// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Thu Jun 27 02:51:32 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383, new_n384, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067_1, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095, new_n1096,
    new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269_1, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333_1, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355, new_n1356,
    new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471_1,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1, new_n2432,
    new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1, new_n2510,
    new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3053, new_n3054, new_n3055, new_n3056, new_n3057,
    new_n3058, new_n3059, new_n3060, new_n3061, new_n3062, new_n3063,
    new_n3064, new_n3065, new_n3066, new_n3067, new_n3068, new_n3069,
    new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074, new_n3075,
    new_n3076, new_n3077, new_n3078, new_n3079, new_n3080, new_n3081,
    new_n3082, new_n3083, new_n3084, new_n3085, new_n3086, new_n3087,
    new_n3088, new_n3089, new_n3090, new_n3091, new_n3092, new_n3093,
    new_n3094, new_n3095, new_n3096, new_n3097, new_n3098, new_n3099,
    new_n3100, new_n3101, new_n3102, new_n3103, new_n3104, new_n3105,
    new_n3106, new_n3107, new_n3108, new_n3109, new_n3110, new_n3111,
    new_n3112, new_n3113, new_n3114, new_n3115, new_n3116, new_n3117,
    new_n3118, new_n3119, new_n3120, new_n3121, new_n3122, new_n3123,
    new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128, new_n3129,
    new_n3130, new_n3131, new_n3132, new_n3133, new_n3134, new_n3135,
    new_n3136, new_n3137, new_n3138, new_n3139, new_n3140, new_n3141,
    new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1, new_n3147,
    new_n3148, new_n3149, new_n3150, new_n3151, new_n3152, new_n3153,
    new_n3154, new_n3155, new_n3156, new_n3157, new_n3158, new_n3159,
    new_n3160, new_n3161, new_n3162, new_n3163, new_n3164, new_n3165,
    new_n3166, new_n3167, new_n3168, new_n3169, new_n3170, new_n3171,
    new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176, new_n3177,
    new_n3178, new_n3179, new_n3180, new_n3181, new_n3182, new_n3183,
    new_n3184, new_n3185, new_n3186, new_n3187, new_n3188, new_n3189,
    new_n3190, new_n3191, new_n3192, new_n3193, new_n3194, new_n3195,
    new_n3196, new_n3197, new_n3198, new_n3199, new_n3200, new_n3201,
    new_n3202, new_n3203, new_n3204, new_n3205, new_n3206, new_n3207,
    new_n3208, new_n3209, new_n3210, new_n3211, new_n3212, new_n3213,
    new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218, new_n3219,
    new_n3220, new_n3221, new_n3222, new_n3223, new_n3224, new_n3225,
    new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1, new_n3231,
    new_n3232, new_n3233, new_n3234, new_n3235, new_n3236, new_n3237,
    new_n3238, new_n3239, new_n3240, new_n3241, new_n3242, new_n3243,
    new_n3244, new_n3245, new_n3246, new_n3247, new_n3248, new_n3249,
    new_n3250, new_n3251, new_n3252, new_n3253, new_n3254, new_n3255,
    new_n3256, new_n3257, new_n3258, new_n3259, new_n3260, new_n3261,
    new_n3262, new_n3263, new_n3264, new_n3265, new_n3266, new_n3267,
    new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1, new_n3273,
    new_n3274, new_n3275, new_n3276, new_n3277, new_n3278, new_n3279,
    new_n3280, new_n3281, new_n3282, new_n3283, new_n3284, new_n3285,
    new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290, new_n3291,
    new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297,
    new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303,
    new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309,
    new_n3310, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321,
    new_n3322, new_n3323, new_n3324, new_n3325, new_n3326, new_n3327,
    new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339_1,
    new_n3340, new_n3341, new_n3342_1, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754_1,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3892, new_n3893,
    new_n3894, new_n3895, new_n3896, new_n3897, new_n3898, new_n3899,
    new_n3900, new_n3901, new_n3902, new_n3903, new_n3904, new_n3905,
    new_n3906, new_n3907, new_n3908, new_n3909, new_n3910, new_n3911,
    new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917,
    new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923,
    new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929,
    new_n3930, new_n3931, new_n3932_1, new_n3933, new_n3934, new_n3935,
    new_n3936, new_n3937, new_n3938, new_n3939, new_n3940, new_n3941,
    new_n3942, new_n3943, new_n3944, new_n3945, new_n3946, new_n3947,
    new_n3948, new_n3949, new_n3950, new_n3951, new_n3952, new_n3953,
    new_n3954, new_n3955, new_n3956, new_n3957, new_n3958, new_n3959,
    new_n3960, new_n3961, new_n3962, new_n3963, new_n3964, new_n3965,
    new_n3966, new_n3967, new_n3968, new_n3969, new_n3970, new_n3971,
    new_n3972, new_n3973, new_n3974, new_n3975, new_n3976, new_n3977,
    new_n3978, new_n3979, new_n3980, new_n3981, new_n3982, new_n3983,
    new_n3984, new_n3985, new_n3986_1, new_n3987, new_n3988, new_n3989,
    new_n3990, new_n3991, new_n3992_1, new_n3993, new_n3994, new_n3995,
    new_n3996, new_n3997, new_n3998, new_n3999, new_n4000, new_n4001,
    new_n4002, new_n4003, new_n4004, new_n4005_1, new_n4006, new_n4007,
    new_n4008, new_n4009, new_n4010, new_n4011, new_n4012, new_n4013,
    new_n4014, new_n4015, new_n4016, new_n4017, new_n4018, new_n4019,
    new_n4020, new_n4021, new_n4022, new_n4023, new_n4024, new_n4025,
    new_n4026, new_n4027, new_n4028, new_n4029, new_n4030, new_n4031,
    new_n4032, new_n4033, new_n4034, new_n4035, new_n4036, new_n4037,
    new_n4038, new_n4039, new_n4040, new_n4041, new_n4042, new_n4043,
    new_n4044, new_n4045, new_n4046, new_n4047, new_n4048, new_n4049,
    new_n4050, new_n4051, new_n4052, new_n4053, new_n4054, new_n4055,
    new_n4056, new_n4057, new_n4058, new_n4059, new_n4060, new_n4061,
    new_n4062, new_n4063, new_n4064, new_n4065, new_n4066, new_n4067,
    new_n4068, new_n4069, new_n4070, new_n4071, new_n4072, new_n4073,
    new_n4074, new_n4075, new_n4076, new_n4077, new_n4078, new_n4079,
    new_n4080, new_n4081, new_n4082, new_n4083, new_n4084, new_n4085,
    new_n4086_1, new_n4087, new_n4088_1, new_n4089, new_n4090, new_n4091,
    new_n4092, new_n4093, new_n4094_1, new_n4095, new_n4096, new_n4097,
    new_n4098, new_n4099, new_n4100, new_n4101, new_n4102, new_n4103,
    new_n4104, new_n4105, new_n4106, new_n4107, new_n4108, new_n4109,
    new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119, new_n4120, new_n4121,
    new_n4122, new_n4123, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141_1, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155_1, new_n4156, new_n4157,
    new_n4158, new_n4159_1, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187_1,
    new_n4188, new_n4189_1, new_n4190_1, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203_1, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4220,
    new_n4222, new_n4223, new_n4224, new_n4225, new_n4226_1, new_n4227,
    new_n4228, new_n4229, new_n4230_1, new_n4231, new_n4232, new_n4233,
    new_n4234, new_n4235, new_n4236, new_n4237, new_n4238, new_n4239,
    new_n4240, new_n4241, new_n4242, new_n4243, new_n4244, new_n4245,
    new_n4246, new_n4247, new_n4248, new_n4249, new_n4250, new_n4251,
    new_n4252, new_n4253, new_n4254, new_n4255, new_n4256, new_n4257,
    new_n4258, new_n4259, new_n4260, new_n4261, new_n4262, new_n4263,
    new_n4264, new_n4265, new_n4266, new_n4267, new_n4268, new_n4269,
    new_n4270, new_n4271, new_n4272, new_n4273, new_n4274, new_n4275,
    new_n4276, new_n4277, new_n4278, new_n4279, new_n4280, new_n4281,
    new_n4282, new_n4283, new_n4284, new_n4285, new_n4286, new_n4287,
    new_n4288, new_n4289, new_n4290, new_n4291, new_n4292, new_n4293,
    new_n4294, new_n4295, new_n4296, new_n4297, new_n4298, new_n4299,
    new_n4300_1, new_n4301, new_n4302, new_n4303, new_n4304, new_n4305,
    new_n4306, new_n4307, new_n4308, new_n4309, new_n4310, new_n4311,
    new_n4312_1, new_n4313, new_n4314, new_n4315, new_n4316, new_n4317,
    new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4324, new_n4325, new_n4326_1, new_n4327, new_n4328, new_n4329,
    new_n4330, new_n4331, new_n4332, new_n4333_1, new_n4334, new_n4335,
    new_n4336, new_n4337, new_n4338, new_n4339, new_n4340, new_n4341,
    new_n4342, new_n4343, new_n4344, new_n4345, new_n4346, new_n4347,
    new_n4348, new_n4349, new_n4350, new_n4351, new_n4352, new_n4353,
    new_n4354, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359,
    new_n4360, new_n4361, new_n4362, new_n4363, new_n4364, new_n4365,
    new_n4366, new_n4367, new_n4368, new_n4369, new_n4370_1, new_n4371,
    new_n4372, new_n4373, new_n4374, new_n4375, new_n4376, new_n4377,
    new_n4378_1, new_n4379, new_n4380, new_n4381, new_n4382, new_n4383,
    new_n4384, new_n4385, new_n4386, new_n4387, new_n4388, new_n4389,
    new_n4390, new_n4391, new_n4392, new_n4393, new_n4394, new_n4395,
    new_n4396, new_n4397_1, new_n4398, new_n4399, new_n4400, new_n4401,
    new_n4402, new_n4403, new_n4404, new_n4405, new_n4406, new_n4407,
    new_n4408, new_n4409, new_n4410, new_n4411, new_n4412, new_n4413,
    new_n4414, new_n4415, new_n4416, new_n4417, new_n4418, new_n4419,
    new_n4420, new_n4421, new_n4422, new_n4423, new_n4424, new_n4425,
    new_n4426, new_n4427, new_n4428, new_n4429, new_n4430, new_n4431,
    new_n4432, new_n4433, new_n4434, new_n4435, new_n4436_1, new_n4437,
    new_n4438, new_n4439, new_n4440, new_n4441, new_n4442, new_n4443,
    new_n4444, new_n4445, new_n4446, new_n4447, new_n4448, new_n4449,
    new_n4450, new_n4451, new_n4452, new_n4453, new_n4454, new_n4455,
    new_n4456, new_n4457, new_n4458, new_n4459, new_n4460, new_n4461,
    new_n4462, new_n4463, new_n4464, new_n4465, new_n4466, new_n4467,
    new_n4468, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473,
    new_n4474, new_n4475, new_n4476, new_n4477, new_n4478, new_n4479,
    new_n4480, new_n4481, new_n4482, new_n4483, new_n4484, new_n4485,
    new_n4486, new_n4487, new_n4488, new_n4489, new_n4490, new_n4491,
    new_n4492, new_n4493, new_n4494, new_n4495, new_n4496, new_n4497,
    new_n4498, new_n4499_1, new_n4500, new_n4501, new_n4502, new_n4503,
    new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509,
    new_n4510, new_n4511, new_n4512, new_n4513, new_n4514, new_n4515,
    new_n4516_1, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521,
    new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527,
    new_n4528, new_n4529, new_n4530, new_n4531, new_n4532, new_n4533,
    new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539,
    new_n4540, new_n4541, new_n4542, new_n4543, new_n4544, new_n4545,
    new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551,
    new_n4552, new_n4553_1, new_n4554, new_n4555, new_n4556, new_n4557,
    new_n4558, new_n4559, new_n4560, new_n4561, new_n4562, new_n4563,
    new_n4564, new_n4565, new_n4566, new_n4567, new_n4568, new_n4569,
    new_n4570, new_n4571, new_n4572, new_n4573, new_n4574, new_n4575,
    new_n4576, new_n4577, new_n4578, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599,
    new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605,
    new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611,
    new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617,
    new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623,
    new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634_1, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686_1, new_n4687, new_n4688, new_n4689_1,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733_1, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757_1, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805_1, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817_1, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826_1, new_n4827,
    new_n4828_1, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212_1,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314_1,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1, new_n5320_1,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5497, new_n5498, new_n5499, new_n5500, new_n5501,
    new_n5502, new_n5503, new_n5504, new_n5505, new_n5506, new_n5507,
    new_n5508, new_n5509, new_n5510, new_n5511, new_n5512, new_n5513,
    new_n5514, new_n5515, new_n5516, new_n5517, new_n5518, new_n5519,
    new_n5520, new_n5521, new_n5522, new_n5523, new_n5524, new_n5525,
    new_n5526, new_n5527, new_n5528, new_n5529, new_n5530, new_n5531,
    new_n5532, new_n5533, new_n5534, new_n5535, new_n5536, new_n5537,
    new_n5538, new_n5539, new_n5540, new_n5541, new_n5542, new_n5543,
    new_n5544, new_n5545, new_n5546, new_n5547, new_n5548, new_n5549,
    new_n5550, new_n5551, new_n5552, new_n5553, new_n5554, new_n5555,
    new_n5556, new_n5557, new_n5558, new_n5559, new_n5560, new_n5561,
    new_n5562, new_n5563, new_n5564, new_n5565, new_n5566, new_n5567,
    new_n5568, new_n5569, new_n5570, new_n5571, new_n5572, new_n5573,
    new_n5574, new_n5575, new_n5576, new_n5577, new_n5578, new_n5579_1,
    new_n5580, new_n5581, new_n5582, new_n5583, new_n5584, new_n5585,
    new_n5586, new_n5587, new_n5588, new_n5589, new_n5590, new_n5591,
    new_n5592, new_n5593, new_n5594, new_n5595, new_n5596, new_n5597,
    new_n5598, new_n5599, new_n5600, new_n5601, new_n5602, new_n5603,
    new_n5604, new_n5605, new_n5606, new_n5607, new_n5608, new_n5609,
    new_n5610, new_n5611, new_n5612, new_n5613, new_n5614, new_n5615,
    new_n5616, new_n5617, new_n5618, new_n5619, new_n5620, new_n5621,
    new_n5622, new_n5623, new_n5624, new_n5625, new_n5626, new_n5627,
    new_n5628, new_n5629, new_n5630, new_n5631, new_n5632, new_n5633,
    new_n5634, new_n5635, new_n5636, new_n5637, new_n5638, new_n5639,
    new_n5640, new_n5641_1, new_n5642, new_n5643, new_n5644, new_n5645_1,
    new_n5646, new_n5647, new_n5648, new_n5649, new_n5650, new_n5651,
    new_n5652, new_n5653, new_n5654, new_n5655, new_n5656, new_n5657,
    new_n5658, new_n5659, new_n5660, new_n5661, new_n5662, new_n5663,
    new_n5664, new_n5665, new_n5666, new_n5667, new_n5668, new_n5669,
    new_n5670_1, new_n5671, new_n5672, new_n5673, new_n5674, new_n5675,
    new_n5676, new_n5677, new_n5678, new_n5679, new_n5680, new_n5681,
    new_n5682, new_n5683, new_n5684, new_n5685, new_n5686, new_n5687,
    new_n5688, new_n5689, new_n5690, new_n5691, new_n5692, new_n5693_1,
    new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698, new_n5699,
    new_n5700, new_n5701, new_n5702, new_n5703, new_n5704, new_n5705,
    new_n5706, new_n5707, new_n5708, new_n5709, new_n5710, new_n5711,
    new_n5712, new_n5713, new_n5714, new_n5715, new_n5716, new_n5717,
    new_n5718, new_n5719, new_n5720, new_n5721, new_n5722, new_n5723,
    new_n5724, new_n5725, new_n5726, new_n5727, new_n5728, new_n5729,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759,
    new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777,
    new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783,
    new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789,
    new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795,
    new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814_1,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857_1, new_n5858, new_n5859, new_n5860_1, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934_1,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964_1,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5994, new_n5995,
    new_n5996, new_n5997, new_n5998, new_n5999, new_n6000, new_n6001,
    new_n6002, new_n6003, new_n6004, new_n6005, new_n6006, new_n6007,
    new_n6008, new_n6009, new_n6010, new_n6011, new_n6012, new_n6013,
    new_n6014, new_n6015, new_n6016_1, new_n6017, new_n6018, new_n6019,
    new_n6020, new_n6021, new_n6022, new_n6023, new_n6024, new_n6025,
    new_n6026, new_n6027, new_n6030, new_n6031, new_n6032, new_n6033,
    new_n6034, new_n6035, new_n6036, new_n6037, new_n6038_1, new_n6039,
    new_n6040, new_n6041, new_n6042, new_n6043, new_n6044, new_n6045,
    new_n6046, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051,
    new_n6052, new_n6053, new_n6054, new_n6055, new_n6056, new_n6057,
    new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063,
    new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069,
    new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075,
    new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081,
    new_n6082, new_n6083, new_n6084, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089_1, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104, new_n6105,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126_1, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153,
    new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159,
    new_n6160, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165,
    new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171,
    new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189,
    new_n6190, new_n6191, new_n6192_1, new_n6193, new_n6194, new_n6195,
    new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201,
    new_n6202, new_n6203, new_n6204, new_n6205, new_n6206, new_n6207,
    new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213,
    new_n6214, new_n6215, new_n6216, new_n6217, new_n6218, new_n6219,
    new_n6220, new_n6221, new_n6222, new_n6223, new_n6224, new_n6225,
    new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231,
    new_n6232, new_n6233, new_n6234, new_n6235, new_n6236, new_n6237,
    new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243,
    new_n6244, new_n6245, new_n6246, new_n6247, new_n6248, new_n6249,
    new_n6250, new_n6251, new_n6252, new_n6253, new_n6254_1, new_n6255,
    new_n6256, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261,
    new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267,
    new_n6268, new_n6269, new_n6270, new_n6271, new_n6272, new_n6273_1,
    new_n6274, new_n6275, new_n6276, new_n6277, new_n6278, new_n6279,
    new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285,
    new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291,
    new_n6292, new_n6293, new_n6294_1, new_n6295, new_n6296, new_n6297,
    new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303,
    new_n6304, new_n6305, new_n6306, new_n6307, new_n6308, new_n6309,
    new_n6310, new_n6311, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323, new_n6324, new_n6325, new_n6326, new_n6327,
    new_n6328, new_n6329, new_n6330, new_n6331, new_n6332, new_n6333,
    new_n6334, new_n6335, new_n6336, new_n6337, new_n6338, new_n6339,
    new_n6340, new_n6341, new_n6342, new_n6343, new_n6344, new_n6345,
    new_n6346, new_n6347, new_n6348, new_n6349, new_n6350, new_n6351,
    new_n6352, new_n6353, new_n6354, new_n6355, new_n6356, new_n6357,
    new_n6358_1, new_n6359_1, new_n6360, new_n6361, new_n6362, new_n6363,
    new_n6364, new_n6365, new_n6366, new_n6367, new_n6368, new_n6369,
    new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375,
    new_n6376, new_n6377, new_n6378, new_n6379, new_n6380, new_n6381,
    new_n6382, new_n6383, new_n6384, new_n6385, new_n6386, new_n6387,
    new_n6388, new_n6389, new_n6390, new_n6391, new_n6392, new_n6393,
    new_n6394, new_n6395, new_n6396, new_n6397, new_n6398, new_n6399,
    new_n6400, new_n6401, new_n6402, new_n6403, new_n6404, new_n6405,
    new_n6406, new_n6407, new_n6408, new_n6409, new_n6410, new_n6411,
    new_n6412, new_n6413, new_n6414, new_n6415, new_n6416, new_n6417,
    new_n6418, new_n6419, new_n6420, new_n6421, new_n6422, new_n6423,
    new_n6424, new_n6425, new_n6426, new_n6427, new_n6428, new_n6429_1,
    new_n6430, new_n6431_1, new_n6432, new_n6433, new_n6434, new_n6435,
    new_n6436, new_n6437, new_n6438, new_n6439, new_n6440, new_n6441_1,
    new_n6442, new_n6443, new_n6444, new_n6445_1, new_n6446, new_n6447,
    new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453,
    new_n6454, new_n6455, new_n6456, new_n6457, new_n6458, new_n6459,
    new_n6460, new_n6461, new_n6462, new_n6463, new_n6464, new_n6465,
    new_n6466, new_n6467, new_n6468, new_n6469, new_n6470, new_n6471,
    new_n6472, new_n6473, new_n6474, new_n6475, new_n6476, new_n6477,
    new_n6478, new_n6479, new_n6480, new_n6481, new_n6484, new_n6485,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502, new_n6503,
    new_n6504, new_n6505, new_n6506, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513, new_n6514, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556, new_n6557,
    new_n6558, new_n6559, new_n6560, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576, new_n6577, new_n6578_1, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587,
    new_n6588, new_n6589, new_n6590, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604_1, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611_1,
    new_n6612, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629,
    new_n6630, new_n6631, new_n6632, new_n6633, new_n6634, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6645_1, new_n6646, new_n6647,
    new_n6648, new_n6649, new_n6650, new_n6651, new_n6652, new_n6653,
    new_n6654, new_n6655, new_n6656, new_n6657, new_n6658, new_n6659,
    new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665,
    new_n6666, new_n6667, new_n6668, new_n6669, new_n6670, new_n6671,
    new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684, new_n6685, new_n6686, new_n6687_1, new_n6688, new_n6689_1,
    new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703_1, new_n6704, new_n6705, new_n6706, new_n6707,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742_1, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770_1, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776_1, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797_1,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806_1, new_n6807, new_n6808, new_n6809_1,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822_1, new_n6823, new_n6824, new_n6825, new_n6826_1, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6860_1, new_n6861, new_n6862, new_n6863,
    new_n6864, new_n6865, new_n6866, new_n6867, new_n6868, new_n6869,
    new_n6870, new_n6871, new_n6872, new_n6873, new_n6874, new_n6875,
    new_n6876, new_n6877_1, new_n6878, new_n6879, new_n6880, new_n6881,
    new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887,
    new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893,
    new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899,
    new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905,
    new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911,
    new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941,
    new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947,
    new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986_1, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013,
    new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019,
    new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025,
    new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031,
    new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7132,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159_1, new_n7160_1, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193_1,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265_1,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270_1, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294_1, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320_1, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523_1,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7805, new_n7806, new_n7807, new_n7808, new_n7809,
    new_n7810, new_n7811, new_n7812, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946_1,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964,
    new_n7965_1, new_n7966_1, new_n7967, new_n7968, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981_1, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028_1, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065_1, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100_1, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138_1,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202_1, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236_1, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276_1,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303_1, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336_1,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384_1,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398_1, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433_1, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476_1, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595_1, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665_1, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717_1,
    new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759_1,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819_1,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927,
    new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933,
    new_n8934, new_n8935, new_n8936, new_n8937, new_n8938, new_n8939,
    new_n8940, new_n8941, new_n8942, new_n8943, new_n8944, new_n8945,
    new_n8946, new_n8947, new_n8948, new_n8949, new_n8950, new_n8951,
    new_n8952, new_n8953, new_n8954, new_n8955, new_n8956, new_n8957,
    new_n8958, new_n8959, new_n8960, new_n8961, new_n8962, new_n8963,
    new_n8964, new_n8965, new_n8966, new_n8967, new_n8968, new_n8969,
    new_n8970, new_n8971, new_n8972, new_n8973, new_n8974, new_n8975,
    new_n8976, new_n8977, new_n8978, new_n8979, new_n8980, new_n8981,
    new_n8982, new_n8983, new_n8984, new_n8985, new_n8986, new_n8987,
    new_n8988, new_n8989, new_n8990, new_n8991, new_n8992, new_n8993,
    new_n8994, new_n8995, new_n8996, new_n8997, new_n8998, new_n8999,
    new_n9000, new_n9001, new_n9002, new_n9003, new_n9004, new_n9005,
    new_n9006, new_n9007, new_n9008, new_n9009, new_n9010, new_n9011,
    new_n9012, new_n9013, new_n9014, new_n9015, new_n9016, new_n9017,
    new_n9018, new_n9019, new_n9020, new_n9021, new_n9022, new_n9023,
    new_n9024, new_n9025, new_n9026, new_n9027, new_n9028, new_n9029,
    new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035,
    new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041,
    new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047,
    new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053,
    new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059,
    new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065,
    new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071,
    new_n9072, new_n9073, new_n9074, new_n9075, new_n9076, new_n9077,
    new_n9078, new_n9079, new_n9080_1, new_n9081, new_n9082, new_n9083,
    new_n9084, new_n9085, new_n9086, new_n9087, new_n9088, new_n9089,
    new_n9090, new_n9091, new_n9092, new_n9093, new_n9094, new_n9095,
    new_n9096, new_n9097, new_n9098, new_n9099, new_n9100, new_n9101,
    new_n9102, new_n9103, new_n9104, new_n9105, new_n9106, new_n9107,
    new_n9108, new_n9109, new_n9110, new_n9111_1, new_n9112, new_n9113,
    new_n9114, new_n9115, new_n9116, new_n9117, new_n9118, new_n9119,
    new_n9120, new_n9121, new_n9122, new_n9123, new_n9124, new_n9125,
    new_n9126, new_n9127, new_n9128, new_n9129, new_n9130, new_n9131,
    new_n9132, new_n9133, new_n9134, new_n9135, new_n9136, new_n9137_1,
    new_n9138, new_n9139, new_n9140, new_n9141, new_n9142, new_n9143,
    new_n9144, new_n9145, new_n9146, new_n9147, new_n9148, new_n9149,
    new_n9150, new_n9151, new_n9152, new_n9153, new_n9154, new_n9155,
    new_n9156, new_n9157, new_n9158, new_n9159, new_n9160, new_n9161,
    new_n9162, new_n9163, new_n9164, new_n9165, new_n9166, new_n9167,
    new_n9168, new_n9169, new_n9170, new_n9171, new_n9172, new_n9173,
    new_n9174, new_n9175, new_n9176, new_n9177, new_n9178, new_n9179,
    new_n9180, new_n9181, new_n9182, new_n9183, new_n9184, new_n9185,
    new_n9186, new_n9187, new_n9188, new_n9189_1, new_n9190, new_n9191,
    new_n9192, new_n9193, new_n9194, new_n9195_1, new_n9196, new_n9197,
    new_n9198, new_n9199, new_n9200, new_n9201, new_n9202, new_n9203,
    new_n9204, new_n9205, new_n9206, new_n9207, new_n9208, new_n9209,
    new_n9210, new_n9211, new_n9212, new_n9213, new_n9214, new_n9215,
    new_n9216, new_n9217, new_n9218, new_n9219, new_n9220, new_n9221,
    new_n9222, new_n9223, new_n9224, new_n9225, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241_1, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387_1, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400_1, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9456, new_n9457_1,
    new_n9458, new_n9459, new_n9460, new_n9461, new_n9462, new_n9463,
    new_n9464, new_n9465, new_n9466, new_n9467, new_n9468, new_n9469,
    new_n9470, new_n9471, new_n9472, new_n9473, new_n9474, new_n9475,
    new_n9476, new_n9477, new_n9478, new_n9479, new_n9480, new_n9481,
    new_n9482, new_n9483, new_n9484, new_n9485, new_n9486, new_n9487,
    new_n9488, new_n9489, new_n9490, new_n9491, new_n9492, new_n9493,
    new_n9494, new_n9495, new_n9496, new_n9497, new_n9498, new_n9499,
    new_n9500, new_n9501, new_n9502, new_n9503, new_n9504, new_n9505,
    new_n9506, new_n9507, new_n9508, new_n9509, new_n9510, new_n9511,
    new_n9512, new_n9513, new_n9514, new_n9515, new_n9516, new_n9517,
    new_n9518, new_n9519, new_n9520, new_n9521, new_n9522, new_n9523,
    new_n9524, new_n9525, new_n9526, new_n9527, new_n9528, new_n9529,
    new_n9530, new_n9531, new_n9532, new_n9533, new_n9534, new_n9535,
    new_n9536, new_n9537, new_n9538, new_n9539, new_n9540, new_n9541,
    new_n9542, new_n9543, new_n9544, new_n9545, new_n9546, new_n9547,
    new_n9548, new_n9549, new_n9550, new_n9551, new_n9552, new_n9553,
    new_n9554, new_n9555, new_n9556, new_n9557, new_n9558, new_n9559,
    new_n9560, new_n9561, new_n9562, new_n9563, new_n9564, new_n9565,
    new_n9566, new_n9567, new_n9568, new_n9569, new_n9570, new_n9571_1,
    new_n9572, new_n9573, new_n9574, new_n9575, new_n9576, new_n9577,
    new_n9578_1, new_n9579, new_n9580, new_n9581, new_n9582, new_n9583_1,
    new_n9584, new_n9585, new_n9586, new_n9587, new_n9588, new_n9589,
    new_n9590, new_n9591, new_n9592, new_n9593, new_n9594, new_n9595,
    new_n9596, new_n9597, new_n9598, new_n9599, new_n9600, new_n9601,
    new_n9602, new_n9603, new_n9604, new_n9605, new_n9606, new_n9607,
    new_n9608, new_n9609, new_n9610, new_n9611, new_n9612, new_n9613,
    new_n9614, new_n9615, new_n9616, new_n9617, new_n9618, new_n9619,
    new_n9620, new_n9621, new_n9622, new_n9623, new_n9624, new_n9625,
    new_n9626, new_n9627, new_n9628, new_n9629, new_n9630, new_n9631,
    new_n9632, new_n9633, new_n9634, new_n9635, new_n9636, new_n9637_1,
    new_n9638, new_n9639, new_n9640_1, new_n9641, new_n9642, new_n9643,
    new_n9644, new_n9645, new_n9646, new_n9647, new_n9648, new_n9649,
    new_n9650, new_n9651, new_n9652, new_n9653, new_n9654, new_n9655,
    new_n9656, new_n9657, new_n9658, new_n9659, new_n9660, new_n9661,
    new_n9662, new_n9663, new_n9664, new_n9665, new_n9666, new_n9667,
    new_n9668, new_n9669, new_n9670, new_n9671, new_n9672, new_n9673,
    new_n9674, new_n9675, new_n9676, new_n9677, new_n9678, new_n9679,
    new_n9680, new_n9681, new_n9682, new_n9683, new_n9684, new_n9685,
    new_n9686, new_n9687, new_n9688, new_n9689, new_n9690, new_n9691,
    new_n9692, new_n9693, new_n9694, new_n9695, new_n9696, new_n9697,
    new_n9698, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703,
    new_n9704, new_n9705, new_n9706_1, new_n9707, new_n9708, new_n9709,
    new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715,
    new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725_1, new_n9726, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9738, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753, new_n9754, new_n9755, new_n9756_1, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763_1,
    new_n9764, new_n9765, new_n9766, new_n9767_1, new_n9768, new_n9769,
    new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799,
    new_n9800, new_n9801, new_n9802, new_n9803, new_n9804, new_n9805,
    new_n9806, new_n9807, new_n9808, new_n9809, new_n9810, new_n9811,
    new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817,
    new_n9818, new_n9819, new_n9820_1, new_n9821, new_n9822, new_n9823,
    new_n9824, new_n9825, new_n9826, new_n9827, new_n9828, new_n9829,
    new_n9830, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835,
    new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841,
    new_n9842, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889,
    new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920_1, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938_1, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956_1, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10006, new_n10007, new_n10008, new_n10009,
    new_n10010, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015,
    new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10022_1, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038,
    new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044,
    new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050,
    new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056,
    new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080,
    new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086,
    new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174_1, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217_1, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223_1, new_n10224, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10252, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259,
    new_n10260, new_n10261, new_n10262, new_n10263, new_n10264, new_n10265,
    new_n10266, new_n10267, new_n10268, new_n10269, new_n10270, new_n10271,
    new_n10272, new_n10273, new_n10274, new_n10275, new_n10276, new_n10277,
    new_n10278_1, new_n10279, new_n10280, new_n10281, new_n10282,
    new_n10283, new_n10284, new_n10285, new_n10286, new_n10287, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300,
    new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306,
    new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312,
    new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318,
    new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326, new_n10327_1, new_n10328, new_n10329,
    new_n10330, new_n10331, new_n10332, new_n10333, new_n10334, new_n10335,
    new_n10336, new_n10337, new_n10338, new_n10339, new_n10340, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345, new_n10346, new_n10347,
    new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10382, new_n10383, new_n10384,
    new_n10385, new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391_1, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439_1, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451_1, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476_1,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510_1, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545_1, new_n10546,
    new_n10547_1, new_n10548, new_n10549, new_n10550, new_n10551,
    new_n10552, new_n10553, new_n10554, new_n10555, new_n10556, new_n10557,
    new_n10558, new_n10559, new_n10560, new_n10561, new_n10562, new_n10563,
    new_n10564, new_n10565, new_n10566, new_n10567, new_n10568, new_n10569,
    new_n10570, new_n10571, new_n10572, new_n10573, new_n10574, new_n10575,
    new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589_1, new_n10590, new_n10591, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616,
    new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622,
    new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628,
    new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644_1, new_n10645,
    new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651,
    new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678_1, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685_1,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695_1, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789_1, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848_1, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898_1, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913_1,
    new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10928_1, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949_1, new_n10950, new_n10951, new_n10952, new_n10953,
    new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959,
    new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965_1, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10988, new_n10989, new_n10990_1, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023_1, new_n11024, new_n11025, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045,
    new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051,
    new_n11052, new_n11053, new_n11054, new_n11055, new_n11056, new_n11057,
    new_n11058, new_n11059, new_n11060, new_n11061, new_n11062, new_n11063,
    new_n11064, new_n11065, new_n11066, new_n11067, new_n11068, new_n11069,
    new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11095, new_n11096, new_n11097, new_n11098, new_n11099,
    new_n11100, new_n11101, new_n11102, new_n11103, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120, new_n11121, new_n11122, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129,
    new_n11130, new_n11131, new_n11132, new_n11133, new_n11134, new_n11135,
    new_n11136, new_n11137, new_n11138, new_n11139, new_n11140, new_n11141,
    new_n11142, new_n11143, new_n11144, new_n11145, new_n11146, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153_1, new_n11154, new_n11155, new_n11156, new_n11157,
    new_n11158, new_n11159, new_n11160, new_n11161, new_n11162, new_n11163,
    new_n11164, new_n11165, new_n11166, new_n11167, new_n11168, new_n11169,
    new_n11170, new_n11171, new_n11172, new_n11173, new_n11174, new_n11175,
    new_n11176, new_n11177, new_n11178, new_n11179, new_n11180, new_n11181,
    new_n11182, new_n11183, new_n11184, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201, new_n11202, new_n11203, new_n11204, new_n11205,
    new_n11206, new_n11207, new_n11208, new_n11213, new_n11216_1,
    new_n11218, new_n11220, new_n11223, new_n11225, new_n11226, new_n11227,
    new_n11228, new_n11229, new_n11230, new_n11231, new_n11232, new_n11233,
    new_n11234, new_n11235, new_n11236, new_n11237, new_n11238, new_n11239,
    new_n11240, new_n11241, new_n11242, new_n11243, new_n11244, new_n11245,
    new_n11246, new_n11247, new_n11248, new_n11249, new_n11250, new_n11251,
    new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257_1, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311_1, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326_1, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407_1,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423_1, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478_1, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536_1, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11554,
    new_n11555, new_n11556, new_n11557, new_n11558, new_n11559, new_n11560,
    new_n11561, new_n11562, new_n11563, new_n11564, new_n11565, new_n11566,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584,
    new_n11585, new_n11586, new_n11587, new_n11588, new_n11589, new_n11590,
    new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596,
    new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602,
    new_n11603, new_n11604, new_n11605, new_n11606, new_n11607, new_n11608,
    new_n11609, new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615, new_n11616, new_n11617, new_n11618, new_n11619, new_n11620,
    new_n11621, new_n11622, new_n11623, new_n11624, new_n11625, new_n11626,
    new_n11627, new_n11628, new_n11629, new_n11630, new_n11631, new_n11632,
    new_n11633, new_n11634, new_n11635, new_n11636, new_n11637, new_n11638,
    new_n11639, new_n11640, new_n11641, new_n11642, new_n11643, new_n11644,
    new_n11645, new_n11646, new_n11647, new_n11648, new_n11649, new_n11650,
    new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656,
    new_n11657, new_n11658, new_n11659, new_n11660, new_n11661,
    new_n11662_1, new_n11663, new_n11664, new_n11665, new_n11666,
    new_n11667, new_n11668, new_n11669, new_n11670, new_n11671, new_n11672,
    new_n11673, new_n11674, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682, new_n11683, new_n11684,
    new_n11685, new_n11686, new_n11687, new_n11688, new_n11689, new_n11690,
    new_n11691, new_n11692, new_n11693, new_n11694, new_n11695, new_n11696,
    new_n11697, new_n11698, new_n11699, new_n11700, new_n11701, new_n11702,
    new_n11703, new_n11704, new_n11705, new_n11706, new_n11707_1,
    new_n11708, new_n11709, new_n11710, new_n11711, new_n11712, new_n11713,
    new_n11714, new_n11715, new_n11716, new_n11717, new_n11718, new_n11719,
    new_n11720, new_n11721, new_n11722, new_n11723, new_n11724, new_n11725,
    new_n11726, new_n11727, new_n11728_1, new_n11729, new_n11730,
    new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11745, new_n11747, new_n11749,
    new_n11751, new_n11752, new_n11753, new_n11754, new_n11755_1,
    new_n11756, new_n11757_1, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780_1, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11790, new_n11791_1, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11817, new_n11818,
    new_n11819, new_n11820, new_n11821_1, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876_1,
    new_n11877_1, new_n11878, new_n11879, new_n11880, new_n11881,
    new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887,
    new_n11888, new_n11889, new_n11890, new_n11891, new_n11892_1,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917_1, new_n11918, new_n11919_1, new_n11920, new_n11921,
    new_n11922_1, new_n11923, new_n11924, new_n11925, new_n11926,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956,
    new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962,
    new_n11963, new_n11964, new_n11965, new_n11966, new_n11967_1,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999_1, new_n12000_1, new_n12001, new_n12002,
    new_n12003, new_n12004, new_n12005_1, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014_1, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020_1, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025_1, new_n12026, new_n12027, new_n12028,
    new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044_1, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069_1, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076_1, new_n12077, new_n12078,
    new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12108, new_n12110, new_n12115,
    new_n12119, new_n12122, new_n12123, new_n12124, new_n12125, new_n12126,
    new_n12127, new_n12128, new_n12129, new_n12130, new_n12131, new_n12132,
    new_n12133, new_n12134, new_n12135, new_n12136, new_n12137, new_n12138,
    new_n12139, new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145_1, new_n12146, new_n12147, new_n12148, new_n12149,
    new_n12150, new_n12151, new_n12152, new_n12153, new_n12154, new_n12155,
    new_n12156, new_n12157, new_n12158, new_n12159, new_n12160, new_n12161,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173,
    new_n12174, new_n12175, new_n12176, new_n12177, new_n12178, new_n12179,
    new_n12180, new_n12181, new_n12182, new_n12183, new_n12184, new_n12185,
    new_n12186, new_n12187, new_n12188, new_n12189, new_n12190, new_n12191,
    new_n12192, new_n12193, new_n12194, new_n12195, new_n12196, new_n12197,
    new_n12198, new_n12199, new_n12200, new_n12201, new_n12202, new_n12203,
    new_n12204, new_n12205, new_n12206, new_n12207, new_n12208, new_n12209,
    new_n12210, new_n12211, new_n12212, new_n12213, new_n12214, new_n12215,
    new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221_1, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247_1, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299_1, new_n12300, new_n12301,
    new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12308,
    new_n12310, new_n12311, new_n12312, new_n12313, new_n12314, new_n12315,
    new_n12316, new_n12317, new_n12318, new_n12319, new_n12320, new_n12321,
    new_n12322, new_n12323, new_n12324, new_n12325, new_n12326, new_n12327,
    new_n12328, new_n12329, new_n12330, new_n12331, new_n12332, new_n12333,
    new_n12334, new_n12335, new_n12336, new_n12337, new_n12338, new_n12339,
    new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12354, new_n12355, new_n12356, new_n12357,
    new_n12358, new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364, new_n12365, new_n12366, new_n12367, new_n12368, new_n12369,
    new_n12370, new_n12371, new_n12372, new_n12373, new_n12374, new_n12375,
    new_n12376, new_n12377, new_n12378, new_n12379, new_n12380, new_n12381,
    new_n12382, new_n12383, new_n12384, new_n12385, new_n12386, new_n12387,
    new_n12388, new_n12389, new_n12390, new_n12391_1, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404,
    new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444_1, new_n12445,
    new_n12446, new_n12447, new_n12448, new_n12449, new_n12450, new_n12451,
    new_n12452, new_n12453, new_n12454, new_n12455, new_n12456, new_n12457,
    new_n12458, new_n12459, new_n12460, new_n12461, new_n12462, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467, new_n12468, new_n12469,
    new_n12470, new_n12471, new_n12472, new_n12473, new_n12474, new_n12475,
    new_n12476, new_n12477, new_n12478, new_n12479, new_n12480, new_n12481,
    new_n12482, new_n12483, new_n12484, new_n12485, new_n12486, new_n12487,
    new_n12488, new_n12489_1, new_n12490, new_n12491, new_n12492,
    new_n12493, new_n12500, new_n12502, new_n12503, new_n12505, new_n12508,
    new_n12510, new_n12511_1, new_n12512, new_n12513, new_n12514,
    new_n12515, new_n12516, new_n12517, new_n12518, new_n12519, new_n12520,
    new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526,
    new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544,
    new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550,
    new_n12551, new_n12552, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561, new_n12562,
    new_n12563, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591_1,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626, new_n12627,
    new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648_1, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12695,
    new_n12699, new_n12702, new_n12707, new_n12708, new_n12709_1,
    new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715,
    new_n12716, new_n12717, new_n12718, new_n12719, new_n12720_1,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753_1, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777_1, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807_1,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12896, new_n12899, new_n12901, new_n12903,
    new_n12906, new_n12908;
nand_5 g00000(n6687, n6038, new_n377);
not_8  g00001(new_n377, new_n378);
nand_5 g00002(n8336, n7354, new_n379);
nand_5 g00003(n11222, n8028, new_n380);
nand_5 g00004(n12069, n1564, new_n381_1);
xor_4  g00005(new_n381_1, new_n380, new_n382);
not_8  g00006(new_n382, new_n383);
xor_4  g00007(new_n383, new_n379, new_n384);
xor_4  g00008(new_n384, new_n378, n112);
nand_5 g00009(n12720, n4312, new_n386);
nand_5 g00010(n12025, n6038, new_n387);
nand_5 g00011(n12705, n2509, new_n388);
xor_4  g00012(new_n388, new_n387, new_n389);
not_8  g00013(new_n389, new_n390);
xor_4  g00014(new_n390, new_n386, new_n391);
nand_5 g00015(n12705, n6038, new_n392);
nand_5 g00016(n12720, n1097, new_n393);
and_5  g00017(new_n393, new_n392, new_n394);
nand_5 g00018(n4312, n2509, new_n395);
not_8  g00019(new_n395, new_n396);
xor_4  g00020(new_n393, new_n392, new_n397_1);
not_8  g00021(new_n397_1, new_n398);
nor_5  g00022(new_n398, new_n396, new_n399);
or_5   g00023(new_n399, new_n394, new_n400);
not_8  g00024(new_n400, new_n401);
xor_4  g00025(new_n401, new_n391, new_n402);
nand_5 g00026(n2508, n1097, new_n403);
nand_5 g00027(n5964, n2585, new_n404);
xor_4  g00028(new_n404, new_n403, new_n405_1);
xor_4  g00029(new_n405_1, new_n402, new_n406);
nand_5 g00030(n5964, n2508, new_n407);
xor_4  g00031(new_n398, new_n396, new_n408);
and_5  g00032(new_n408, new_n407, new_n409);
xor_4  g00033(new_n408, new_n407, new_n410);
not_8  g00034(new_n410, new_n411);
nand_5 g00035(n6038, n4312, new_n412);
nand_5 g00036(n12720, n5964, new_n413);
and_5  g00037(new_n413, new_n412, new_n414);
nor_5  g00038(new_n413, new_n412, new_n415);
nand_5 g00039(n2509, n1097, new_n416);
not_8  g00040(new_n416, new_n417);
nor_5  g00041(new_n417, new_n415, new_n418);
nor_5  g00042(new_n418, new_n414, new_n419);
nor_5  g00043(new_n419, new_n411, new_n420);
or_5   g00044(new_n420, new_n409, new_n421);
not_8  g00045(new_n421, new_n422);
xor_4  g00046(new_n422, new_n406, new_n423);
nand_5 g00047(n5305, n2585, new_n424);
not_8  g00048(new_n424, new_n425);
xor_4  g00049(new_n419, new_n411, new_n426);
not_8  g00050(new_n426, new_n427);
nor_5  g00051(new_n427, new_n425, new_n428);
xor_4  g00052(new_n427, new_n425, new_n429);
nand_5 g00053(n5305, n2508, new_n430);
nand_5 g00054(n6038, n1097, new_n431);
nand_5 g00055(n12720, n5305, new_n432);
nor_5  g00056(new_n432, new_n431, new_n433);
and_5  g00057(new_n432, new_n431, new_n434);
nand_5 g00058(n5964, n2509, new_n435);
or_5   g00059(new_n435, new_n434, new_n436);
not_8  g00060(new_n436, new_n437);
nor_5  g00061(new_n437, new_n433, new_n438);
nor_5  g00062(new_n438, new_n430, new_n439);
xor_4  g00063(new_n438, new_n430, new_n440);
xor_4  g00064(new_n413, new_n412, new_n441);
xor_4  g00065(new_n441, new_n417, new_n442);
and_5  g00066(new_n442, new_n440, new_n443);
or_5   g00067(new_n443, new_n439, new_n444);
not_8  g00068(new_n444, new_n445);
and_5  g00069(new_n445, new_n429, new_n446);
or_5   g00070(new_n446, new_n428, new_n447_1);
not_8  g00071(new_n447_1, new_n448);
nand_5 g00072(new_n448, new_n423, new_n449);
nor_5  g00073(new_n390, new_n386, new_n450);
and_5  g00074(new_n401, new_n391, new_n451);
or_5   g00075(new_n451, new_n450, new_n452);
not_8  g00076(new_n452, new_n453);
nand_5 g00077(n5964, n4005, new_n454);
nand_5 g00078(n2585, n1097, new_n455);
nand_5 g00079(n12706, n5305, new_n456);
xor_4  g00080(new_n456, new_n455, new_n457);
xor_4  g00081(new_n457, new_n454, new_n458);
xor_4  g00082(new_n458, new_n453, new_n459);
or_5   g00083(new_n388, new_n387, new_n460);
not_8  g00084(new_n460, new_n461);
nand_5 g00085(n4312, n2508, new_n462);
not_8  g00086(new_n462, new_n463);
xor_4  g00087(new_n463, new_n461, new_n464);
nand_5 g00088(n12025, n2509, new_n465);
nand_5 g00089(n12720, n12705, new_n466);
nand_5 g00090(n11257, n6038, new_n467);
xor_4  g00091(new_n467, new_n466, new_n468);
not_8  g00092(new_n468, new_n469);
xor_4  g00093(new_n469, new_n465, new_n470);
xor_4  g00094(new_n470, new_n464, new_n471);
xor_4  g00095(new_n471, new_n459, new_n472);
not_8  g00096(new_n472, new_n473);
and_5  g00097(new_n405_1, new_n402, new_n474);
or_5   g00098(new_n404, new_n403, new_n475);
nand_5 g00099(new_n422, new_n406, new_n476);
xor_4  g00100(new_n476, new_n475, new_n477);
nor_5  g00101(new_n477, new_n474, new_n478);
xor_4  g00102(new_n478, new_n473, new_n479);
not_8  g00103(new_n479, new_n480);
xor_4  g00104(new_n480, new_n449, new_n481);
not_8  g00105(new_n481, new_n482);
nand_5 g00106(n5305, n4005, new_n483);
not_8  g00107(new_n483, new_n484);
xor_4  g00108(new_n448, new_n423, new_n485);
and_5  g00109(new_n485, new_n484, new_n486);
nor_5  g00110(new_n485, new_n484, new_n487);
xor_4  g00111(new_n442, new_n440, new_n488);
not_8  g00112(new_n488, new_n489);
xor_4  g00113(new_n432, new_n431, new_n490);
nand_5 g00114(n6038, n5964, new_n491);
nand_5 g00115(n5305, n2509, new_n492);
or_5   g00116(new_n492, new_n491, new_n493);
or_5   g00117(new_n493, new_n490, new_n494);
or_5   g00118(new_n494, new_n489, new_n495);
xor_4  g00119(new_n445, new_n429, new_n496);
or_5   g00120(new_n496, new_n495, new_n497);
nor_5  g00121(new_n497, new_n487, new_n498);
nor_5  g00122(new_n498, new_n486, new_n499);
xor_4  g00123(new_n499, new_n482, new_n500);
nand_5 g00124(n8759, n5105, new_n501);
nand_5 g00125(n12299, n7354, new_n502);
nand_5 g00126(n8759, n1209, new_n503_1);
nand_5 g00127(new_n503_1, new_n502, new_n504);
not_8  g00128(new_n504, new_n505);
nor_5  g00129(new_n503_1, new_n502, new_n506);
nand_5 g00130(n7500, n6776, new_n507);
not_8  g00131(new_n507, new_n508);
nor_5  g00132(new_n508, new_n506, new_n509);
nor_5  g00133(new_n509, new_n505, new_n510);
not_8  g00134(new_n510, new_n511);
xor_4  g00135(new_n511, new_n501, new_n512);
nand_5 g00136(n12299, n7500, new_n513);
nand_5 g00137(n7436, n7354, new_n514);
nand_5 g00138(n6776, n1209, new_n515);
xor_4  g00139(new_n515, new_n514, new_n516);
not_8  g00140(new_n516, new_n517);
xor_4  g00141(new_n517, new_n513, new_n518);
xor_4  g00142(new_n518, new_n512, new_n519);
and_5  g00143(n8759, n7354, new_n520);
or_5   g00144(new_n520, new_n507, new_n521_1);
not_8  g00145(new_n521_1, new_n522);
nor_5  g00146(new_n522, new_n504, new_n523);
or_5   g00147(new_n523, new_n506, new_n524);
not_8  g00148(new_n524, new_n525);
or_5   g00149(new_n525, new_n507, new_n526);
not_8  g00150(new_n526, new_n527);
nand_5 g00151(new_n527, new_n519, new_n528);
nand_5 g00152(n8759, n4141, new_n529);
nand_5 g00153(n6776, n5105, new_n530);
not_8  g00154(new_n530, new_n531);
and_5  g00155(new_n515, new_n514, new_n532);
not_8  g00156(new_n513, new_n533_1);
nor_5  g00157(new_n517, new_n533_1, new_n534);
or_5   g00158(new_n534, new_n532, new_n535);
not_8  g00159(new_n535, new_n536);
xor_4  g00160(new_n536, new_n531, new_n537);
nand_5 g00161(n7500, n7436, new_n538);
nand_5 g00162(n12299, n1209, new_n539);
nand_5 g00163(n8276, n7354, new_n540);
xor_4  g00164(new_n540, new_n539, new_n541);
not_8  g00165(new_n541, new_n542);
xor_4  g00166(new_n542, new_n538, new_n543);
xor_4  g00167(new_n543, new_n537, new_n544);
not_8  g00168(new_n544, new_n545);
xor_4  g00169(new_n545, new_n529, new_n546);
nor_5  g00170(new_n511, new_n501, new_n547);
and_5  g00171(new_n518, new_n512, new_n548);
or_5   g00172(new_n548, new_n547, new_n549);
xor_4  g00173(new_n549, new_n546, new_n550);
not_8  g00174(new_n550, new_n551);
or_5   g00175(new_n551, new_n528, new_n552);
not_8  g00176(new_n552, new_n553);
nand_5 g00177(n8759, n4928, new_n554);
nand_5 g00178(n7436, n1209, new_n555);
nand_5 g00179(n8276, n7500, new_n556);
nand_5 g00180(n9241, n7354, new_n557);
xor_4  g00181(new_n557, new_n556, new_n558);
not_8  g00182(new_n558, new_n559);
xor_4  g00183(new_n559, new_n555, new_n560);
and_5  g00184(new_n540, new_n539, new_n561);
not_8  g00185(new_n538, new_n562);
nor_5  g00186(new_n542, new_n562, new_n563);
or_5   g00187(new_n563, new_n561, new_n564);
not_8  g00188(new_n564, new_n565);
xor_4  g00189(new_n565, new_n560, new_n566);
nand_5 g00190(n6776, n4141, new_n567);
nand_5 g00191(n12299, n5105, new_n568);
xor_4  g00192(new_n568, new_n567, new_n569);
xor_4  g00193(new_n569, new_n566, new_n570);
not_8  g00194(new_n570, new_n571);
and_5  g00195(new_n536, new_n531, new_n572);
and_5  g00196(new_n543, new_n537, new_n573);
nor_5  g00197(new_n573, new_n572, new_n574);
xor_4  g00198(new_n574, new_n571, new_n575);
not_8  g00199(new_n575, new_n576);
nor_5  g00200(new_n545, new_n529, new_n577);
and_5  g00201(new_n549, new_n546, new_n578);
nor_5  g00202(new_n578, new_n577, new_n579);
xor_4  g00203(new_n579, new_n576, new_n580);
not_8  g00204(new_n580, new_n581);
xor_4  g00205(new_n581, new_n554, new_n582);
xor_4  g00206(new_n582, new_n553, new_n583);
xor_4  g00207(new_n551, new_n528, new_n584);
xor_4  g00208(new_n526, new_n519, new_n585);
not_8  g00209(new_n585, new_n586);
nand_5 g00210(n5331, n1564, new_n587);
nand_5 g00211(n8028, n7965, new_n588);
xnor_4 g00212(new_n588, new_n587, new_n589);
not_8  g00213(new_n589, new_n590);
nand_5 g00214(new_n590, new_n520, new_n591);
nand_5 g00215(n7354, n6776, new_n592);
and_5  g00216(n8759, n7500, new_n593);
xor_4  g00217(new_n593, new_n592, new_n594);
and_5  g00218(new_n594, new_n591, new_n595);
or_5   g00219(new_n588, new_n587, new_n596);
nand_5 g00220(n5331, n1512, new_n597);
and_5  g00221(n8476, n1564, new_n598);
xor_4  g00222(new_n598, new_n597, new_n599);
not_8  g00223(new_n599, new_n600);
xor_4  g00224(new_n600, new_n596, new_n601);
nand_5 g00225(n8028, n7388, new_n602);
and_5  g00226(n10848, n7965, new_n603);
xor_4  g00227(new_n603, new_n602, new_n604);
xor_4  g00228(new_n604, new_n601, new_n605);
and_5  g00229(n7354, n6776, new_n606);
xor_4  g00230(new_n593, new_n606, new_n607);
xor_4  g00231(new_n607, new_n591, new_n608);
nor_5  g00232(new_n608, new_n605, new_n609);
or_5   g00233(new_n609, new_n595, new_n610);
not_8  g00234(new_n610, new_n611);
or_5   g00235(new_n521_1, new_n505, new_n612);
and_5  g00236(new_n612, new_n525, new_n613);
nor_5  g00237(new_n613, new_n611, new_n614);
not_8  g00238(new_n588, new_n615_1);
nand_5 g00239(n10848, n7388, new_n616);
or_5   g00240(new_n616, new_n615_1, new_n617);
not_8  g00241(new_n617, new_n618);
and_5  g00242(n11892, n8028, new_n619);
and_5  g00243(n7965, n1980, new_n620);
nor_5  g00244(new_n620, new_n619, new_n621);
nand_5 g00245(n11892, n1980, new_n622);
nor_5  g00246(new_n622, new_n588, new_n623);
nor_5  g00247(new_n623, new_n621, new_n624);
or_5   g00248(new_n624, new_n618, new_n625);
not_8  g00249(new_n625, new_n626);
nor_5  g00250(new_n621, new_n617, new_n627);
or_5   g00251(new_n627, new_n626, new_n628);
not_8  g00252(new_n587, new_n629);
nand_5 g00253(n8476, n1512, new_n630);
or_5   g00254(new_n630, new_n629, new_n631);
nand_5 g00255(n2530, n1564, new_n632);
nand_5 g00256(n5331, n533, new_n633);
nand_5 g00257(new_n633, new_n632, new_n634);
not_8  g00258(new_n634, new_n635);
and_5  g00259(new_n635, new_n631, new_n636);
nor_5  g00260(new_n633, new_n632, new_n637);
or_5   g00261(new_n637, new_n636, new_n638);
not_8  g00262(new_n638, new_n639);
or_5   g00263(new_n635, new_n631, new_n640);
nand_5 g00264(new_n640, new_n639, new_n641);
xnor_4 g00265(new_n641, new_n628, new_n642);
nor_5  g00266(new_n599, new_n596, new_n643);
nor_5  g00267(new_n604, new_n601, new_n644);
nor_5  g00268(new_n644, new_n643, new_n645);
xor_4  g00269(new_n645, new_n642, new_n646);
and_5  g00270(new_n613, new_n611, new_n647);
or_5   g00271(new_n647, new_n614, new_n648);
nor_5  g00272(new_n648, new_n646, new_n649);
nor_5  g00273(new_n649, new_n614, new_n650);
nor_5  g00274(new_n650, new_n586, new_n651);
nand_5 g00275(n5331, n2802, new_n652);
not_8  g00276(new_n630, new_n653);
nor_5  g00277(new_n637, new_n653, new_n654);
nor_5  g00278(new_n654, new_n635, new_n655);
not_8  g00279(new_n655, new_n656);
xor_4  g00280(new_n656, new_n652, new_n657);
nand_5 g00281(n2530, n1512, new_n658_1);
nand_5 g00282(n12648, n1564, new_n659);
nand_5 g00283(n8476, n533, new_n660);
xnor_4 g00284(new_n660, new_n659, new_n661);
not_8  g00285(new_n661, new_n662);
xor_4  g00286(new_n662, new_n658_1, new_n663);
xor_4  g00287(new_n663, new_n657, new_n664);
nor_5  g00288(new_n639, new_n630, new_n665);
xor_4  g00289(new_n665, new_n664, new_n666);
not_8  g00290(new_n666, new_n667);
nand_5 g00291(n7965, n7294, new_n668);
not_8  g00292(new_n616, new_n669);
nor_5  g00293(new_n623, new_n669, new_n670);
nor_5  g00294(new_n670, new_n621, new_n671_1);
not_8  g00295(new_n671_1, new_n672);
xor_4  g00296(new_n672, new_n668, new_n673);
nand_5 g00297(n11892, n10848, new_n674);
not_8  g00298(new_n674, new_n675);
nand_5 g00299(n7388, n1980, new_n676);
nand_5 g00300(n8028, n2393, new_n677);
xor_4  g00301(new_n677, new_n676, new_n678);
xor_4  g00302(new_n678, new_n675, new_n679);
xor_4  g00303(new_n679, new_n673, new_n680);
and_5  g00304(new_n626, new_n669, new_n681);
xor_4  g00305(new_n681, new_n680, new_n682);
xor_4  g00306(new_n682, new_n667, new_n683);
nor_5  g00307(new_n641, new_n628, new_n684);
nor_5  g00308(new_n645, new_n642, new_n685);
or_5   g00309(new_n685, new_n684, new_n686);
not_8  g00310(new_n686, new_n687);
xnor_4 g00311(new_n687, new_n683, new_n688);
xor_4  g00312(new_n650, new_n586, new_n689);
not_8  g00313(new_n689, new_n690);
nor_5  g00314(new_n690, new_n688, new_n691);
nor_5  g00315(new_n691, new_n651, new_n692);
nor_5  g00316(new_n692, new_n584, new_n693);
nand_5 g00317(new_n681, new_n680, new_n694);
or_5   g00318(new_n672, new_n668, new_n695);
nand_5 g00319(new_n679, new_n673, new_n696);
nand_5 g00320(new_n696, new_n695, new_n697);
nand_5 g00321(n12704, n7965, new_n698);
not_8  g00322(new_n698, new_n699);
nand_5 g00323(n7388, n7294, new_n700);
not_8  g00324(new_n700, new_n701);
and_5  g00325(new_n677, new_n676, new_n702);
nor_5  g00326(new_n677, new_n676, new_n703);
nor_5  g00327(new_n703, new_n675, new_n704);
or_5   g00328(new_n704, new_n702, new_n705);
not_8  g00329(new_n705, new_n706);
and_5  g00330(new_n706, new_n701, new_n707);
nor_5  g00331(new_n706, new_n701, new_n708);
or_5   g00332(new_n708, new_n707, new_n709);
nand_5 g00333(n10848, n2393, new_n710);
not_8  g00334(new_n710, new_n711);
nand_5 g00335(n8028, n5860, new_n712);
xor_4  g00336(new_n712, new_n622, new_n713);
xor_4  g00337(new_n713, new_n711, new_n714);
not_8  g00338(new_n714, new_n715);
xor_4  g00339(new_n715, new_n709, new_n716);
xor_4  g00340(new_n716, new_n699, new_n717);
xor_4  g00341(new_n717, new_n697, new_n718);
not_8  g00342(new_n718, new_n719);
xor_4  g00343(new_n719, new_n694, new_n720);
not_8  g00344(new_n720, new_n721);
not_8  g00345(new_n665, new_n722);
or_5   g00346(new_n722, new_n664, new_n723);
nand_5 g00347(n6806, n5331, new_n724);
nand_5 g00348(n8476, n2802, new_n725);
not_8  g00349(new_n725, new_n726);
and_5  g00350(new_n660, new_n659, new_n727);
and_5  g00351(new_n662, new_n658_1, new_n728);
or_5   g00352(new_n728, new_n727, new_n729);
not_8  g00353(new_n729, new_n730);
xor_4  g00354(new_n730, new_n726, new_n731);
nand_5 g00355(n12648, n1512, new_n732);
nand_5 g00356(n2530, n533, new_n733);
nand_5 g00357(n10545, n1564, new_n734);
xor_4  g00358(new_n734, new_n733, new_n735);
not_8  g00359(new_n735, new_n736);
xor_4  g00360(new_n736, new_n732, new_n737);
xor_4  g00361(new_n737, new_n731, new_n738);
not_8  g00362(new_n738, new_n739);
xor_4  g00363(new_n739, new_n724, new_n740);
or_5   g00364(new_n656, new_n652, new_n741);
not_8  g00365(new_n741, new_n742);
not_8  g00366(new_n658_1, new_n743);
xor_4  g00367(new_n662, new_n743, new_n744);
and_5  g00368(new_n744, new_n657, new_n745);
or_5   g00369(new_n745, new_n742, new_n746);
xor_4  g00370(new_n746, new_n740, new_n747);
not_8  g00371(new_n747, new_n748);
xor_4  g00372(new_n748, new_n723, new_n749);
nor_5  g00373(new_n682, new_n667, new_n750);
and_5  g00374(new_n687, new_n683, new_n751);
nor_5  g00375(new_n751, new_n750, new_n752);
xor_4  g00376(new_n752, new_n749, new_n753_1);
not_8  g00377(new_n753_1, new_n754);
xor_4  g00378(new_n754, new_n721, new_n755);
xor_4  g00379(new_n692, new_n584, new_n756);
not_8  g00380(new_n756, new_n757);
nor_5  g00381(new_n757, new_n755, new_n758);
nor_5  g00382(new_n758, new_n693, new_n759);
xor_4  g00383(new_n759, new_n583, new_n760);
not_8  g00384(new_n760, new_n761);
nor_5  g00385(new_n752, new_n749, new_n762);
nor_5  g00386(new_n754, new_n720, new_n763);
or_5   g00387(new_n763, new_n762, new_n764);
or_5   g00388(new_n748, new_n723, new_n765);
nand_5 g00389(n5331, n5069, new_n766);
nand_5 g00390(n12648, n533, new_n767);
nand_5 g00391(n10545, n1512, new_n768);
nand_5 g00392(n7690, n1564, new_n769);
xor_4  g00393(new_n769, new_n768, new_n770);
not_8  g00394(new_n770, new_n771);
xor_4  g00395(new_n771, new_n767, new_n772);
and_5  g00396(new_n734, new_n733, new_n773);
not_8  g00397(new_n732, new_n774);
nor_5  g00398(new_n736, new_n774, new_n775);
or_5   g00399(new_n775, new_n773, new_n776);
not_8  g00400(new_n776, new_n777);
xor_4  g00401(new_n777, new_n772, new_n778);
nand_5 g00402(n8476, n6806, new_n779);
nand_5 g00403(n2802, n2530, new_n780);
xor_4  g00404(new_n780, new_n779, new_n781);
xor_4  g00405(new_n781, new_n778, new_n782);
not_8  g00406(new_n782, new_n783_1);
and_5  g00407(new_n730, new_n726, new_n784);
and_5  g00408(new_n737, new_n731, new_n785);
nor_5  g00409(new_n785, new_n784, new_n786);
xor_4  g00410(new_n786, new_n783_1, new_n787);
not_8  g00411(new_n787, new_n788);
nor_5  g00412(new_n739, new_n724, new_n789);
and_5  g00413(new_n746, new_n740, new_n790);
nor_5  g00414(new_n790, new_n789, new_n791);
xor_4  g00415(new_n791, new_n788, new_n792);
not_8  g00416(new_n792, new_n793);
xor_4  g00417(new_n793, new_n766, new_n794);
xor_4  g00418(new_n794, new_n765, new_n795);
xor_4  g00419(new_n795, new_n764, new_n796);
not_8  g00420(new_n796, new_n797);
or_5   g00421(new_n719, new_n694, new_n798);
nand_5 g00422(n7965, n5814, new_n799);
not_8  g00423(new_n799, new_n800);
nand_5 g00424(n2393, n1980, new_n801);
nand_5 g00425(n8028, n3986, new_n802);
nand_5 g00426(n10848, n5860, new_n803);
xor_4  g00427(new_n803, new_n802, new_n804);
not_8  g00428(new_n804, new_n805);
xor_4  g00429(new_n805, new_n801, new_n806_1);
and_5  g00430(new_n712, new_n622, new_n807);
nor_5  g00431(new_n712, new_n622, new_n808);
nor_5  g00432(new_n808, new_n711, new_n809);
or_5   g00433(new_n809, new_n807, new_n810);
not_8  g00434(new_n810, new_n811);
xor_4  g00435(new_n811, new_n806_1, new_n812);
nand_5 g00436(n12704, n7388, new_n813);
nand_5 g00437(n11892, n7294, new_n814);
xor_4  g00438(new_n814, new_n813, new_n815);
xor_4  g00439(new_n815, new_n812, new_n816);
not_8  g00440(new_n816, new_n817);
nor_5  g00441(new_n715, new_n709, new_n818);
nor_5  g00442(new_n818, new_n707, new_n819);
xor_4  g00443(new_n819, new_n817, new_n820);
nor_5  g00444(new_n716, new_n699, new_n821);
and_5  g00445(new_n716, new_n699, new_n822);
nor_5  g00446(new_n822, new_n697, new_n823);
or_5   g00447(new_n823, new_n821, new_n824);
not_8  g00448(new_n824, new_n825);
xor_4  g00449(new_n825, new_n820, new_n826);
xor_4  g00450(new_n826, new_n800, new_n827);
xor_4  g00451(new_n827, new_n798, new_n828);
not_8  g00452(new_n828, new_n829);
xor_4  g00453(new_n829, new_n797, new_n830);
not_8  g00454(new_n830, new_n831);
xor_4  g00455(new_n831, new_n761, new_n832);
xor_4  g00456(new_n485, new_n484, new_n833);
xor_4  g00457(new_n833, new_n497, new_n834);
nor_5  g00458(new_n834, new_n832, new_n835);
xor_4  g00459(new_n496, new_n495, new_n836);
not_8  g00460(new_n836, new_n837_1);
xor_4  g00461(new_n757, new_n755, new_n838);
nor_5  g00462(new_n838, new_n837_1, new_n839);
xor_4  g00463(new_n838, new_n836, new_n840);
xor_4  g00464(new_n494, new_n489, new_n841);
not_8  g00465(new_n841, new_n842);
xor_4  g00466(new_n690, new_n688, new_n843);
or_5   g00467(new_n843, new_n842, new_n844_1);
not_8  g00468(new_n646, new_n845);
xor_4  g00469(new_n648, new_n845, new_n846);
not_8  g00470(new_n435, new_n847);
nand_5 g00471(n6038, n5305, new_n848);
and_5  g00472(new_n848, new_n847, new_n849);
nor_5  g00473(new_n849, new_n490, new_n850);
and_5  g00474(new_n848, new_n437, new_n851);
nor_5  g00475(new_n851, new_n850, new_n852);
nor_5  g00476(new_n852, new_n846, new_n853);
xor_4  g00477(new_n852, new_n846, new_n854);
not_8  g00478(new_n854, new_n855);
not_8  g00479(new_n848, new_n856);
xor_4  g00480(new_n590, new_n520, new_n857);
nand_5 g00481(new_n857, new_n856, new_n858);
xnor_4 g00482(new_n492, new_n491, new_n859);
and_5  g00483(new_n859, new_n858, new_n860);
not_8  g00484(new_n608, new_n861);
xor_4  g00485(new_n861, new_n605, new_n862);
xor_4  g00486(new_n859, new_n858, new_n863);
not_8  g00487(new_n863, new_n864);
nor_5  g00488(new_n864, new_n862, new_n865);
or_5   g00489(new_n865, new_n860, new_n866);
not_8  g00490(new_n866, new_n867);
nor_5  g00491(new_n867, new_n855, new_n868);
or_5   g00492(new_n868, new_n853, new_n869);
xor_4  g00493(new_n843, new_n841, new_n870);
or_5   g00494(new_n870, new_n869, new_n871);
and_5  g00495(new_n871, new_n844_1, new_n872);
nor_5  g00496(new_n872, new_n840, new_n873);
nor_5  g00497(new_n873, new_n839, new_n874);
not_8  g00498(new_n834, new_n875);
xor_4  g00499(new_n875, new_n832, new_n876);
nor_5  g00500(new_n876, new_n874, new_n877);
nor_5  g00501(new_n877, new_n835, new_n878);
xor_4  g00502(new_n878, new_n500, new_n879);
not_8  g00503(new_n879, new_n880);
or_5   g00504(new_n579, new_n576, new_n881);
not_8  g00505(new_n881, new_n882);
nor_5  g00506(new_n559, new_n555, new_n883);
and_5  g00507(new_n565, new_n560, new_n884);
or_5   g00508(new_n884, new_n883, new_n885);
not_8  g00509(new_n885, new_n886);
nand_5 g00510(n6776, n4928, new_n887);
not_8  g00511(new_n887, new_n888);
nand_5 g00512(n12299, n4141, new_n889);
nand_5 g00513(n8759, n8236, new_n890);
xor_4  g00514(new_n890, new_n889, new_n891);
not_8  g00515(new_n891, new_n892);
xor_4  g00516(new_n892, new_n888, new_n893);
xor_4  g00517(new_n893, new_n886, new_n894);
or_5   g00518(new_n557, new_n556, new_n895);
not_8  g00519(new_n895, new_n896);
nand_5 g00520(n7436, n5105, new_n897);
not_8  g00521(new_n897, new_n898);
xor_4  g00522(new_n898, new_n896, new_n899);
and_5  g00523(n9241, n7500, new_n900);
nand_5 g00524(n8276, n1209, new_n901);
nand_5 g00525(n10510, n7354, new_n902);
xor_4  g00526(new_n902, new_n901, new_n903);
xor_4  g00527(new_n903, new_n900, new_n904);
xor_4  g00528(new_n904, new_n899, new_n905);
xor_4  g00529(new_n905, new_n894, new_n906);
not_8  g00530(new_n906, new_n907);
and_5  g00531(new_n569, new_n566, new_n908);
or_5   g00532(new_n568, new_n567, new_n909);
not_8  g00533(new_n909, new_n910);
or_5   g00534(new_n574, new_n571, new_n911_1);
not_8  g00535(new_n911_1, new_n912);
xor_4  g00536(new_n912, new_n910, new_n913);
nor_5  g00537(new_n913, new_n908, new_n914);
xor_4  g00538(new_n914, new_n907, new_n915);
not_8  g00539(new_n915, new_n916);
xnor_4 g00540(new_n916, new_n882, new_n917);
not_8  g00541(new_n917, new_n918);
nor_5  g00542(new_n581, new_n554, new_n919);
and_5  g00543(new_n582, new_n553, new_n920);
nor_5  g00544(new_n920, new_n919, new_n921);
xor_4  g00545(new_n921, new_n918, new_n922);
not_8  g00546(new_n922, new_n923);
or_5   g00547(new_n791, new_n788, new_n924);
not_8  g00548(new_n924, new_n925);
nor_5  g00549(new_n771, new_n767, new_n926);
and_5  g00550(new_n777, new_n772, new_n927);
or_5   g00551(new_n927, new_n926, new_n928);
not_8  g00552(new_n928, new_n929);
nand_5 g00553(n8476, n5069, new_n930);
not_8  g00554(new_n930, new_n931);
nand_5 g00555(n6806, n2530, new_n932);
nand_5 g00556(n12044, n5331, new_n933);
xor_4  g00557(new_n933, new_n932, new_n934);
not_8  g00558(new_n934, new_n935);
xor_4  g00559(new_n935, new_n931, new_n936);
xor_4  g00560(new_n936, new_n929, new_n937);
or_5   g00561(new_n769, new_n768, new_n938);
not_8  g00562(new_n938, new_n939);
nand_5 g00563(n12648, n2802, new_n940);
not_8  g00564(new_n940, new_n941);
xor_4  g00565(new_n941, new_n939, new_n942);
nand_5 g00566(n7690, n1512, new_n943);
nand_5 g00567(n10545, n533, new_n944);
nand_5 g00568(n3616, n1564, new_n945);
xor_4  g00569(new_n945, new_n944, new_n946);
not_8  g00570(new_n946, new_n947);
xor_4  g00571(new_n947, new_n943, new_n948);
xor_4  g00572(new_n948, new_n942, new_n949);
xor_4  g00573(new_n949, new_n937, new_n950);
not_8  g00574(new_n950, new_n951);
and_5  g00575(new_n781, new_n778, new_n952);
or_5   g00576(new_n780, new_n779, new_n953);
not_8  g00577(new_n953, new_n954);
or_5   g00578(new_n786, new_n783_1, new_n955);
not_8  g00579(new_n955, new_n956);
xor_4  g00580(new_n956, new_n954, new_n957);
nor_5  g00581(new_n957, new_n952, new_n958);
xor_4  g00582(new_n958, new_n951, new_n959);
not_8  g00583(new_n959, new_n960);
xnor_4 g00584(new_n960, new_n925, new_n961);
not_8  g00585(new_n961, new_n962);
nor_5  g00586(new_n793, new_n766, new_n963);
and_5  g00587(new_n793, new_n766, new_n964);
nor_5  g00588(new_n964, new_n765, new_n965);
nor_5  g00589(new_n965, new_n963, new_n966);
xor_4  g00590(new_n966, new_n962, new_n967);
not_8  g00591(new_n967, new_n968);
nand_5 g00592(new_n825, new_n820, new_n969);
nor_5  g00593(new_n805, new_n801, new_n970);
and_5  g00594(new_n811, new_n806_1, new_n971);
or_5   g00595(new_n971, new_n970, new_n972);
nand_5 g00596(n7388, n5814, new_n973);
not_8  g00597(new_n973, new_n974);
nand_5 g00598(n12704, n11892, new_n975);
nand_5 g00599(n7965, n4903, new_n976);
xor_4  g00600(new_n976, new_n975, new_n977);
not_8  g00601(new_n977, new_n978);
xor_4  g00602(new_n978, new_n974, new_n979);
not_8  g00603(new_n979, new_n980);
xor_4  g00604(new_n980, new_n972, new_n981);
or_5   g00605(new_n803, new_n802, new_n982);
not_8  g00606(new_n982, new_n983);
nand_5 g00607(n7294, n2393, new_n984);
not_8  g00608(new_n984, new_n985);
xor_4  g00609(new_n985, new_n983, new_n986);
nand_5 g00610(n10848, n3986, new_n987);
nand_5 g00611(n5860, n1980, new_n988);
nand_5 g00612(n8028, n5857, new_n989);
xor_4  g00613(new_n989, new_n988, new_n990);
not_8  g00614(new_n990, new_n991);
xor_4  g00615(new_n991, new_n987, new_n992_1);
xor_4  g00616(new_n992_1, new_n986, new_n993);
xor_4  g00617(new_n993, new_n981, new_n994);
not_8  g00618(new_n994, new_n995);
nand_5 g00619(new_n815, new_n812, new_n996_1);
or_5   g00620(new_n814, new_n813, new_n997);
or_5   g00621(new_n819, new_n817, new_n998);
not_8  g00622(new_n998, new_n999);
xor_4  g00623(new_n999, new_n997, new_n1000);
and_5  g00624(new_n1000, new_n996_1, new_n1001);
xor_4  g00625(new_n1001, new_n995, new_n1002);
xnor_4 g00626(new_n1002, new_n969, new_n1003);
nor_5  g00627(new_n826, new_n800, new_n1004);
not_8  g00628(new_n798, new_n1005);
and_5  g00629(new_n826, new_n800, new_n1006);
nor_5  g00630(new_n1006, new_n1005, new_n1007);
or_5   g00631(new_n1007, new_n1004, new_n1008);
not_8  g00632(new_n1008, new_n1009);
xnor_4 g00633(new_n1009, new_n1003, new_n1010);
xor_4  g00634(new_n1010, new_n968, new_n1011);
or_5   g00635(new_n795, new_n764, new_n1012);
not_8  g00636(new_n1012, new_n1013);
nand_5 g00637(new_n795, new_n764, new_n1014);
and_5  g00638(new_n829, new_n1014, new_n1015);
or_5   g00639(new_n1015, new_n1013, new_n1016);
not_8  g00640(new_n1016, new_n1017);
xor_4  g00641(new_n1017, new_n1011, new_n1018);
xor_4  g00642(new_n1018, new_n923, new_n1019);
nor_5  g00643(new_n759, new_n583, new_n1020_1);
nor_5  g00644(new_n831, new_n761, new_n1021);
or_5   g00645(new_n1021, new_n1020_1, new_n1022);
xor_4  g00646(new_n1022, new_n1019, new_n1023);
not_8  g00647(new_n1023, new_n1024);
nand_5 g00648(new_n1024, new_n880, new_n1025);
or_5   g00649(new_n1024, new_n880, new_n1026);
and_5  g00650(new_n1026, new_n1025, n226);
nand_5 g00651(n5305, n4634, new_n1028);
not_8  g00652(new_n1028, new_n1029);
and_5  g00653(n10223, n5305, new_n1030);
and_5  g00654(n7265, n1097, new_n1031);
nor_5  g00655(new_n1031, new_n1030, new_n1032);
nand_5 g00656(n7265, n5305, new_n1033);
nand_5 g00657(n10223, n1097, new_n1034);
nor_5  g00658(new_n1034, new_n1033, new_n1035);
nand_5 g00659(n5964, n2879, new_n1036);
not_8  g00660(new_n1036, new_n1037);
nor_5  g00661(new_n1037, new_n1035, new_n1038);
or_5   g00662(new_n1038, new_n1032, new_n1039);
not_8  g00663(new_n1039, new_n1040);
and_5  g00664(new_n1040, new_n1029, new_n1041);
nor_5  g00665(new_n1040, new_n1029, new_n1042);
or_5   g00666(new_n1042, new_n1041, new_n1043);
nand_5 g00667(n2879, n1097, new_n1044);
not_8  g00668(new_n1044, new_n1045);
nand_5 g00669(n10223, n5964, new_n1046);
nand_5 g00670(n7265, n4312, new_n1047);
xor_4  g00671(new_n1047, new_n1046, new_n1048);
xor_4  g00672(new_n1048, new_n1045, new_n1049);
not_8  g00673(new_n1049, new_n1050);
xor_4  g00674(new_n1050, new_n1043, new_n1051);
not_8  g00675(new_n1033, new_n1052);
or_5   g00676(new_n1036, new_n1052, new_n1053);
not_8  g00677(new_n1053, new_n1054);
nor_5  g00678(new_n1035, new_n1032, new_n1055);
or_5   g00679(new_n1055, new_n1054, new_n1056);
not_8  g00680(new_n1056, new_n1057);
nand_5 g00681(new_n1057, new_n1037, new_n1058);
not_8  g00682(new_n1058, new_n1059);
xor_4  g00683(new_n1059, new_n1051, new_n1060);
not_8  g00684(new_n1060, new_n1061);
nor_5  g00685(new_n1053, new_n1032, new_n1062);
or_5   g00686(new_n1062, new_n1057, new_n1063);
nand_5 g00687(n8759, n7946, new_n1064);
not_8  g00688(new_n1064, new_n1065);
nand_5 g00689(n5331, n2558, new_n1066);
nand_5 g00690(n9763, n7965, new_n1067_1);
xnor_4 g00691(new_n1067_1, new_n1066, new_n1068);
not_8  g00692(new_n1068, new_n1069);
nand_5 g00693(new_n1069, new_n1065, new_n1070);
and_5  g00694(n7946, n6776, new_n1071);
and_5  g00695(n8759, n2024, new_n1072);
xor_4  g00696(new_n1072, new_n1071, new_n1073);
not_8  g00697(new_n1073, new_n1074);
nor_5  g00698(new_n1074, new_n1070, new_n1075);
or_5   g00699(new_n1067_1, new_n1066, new_n1076);
and_5  g00700(n9111, n7965, new_n1077);
and_5  g00701(n9763, n7388, new_n1078);
xor_4  g00702(new_n1078, new_n1077, new_n1079);
xor_4  g00703(new_n1079, new_n1076, new_n1080);
not_8  g00704(new_n1080, new_n1081);
and_5  g00705(n5331, n2498, new_n1082);
and_5  g00706(n8476, n2558, new_n1083);
xnor_4 g00707(new_n1083, new_n1082, new_n1084);
xor_4  g00708(new_n1084, new_n1081, new_n1085);
xor_4  g00709(new_n1073, new_n1070, new_n1086);
nor_5  g00710(new_n1086, new_n1085, new_n1087);
nor_5  g00711(new_n1087, new_n1075, new_n1088);
not_8  g00712(new_n1088, new_n1089);
nand_5 g00713(n6776, n2024, new_n1090);
or_5   g00714(new_n1090, new_n1065, new_n1091);
nand_5 g00715(n12299, n7946, new_n1092);
nand_5 g00716(n9189, n8759, new_n1093);
xnor_4 g00717(new_n1093, new_n1092, new_n1094_1);
and_5  g00718(new_n1094_1, new_n1091, new_n1095);
and_5  g00719(new_n1093, new_n1092, new_n1096);
nor_5  g00720(new_n1096, new_n1091, new_n1097_1);
or_5   g00721(new_n1097_1, new_n1095, new_n1098);
xor_4  g00722(new_n1098, new_n1089, new_n1099);
not_8  g00723(new_n1076, new_n1100);
nor_5  g00724(new_n1079, new_n1100, new_n1101);
and_5  g00725(new_n1084, new_n1081, new_n1102);
or_5   g00726(new_n1102, new_n1101, new_n1103);
and_5  g00727(n9111, n7388, new_n1104);
and_5  g00728(new_n1104, new_n1067_1, new_n1105);
nand_5 g00729(n11892, n3342, new_n1106);
nor_5  g00730(new_n1106, new_n1067_1, new_n1107);
and_5  g00731(n11892, n9763, new_n1108);
and_5  g00732(n7965, n3342, new_n1109);
nor_5  g00733(new_n1109, new_n1108, new_n1110);
nor_5  g00734(new_n1110, new_n1107, new_n1111);
or_5   g00735(new_n1111, new_n1105, new_n1112);
not_8  g00736(new_n1112, new_n1113);
not_8  g00737(new_n1105, new_n1114);
nor_5  g00738(new_n1110, new_n1114, new_n1115);
or_5   g00739(new_n1115, new_n1113, new_n1116);
xor_4  g00740(new_n1116, new_n1103, new_n1117);
and_5  g00741(n8476, n2498, new_n1118);
nand_5 g00742(new_n1118, new_n1066, new_n1119);
and_5  g00743(n2558, n2530, new_n1120);
and_5  g00744(n5579, n5331, new_n1121);
nor_5  g00745(new_n1121, new_n1120, new_n1122);
not_8  g00746(new_n1122, new_n1123);
nor_5  g00747(new_n1123, new_n1119, new_n1124);
nand_5 g00748(n5579, n2530, new_n1125);
nor_5  g00749(new_n1125, new_n1066, new_n1126);
or_5   g00750(new_n1126, new_n1122, new_n1127);
not_8  g00751(new_n1127, new_n1128);
and_5  g00752(new_n1128, new_n1119, new_n1129);
or_5   g00753(new_n1129, new_n1124, new_n1130);
not_8  g00754(new_n1130, new_n1131);
xor_4  g00755(new_n1131, new_n1117, new_n1132);
not_8  g00756(new_n1132, new_n1133);
xor_4  g00757(new_n1133, new_n1099, new_n1134);
or_5   g00758(new_n1134, new_n1063, new_n1135);
xor_4  g00759(new_n1069, new_n1065, new_n1136_1);
nand_5 g00760(new_n1136_1, new_n1052, new_n1137);
nand_5 g00761(n7265, n5964, new_n1138_1);
and_5  g00762(n5305, n2879, new_n1139);
xor_4  g00763(new_n1139, new_n1138_1, new_n1140);
and_5  g00764(new_n1140, new_n1137, new_n1141);
xor_4  g00765(new_n1086, new_n1085, new_n1142);
xor_4  g00766(new_n1140, new_n1137, new_n1143);
not_8  g00767(new_n1143, new_n1144);
nor_5  g00768(new_n1144, new_n1142, new_n1145);
or_5   g00769(new_n1145, new_n1141, new_n1146);
not_8  g00770(new_n1146, new_n1147);
not_8  g00771(new_n1063, new_n1148);
xor_4  g00772(new_n1134, new_n1148, new_n1149);
not_8  g00773(new_n1149, new_n1150);
nand_5 g00774(new_n1150, new_n1147, new_n1151);
and_5  g00775(new_n1151, new_n1135, new_n1152);
xor_4  g00776(new_n1152, new_n1061, new_n1153);
not_8  g00777(new_n1153, new_n1154);
nand_5 g00778(n8759, n2522, new_n1155);
not_8  g00779(new_n1155, new_n1156);
not_8  g00780(new_n1090, new_n1157);
nor_5  g00781(new_n1093, new_n1092, new_n1158);
nor_5  g00782(new_n1158, new_n1157, new_n1159);
nor_5  g00783(new_n1159, new_n1096, new_n1160);
not_8  g00784(new_n1160, new_n1161);
xor_4  g00785(new_n1161, new_n1156, new_n1162);
nand_5 g00786(n12299, n2024, new_n1163);
not_8  g00787(new_n1163, new_n1164);
nand_5 g00788(n7946, n7436, new_n1165);
nand_5 g00789(n9189, n6776, new_n1166);
xor_4  g00790(new_n1166, new_n1165, new_n1167);
xor_4  g00791(new_n1167, new_n1164, new_n1168);
not_8  g00792(new_n1168, new_n1169);
xor_4  g00793(new_n1169, new_n1162, new_n1170);
not_8  g00794(new_n1095, new_n1171);
or_5   g00795(new_n1171, new_n1090, new_n1172);
not_8  g00796(new_n1172, new_n1173);
xor_4  g00797(new_n1173, new_n1170, new_n1174);
not_8  g00798(new_n1174, new_n1175);
not_8  g00799(new_n1098, new_n1176);
nor_5  g00800(new_n1176, new_n1089, new_n1177);
nor_5  g00801(new_n1133, new_n1099, new_n1178);
or_5   g00802(new_n1178, new_n1177, new_n1179);
not_8  g00803(new_n1179, new_n1180);
xor_4  g00804(new_n1180, new_n1175, new_n1181);
nand_5 g00805(n5331, n521, new_n1182);
not_8  g00806(new_n1182, new_n1183);
nor_5  g00807(new_n1126, new_n1118, new_n1184);
or_5   g00808(new_n1184, new_n1122, new_n1185);
not_8  g00809(new_n1185, new_n1186);
and_5  g00810(new_n1186, new_n1183, new_n1187);
nor_5  g00811(new_n1186, new_n1183, new_n1188);
or_5   g00812(new_n1188, new_n1187, new_n1189);
and_5  g00813(n2530, n2498, new_n1190);
not_8  g00814(new_n1190, new_n1191);
nand_5 g00815(n12648, n2558, new_n1192);
and_5  g00816(n8476, n5579, new_n1193);
xor_4  g00817(new_n1193, new_n1192, new_n1194);
not_8  g00818(new_n1194, new_n1195);
xor_4  g00819(new_n1195, new_n1191, new_n1196);
xor_4  g00820(new_n1196, new_n1189, new_n1197);
nand_5 g00821(new_n1083, new_n1082, new_n1198_1);
or_5   g00822(new_n1128, new_n1198_1, new_n1199_1);
not_8  g00823(new_n1199_1, new_n1200);
xor_4  g00824(new_n1200, new_n1197, new_n1201);
nand_5 g00825(n7965, n806, new_n1202);
nand_5 g00826(n9111, n7388, new_n1203);
nor_5  g00827(new_n1110, new_n1203, new_n1204);
nor_5  g00828(new_n1204, new_n1107, new_n1205);
xor_4  g00829(new_n1205, new_n1202, new_n1206);
not_8  g00830(new_n1206, new_n1207);
and_5  g00831(n11892, n9111, new_n1208);
not_8  g00832(new_n1208, new_n1209_1);
nand_5 g00833(n9763, n2393, new_n1210);
and_5  g00834(n7388, n3342, new_n1211);
xor_4  g00835(new_n1211, new_n1210, new_n1212);
not_8  g00836(new_n1212, new_n1213);
xor_4  g00837(new_n1213, new_n1209_1, new_n1214);
nor_5  g00838(new_n1214, new_n1207, new_n1215);
and_5  g00839(new_n1214, new_n1207, new_n1216);
or_5   g00840(new_n1216, new_n1215, new_n1217);
and_5  g00841(new_n1113, new_n1104, new_n1218);
xnor_4 g00842(new_n1218, new_n1217, new_n1219);
xor_4  g00843(new_n1219, new_n1201, new_n1220);
not_8  g00844(new_n1220, new_n1221);
and_5  g00845(new_n1116, new_n1103, new_n1222);
and_5  g00846(new_n1131, new_n1117, new_n1223);
nor_5  g00847(new_n1223, new_n1222, new_n1224);
xor_4  g00848(new_n1224, new_n1221, new_n1225);
xor_4  g00849(new_n1225, new_n1181, new_n1226);
xnor_4 g00850(new_n1226, new_n1154, n381);
nand_5 g00851(n7862, n6038, new_n1228);
not_8  g00852(new_n1228, new_n1229);
nand_5 g00853(n7354, n6877, new_n1230);
nand_5 g00854(n4805, n1564, new_n1231);
nand_5 g00855(n8028, n7236, new_n1232);
xor_4  g00856(new_n1232, new_n1231, new_n1233);
not_8  g00857(new_n1233, new_n1234);
xor_4  g00858(new_n1234, new_n1230, new_n1235);
xor_4  g00859(new_n1235, new_n1229, n397);
nand_5 g00860(n6687, n4370, new_n1237);
not_8  g00861(new_n1237, new_n1238);
nand_5 g00862(n11407, n4189, new_n1239);
nand_5 g00863(n11877, n6687, new_n1240);
nand_5 g00864(new_n1240, new_n1239, new_n1241);
not_8  g00865(new_n1241, new_n1242);
nor_5  g00866(new_n1240, new_n1239, new_n1243);
nand_5 g00867(n5212, n2564, new_n1244);
not_8  g00868(new_n1244, new_n1245);
nor_5  g00869(new_n1245, new_n1243, new_n1246);
nor_5  g00870(new_n1246, new_n1242, new_n1247);
not_8  g00871(new_n1247, new_n1248);
xor_4  g00872(new_n1248, new_n1238, new_n1249);
nand_5 g00873(n5212, n4189, new_n1250);
not_8  g00874(new_n1250, new_n1251);
nand_5 g00875(n11407, n6770, new_n1252);
nand_5 g00876(n11877, n2564, new_n1253);
xor_4  g00877(new_n1253, new_n1252, new_n1254);
not_8  g00878(new_n1254, new_n1255);
xor_4  g00879(new_n1255, new_n1251, new_n1256);
xor_4  g00880(new_n1256, new_n1249, new_n1257);
nand_5 g00881(n11407, n6687, new_n1258);
not_8  g00882(new_n1258, new_n1259);
or_5   g00883(new_n1259, new_n1244, new_n1260);
and_5  g00884(new_n1260, new_n1242, new_n1261);
or_5   g00885(new_n1261, new_n1243, new_n1262);
not_8  g00886(new_n1262, new_n1263);
or_5   g00887(new_n1263, new_n1244, new_n1264);
xor_4  g00888(new_n1264, new_n1257, new_n1265);
not_8  g00889(new_n1265, new_n1266);
nand_5 g00890(n12709, n8336, new_n1267);
not_8  g00891(new_n1267, new_n1268);
nand_5 g00892(n11222, n10990, new_n1269_1);
nand_5 g00893(n12489, n12069, new_n1270);
xnor_4 g00894(new_n1270, new_n1269_1, new_n1271);
not_8  g00895(new_n1271, new_n1272);
nand_5 g00896(new_n1272, new_n1268, new_n1273);
nand_5 g00897(n11728, n8336, new_n1274);
and_5  g00898(n12709, n10928, new_n1275);
xor_4  g00899(new_n1275, new_n1274, new_n1276);
and_5  g00900(new_n1276, new_n1273, new_n1277);
or_5   g00901(new_n1270, new_n1269_1, new_n1278);
nand_5 g00902(n11222, n5760, new_n1279);
and_5  g00903(n11153, n10990, new_n1280);
xor_4  g00904(new_n1280, new_n1279, new_n1281);
not_8  g00905(new_n1281, new_n1282);
xor_4  g00906(new_n1282, new_n1278, new_n1283);
nand_5 g00907(n12069, n7159, new_n1284);
and_5  g00908(n12489, n12391, new_n1285);
xor_4  g00909(new_n1285, new_n1284, new_n1286);
xor_4  g00910(new_n1286, new_n1283, new_n1287);
and_5  g00911(n11728, n8336, new_n1288);
xor_4  g00912(new_n1275, new_n1288, new_n1289);
xor_4  g00913(new_n1289, new_n1273, new_n1290);
nor_5  g00914(new_n1290, new_n1287, new_n1291);
or_5   g00915(new_n1291, new_n1277, new_n1292);
not_8  g00916(new_n1292, new_n1293);
nand_5 g00917(n11728, n10928, new_n1294);
not_8  g00918(new_n1294, new_n1295);
and_5  g00919(new_n1295, new_n1267, new_n1296);
nand_5 g00920(n6986, n6429, new_n1297);
nor_5  g00921(new_n1297, new_n1267, new_n1298);
and_5  g00922(n12709, n6986, new_n1299);
and_5  g00923(n8336, n6429, new_n1300);
nor_5  g00924(new_n1300, new_n1299, new_n1301);
nor_5  g00925(new_n1301, new_n1298, new_n1302);
nor_5  g00926(new_n1302, new_n1296, new_n1303);
not_8  g00927(new_n1303, new_n1304);
or_5   g00928(new_n1300, new_n1299, new_n1305);
nand_5 g00929(new_n1305, new_n1296, new_n1306);
and_5  g00930(new_n1306, new_n1304, new_n1307);
and_5  g00931(new_n1307, new_n1293, new_n1308);
nor_5  g00932(new_n1307, new_n1293, new_n1309);
or_5   g00933(new_n1309, new_n1308, new_n1310);
not_8  g00934(new_n1270, new_n1311);
nand_5 g00935(n12391, n7159, new_n1312);
or_5   g00936(new_n1312, new_n1311, new_n1313);
nand_5 g00937(n12489, n7891, new_n1314);
nand_5 g00938(n12777, n12069, new_n1315);
nand_5 g00939(new_n1315, new_n1314, new_n1316);
not_8  g00940(new_n1316, new_n1317);
and_5  g00941(new_n1317, new_n1313, new_n1318);
nor_5  g00942(new_n1315, new_n1314, new_n1319);
or_5   g00943(new_n1319, new_n1318, new_n1320);
not_8  g00944(new_n1320, new_n1321);
or_5   g00945(new_n1317, new_n1313, new_n1322);
nand_5 g00946(new_n1322, new_n1321, new_n1323);
not_8  g00947(new_n1269_1, new_n1324);
nand_5 g00948(n11153, n5760, new_n1325);
or_5   g00949(new_n1325, new_n1324, new_n1326);
nand_5 g00950(n10990, n5314, new_n1327);
nand_5 g00951(n11222, n1478, new_n1328);
xnor_4 g00952(new_n1328, new_n1327, new_n1329);
and_5  g00953(new_n1329, new_n1326, new_n1330);
and_5  g00954(new_n1328, new_n1327, new_n1331);
nor_5  g00955(new_n1331, new_n1326, new_n1332);
or_5   g00956(new_n1332, new_n1330, new_n1333_1);
not_8  g00957(new_n1333_1, new_n1334);
xor_4  g00958(new_n1334, new_n1323, new_n1335);
nor_5  g00959(new_n1281, new_n1278, new_n1336);
nor_5  g00960(new_n1286, new_n1283, new_n1337);
nor_5  g00961(new_n1337, new_n1336, new_n1338);
xor_4  g00962(new_n1338, new_n1335, new_n1339);
xor_4  g00963(new_n1339, new_n1310, new_n1340);
or_5   g00964(new_n1260, new_n1242, new_n1341);
nand_5 g00965(new_n1341, new_n1263, new_n1342);
and_5  g00966(new_n1342, new_n1340, new_n1343);
and_5  g00967(new_n1341, new_n1263, new_n1344);
xor_4  g00968(new_n1344, new_n1340, new_n1345);
not_8  g00969(new_n1345, new_n1346);
xor_4  g00970(new_n1272, new_n1268, new_n1347);
nand_5 g00971(new_n1347, new_n1259, new_n1348);
nand_5 g00972(n11407, n2564, new_n1349);
and_5  g00973(n6687, n5212, new_n1350);
xor_4  g00974(new_n1350, new_n1349, new_n1351);
and_5  g00975(new_n1351, new_n1348, new_n1352);
not_8  g00976(new_n1290, new_n1353_1);
xor_4  g00977(new_n1353_1, new_n1287, new_n1354);
xor_4  g00978(new_n1351, new_n1348, new_n1355);
not_8  g00979(new_n1355, new_n1356);
nor_5  g00980(new_n1356, new_n1354, new_n1357_1);
or_5   g00981(new_n1357_1, new_n1352, new_n1358);
and_5  g00982(new_n1358, new_n1346, new_n1359);
or_5   g00983(new_n1359, new_n1343, new_n1360);
not_8  g00984(new_n1360, new_n1361);
xor_4  g00985(new_n1361, new_n1266, new_n1362);
nand_5 g00986(n8819, n8336, new_n1363);
nand_5 g00987(n11728, n6986, new_n1364);
not_8  g00988(new_n1364, new_n1365);
nand_5 g00989(n10928, n6429, new_n1366);
nand_5 g00990(n12709, n2226, new_n1367);
xor_4  g00991(new_n1367, new_n1366, new_n1368);
xor_4  g00992(new_n1368, new_n1365, new_n1369);
not_8  g00993(new_n1369, new_n1370);
xor_4  g00994(new_n1370, new_n1363, new_n1371);
nor_5  g00995(new_n1301, new_n1294, new_n1372);
or_5   g00996(new_n1372, new_n1298, new_n1373);
xor_4  g00997(new_n1373, new_n1371, new_n1374);
not_8  g00998(new_n1374, new_n1375);
or_5   g00999(new_n1304, new_n1294, new_n1376);
xor_4  g01000(new_n1376, new_n1375, new_n1377);
nand_5 g01001(n12069, n6254, new_n1378);
not_8  g01002(new_n1312, new_n1379);
nor_5  g01003(new_n1319, new_n1379, new_n1380);
nor_5  g01004(new_n1380, new_n1317, new_n1381);
not_8  g01005(new_n1381, new_n1382);
xor_4  g01006(new_n1382, new_n1378, new_n1383);
nand_5 g01007(n12489, n7160, new_n1384);
nand_5 g01008(n12777, n12391, new_n1385);
nand_5 g01009(n7891, n7159, new_n1386);
xor_4  g01010(new_n1386, new_n1385, new_n1387);
not_8  g01011(new_n1387, new_n1388);
xor_4  g01012(new_n1388, new_n1384, new_n1389);
xor_4  g01013(new_n1389, new_n1383, new_n1390);
nor_5  g01014(new_n1321, new_n1312, new_n1391);
xor_4  g01015(new_n1391, new_n1390, new_n1392);
nand_5 g01016(n11791, n11222, new_n1393);
not_8  g01017(new_n1393, new_n1394);
not_8  g01018(new_n1325, new_n1395);
nor_5  g01019(new_n1328, new_n1327, new_n1396);
nor_5  g01020(new_n1396, new_n1395, new_n1397);
nor_5  g01021(new_n1397, new_n1331, new_n1398);
not_8  g01022(new_n1398, new_n1399);
xor_4  g01023(new_n1399, new_n1394, new_n1400);
nand_5 g01024(n5760, n5314, new_n1401);
not_8  g01025(new_n1401, new_n1402);
nand_5 g01026(n10990, n996, new_n1403);
nand_5 g01027(n11153, n1478, new_n1404);
xor_4  g01028(new_n1404, new_n1403, new_n1405);
not_8  g01029(new_n1405, new_n1406);
xor_4  g01030(new_n1406, new_n1402, new_n1407);
xor_4  g01031(new_n1407, new_n1400, new_n1408);
not_8  g01032(new_n1330, new_n1409);
nor_5  g01033(new_n1409, new_n1325, new_n1410);
xor_4  g01034(new_n1410, new_n1408, new_n1411);
xor_4  g01035(new_n1411, new_n1392, new_n1412);
not_8  g01036(new_n1412, new_n1413);
nor_5  g01037(new_n1333_1, new_n1323, new_n1414);
nor_5  g01038(new_n1338, new_n1335, new_n1415);
or_5   g01039(new_n1415, new_n1414, new_n1416);
not_8  g01040(new_n1416, new_n1417);
xnor_4 g01041(new_n1417, new_n1413, new_n1418);
xor_4  g01042(new_n1418, new_n1377, new_n1419);
nor_5  g01043(new_n1339, new_n1310, new_n1420);
or_5   g01044(new_n1420, new_n1309, new_n1421);
not_8  g01045(new_n1421, new_n1422);
xor_4  g01046(new_n1422, new_n1419, new_n1423);
xnor_4 g01047(new_n1423, new_n1362, n658);
nand_5 g01048(n7862, n2585, new_n1425);
not_8  g01049(new_n1425, new_n1426);
and_5  g01050(n2508, n1333, new_n1427);
nand_5 g01051(n11757, n6038, new_n1428);
nand_5 g01052(n12720, n1333, new_n1429);
and_5  g01053(new_n1429, new_n1428, new_n1430);
nor_5  g01054(new_n1429, new_n1428, new_n1431);
nand_5 g01055(n3172, n2509, new_n1432);
not_8  g01056(new_n1432, new_n1433);
nor_5  g01057(new_n1433, new_n1431, new_n1434);
or_5   g01058(new_n1434, new_n1430, new_n1435);
not_8  g01059(new_n1435, new_n1436);
and_5  g01060(new_n1436, new_n1427, new_n1437);
nor_5  g01061(new_n1436, new_n1427, new_n1438);
or_5   g01062(new_n1438, new_n1437, new_n1439);
nand_5 g01063(n11757, n2509, new_n1440);
not_8  g01064(new_n1440, new_n1441);
nand_5 g01065(n6038, n5240, new_n1442);
nand_5 g01066(n12720, n3172, new_n1443);
xor_4  g01067(new_n1443, new_n1442, new_n1444);
not_8  g01068(new_n1444, new_n1445);
xor_4  g01069(new_n1445, new_n1441, new_n1446);
xor_4  g01070(new_n1446, new_n1439, new_n1447);
nor_5  g01071(new_n1447, new_n1426, new_n1448);
xor_4  g01072(new_n1447, new_n1426, new_n1449);
not_8  g01073(new_n1449, new_n1450);
nand_5 g01074(n7862, n2508, new_n1451);
nand_5 g01075(n2509, n1333, new_n1452);
nand_5 g01076(n6038, n3172, new_n1453);
nand_5 g01077(n12720, n7862, new_n1454);
and_5  g01078(new_n1454, new_n1453, new_n1455);
or_5   g01079(new_n1455, new_n1452, new_n1456);
not_8  g01080(new_n1456, new_n1457);
nor_5  g01081(new_n1454, new_n1453, new_n1458);
nor_5  g01082(new_n1458, new_n1457, new_n1459);
nor_5  g01083(new_n1459, new_n1451, new_n1460);
xor_4  g01084(new_n1459, new_n1451, new_n1461);
xor_4  g01085(new_n1429, new_n1428, new_n1462);
xor_4  g01086(new_n1462, new_n1433, new_n1463);
and_5  g01087(new_n1463, new_n1461, new_n1464);
or_5   g01088(new_n1464, new_n1460, new_n1465);
nor_5  g01089(new_n1465, new_n1450, new_n1466);
or_5   g01090(new_n1466, new_n1448, new_n1467);
not_8  g01091(new_n1467, new_n1468);
nand_5 g01092(n12720, n11757, new_n1469);
nand_5 g01093(n5240, n2509, new_n1470);
nand_5 g01094(n11821, n6038, new_n1471_1);
xor_4  g01095(new_n1471_1, new_n1470, new_n1472);
not_8  g01096(new_n1472, new_n1473);
xor_4  g01097(new_n1473, new_n1469, new_n1474);
and_5  g01098(new_n1443, new_n1442, new_n1475);
nor_5  g01099(new_n1445, new_n1441, new_n1476);
or_5   g01100(new_n1476, new_n1475, new_n1477);
not_8  g01101(new_n1477, new_n1478_1);
xor_4  g01102(new_n1478_1, new_n1474, new_n1479);
nor_5  g01103(new_n1446, new_n1439, new_n1480);
or_5   g01104(new_n1480, new_n1437, new_n1481);
not_8  g01105(new_n1481, new_n1482);
nand_5 g01106(n2585, n1333, new_n1483);
nand_5 g01107(n3172, n2508, new_n1484);
xor_4  g01108(new_n1484, new_n1483, new_n1485);
not_8  g01109(new_n1485, new_n1486);
xor_4  g01110(new_n1486, new_n1482, new_n1487);
xor_4  g01111(new_n1487, new_n1479, new_n1488);
nand_5 g01112(new_n1488, new_n1468, new_n1489);
nor_5  g01113(new_n1486, new_n1482, new_n1490);
or_5   g01114(new_n1484, new_n1483, new_n1491);
not_8  g01115(new_n1479, new_n1492);
and_5  g01116(new_n1486, new_n1482, new_n1493);
or_5   g01117(new_n1493, new_n1492, new_n1494);
xor_4  g01118(new_n1494, new_n1491, new_n1495);
or_5   g01119(new_n1495, new_n1490, new_n1496);
not_8  g01120(new_n1496, new_n1497);
or_5   g01121(new_n1471_1, new_n1470, new_n1498);
not_8  g01122(new_n1498, new_n1499);
nand_5 g01123(n11757, n2508, new_n1500);
not_8  g01124(new_n1500, new_n1501);
xor_4  g01125(new_n1501, new_n1499, new_n1502);
nand_5 g01126(n11821, n2509, new_n1503);
nand_5 g01127(n12720, n5240, new_n1504);
nand_5 g01128(n9080, n6038, new_n1505);
xor_4  g01129(new_n1505, new_n1504, new_n1506);
not_8  g01130(new_n1506, new_n1507);
xor_4  g01131(new_n1507, new_n1503, new_n1508);
xor_4  g01132(new_n1508, new_n1502, new_n1509);
not_8  g01133(new_n1509, new_n1510_1);
nor_5  g01134(new_n1473, new_n1469, new_n1511);
and_5  g01135(new_n1478_1, new_n1474, new_n1512_1);
or_5   g01136(new_n1512_1, new_n1511, new_n1513);
not_8  g01137(new_n1513, new_n1514);
nand_5 g01138(n4005, n1333, new_n1515);
nand_5 g01139(n3172, n2585, new_n1516);
nand_5 g01140(n12706, n7862, new_n1517);
xor_4  g01141(new_n1517, new_n1516, new_n1518);
xor_4  g01142(new_n1518, new_n1515, new_n1519);
xor_4  g01143(new_n1519, new_n1514, new_n1520);
xor_4  g01144(new_n1520, new_n1510_1, new_n1521);
xor_4  g01145(new_n1521, new_n1497, new_n1522);
xor_4  g01146(new_n1522, new_n1489, new_n1523_1);
nand_5 g01147(n7862, n4005, new_n1524);
not_8  g01148(new_n1524, new_n1525);
xor_4  g01149(new_n1488, new_n1468, new_n1526);
and_5  g01150(new_n1526, new_n1525, new_n1527);
xor_4  g01151(new_n1463, new_n1461, new_n1528);
not_8  g01152(new_n1528, new_n1529);
xor_4  g01153(new_n1454, new_n1453, new_n1530);
nand_5 g01154(n6038, n1333, new_n1531);
nand_5 g01155(n7862, n2509, new_n1532);
or_5   g01156(new_n1532, new_n1531, new_n1533);
or_5   g01157(new_n1533, new_n1530, new_n1534);
or_5   g01158(new_n1534, new_n1529, new_n1535);
not_8  g01159(new_n1465, new_n1536);
xnor_4 g01160(new_n1536, new_n1450, new_n1537);
or_5   g01161(new_n1537, new_n1535, new_n1538);
xor_4  g01162(new_n1526, new_n1525, new_n1539);
not_8  g01163(new_n1539, new_n1540);
nor_5  g01164(new_n1540, new_n1538, new_n1541);
nor_5  g01165(new_n1541, new_n1527, new_n1542);
xor_4  g01166(new_n1542, new_n1523_1, new_n1543);
not_8  g01167(new_n1543, new_n1544);
nand_5 g01168(n6877, n5105, new_n1545);
and_5  g01169(n6877, n1209, new_n1546);
and_5  g01170(n7354, n2464, new_n1547);
and_5  g01171(new_n1547, new_n1546, new_n1548);
nor_5  g01172(new_n1547, new_n1546, new_n1549);
not_8  g01173(new_n1549, new_n1550);
and_5  g01174(n9400, n7500, new_n1551);
and_5  g01175(new_n1551, new_n1550, new_n1552);
nor_5  g01176(new_n1552, new_n1548, new_n1553);
xor_4  g01177(new_n1553, new_n1545, new_n1554);
not_8  g01178(new_n1554, new_n1555);
nand_5 g01179(n7500, n2464, new_n1556);
not_8  g01180(new_n1556, new_n1557);
nand_5 g01181(n9400, n1209, new_n1558);
nand_5 g01182(n11311, n7354, new_n1559);
xor_4  g01183(new_n1559, new_n1558, new_n1560);
xor_4  g01184(new_n1560, new_n1557, new_n1561);
not_8  g01185(new_n1561, new_n1562);
xor_4  g01186(new_n1562, new_n1555, new_n1563);
xor_4  g01187(new_n1547, new_n1546, new_n1564_1);
nand_5 g01188(n9400, n7354, new_n1565);
nand_5 g01189(n7500, n6877, new_n1566);
or_5   g01190(new_n1566, new_n1565, new_n1567);
or_5   g01191(new_n1567, new_n1564_1, new_n1568);
not_8  g01192(new_n1568, new_n1569);
nand_5 g01193(new_n1569, new_n1563, new_n1570);
nand_5 g01194(n11311, n7500, new_n1571);
not_8  g01195(new_n1571, new_n1572);
nand_5 g01196(n2464, n1209, new_n1573);
nand_5 g01197(n7354, n4187, new_n1574);
xor_4  g01198(new_n1574, new_n1573, new_n1575);
not_8  g01199(new_n1575, new_n1576_1);
xor_4  g01200(new_n1576_1, new_n1572, new_n1577);
nand_5 g01201(n9400, n5105, new_n1578);
not_8  g01202(new_n1578, new_n1579);
and_5  g01203(new_n1559, new_n1558, new_n1580);
nor_5  g01204(new_n1559, new_n1558, new_n1581);
nor_5  g01205(new_n1581, new_n1557, new_n1582);
or_5   g01206(new_n1582, new_n1580, new_n1583);
not_8  g01207(new_n1583, new_n1584);
and_5  g01208(new_n1584, new_n1579, new_n1585);
nor_5  g01209(new_n1584, new_n1579, new_n1586);
or_5   g01210(new_n1586, new_n1585, new_n1587);
xor_4  g01211(new_n1587, new_n1577, new_n1588);
not_8  g01212(new_n1588, new_n1589);
nand_5 g01213(n6877, n4141, new_n1590);
nor_5  g01214(new_n1553, new_n1545, new_n1591);
nor_5  g01215(new_n1562, new_n1555, new_n1592);
or_5   g01216(new_n1592, new_n1591, new_n1593);
not_8  g01217(new_n1593, new_n1594);
xor_4  g01218(new_n1594, new_n1590, new_n1595);
xor_4  g01219(new_n1595, new_n1589, new_n1596);
or_5   g01220(new_n1596, new_n1570, new_n1597);
not_8  g01221(new_n1597, new_n1598);
nand_5 g01222(n6877, n4928, new_n1599);
not_8  g01223(new_n1599, new_n1600);
and_5  g01224(new_n1594, new_n1590, new_n1601);
and_5  g01225(new_n1595, new_n1589, new_n1602);
or_5   g01226(new_n1602, new_n1601, new_n1603);
not_8  g01227(new_n1603, new_n1604);
nand_5 g01228(n11311, n1209, new_n1605);
nand_5 g01229(n7500, n4187, new_n1606);
nand_5 g01230(n7354, n4203, new_n1607);
xor_4  g01231(new_n1607, new_n1606, new_n1608);
not_8  g01232(new_n1608, new_n1609);
xor_4  g01233(new_n1609, new_n1605, new_n1610);
and_5  g01234(new_n1574, new_n1573, new_n1611);
nor_5  g01235(new_n1576_1, new_n1572, new_n1612);
or_5   g01236(new_n1612, new_n1611, new_n1613);
not_8  g01237(new_n1613, new_n1614);
xor_4  g01238(new_n1614, new_n1610, new_n1615);
nor_5  g01239(new_n1587, new_n1577, new_n1616);
or_5   g01240(new_n1616, new_n1585, new_n1617);
not_8  g01241(new_n1617, new_n1618);
nand_5 g01242(n9400, n4141, new_n1619);
nand_5 g01243(n5105, n2464, new_n1620);
xor_4  g01244(new_n1620, new_n1619, new_n1621);
not_8  g01245(new_n1621, new_n1622);
xor_4  g01246(new_n1622, new_n1618, new_n1623);
xor_4  g01247(new_n1623, new_n1615, new_n1624);
xor_4  g01248(new_n1624, new_n1604, new_n1625);
xor_4  g01249(new_n1625, new_n1600, new_n1626);
xor_4  g01250(new_n1626, new_n1598, new_n1627);
not_8  g01251(new_n1627, new_n1628);
nand_5 g01252(n7294, n7236, new_n1629);
not_8  g01253(new_n1629, new_n1630);
nand_5 g01254(n10848, n3992, new_n1631);
nand_5 g01255(n8384, n8028, new_n1632);
nand_5 g01256(n7236, n1980, new_n1633);
and_5  g01257(new_n1633, new_n1632, new_n1634);
nor_5  g01258(new_n1634, new_n1631, new_n1635);
not_8  g01259(new_n1635, new_n1636);
or_5   g01260(new_n1633, new_n1632, new_n1637);
and_5  g01261(new_n1637, new_n1636, new_n1638);
xor_4  g01262(new_n1638, new_n1630, new_n1639);
nand_5 g01263(n8028, n6358, new_n1640);
nand_5 g01264(n10848, n8384, new_n1641);
nand_5 g01265(n3992, n1980, new_n1642);
xnor_4 g01266(new_n1642, new_n1641, new_n1643);
not_8  g01267(new_n1643, new_n1644);
xor_4  g01268(new_n1644, new_n1640, new_n1645);
xor_4  g01269(new_n1645, new_n1639, new_n1646);
not_8  g01270(new_n1646, new_n1647);
xor_4  g01271(new_n1633, new_n1632, new_n1648);
nand_5 g01272(n10848, n7236, new_n1649);
nand_5 g01273(n8028, n3992, new_n1650);
or_5   g01274(new_n1650, new_n1649, new_n1651);
or_5   g01275(new_n1651, new_n1648, new_n1652);
or_5   g01276(new_n1652, new_n1647, new_n1653);
nand_5 g01277(n10848, n6358, new_n1654);
not_8  g01278(new_n1654, new_n1655);
nand_5 g01279(n8384, n1980, new_n1656);
nand_5 g01280(n8028, n5198, new_n1657);
xor_4  g01281(new_n1657, new_n1656, new_n1658_1);
not_8  g01282(new_n1658_1, new_n1659);
xor_4  g01283(new_n1659, new_n1655, new_n1660);
not_8  g01284(new_n1660, new_n1661);
nand_5 g01285(n7294, n3992, new_n1662);
not_8  g01286(new_n1662, new_n1663);
and_5  g01287(new_n1642, new_n1641, new_n1664);
and_5  g01288(new_n1644, new_n1640, new_n1665);
or_5   g01289(new_n1665, new_n1664, new_n1666);
not_8  g01290(new_n1666, new_n1667);
xor_4  g01291(new_n1667, new_n1663, new_n1668);
xor_4  g01292(new_n1668, new_n1661, new_n1669);
nand_5 g01293(n12704, n7236, new_n1670);
nor_5  g01294(new_n1638, new_n1629, new_n1671);
nor_5  g01295(new_n1645, new_n1639, new_n1672);
nor_5  g01296(new_n1672, new_n1671, new_n1673);
not_8  g01297(new_n1673, new_n1674);
xor_4  g01298(new_n1674, new_n1670, new_n1675);
xor_4  g01299(new_n1675, new_n1669, new_n1676);
or_5   g01300(new_n1676, new_n1653, new_n1677);
nand_5 g01301(n7236, n5814, new_n1678);
not_8  g01302(new_n1678, new_n1679);
and_5  g01303(new_n1667, new_n1663, new_n1680);
and_5  g01304(new_n1668, new_n1661, new_n1681);
or_5   g01305(new_n1681, new_n1680, new_n1682);
not_8  g01306(new_n1682, new_n1683);
nand_5 g01307(n8384, n7294, new_n1684);
nand_5 g01308(n12704, n3992, new_n1685);
xor_4  g01309(new_n1685, new_n1684, new_n1686);
not_8  g01310(new_n1686, new_n1687);
xor_4  g01311(new_n1687, new_n1683, new_n1688);
nand_5 g01312(n6358, n1980, new_n1689);
not_8  g01313(new_n1689, new_n1690);
and_5  g01314(new_n1657, new_n1656, new_n1691);
nor_5  g01315(new_n1659, new_n1655, new_n1692);
nor_5  g01316(new_n1692, new_n1691, new_n1693);
xor_4  g01317(new_n1693, new_n1690, new_n1694);
not_8  g01318(new_n1694, new_n1695);
nand_5 g01319(n10848, n5198, new_n1696);
nand_5 g01320(n8028, n1471, new_n1697);
xnor_4 g01321(new_n1697, new_n1696, new_n1698);
xor_4  g01322(new_n1698, new_n1695, new_n1699);
xor_4  g01323(new_n1699, new_n1688, new_n1700);
not_8  g01324(new_n1670, new_n1701);
nor_5  g01325(new_n1674, new_n1701, new_n1702);
nor_5  g01326(new_n1675, new_n1669, new_n1703);
or_5   g01327(new_n1703, new_n1702, new_n1704);
not_8  g01328(new_n1704, new_n1705);
xor_4  g01329(new_n1705, new_n1700, new_n1706);
xor_4  g01330(new_n1706, new_n1679, new_n1707);
not_8  g01331(new_n1707, new_n1708);
xor_4  g01332(new_n1708, new_n1677, new_n1709);
nand_5 g01333(n4805, n2802, new_n1710);
and_5  g01334(n5283, n1564, new_n1711);
and_5  g01335(n4805, n533, new_n1712);
and_5  g01336(new_n1712, new_n1711, new_n1713);
nor_5  g01337(new_n1712, new_n1711, new_n1714);
nand_5 g01338(n11478, n1512, new_n1715);
or_5   g01339(new_n1715, new_n1714, new_n1716);
not_8  g01340(new_n1716, new_n1717);
nor_5  g01341(new_n1717, new_n1713, new_n1718);
xor_4  g01342(new_n1718, new_n1710, new_n1719);
nand_5 g01343(n1564, n137, new_n1720);
nand_5 g01344(n5283, n1512, new_n1721);
nand_5 g01345(n11478, n533, new_n1722);
xnor_4 g01346(new_n1722, new_n1721, new_n1723);
not_8  g01347(new_n1723, new_n1724);
xor_4  g01348(new_n1724, new_n1720, new_n1725);
xor_4  g01349(new_n1725, new_n1719, new_n1726);
not_8  g01350(new_n1726, new_n1727);
xor_4  g01351(new_n1712, new_n1711, new_n1728);
and_5  g01352(n4805, n1512, new_n1729);
and_5  g01353(n11478, n1564, new_n1730);
nand_5 g01354(new_n1730, new_n1729, new_n1731);
or_5   g01355(new_n1731, new_n1728, new_n1732);
not_8  g01356(new_n1732, new_n1733);
nand_5 g01357(new_n1733, new_n1727, new_n1734);
nand_5 g01358(n6806, n4805, new_n1735);
not_8  g01359(new_n1735, new_n1736);
nand_5 g01360(n11478, n2802, new_n1737);
and_5  g01361(new_n1722, new_n1721, new_n1738);
and_5  g01362(new_n1724, new_n1720, new_n1739);
or_5   g01363(new_n1739, new_n1738, new_n1740);
not_8  g01364(new_n1740, new_n1741);
xor_4  g01365(new_n1741, new_n1737, new_n1742);
nand_5 g01366(n1512, n137, new_n1743);
not_8  g01367(new_n1743, new_n1744);
nand_5 g01368(n5283, n533, new_n1745);
nand_5 g01369(n6294, n1564, new_n1746);
xor_4  g01370(new_n1746, new_n1745, new_n1747);
not_8  g01371(new_n1747, new_n1748);
xor_4  g01372(new_n1748, new_n1744, new_n1749);
xor_4  g01373(new_n1749, new_n1742, new_n1750);
xor_4  g01374(new_n1750, new_n1736, new_n1751);
not_8  g01375(new_n1751, new_n1752);
nor_5  g01376(new_n1718, new_n1710, new_n1753);
not_8  g01377(new_n1720, new_n1754);
xor_4  g01378(new_n1724, new_n1754, new_n1755);
and_5  g01379(new_n1755, new_n1719, new_n1756);
or_5   g01380(new_n1756, new_n1753, new_n1757);
not_8  g01381(new_n1757, new_n1758);
xnor_4 g01382(new_n1758, new_n1752, new_n1759);
nor_5  g01383(new_n1759, new_n1734, new_n1760);
not_8  g01384(new_n1760, new_n1761);
nand_5 g01385(n5069, n4805, new_n1762);
not_8  g01386(new_n1762, new_n1763);
nand_5 g01387(n533, n137, new_n1764);
nand_5 g01388(n6294, n1512, new_n1765);
nand_5 g01389(n6797, n1564, new_n1766);
xor_4  g01390(new_n1766, new_n1765, new_n1767);
not_8  g01391(new_n1767, new_n1768);
xor_4  g01392(new_n1768, new_n1764, new_n1769);
and_5  g01393(new_n1746, new_n1745, new_n1770);
nor_5  g01394(new_n1748, new_n1744, new_n1771);
or_5   g01395(new_n1771, new_n1770, new_n1772);
not_8  g01396(new_n1772, new_n1773);
xor_4  g01397(new_n1773, new_n1769, new_n1774);
nand_5 g01398(n11478, n6806, new_n1775);
nand_5 g01399(n5283, n2802, new_n1776);
xor_4  g01400(new_n1776, new_n1775, new_n1777);
xor_4  g01401(new_n1777, new_n1774, new_n1778);
not_8  g01402(new_n1778, new_n1779);
not_8  g01403(new_n1737, new_n1780);
and_5  g01404(new_n1741, new_n1780, new_n1781);
nor_5  g01405(new_n1749, new_n1742, new_n1782);
nor_5  g01406(new_n1782, new_n1781, new_n1783);
xor_4  g01407(new_n1783, new_n1779, new_n1784);
nor_5  g01408(new_n1750, new_n1736, new_n1785);
nor_5  g01409(new_n1757, new_n1752, new_n1786);
or_5   g01410(new_n1786, new_n1785, new_n1787);
not_8  g01411(new_n1787, new_n1788);
xor_4  g01412(new_n1788, new_n1784, new_n1789);
xor_4  g01413(new_n1789, new_n1763, new_n1790);
not_8  g01414(new_n1790, new_n1791);
xor_4  g01415(new_n1791, new_n1761, new_n1792);
xor_4  g01416(new_n1792, new_n1709, new_n1793);
not_8  g01417(new_n1793, new_n1794);
xor_4  g01418(new_n1676, new_n1653, new_n1795);
xor_4  g01419(new_n1732, new_n1727, new_n1796);
not_8  g01420(new_n1652, new_n1797);
xor_4  g01421(new_n1797, new_n1647, new_n1798_1);
and_5  g01422(new_n1798_1, new_n1796, new_n1799);
or_5   g01423(new_n1232, new_n1231, new_n1800);
not_8  g01424(new_n1800, new_n1801);
xor_4  g01425(new_n1730, new_n1729, new_n1802);
nor_5  g01426(new_n1802, new_n1801, new_n1803);
xor_4  g01427(new_n1802, new_n1800, new_n1804);
not_8  g01428(new_n1804, new_n1805);
xnor_4 g01429(new_n1650, new_n1649, new_n1806);
and_5  g01430(new_n1806, new_n1805, new_n1807);
or_5   g01431(new_n1807, new_n1803, new_n1808);
not_8  g01432(new_n1715, new_n1809);
and_5  g01433(new_n1809, new_n1231, new_n1810);
nor_5  g01434(new_n1810, new_n1728, new_n1811);
and_5  g01435(new_n1717, new_n1231, new_n1812);
or_5   g01436(new_n1812, new_n1811, new_n1813);
and_5  g01437(new_n1813, new_n1808, new_n1814);
nor_5  g01438(new_n1812, new_n1811, new_n1815);
xor_4  g01439(new_n1815, new_n1808, new_n1816);
not_8  g01440(new_n1816, new_n1817);
not_8  g01441(new_n1631, new_n1818);
and_5  g01442(new_n1818, new_n1232, new_n1819);
nor_5  g01443(new_n1819, new_n1648, new_n1820);
not_8  g01444(new_n1232, new_n1821);
nor_5  g01445(new_n1636, new_n1821, new_n1822);
or_5   g01446(new_n1822, new_n1820, new_n1823);
and_5  g01447(new_n1823, new_n1817, new_n1824);
or_5   g01448(new_n1824, new_n1814, new_n1825);
not_8  g01449(new_n1825, new_n1826);
xor_4  g01450(new_n1798_1, new_n1796, new_n1827);
not_8  g01451(new_n1827, new_n1828);
nor_5  g01452(new_n1828, new_n1826, new_n1829);
nor_5  g01453(new_n1829, new_n1799, new_n1830);
nor_5  g01454(new_n1830, new_n1795, new_n1831);
xor_4  g01455(new_n1758, new_n1752, new_n1832);
xor_4  g01456(new_n1832, new_n1734, new_n1833);
not_8  g01457(new_n1833, new_n1834);
xor_4  g01458(new_n1830, new_n1795, new_n1835_1);
not_8  g01459(new_n1835_1, new_n1836);
nor_5  g01460(new_n1836, new_n1834, new_n1837);
nor_5  g01461(new_n1837, new_n1831, new_n1838);
xor_4  g01462(new_n1838, new_n1794, new_n1839);
and_5  g01463(new_n1839, new_n1628, new_n1840);
xor_4  g01464(new_n1839, new_n1628, new_n1841);
not_8  g01465(new_n1841, new_n1842);
xor_4  g01466(new_n1596, new_n1570, new_n1843);
not_8  g01467(new_n1843, new_n1844);
xor_4  g01468(new_n1836, new_n1834, new_n1845);
nor_5  g01469(new_n1845, new_n1844, new_n1846);
xor_4  g01470(new_n1845, new_n1843, new_n1847_1);
xor_4  g01471(new_n1569, new_n1563, new_n1848);
not_8  g01472(new_n1848, new_n1849);
xor_4  g01473(new_n1828, new_n1826, new_n1850);
nor_5  g01474(new_n1850, new_n1849, new_n1851);
xor_4  g01475(new_n1850, new_n1848, new_n1852);
xor_4  g01476(new_n1823, new_n1817, new_n1853);
nand_5 g01477(new_n1551, new_n1230, new_n1854);
nor_5  g01478(new_n1854, new_n1550, new_n1855);
not_8  g01479(new_n1564_1, new_n1856);
not_8  g01480(new_n1854, new_n1857);
nor_5  g01481(new_n1857, new_n1856, new_n1858);
nor_5  g01482(new_n1858, new_n1855, new_n1859);
nor_5  g01483(new_n1859, new_n1853, new_n1860);
xor_4  g01484(new_n1859, new_n1853, new_n1861);
xor_4  g01485(new_n1806, new_n1805, new_n1862);
xor_4  g01486(new_n1566, new_n1565, new_n1863);
not_8  g01487(new_n1863, new_n1864);
nor_5  g01488(new_n1864, new_n1862, new_n1865);
or_5   g01489(new_n1234, new_n1230, new_n1866);
not_8  g01490(new_n1866, new_n1867);
xor_4  g01491(new_n1864, new_n1862, new_n1868);
and_5  g01492(new_n1868, new_n1867, new_n1869);
or_5   g01493(new_n1869, new_n1865, new_n1870);
and_5  g01494(new_n1870, new_n1861, new_n1871);
nor_5  g01495(new_n1871, new_n1860, new_n1872);
nor_5  g01496(new_n1872, new_n1852, new_n1873);
nor_5  g01497(new_n1873, new_n1851, new_n1874);
nor_5  g01498(new_n1874, new_n1847_1, new_n1875);
or_5   g01499(new_n1875, new_n1846, new_n1876);
nor_5  g01500(new_n1876, new_n1842, new_n1877);
or_5   g01501(new_n1877, new_n1840, new_n1878);
not_8  g01502(new_n1878, new_n1879);
nand_5 g01503(new_n1624, new_n1604, new_n1880);
nor_5  g01504(new_n1609, new_n1605, new_n1881);
and_5  g01505(new_n1614, new_n1610, new_n1882);
or_5   g01506(new_n1882, new_n1881, new_n1883);
not_8  g01507(new_n1883, new_n1884);
nand_5 g01508(n9400, n4928, new_n1885);
nand_5 g01509(n4141, n2464, new_n1886);
nand_5 g01510(n8236, n6877, new_n1887);
xor_4  g01511(new_n1887, new_n1886, new_n1888);
xor_4  g01512(new_n1888, new_n1885, new_n1889);
xor_4  g01513(new_n1889, new_n1884, new_n1890);
or_5   g01514(new_n1607, new_n1606, new_n1891);
not_8  g01515(new_n1891, new_n1892);
nand_5 g01516(n11311, n5105, new_n1893);
not_8  g01517(new_n1893, new_n1894);
xor_4  g01518(new_n1894, new_n1892, new_n1895);
nand_5 g01519(n7500, n4203, new_n1896);
nand_5 g01520(n4187, n1209, new_n1897);
nand_5 g01521(n12753, n7354, new_n1898);
xor_4  g01522(new_n1898, new_n1897, new_n1899);
not_8  g01523(new_n1899, new_n1900);
xor_4  g01524(new_n1900, new_n1896, new_n1901);
xor_4  g01525(new_n1901, new_n1895, new_n1902);
xor_4  g01526(new_n1902, new_n1890, new_n1903);
not_8  g01527(new_n1903, new_n1904);
nor_5  g01528(new_n1622, new_n1618, new_n1905);
or_5   g01529(new_n1620, new_n1619, new_n1906_1);
not_8  g01530(new_n1615, new_n1907);
and_5  g01531(new_n1622, new_n1618, new_n1908);
or_5   g01532(new_n1908, new_n1907, new_n1909);
xor_4  g01533(new_n1909, new_n1906_1, new_n1910);
nor_5  g01534(new_n1910, new_n1905, new_n1911);
xor_4  g01535(new_n1911, new_n1904, new_n1912);
not_8  g01536(new_n1912, new_n1913);
nor_5  g01537(new_n1913, new_n1880, new_n1914);
and_5  g01538(new_n1913, new_n1880, new_n1915);
or_5   g01539(new_n1915, new_n1914, new_n1916);
and_5  g01540(new_n1625, new_n1600, new_n1917);
and_5  g01541(new_n1626, new_n1598, new_n1918);
nor_5  g01542(new_n1918, new_n1917, new_n1919);
xor_4  g01543(new_n1919, new_n1916, new_n1920);
nand_5 g01544(new_n1705, new_n1700, new_n1921);
nor_5  g01545(new_n1693, new_n1690, new_n1922);
xor_4  g01546(new_n1697, new_n1696, new_n1923);
nor_5  g01547(new_n1923, new_n1695, new_n1924);
or_5   g01548(new_n1924, new_n1922, new_n1925);
nand_5 g01549(n5814, n3992, new_n1926);
not_8  g01550(new_n1926, new_n1927);
nand_5 g01551(n12704, n8384, new_n1928);
nand_5 g01552(n7236, n4903, new_n1929);
xor_4  g01553(new_n1929, new_n1928, new_n1930);
not_8  g01554(new_n1930, new_n1931);
xor_4  g01555(new_n1931, new_n1927, new_n1932);
not_8  g01556(new_n1932, new_n1933);
xor_4  g01557(new_n1933, new_n1925, new_n1934);
not_8  g01558(new_n1934, new_n1935);
or_5   g01559(new_n1697, new_n1696, new_n1936);
nand_5 g01560(n7294, n6358, new_n1937);
not_8  g01561(new_n1937, new_n1938);
xor_4  g01562(new_n1938, new_n1936, new_n1939);
nand_5 g01563(n10848, n1471, new_n1940);
not_8  g01564(new_n1940, new_n1941);
nand_5 g01565(n5198, n1980, new_n1942);
nand_5 g01566(n8028, n7646, new_n1943);
xor_4  g01567(new_n1943, new_n1942, new_n1944);
not_8  g01568(new_n1944, new_n1945);
xor_4  g01569(new_n1945, new_n1941, new_n1946);
xor_4  g01570(new_n1946, new_n1939, new_n1947);
xnor_4 g01571(new_n1947, new_n1935, new_n1948);
nor_5  g01572(new_n1687, new_n1683, new_n1949);
or_5   g01573(new_n1685, new_n1684, new_n1950);
not_8  g01574(new_n1950, new_n1951);
and_5  g01575(new_n1699, new_n1688, new_n1952);
xor_4  g01576(new_n1952, new_n1951, new_n1953);
nor_5  g01577(new_n1953, new_n1949, new_n1954);
xor_4  g01578(new_n1954, new_n1948, new_n1955);
not_8  g01579(new_n1955, new_n1956);
xor_4  g01580(new_n1956, new_n1921, new_n1957);
not_8  g01581(new_n1957, new_n1958);
and_5  g01582(new_n1706, new_n1679, new_n1959);
nor_5  g01583(new_n1708, new_n1677, new_n1960);
nor_5  g01584(new_n1960, new_n1959, new_n1961);
xor_4  g01585(new_n1961, new_n1958, new_n1962);
not_8  g01586(new_n1962, new_n1963);
and_5  g01587(new_n1789, new_n1763, new_n1964);
nor_5  g01588(new_n1791, new_n1761, new_n1965);
or_5   g01589(new_n1965, new_n1964, new_n1966);
not_8  g01590(new_n1966, new_n1967);
nand_5 g01591(new_n1788, new_n1784, new_n1968);
nor_5  g01592(new_n1768, new_n1764, new_n1969);
and_5  g01593(new_n1773, new_n1769, new_n1970);
or_5   g01594(new_n1970, new_n1969, new_n1971);
not_8  g01595(new_n1971, new_n1972);
nand_5 g01596(n11478, n5069, new_n1973);
nand_5 g01597(n6806, n5283, new_n1974);
nand_5 g01598(n12044, n4805, new_n1975);
xor_4  g01599(new_n1975, new_n1974, new_n1976);
xor_4  g01600(new_n1976, new_n1973, new_n1977);
xor_4  g01601(new_n1977, new_n1972, new_n1978);
or_5   g01602(new_n1766, new_n1765, new_n1979);
not_8  g01603(new_n1979, new_n1980_1);
nand_5 g01604(n2802, n137, new_n1981);
not_8  g01605(new_n1981, new_n1982);
xor_4  g01606(new_n1982, new_n1980_1, new_n1983);
nand_5 g01607(n6797, n1512, new_n1984);
nand_5 g01608(n6294, n533, new_n1985);
nand_5 g01609(n3146, n1564, new_n1986);
xor_4  g01610(new_n1986, new_n1985, new_n1987);
not_8  g01611(new_n1987, new_n1988);
xor_4  g01612(new_n1988, new_n1984, new_n1989);
xor_4  g01613(new_n1989, new_n1983, new_n1990);
xor_4  g01614(new_n1990, new_n1978, new_n1991);
not_8  g01615(new_n1991, new_n1992);
and_5  g01616(new_n1777, new_n1774, new_n1993);
or_5   g01617(new_n1776, new_n1775, new_n1994);
not_8  g01618(new_n1994, new_n1995);
or_5   g01619(new_n1783, new_n1779, new_n1996);
not_8  g01620(new_n1996, new_n1997);
xor_4  g01621(new_n1997, new_n1995, new_n1998);
nor_5  g01622(new_n1998, new_n1993, new_n1999);
xor_4  g01623(new_n1999, new_n1992, new_n2000);
not_8  g01624(new_n2000, new_n2001);
xnor_4 g01625(new_n2001, new_n1968, new_n2002);
not_8  g01626(new_n2002, new_n2003);
xor_4  g01627(new_n2003, new_n1967, new_n2004);
xor_4  g01628(new_n2004, new_n1963, new_n2005);
nor_5  g01629(new_n1792, new_n1709, new_n2006);
nor_5  g01630(new_n1838, new_n1794, new_n2007);
or_5   g01631(new_n2007, new_n2006, new_n2008);
xor_4  g01632(new_n2008, new_n2005, new_n2009);
not_8  g01633(new_n2009, new_n2010);
xor_4  g01634(new_n2010, new_n1920, new_n2011);
xnor_4 g01635(new_n2011, new_n1879, new_n2012);
nor_5  g01636(new_n2012, new_n1544, new_n2013);
xor_4  g01637(new_n2012, new_n1543, new_n2014);
xor_4  g01638(new_n1540, new_n1538, new_n2015);
not_8  g01639(new_n2015, new_n2016);
not_8  g01640(new_n1876, new_n2017);
xnor_4 g01641(new_n2017, new_n1842, new_n2018);
nor_5  g01642(new_n2018, new_n2016, new_n2019);
xor_4  g01643(new_n1537, new_n1535, new_n2020);
xor_4  g01644(new_n1874, new_n1847_1, new_n2021);
nor_5  g01645(new_n2021, new_n2020, new_n2022);
xor_4  g01646(new_n2021, new_n2020, new_n2023);
not_8  g01647(new_n2023, new_n2024_1);
xor_4  g01648(new_n1534, new_n1529, new_n2025);
xor_4  g01649(new_n1872, new_n1852, new_n2026);
nor_5  g01650(new_n2026, new_n2025, new_n2027);
xor_4  g01651(new_n1870, new_n1861, new_n2028);
not_8  g01652(new_n2028, new_n2029);
not_8  g01653(new_n1452, new_n2030);
and_5  g01654(new_n2030, new_n1228, new_n2031);
nor_5  g01655(new_n2031, new_n1530, new_n2032);
and_5  g01656(new_n1457, new_n1228, new_n2033);
or_5   g01657(new_n2033, new_n2032, new_n2034);
and_5  g01658(new_n2034, new_n2029, new_n2035);
xor_4  g01659(new_n2034, new_n2029, new_n2036);
nand_5 g01660(new_n1235, new_n1229, new_n2037);
xnor_4 g01661(new_n1532, new_n1531, new_n2038);
and_5  g01662(new_n2038, new_n2037, new_n2039);
xor_4  g01663(new_n1868, new_n1867, new_n2040);
xor_4  g01664(new_n2038, new_n2037, new_n2041);
not_8  g01665(new_n2041, new_n2042);
nor_5  g01666(new_n2042, new_n2040, new_n2043);
or_5   g01667(new_n2043, new_n2039, new_n2044);
and_5  g01668(new_n2044, new_n2036, new_n2045);
or_5   g01669(new_n2045, new_n2035, new_n2046);
not_8  g01670(new_n2046, new_n2047);
xor_4  g01671(new_n2026, new_n2025, new_n2048);
not_8  g01672(new_n2048, new_n2049);
nor_5  g01673(new_n2049, new_n2047, new_n2050);
or_5   g01674(new_n2050, new_n2027, new_n2051);
not_8  g01675(new_n2051, new_n2052);
nor_5  g01676(new_n2052, new_n2024_1, new_n2053);
or_5   g01677(new_n2053, new_n2022, new_n2054);
xor_4  g01678(new_n2018, new_n2016, new_n2055);
not_8  g01679(new_n2055, new_n2056);
nor_5  g01680(new_n2056, new_n2054, new_n2057);
nor_5  g01681(new_n2057, new_n2019, new_n2058);
nor_5  g01682(new_n2058, new_n2014, new_n2059);
or_5   g01683(new_n2059, new_n2013, new_n2060);
nor_5  g01684(new_n2010, new_n1920, new_n2061);
and_5  g01685(new_n2011, new_n1878, new_n2062);
nor_5  g01686(new_n2062, new_n2061, new_n2063);
and_5  g01687(new_n2004, new_n1963, new_n2064);
and_5  g01688(new_n2008, new_n2005, new_n2065);
nor_5  g01689(new_n2065, new_n2064, new_n2066);
not_8  g01690(new_n1489, new_n2067);
and_5  g01691(new_n1522, new_n2067, new_n2068);
nor_5  g01692(new_n1542, new_n1523_1, new_n2069);
nor_5  g01693(new_n2069, new_n2068, new_n2070);
nor_5  g01694(new_n1956, new_n1921, new_n2071);
nor_5  g01695(new_n1961, new_n1958, new_n2072);
nor_5  g01696(new_n2072, new_n2071, new_n2073);
xor_4  g01697(new_n2073, new_n2070, new_n2074);
and_5  g01698(new_n1952, new_n1951, new_n2075);
nor_5  g01699(new_n1954, new_n1948, new_n2076);
nor_5  g01700(new_n2076, new_n2075, new_n2077);
and_5  g01701(new_n1982, new_n1980_1, new_n2078);
and_5  g01702(new_n1989, new_n1983, new_n2079);
nor_5  g01703(new_n2079, new_n2078, new_n2080);
and_5  g01704(n7862, n615, new_n2081);
nand_5 g01705(n4903, n3992, new_n2082);
and_5  g01706(n6806, n137, new_n2083);
xor_4  g01707(new_n2083, new_n2082, new_n2084);
xor_4  g01708(new_n2084, new_n2081, new_n2085);
xor_4  g01709(new_n2085, new_n2080, new_n2086);
nand_5 g01710(n6797, n533, new_n2087_1);
and_5  g01711(n8384, n5814, new_n2088);
xor_4  g01712(new_n2088, new_n2087_1, new_n2089);
nand_5 g01713(n12044, n11478, new_n2090);
and_5  g01714(n7294, n5198, new_n2091);
xor_4  g01715(new_n2091, new_n2090, new_n2092);
xor_4  g01716(new_n2092, new_n2089, new_n2093);
nor_5  g01717(new_n1975, new_n1974, new_n2094);
and_5  g01718(new_n1975, new_n1974, new_n2095);
nor_5  g01719(new_n2095, new_n1973, new_n2096_1);
nor_5  g01720(new_n2096_1, new_n2094, new_n2097);
xor_4  g01721(new_n2097, new_n2093, new_n2098);
nand_5 g01722(n10174, n7354, new_n2099);
nand_5 g01723(n4928, n2464, new_n2100);
and_5  g01724(n11311, n4141, new_n2101);
xor_4  g01725(new_n2101, new_n2100, new_n2102);
and_5  g01726(n4005, n3172, new_n2103);
and_5  g01727(n7236, n1906, new_n2104);
xor_4  g01728(new_n2104, new_n2103, new_n2105);
xor_4  g01729(new_n2105, new_n2102, new_n2106);
xor_4  g01730(new_n2106, new_n2099, new_n2107);
xor_4  g01731(new_n2107, new_n2098, new_n2108);
xor_4  g01732(new_n2108, new_n2086, new_n2109);
xor_4  g01733(new_n2109, new_n2077, new_n2110);
and_5  g01734(new_n1932, new_n1925, new_n2111);
nor_5  g01735(new_n1947, new_n1934, new_n2112);
or_5   g01736(new_n2112, new_n2111, new_n2113);
and_5  g01737(n9080, n2509, new_n2114);
and_5  g01738(new_n1505, new_n1504, new_n2115);
not_8  g01739(new_n1503, new_n2116);
nor_5  g01740(new_n1507, new_n2116, new_n2117);
or_5   g01741(new_n2117, new_n2115, new_n2118);
and_5  g01742(n5240, n2508, new_n2119);
nand_5 g01743(n11757, n2585, new_n2120);
and_5  g01744(n12706, n1333, new_n2121);
xor_4  g01745(new_n2121, new_n2120, new_n2122);
xor_4  g01746(new_n2122, new_n2119, new_n2123);
xor_4  g01747(new_n2123, new_n2118, new_n2124);
xor_4  g01748(new_n2124, new_n2114, new_n2125);
xor_4  g01749(new_n2125, new_n2113, new_n2126);
xor_4  g01750(new_n2126, new_n2110, new_n2127);
nor_5  g01751(new_n1909, new_n1906_1, new_n2128);
nor_5  g01752(new_n1911, new_n1904, new_n2129);
or_5   g01753(new_n2129, new_n2128, new_n2130);
nor_5  g01754(new_n1494, new_n1491, new_n2131_1);
nor_5  g01755(new_n1521, new_n1497, new_n2132);
nor_5  g01756(new_n2132, new_n2131_1, new_n2133);
xor_4  g01757(new_n2133, new_n2130, new_n2134);
nand_5 g01758(new_n1889, new_n1884, new_n2135);
not_8  g01759(new_n1902, new_n2136);
nand_5 g01760(new_n2136, new_n1890, new_n2137);
nand_5 g01761(new_n2137, new_n2135, new_n2138);
and_5  g01762(n12704, n6358, new_n2139);
and_5  g01763(n3146, n1512, new_n2140);
xor_4  g01764(new_n2140, new_n2139, new_n2141);
and_5  g01765(n5105, n4187, new_n2142);
and_5  g01766(n6294, n2802, new_n2143);
xor_4  g01767(new_n2143, new_n2142, new_n2144);
and_5  g01768(n9400, n8236, new_n2145);
and_5  g01769(n1980, n1471, new_n2146);
xor_4  g01770(new_n2146, new_n2145, new_n2147);
xor_4  g01771(new_n2147, new_n2144, new_n2148);
xor_4  g01772(new_n2148, new_n2141, new_n2149);
nand_5 g01773(n12720, n11821, new_n2150);
and_5  g01774(n4938, n1564, new_n2151);
and_5  g01775(n5694, n4805, new_n2152);
xor_4  g01776(new_n2152, new_n2151, new_n2153);
xor_4  g01777(new_n2153, new_n2150, new_n2154);
xor_4  g01778(new_n2154, new_n2149, new_n2155);
and_5  g01779(new_n1929, new_n1928, new_n2156);
nor_5  g01780(new_n1931, new_n1927, new_n2157);
nor_5  g01781(new_n2157, new_n2156, new_n2158);
and_5  g01782(new_n1501, new_n1499, new_n2159);
and_5  g01783(new_n1508, new_n1502, new_n2160);
nor_5  g01784(new_n2160, new_n2159, new_n2161);
xor_4  g01785(new_n2161, new_n2158, new_n2162);
xor_4  g01786(new_n2162, new_n2155, new_n2163);
xor_4  g01787(new_n2163, new_n2138, new_n2164);
and_5  g01788(new_n1997, new_n1995, new_n2165);
nor_5  g01789(new_n1999, new_n1992, new_n2166);
or_5   g01790(new_n2166, new_n2165, new_n2167);
nand_5 g01791(new_n1977, new_n1972, new_n2168);
not_8  g01792(new_n1990, new_n2169);
nand_5 g01793(new_n2169, new_n1978, new_n2170);
nand_5 g01794(new_n2170, new_n2168, new_n2171);
nor_5  g01795(new_n1937, new_n1936, new_n2172);
nor_5  g01796(new_n1946, new_n1939, new_n2173);
or_5   g01797(new_n2173, new_n2172, new_n2174);
nand_5 g01798(n4203, n1209, new_n2175);
nand_5 g01799(n6826, n6038, new_n2176);
and_5  g01800(n5283, n5069, new_n2177);
xor_4  g01801(new_n2177, new_n2176, new_n2178);
xor_4  g01802(new_n2178, new_n2175, new_n2179);
xor_4  g01803(new_n2179, new_n2174, new_n2180);
and_5  g01804(new_n1986, new_n1985, new_n2181);
not_8  g01805(new_n1984, new_n2182);
nor_5  g01806(new_n1988, new_n2182, new_n2183);
or_5   g01807(new_n2183, new_n2181, new_n2184);
and_5  g01808(new_n1943, new_n1942, new_n2185);
nor_5  g01809(new_n1945, new_n1941, new_n2186);
or_5   g01810(new_n2186, new_n2185, new_n2187);
nor_5  g01811(new_n1887, new_n1886, new_n2188);
and_5  g01812(new_n1887, new_n1886, new_n2189);
nor_5  g01813(new_n2189, new_n1885, new_n2190);
nor_5  g01814(new_n2190, new_n2188, new_n2191);
xor_4  g01815(new_n2191, new_n2187, new_n2192);
xor_4  g01816(new_n2192, new_n2184, new_n2193);
xor_4  g01817(new_n2193, new_n2180, new_n2194);
xor_4  g01818(new_n2194, new_n2171, new_n2195);
xor_4  g01819(new_n2195, new_n2167, new_n2196);
xor_4  g01820(new_n2196, new_n2164, new_n2197);
xor_4  g01821(new_n2197, new_n2134, new_n2198);
xor_4  g01822(new_n2198, new_n2127, new_n2199);
xor_4  g01823(new_n2199, new_n2074, new_n2200);
xor_4  g01824(new_n2200, new_n2066, new_n2201);
and_5  g01825(new_n1894, new_n1892, new_n2202);
and_5  g01826(new_n1901, new_n1895, new_n2203);
nor_5  g01827(new_n2203, new_n2202, new_n2204);
nand_5 g01828(n6877, n783, new_n2205);
and_5  g01829(n8028, n4722, new_n2206);
xor_4  g01830(new_n2206, new_n2205, new_n2207);
xor_4  g01831(new_n2207, new_n2204, new_n2208);
nor_5  g01832(new_n1919, new_n1916, new_n2209);
or_5   g01833(new_n2209, new_n1914, new_n2210);
and_5  g01834(n10848, n7646, new_n2211);
xor_4  g01835(new_n2211, new_n2210, new_n2212);
xor_4  g01836(new_n2212, new_n2208, new_n2213);
nor_5  g01837(new_n2001, new_n1968, new_n2214);
nor_5  g01838(new_n2002, new_n1967, new_n2215);
nor_5  g01839(new_n2215, new_n2214, new_n2216);
and_5  g01840(new_n1519, new_n1514, new_n2217);
and_5  g01841(new_n1520, new_n1510_1, new_n2218);
or_5   g01842(new_n2218, new_n2217, new_n2219);
and_5  g01843(new_n1898, new_n1897, new_n2220);
not_8  g01844(new_n1896, new_n2221);
nor_5  g01845(new_n1900, new_n2221, new_n2222);
or_5   g01846(new_n2222, new_n2220, new_n2223);
nand_5 g01847(n12753, n7500, new_n2224);
nor_5  g01848(new_n1517, new_n1516, new_n2225);
and_5  g01849(new_n1517, new_n1516, new_n2226_1);
nor_5  g01850(new_n2226_1, new_n1515, new_n2227);
nor_5  g01851(new_n2227, new_n2225, new_n2228);
xor_4  g01852(new_n2228, new_n2224, new_n2229);
xor_4  g01853(new_n2229, new_n2223, new_n2230);
xor_4  g01854(new_n2230, new_n2219, new_n2231);
xor_4  g01855(new_n2231, new_n2216, new_n2232);
xor_4  g01856(new_n2232, new_n2213, new_n2233);
xor_4  g01857(new_n2233, new_n2201, new_n2234);
xor_4  g01858(new_n2234, new_n2063, new_n2235);
xor_4  g01859(new_n2235, new_n2060, n671);
nand_5 g01860(n11917, n4312, new_n2237);
not_8  g01861(new_n2237, new_n2238);
nand_5 g01862(n12705, n4921, new_n2239);
nand_5 g01863(n12025, n9956, new_n2240);
xor_4  g01864(new_n2240, new_n2239, new_n2241);
xor_4  g01865(new_n2241, new_n2238, new_n2242);
not_8  g01866(new_n2242, new_n2243);
nand_5 g01867(n12705, n9956, new_n2244);
nand_5 g01868(n11917, n1097, new_n2245);
and_5  g01869(new_n2245, new_n2244, new_n2246);
nor_5  g01870(new_n2245, new_n2244, new_n2247);
nand_5 g01871(n4921, n4312, new_n2248);
not_8  g01872(new_n2248, new_n2249);
nor_5  g01873(new_n2249, new_n2247, new_n2250);
nor_5  g01874(new_n2250, new_n2246, new_n2251);
xor_4  g01875(new_n2251, new_n2243, new_n2252);
not_8  g01876(new_n2252, new_n2253_1);
nand_5 g01877(n5964, n2577, new_n2254);
nand_5 g01878(n3842, n1097, new_n2255);
xor_4  g01879(new_n2255, new_n2254, new_n2256);
xor_4  g01880(new_n2256, new_n2253_1, new_n2257);
and_5  g01881(n5964, n3842, new_n2258);
nand_5 g01882(n9956, n4312, new_n2259);
nand_5 g01883(n11917, n5964, new_n2260);
and_5  g01884(new_n2260, new_n2259, new_n2261);
nor_5  g01885(new_n2260, new_n2259, new_n2262);
nand_5 g01886(n4921, n1097, new_n2263);
not_8  g01887(new_n2263, new_n2264);
nor_5  g01888(new_n2264, new_n2262, new_n2265);
or_5   g01889(new_n2265, new_n2261, new_n2266);
not_8  g01890(new_n2266, new_n2267);
and_5  g01891(new_n2267, new_n2258, new_n2268);
nor_5  g01892(new_n2267, new_n2258, new_n2269);
or_5   g01893(new_n2269, new_n2268, new_n2270);
xor_4  g01894(new_n2245, new_n2244, new_n2271);
xor_4  g01895(new_n2271, new_n2248, new_n2272);
nor_5  g01896(new_n2272, new_n2270, new_n2273);
or_5   g01897(new_n2273, new_n2268, new_n2274);
xor_4  g01898(new_n2274, new_n2257, new_n2275);
nand_5 g01899(n5305, n2577, new_n2276);
not_8  g01900(new_n2276, new_n2277);
xor_4  g01901(new_n2272, new_n2270, new_n2278_1);
nor_5  g01902(new_n2278_1, new_n2277, new_n2279);
xor_4  g01903(new_n2278_1, new_n2277, new_n2280);
not_8  g01904(new_n2280, new_n2281);
nand_5 g01905(n5305, n3842, new_n2282);
nand_5 g01906(n9956, n1097, new_n2283);
nand_5 g01907(n11917, n5305, new_n2284);
nor_5  g01908(new_n2284, new_n2283, new_n2285);
and_5  g01909(new_n2284, new_n2283, new_n2286);
nand_5 g01910(n5964, n4921, new_n2287);
nor_5  g01911(new_n2287, new_n2286, new_n2288);
nor_5  g01912(new_n2288, new_n2285, new_n2289);
nor_5  g01913(new_n2289, new_n2282, new_n2290);
xor_4  g01914(new_n2289, new_n2282, new_n2291);
not_8  g01915(new_n2291, new_n2292);
xor_4  g01916(new_n2260, new_n2259, new_n2293);
xor_4  g01917(new_n2293, new_n2263, new_n2294);
nor_5  g01918(new_n2294, new_n2292, new_n2295);
or_5   g01919(new_n2295, new_n2290, new_n2296);
nor_5  g01920(new_n2296, new_n2281, new_n2297);
or_5   g01921(new_n2297, new_n2279, new_n2298);
not_8  g01922(new_n2298, new_n2299);
nand_5 g01923(new_n2299, new_n2275, new_n2300);
nor_5  g01924(new_n2241, new_n2238, new_n2301_1);
nor_5  g01925(new_n2251, new_n2243, new_n2302);
or_5   g01926(new_n2302, new_n2301_1, new_n2303);
not_8  g01927(new_n2303, new_n2304);
nand_5 g01928(n9637, n5964, new_n2305);
not_8  g01929(new_n2305, new_n2306);
nand_5 g01930(n2577, n1097, new_n2307);
nand_5 g01931(n5305, n1835, new_n2308);
xor_4  g01932(new_n2308, new_n2307, new_n2309);
not_8  g01933(new_n2309, new_n2310);
xor_4  g01934(new_n2310, new_n2306, new_n2311);
not_8  g01935(new_n2311, new_n2312);
nor_5  g01936(new_n2312, new_n2304, new_n2313);
and_5  g01937(new_n2312, new_n2304, new_n2314);
or_5   g01938(new_n2314, new_n2313, new_n2315);
or_5   g01939(new_n2240, new_n2239, new_n2316_1);
not_8  g01940(new_n2316_1, new_n2317);
and_5  g01941(n4312, n3842, new_n2318);
xor_4  g01942(new_n2318, new_n2317, new_n2319);
nand_5 g01943(n12025, n4921, new_n2320);
not_8  g01944(new_n2320, new_n2321);
nand_5 g01945(n12705, n11917, new_n2322);
nand_5 g01946(n11257, n9956, new_n2323);
xor_4  g01947(new_n2323, new_n2322, new_n2324);
not_8  g01948(new_n2324, new_n2325);
xor_4  g01949(new_n2325, new_n2321, new_n2326);
xor_4  g01950(new_n2326, new_n2319, new_n2327);
not_8  g01951(new_n2327, new_n2328);
xor_4  g01952(new_n2328, new_n2315, new_n2329);
and_5  g01953(new_n2256, new_n2253_1, new_n2330);
or_5   g01954(new_n2255, new_n2254, new_n2331);
not_8  g01955(new_n2331, new_n2332);
nand_5 g01956(new_n2274, new_n2257, new_n2333);
not_8  g01957(new_n2333, new_n2334);
xor_4  g01958(new_n2334, new_n2332, new_n2335);
nor_5  g01959(new_n2335, new_n2330, new_n2336);
xor_4  g01960(new_n2336, new_n2329, new_n2337);
not_8  g01961(new_n2337, new_n2338);
xor_4  g01962(new_n2338, new_n2300, new_n2339);
not_8  g01963(new_n2339, new_n2340);
nand_5 g01964(n9637, n5305, new_n2341);
not_8  g01965(new_n2341, new_n2342);
xor_4  g01966(new_n2299, new_n2275, new_n2343);
and_5  g01967(new_n2343, new_n2342, new_n2344);
and_5  g01968(new_n2294, new_n2292, new_n2345);
or_5   g01969(new_n2345, new_n2295, new_n2346);
xor_4  g01970(new_n2284, new_n2283, new_n2347_1);
nand_5 g01971(n9956, n5964, new_n2348);
nand_5 g01972(n5305, n4921, new_n2349);
or_5   g01973(new_n2349, new_n2348, new_n2350);
or_5   g01974(new_n2350, new_n2347_1, new_n2351);
or_5   g01975(new_n2351, new_n2346, new_n2352);
xor_4  g01976(new_n2296, new_n2281, new_n2353);
or_5   g01977(new_n2353, new_n2352, new_n2354);
xor_4  g01978(new_n2343, new_n2342, new_n2355);
not_8  g01979(new_n2355, new_n2356);
nor_5  g01980(new_n2356, new_n2354, new_n2357);
nor_5  g01981(new_n2357, new_n2344, new_n2358);
xor_4  g01982(new_n2358, new_n2340, new_n2359);
not_8  g01983(new_n2359, new_n2360);
nand_5 g01984(n8759, n8065, new_n2361);
not_8  g01985(new_n2361, new_n2362);
nand_5 g01986(n7436, n6126, new_n2363);
nand_5 g01987(n9241, n3719, new_n2364);
nand_5 g01988(n8276, n3602, new_n2365);
xor_4  g01989(new_n2365, new_n2364, new_n2366);
not_8  g01990(new_n2366, new_n2367);
xor_4  g01991(new_n2367, new_n2363, new_n2368);
nand_5 g01992(n8276, n3719, new_n2369);
nand_5 g01993(n12299, n6126, new_n2370);
and_5  g01994(new_n2370, new_n2369, new_n2371);
nor_5  g01995(new_n2370, new_n2369, new_n2372);
nand_5 g01996(n7436, n3602, new_n2373);
not_8  g01997(new_n2373, new_n2374);
nor_5  g01998(new_n2374, new_n2372, new_n2375);
or_5   g01999(new_n2375, new_n2371, new_n2376);
not_8  g02000(new_n2376, new_n2377);
xor_4  g02001(new_n2377, new_n2368, new_n2378);
nand_5 g02002(n10439, n6776, new_n2379);
nand_5 g02003(n12299, n8595, new_n2380);
xor_4  g02004(new_n2380, new_n2379, new_n2381);
xor_4  g02005(new_n2381, new_n2378, new_n2382);
nand_5 g02006(n8595, n6776, new_n2383_1);
nand_5 g02007(n7436, n3719, new_n2384);
nand_5 g02008(n6776, n6126, new_n2385);
and_5  g02009(new_n2385, new_n2384, new_n2386);
nor_5  g02010(new_n2385, new_n2384, new_n2387);
nand_5 g02011(n12299, n3602, new_n2388);
not_8  g02012(new_n2388, new_n2389);
nor_5  g02013(new_n2389, new_n2387, new_n2390);
nor_5  g02014(new_n2390, new_n2386, new_n2391);
not_8  g02015(new_n2391, new_n2392);
nor_5  g02016(new_n2392, new_n2383_1, new_n2393_1);
xor_4  g02017(new_n2392, new_n2383_1, new_n2394);
xor_4  g02018(new_n2370, new_n2369, new_n2395);
xor_4  g02019(new_n2395, new_n2374, new_n2396);
and_5  g02020(new_n2396, new_n2394, new_n2397);
or_5   g02021(new_n2397, new_n2393_1, new_n2398);
xor_4  g02022(new_n2398, new_n2382, new_n2399);
nand_5 g02023(n10439, n8759, new_n2400);
not_8  g02024(new_n2400, new_n2401);
xor_4  g02025(new_n2396, new_n2394, new_n2402);
nor_5  g02026(new_n2402, new_n2401, new_n2403);
xor_4  g02027(new_n2402, new_n2401, new_n2404);
not_8  g02028(new_n2404, new_n2405);
nand_5 g02029(n8759, n8595, new_n2406);
and_5  g02030(n12299, n3719, new_n2407);
and_5  g02031(n8759, n6126, new_n2408);
and_5  g02032(new_n2408, new_n2407, new_n2409);
nor_5  g02033(new_n2408, new_n2407, new_n2410);
nand_5 g02034(n6776, n3602, new_n2411);
nor_5  g02035(new_n2411, new_n2410, new_n2412);
nor_5  g02036(new_n2412, new_n2409, new_n2413);
nor_5  g02037(new_n2413, new_n2406, new_n2414);
not_8  g02038(new_n2406, new_n2415);
xor_4  g02039(new_n2413, new_n2415, new_n2416);
not_8  g02040(new_n2416, new_n2417);
xor_4  g02041(new_n2385, new_n2384, new_n2418);
xor_4  g02042(new_n2418, new_n2389, new_n2419);
and_5  g02043(new_n2419, new_n2417, new_n2420);
or_5   g02044(new_n2420, new_n2414, new_n2421);
nor_5  g02045(new_n2421, new_n2405, new_n2422);
or_5   g02046(new_n2422, new_n2403, new_n2423);
not_8  g02047(new_n2423, new_n2424);
xor_4  g02048(new_n2424, new_n2399, new_n2425_1);
and_5  g02049(new_n2425_1, new_n2362, new_n2426);
nor_5  g02050(new_n2419, new_n2417, new_n2427);
or_5   g02051(new_n2427, new_n2420, new_n2428);
xor_4  g02052(new_n2408, new_n2407, new_n2429);
nand_5 g02053(n6776, n3719, new_n2430);
nand_5 g02054(n8759, n3602, new_n2431_1);
or_5   g02055(new_n2431_1, new_n2430, new_n2432);
or_5   g02056(new_n2432, new_n2429, new_n2433_1);
or_5   g02057(new_n2433_1, new_n2428, new_n2434_1);
xor_4  g02058(new_n2421, new_n2405, new_n2435);
or_5   g02059(new_n2435, new_n2434_1, new_n2436);
not_8  g02060(new_n2436, new_n2437);
xor_4  g02061(new_n2425_1, new_n2362, new_n2438);
and_5  g02062(new_n2438, new_n2437, new_n2439);
or_5   g02063(new_n2439, new_n2426, new_n2440);
not_8  g02064(new_n2440, new_n2441);
nand_5 g02065(new_n2424, new_n2399, new_n2442);
nor_5  g02066(new_n2367, new_n2363, new_n2443);
and_5  g02067(new_n2377, new_n2368, new_n2444);
or_5   g02068(new_n2444, new_n2443, new_n2445);
nand_5 g02069(n8065, n6776, new_n2446);
not_8  g02070(new_n2446, new_n2447);
nand_5 g02071(n12299, n10439, new_n2448);
nand_5 g02072(n10391, n8759, new_n2449);
xor_4  g02073(new_n2449, new_n2448, new_n2450);
not_8  g02074(new_n2450, new_n2451);
xor_4  g02075(new_n2451, new_n2447, new_n2452);
not_8  g02076(new_n2452, new_n2453);
xor_4  g02077(new_n2453, new_n2445, new_n2454);
or_5   g02078(new_n2365, new_n2364, new_n2455);
not_8  g02079(new_n2455, new_n2456);
nand_5 g02080(n8595, n7436, new_n2457);
not_8  g02081(new_n2457, new_n2458);
xor_4  g02082(new_n2458, new_n2456, new_n2459);
and_5  g02083(n9241, n3602, new_n2460);
nand_5 g02084(n8276, n6126, new_n2461);
nand_5 g02085(n10510, n3719, new_n2462);
xor_4  g02086(new_n2462, new_n2461, new_n2463);
xor_4  g02087(new_n2463, new_n2460, new_n2464_1);
xor_4  g02088(new_n2464_1, new_n2459, new_n2465);
xor_4  g02089(new_n2465, new_n2454, new_n2466);
not_8  g02090(new_n2466, new_n2467);
and_5  g02091(new_n2381, new_n2378, new_n2468);
or_5   g02092(new_n2380, new_n2379, new_n2469);
not_8  g02093(new_n2469, new_n2470);
nand_5 g02094(new_n2398, new_n2382, new_n2471);
not_8  g02095(new_n2471, new_n2472);
xor_4  g02096(new_n2472, new_n2470, new_n2473);
nor_5  g02097(new_n2473, new_n2468, new_n2474);
xor_4  g02098(new_n2474, new_n2467, new_n2475);
not_8  g02099(new_n2475, new_n2476);
xor_4  g02100(new_n2476, new_n2442, new_n2477);
not_8  g02101(new_n2477, new_n2478);
xor_4  g02102(new_n2478, new_n2441, new_n2479);
not_8  g02103(new_n2479, new_n2480);
nand_5 g02104(n12648, n4826, new_n2481);
nand_5 g02105(n10545, n7733, new_n2482);
nand_5 g02106(n12925, n7690, new_n2483);
xor_4  g02107(new_n2483, new_n2482, new_n2484);
not_8  g02108(new_n2484, new_n2485);
xor_4  g02109(new_n2485, new_n2481, new_n2486);
nand_5 g02110(n12925, n10545, new_n2487);
nand_5 g02111(n4826, n2530, new_n2488);
and_5  g02112(new_n2488, new_n2487, new_n2489);
nand_5 g02113(n12648, n7733, new_n2490);
not_8  g02114(new_n2490, new_n2491);
xor_4  g02115(new_n2488, new_n2487, new_n2492);
not_8  g02116(new_n2492, new_n2493);
nor_5  g02117(new_n2493, new_n2491, new_n2494);
or_5   g02118(new_n2494, new_n2489, new_n2495);
not_8  g02119(new_n2495, new_n2496);
xor_4  g02120(new_n2496, new_n2486, new_n2497);
nand_5 g02121(n8476, n4970, new_n2498_1);
nand_5 g02122(n7610, n2530, new_n2499);
xor_4  g02123(new_n2499, new_n2498_1, new_n2500);
xor_4  g02124(new_n2500, new_n2497, new_n2501);
not_8  g02125(new_n2501, new_n2502);
nand_5 g02126(n8476, n7610, new_n2503);
not_8  g02127(new_n2503, new_n2504);
nand_5 g02128(n12925, n12648, new_n2505);
nand_5 g02129(n8476, n4826, new_n2506);
and_5  g02130(new_n2506, new_n2505, new_n2507_1);
nand_5 g02131(n7733, n2530, new_n2508_1);
not_8  g02132(new_n2508_1, new_n2509_1);
xor_4  g02133(new_n2506, new_n2505, new_n2510);
not_8  g02134(new_n2510, new_n2511);
nor_5  g02135(new_n2511, new_n2509_1, new_n2512_1);
or_5   g02136(new_n2512_1, new_n2507_1, new_n2513);
not_8  g02137(new_n2513, new_n2514);
and_5  g02138(new_n2514, new_n2504, new_n2515_1);
xor_4  g02139(new_n2514, new_n2504, new_n2516);
xor_4  g02140(new_n2493, new_n2490, new_n2517);
and_5  g02141(new_n2517, new_n2516, new_n2518);
nor_5  g02142(new_n2518, new_n2515_1, new_n2519);
xor_4  g02143(new_n2519, new_n2502, new_n2520);
not_8  g02144(new_n2520, new_n2521);
nand_5 g02145(n5331, n4970, new_n2522_1);
nand_5 g02146(n7610, n5331, new_n2523);
not_8  g02147(new_n2523, new_n2524);
nand_5 g02148(n12925, n2530, new_n2525);
nand_5 g02149(n5331, n4826, new_n2526);
nand_5 g02150(new_n2526, new_n2525, new_n2527);
not_8  g02151(new_n2527, new_n2528);
nor_5  g02152(new_n2526, new_n2525, new_n2529);
nand_5 g02153(n8476, n7733, new_n2530_1);
not_8  g02154(new_n2530_1, new_n2531);
nor_5  g02155(new_n2531, new_n2529, new_n2532);
or_5   g02156(new_n2532, new_n2528, new_n2533);
not_8  g02157(new_n2533, new_n2534);
and_5  g02158(new_n2534, new_n2524, new_n2535);
xor_4  g02159(new_n2534, new_n2524, new_n2536);
xor_4  g02160(new_n2511, new_n2508_1, new_n2537);
and_5  g02161(new_n2537, new_n2536, new_n2538);
or_5   g02162(new_n2538, new_n2535, new_n2539);
not_8  g02163(new_n2539, new_n2540);
nand_5 g02164(new_n2540, new_n2522_1, new_n2541);
xor_4  g02165(new_n2517, new_n2516, new_n2542);
not_8  g02166(new_n2522_1, new_n2543);
xor_4  g02167(new_n2540, new_n2543, new_n2544);
or_5   g02168(new_n2544, new_n2542, new_n2545);
and_5  g02169(new_n2545, new_n2541, new_n2546);
not_8  g02170(new_n2546, new_n2547);
or_5   g02171(new_n2547, new_n2521, new_n2548);
and_5  g02172(new_n2500, new_n2497, new_n2549);
or_5   g02173(new_n2499, new_n2498_1, new_n2550);
not_8  g02174(new_n2550, new_n2551_1);
or_5   g02175(new_n2519, new_n2502, new_n2552);
not_8  g02176(new_n2552, new_n2553);
xor_4  g02177(new_n2553, new_n2551_1, new_n2554);
or_5   g02178(new_n2554, new_n2549, new_n2555);
or_5   g02179(new_n2483, new_n2482, new_n2556);
not_8  g02180(new_n2556, new_n2557);
nand_5 g02181(n12648, n7610, new_n2558_1);
not_8  g02182(new_n2558_1, new_n2559);
xor_4  g02183(new_n2559, new_n2557, new_n2560);
nand_5 g02184(n7733, n7690, new_n2561);
nand_5 g02185(n10545, n4826, new_n2562);
nand_5 g02186(n12925, n3616, new_n2563);
xor_4  g02187(new_n2563, new_n2562, new_n2564_1);
not_8  g02188(new_n2564_1, new_n2565);
xor_4  g02189(new_n2565, new_n2561, new_n2566);
xor_4  g02190(new_n2566, new_n2560, new_n2567);
nor_5  g02191(new_n2485, new_n2481, new_n2568);
and_5  g02192(new_n2496, new_n2486, new_n2569);
or_5   g02193(new_n2569, new_n2568, new_n2570);
not_8  g02194(new_n2570, new_n2571);
nand_5 g02195(n8476, n503, new_n2572);
not_8  g02196(new_n2572, new_n2573);
nand_5 g02197(n4970, n2530, new_n2574);
nand_5 g02198(n10965, n5331, new_n2575);
xor_4  g02199(new_n2575, new_n2574, new_n2576);
not_8  g02200(new_n2576, new_n2577_1);
xor_4  g02201(new_n2577_1, new_n2573, new_n2578);
xor_4  g02202(new_n2578, new_n2571, new_n2579);
xor_4  g02203(new_n2579, new_n2567, new_n2580);
xor_4  g02204(new_n2580, new_n2555, new_n2581_1);
not_8  g02205(new_n2581_1, new_n2582);
xor_4  g02206(new_n2582, new_n2548, new_n2583);
not_8  g02207(new_n2583, new_n2584);
nand_5 g02208(n5331, n503, new_n2585_1);
not_8  g02209(new_n2585_1, new_n2586);
xor_4  g02210(new_n2547, new_n2521, new_n2587);
and_5  g02211(new_n2587, new_n2586, new_n2588);
xor_4  g02212(new_n2511, new_n2509_1, new_n2589);
xor_4  g02213(new_n2589, new_n2536, new_n2590);
nand_5 g02214(n12925, n5331, new_n2591);
not_8  g02215(new_n2591, new_n2592);
nor_5  g02216(new_n2592, new_n2530_1, new_n2593);
nor_5  g02217(new_n2593, new_n2527, new_n2594);
or_5   g02218(new_n2594, new_n2529, new_n2595);
not_8  g02219(new_n2595, new_n2596);
or_5   g02220(new_n2596, new_n2530_1, new_n2597);
or_5   g02221(new_n2597, new_n2590, new_n2598);
xor_4  g02222(new_n2544, new_n2542, new_n2599);
or_5   g02223(new_n2599, new_n2598, new_n2600);
not_8  g02224(new_n2600, new_n2601);
xor_4  g02225(new_n2587, new_n2586, new_n2602);
and_5  g02226(new_n2602, new_n2601, new_n2603);
nor_5  g02227(new_n2603, new_n2588, new_n2604);
xor_4  g02228(new_n2604, new_n2584, new_n2605);
not_8  g02229(new_n2605, new_n2606);
nand_5 g02230(n4086, n2393, new_n2607);
nand_5 g02231(n5860, n405, new_n2608);
nand_5 g02232(n8433, n3986, new_n2609);
xor_4  g02233(new_n2609, new_n2608, new_n2610);
not_8  g02234(new_n2610, new_n2611);
xor_4  g02235(new_n2611, new_n2607, new_n2612);
nand_5 g02236(n8433, n5860, new_n2613);
nand_5 g02237(n11892, n4086, new_n2614);
and_5  g02238(new_n2614, new_n2613, new_n2615);
nand_5 g02239(n2393, n405, new_n2616);
not_8  g02240(new_n2616, new_n2617);
xor_4  g02241(new_n2614, new_n2613, new_n2618);
not_8  g02242(new_n2618, new_n2619);
nor_5  g02243(new_n2619, new_n2617, new_n2620);
or_5   g02244(new_n2620, new_n2615, new_n2621);
not_8  g02245(new_n2621, new_n2622);
xor_4  g02246(new_n2622, new_n2612, new_n2623);
nand_5 g02247(n7388, n6611, new_n2624_1);
nand_5 g02248(n11892, n217, new_n2625);
xor_4  g02249(new_n2625, new_n2624_1, new_n2626);
xor_4  g02250(new_n2626, new_n2623, new_n2627);
not_8  g02251(new_n2627, new_n2628);
nand_5 g02252(n7388, n217, new_n2629);
not_8  g02253(new_n2629, new_n2630);
nand_5 g02254(n8433, n2393, new_n2631);
nand_5 g02255(n7388, n4086, new_n2632);
and_5  g02256(new_n2632, new_n2631, new_n2633);
nand_5 g02257(n11892, n405, new_n2634);
xnor_4 g02258(new_n2632, new_n2631, new_n2635);
not_8  g02259(new_n2635, new_n2636);
and_5  g02260(new_n2636, new_n2634, new_n2637);
or_5   g02261(new_n2637, new_n2633, new_n2638);
not_8  g02262(new_n2638, new_n2639);
and_5  g02263(new_n2639, new_n2630, new_n2640);
xor_4  g02264(new_n2639, new_n2630, new_n2641);
xor_4  g02265(new_n2619, new_n2616, new_n2642);
and_5  g02266(new_n2642, new_n2641, new_n2643);
nor_5  g02267(new_n2643, new_n2640, new_n2644);
xor_4  g02268(new_n2644, new_n2628, new_n2645);
not_8  g02269(new_n2645, new_n2646);
nand_5 g02270(n7965, n6611, new_n2647);
xor_4  g02271(new_n2642, new_n2641, new_n2648);
not_8  g02272(new_n2648, new_n2649);
nor_5  g02273(new_n2649, new_n2647, new_n2650);
xor_4  g02274(new_n2649, new_n2647, new_n2651);
nand_5 g02275(n7965, n217, new_n2652);
and_5  g02276(n11892, n8433, new_n2653);
and_5  g02277(n7965, n4086, new_n2654);
and_5  g02278(new_n2654, new_n2653, new_n2655);
nor_5  g02279(new_n2654, new_n2653, new_n2656);
nand_5 g02280(n7388, n405, new_n2657);
nor_5  g02281(new_n2657, new_n2656, new_n2658);
nor_5  g02282(new_n2658, new_n2655, new_n2659);
or_5   g02283(new_n2659, new_n2652, new_n2660);
not_8  g02284(new_n2652, new_n2661);
xor_4  g02285(new_n2659, new_n2661, new_n2662);
not_8  g02286(new_n2662, new_n2663);
not_8  g02287(new_n2634, new_n2664);
xor_4  g02288(new_n2636, new_n2664, new_n2665);
nand_5 g02289(new_n2665, new_n2663, new_n2666);
nand_5 g02290(new_n2666, new_n2660, new_n2667);
and_5  g02291(new_n2667, new_n2651, new_n2668);
nor_5  g02292(new_n2668, new_n2650, new_n2669);
or_5   g02293(new_n2669, new_n2646, new_n2670);
not_8  g02294(new_n2670, new_n2671);
and_5  g02295(new_n2626, new_n2623, new_n2672);
or_5   g02296(new_n2625, new_n2624_1, new_n2673);
not_8  g02297(new_n2673, new_n2674);
or_5   g02298(new_n2644, new_n2628, new_n2675);
not_8  g02299(new_n2675, new_n2676);
xor_4  g02300(new_n2676, new_n2674, new_n2677);
or_5   g02301(new_n2677, new_n2672, new_n2678);
or_5   g02302(new_n2609, new_n2608, new_n2679_1);
not_8  g02303(new_n2679_1, new_n2680);
nand_5 g02304(n2393, n217, new_n2681);
not_8  g02305(new_n2681, new_n2682);
xor_4  g02306(new_n2682, new_n2680, new_n2683);
nand_5 g02307(n3986, n405, new_n2684);
nand_5 g02308(n5860, n4086, new_n2685);
nand_5 g02309(n8433, n5857, new_n2686);
xor_4  g02310(new_n2686, new_n2685, new_n2687);
not_8  g02311(new_n2687, new_n2688);
xor_4  g02312(new_n2688, new_n2684, new_n2689);
xor_4  g02313(new_n2689, new_n2683, new_n2690);
nor_5  g02314(new_n2611, new_n2607, new_n2691);
and_5  g02315(new_n2622, new_n2612, new_n2692);
or_5   g02316(new_n2692, new_n2691, new_n2693);
not_8  g02317(new_n2693, new_n2694);
nand_5 g02318(n11296, n7965, new_n2695);
not_8  g02319(new_n2695, new_n2696);
nand_5 g02320(n11892, n6611, new_n2697);
nand_5 g02321(n7388, n6359, new_n2698);
xor_4  g02322(new_n2698, new_n2697, new_n2699);
not_8  g02323(new_n2699, new_n2700);
xor_4  g02324(new_n2700, new_n2696, new_n2701);
xor_4  g02325(new_n2701, new_n2694, new_n2702);
xor_4  g02326(new_n2702, new_n2690, new_n2703);
xor_4  g02327(new_n2703, new_n2678, new_n2704);
not_8  g02328(new_n2704, new_n2705);
xnor_4 g02329(new_n2705, new_n2671, new_n2706);
not_8  g02330(new_n2706, new_n2707);
nand_5 g02331(n7965, n6359, new_n2708_1);
xor_4  g02332(new_n2669, new_n2646, new_n2709);
not_8  g02333(new_n2709, new_n2710);
nor_5  g02334(new_n2710, new_n2708_1, new_n2711);
or_5   g02335(new_n2665, new_n2663, new_n2712);
and_5  g02336(new_n2712, new_n2666, new_n2713);
xor_4  g02337(new_n2654, new_n2653, new_n2714);
and_5  g02338(n8433, n7388, new_n2715);
and_5  g02339(n7965, n405, new_n2716);
nand_5 g02340(new_n2716, new_n2715, new_n2717);
or_5   g02341(new_n2717, new_n2714, new_n2718);
not_8  g02342(new_n2718, new_n2719);
nand_5 g02343(new_n2719, new_n2713, new_n2720);
xor_4  g02344(new_n2667, new_n2651, new_n2721);
not_8  g02345(new_n2721, new_n2722);
or_5   g02346(new_n2722, new_n2720, new_n2723);
not_8  g02347(new_n2723, new_n2724);
xor_4  g02348(new_n2710, new_n2708_1, new_n2725);
and_5  g02349(new_n2725, new_n2724, new_n2726);
nor_5  g02350(new_n2726, new_n2711, new_n2727);
xor_4  g02351(new_n2727, new_n2707, new_n2728);
not_8  g02352(new_n2728, new_n2729);
xnor_4 g02353(new_n2729, new_n2606, new_n2730);
xor_4  g02354(new_n2602, new_n2600, new_n2731);
not_8  g02355(new_n2731, new_n2732);
xor_4  g02356(new_n2725, new_n2724, new_n2733);
nor_5  g02357(new_n2733, new_n2732, new_n2734);
xor_4  g02358(new_n2722, new_n2720, new_n2735);
xnor_4 g02359(new_n2597, new_n2590, new_n2736);
not_8  g02360(new_n2736, new_n2737);
xor_4  g02361(new_n2719, new_n2713, new_n2738);
nor_5  g02362(new_n2738, new_n2737, new_n2739);
nand_5 g02363(n8433, n7965, new_n2740);
or_5   g02364(new_n2740, new_n2591, new_n2741);
not_8  g02365(new_n2741, new_n2742);
xor_4  g02366(new_n2716, new_n2715, new_n2743);
nor_5  g02367(new_n2743, new_n2742, new_n2744);
xor_4  g02368(new_n2743, new_n2741, new_n2745);
not_8  g02369(new_n2745, new_n2746);
nand_5 g02370(n12925, n8476, new_n2747);
and_5  g02371(n7733, n5331, new_n2748);
xor_4  g02372(new_n2748, new_n2747, new_n2749_1);
and_5  g02373(new_n2749_1, new_n2746, new_n2750);
or_5   g02374(new_n2750, new_n2744, new_n2751);
nand_5 g02375(new_n2593, new_n2527, new_n2752);
nand_5 g02376(new_n2752, new_n2596, new_n2753);
and_5  g02377(new_n2753, new_n2751, new_n2754);
xor_4  g02378(new_n2753, new_n2751, new_n2755);
not_8  g02379(new_n2657, new_n2756);
and_5  g02380(new_n2740, new_n2756, new_n2757);
nor_5  g02381(new_n2757, new_n2714, new_n2758);
or_5   g02382(new_n2654, new_n2653, new_n2759);
and_5  g02383(new_n2757, new_n2759, new_n2760);
or_5   g02384(new_n2760, new_n2758, new_n2761);
and_5  g02385(new_n2761, new_n2755, new_n2762);
or_5   g02386(new_n2762, new_n2754, new_n2763);
xor_4  g02387(new_n2738, new_n2737, new_n2764);
and_5  g02388(new_n2764, new_n2763, new_n2765);
nor_5  g02389(new_n2765, new_n2739, new_n2766);
nor_5  g02390(new_n2766, new_n2735, new_n2767);
xor_4  g02391(new_n2599, new_n2598, new_n2768);
xor_4  g02392(new_n2766, new_n2735, new_n2769);
not_8  g02393(new_n2769, new_n2770);
nor_5  g02394(new_n2770, new_n2768, new_n2771);
or_5   g02395(new_n2771, new_n2767, new_n2772);
xor_4  g02396(new_n2733, new_n2732, new_n2773);
and_5  g02397(new_n2773, new_n2772, new_n2774);
nor_5  g02398(new_n2774, new_n2734, new_n2775);
xor_4  g02399(new_n2775, new_n2730, new_n2776);
xor_4  g02400(new_n2776, new_n2480, new_n2777);
not_8  g02401(new_n2777, new_n2778);
xor_4  g02402(new_n2438, new_n2437, new_n2779);
xor_4  g02403(new_n2773, new_n2772, new_n2780);
not_8  g02404(new_n2780, new_n2781);
nor_5  g02405(new_n2781, new_n2779, new_n2782);
xor_4  g02406(new_n2781, new_n2779, new_n2783);
xor_4  g02407(new_n2435, new_n2434_1, new_n2784);
xnor_4 g02408(new_n2770, new_n2768, new_n2785);
and_5  g02409(new_n2785, new_n2784, new_n2786);
xor_4  g02410(new_n2770, new_n2768, new_n2787);
xor_4  g02411(new_n2787, new_n2784, new_n2788);
xor_4  g02412(new_n2433_1, new_n2428, new_n2789);
not_8  g02413(new_n2789, new_n2790);
not_8  g02414(new_n2763, new_n2791);
xnor_4 g02415(new_n2764, new_n2791, new_n2792);
nor_5  g02416(new_n2792, new_n2790, new_n2793);
xor_4  g02417(new_n2792, new_n2789, new_n2794);
xor_4  g02418(new_n2761, new_n2755, new_n2795);
not_8  g02419(new_n2795, new_n2796);
not_8  g02420(new_n2411, new_n2797);
nand_5 g02421(n8759, n3719, new_n2798);
and_5  g02422(new_n2798, new_n2797, new_n2799);
nor_5  g02423(new_n2799, new_n2429, new_n2800);
or_5   g02424(new_n2408, new_n2407, new_n2801);
and_5  g02425(new_n2799, new_n2801, new_n2802_1);
or_5   g02426(new_n2802_1, new_n2800, new_n2803);
not_8  g02427(new_n2803, new_n2804);
and_5  g02428(new_n2804, new_n2796, new_n2805);
xor_4  g02429(new_n2804, new_n2796, new_n2806);
xor_4  g02430(new_n2749_1, new_n2746, new_n2807);
xor_4  g02431(new_n2431_1, new_n2430, new_n2808);
not_8  g02432(new_n2808, new_n2809);
nor_5  g02433(new_n2809, new_n2807, new_n2810);
xor_4  g02434(new_n2740, new_n2591, new_n2811);
not_8  g02435(new_n2811, new_n2812);
or_5   g02436(new_n2812, new_n2798, new_n2813);
not_8  g02437(new_n2813, new_n2814);
xor_4  g02438(new_n2809, new_n2807, new_n2815);
and_5  g02439(new_n2815, new_n2814, new_n2816);
or_5   g02440(new_n2816, new_n2810, new_n2817);
and_5  g02441(new_n2817, new_n2806, new_n2818_1);
nor_5  g02442(new_n2818_1, new_n2805, new_n2819);
nor_5  g02443(new_n2819, new_n2794, new_n2820);
nor_5  g02444(new_n2820, new_n2793, new_n2821);
nor_5  g02445(new_n2821, new_n2788, new_n2822);
or_5   g02446(new_n2822, new_n2786, new_n2823);
not_8  g02447(new_n2823, new_n2824);
and_5  g02448(new_n2824, new_n2783, new_n2825);
or_5   g02449(new_n2825, new_n2782, new_n2826);
not_8  g02450(new_n2826, new_n2827);
xor_4  g02451(new_n2827, new_n2778, new_n2828);
nor_5  g02452(new_n2828, new_n2360, new_n2829);
xor_4  g02453(new_n2828, new_n2359, new_n2830);
xor_4  g02454(new_n2356, new_n2354, new_n2831);
not_8  g02455(new_n2831, new_n2832);
xor_4  g02456(new_n2824, new_n2783, new_n2833);
nor_5  g02457(new_n2833, new_n2832, new_n2834);
xor_4  g02458(new_n2353, new_n2352, new_n2835);
xor_4  g02459(new_n2821, new_n2788, new_n2836);
nor_5  g02460(new_n2836, new_n2835, new_n2837);
xor_4  g02461(new_n2836, new_n2835, new_n2838);
not_8  g02462(new_n2838, new_n2839);
xor_4  g02463(new_n2351, new_n2346, new_n2840);
xor_4  g02464(new_n2819, new_n2794, new_n2841);
nor_5  g02465(new_n2841, new_n2840, new_n2842);
xor_4  g02466(new_n2817, new_n2806, new_n2843);
not_8  g02467(new_n2843, new_n2844);
not_8  g02468(new_n2287, new_n2845);
nand_5 g02469(n9956, n5305, new_n2846);
and_5  g02470(new_n2846, new_n2845, new_n2847);
nor_5  g02471(new_n2847, new_n2347_1, new_n2848);
nand_5 g02472(new_n2284, new_n2283, new_n2849);
and_5  g02473(new_n2847, new_n2849, new_n2850);
or_5   g02474(new_n2850, new_n2848, new_n2851);
and_5  g02475(new_n2851, new_n2844, new_n2852);
xor_4  g02476(new_n2851, new_n2844, new_n2853);
not_8  g02477(new_n2846, new_n2854);
xor_4  g02478(new_n2812, new_n2798, new_n2855);
nand_5 g02479(new_n2855, new_n2854, new_n2856);
xnor_4 g02480(new_n2349, new_n2348, new_n2857);
and_5  g02481(new_n2857, new_n2856, new_n2858);
xor_4  g02482(new_n2815, new_n2814, new_n2859);
xor_4  g02483(new_n2857, new_n2856, new_n2860);
not_8  g02484(new_n2860, new_n2861);
nor_5  g02485(new_n2861, new_n2859, new_n2862);
or_5   g02486(new_n2862, new_n2858, new_n2863);
and_5  g02487(new_n2863, new_n2853, new_n2864);
or_5   g02488(new_n2864, new_n2852, new_n2865);
not_8  g02489(new_n2865, new_n2866);
xor_4  g02490(new_n2841, new_n2840, new_n2867);
not_8  g02491(new_n2867, new_n2868);
nor_5  g02492(new_n2868, new_n2866, new_n2869);
or_5   g02493(new_n2869, new_n2842, new_n2870);
not_8  g02494(new_n2870, new_n2871);
nor_5  g02495(new_n2871, new_n2839, new_n2872);
or_5   g02496(new_n2872, new_n2837, new_n2873);
xor_4  g02497(new_n2833, new_n2832, new_n2874);
not_8  g02498(new_n2874, new_n2875);
nor_5  g02499(new_n2875, new_n2873, new_n2876);
nor_5  g02500(new_n2876, new_n2834, new_n2877);
nor_5  g02501(new_n2877, new_n2830, new_n2878);
or_5   g02502(new_n2878, new_n2829, new_n2879_1);
nor_5  g02503(new_n2776, new_n2480, new_n2880);
nor_5  g02504(new_n2826, new_n2778, new_n2881);
nor_5  g02505(new_n2881, new_n2880, new_n2882);
and_5  g02506(new_n2559, new_n2557, new_n2883);
and_5  g02507(new_n2566, new_n2560, new_n2884);
or_5   g02508(new_n2884, new_n2883, new_n2885);
and_5  g02509(new_n2563, new_n2562, new_n2886);
not_8  g02510(new_n2561, new_n2887);
nor_5  g02511(new_n2565, new_n2887, new_n2888);
or_5   g02512(new_n2888, new_n2886, new_n2889);
nand_5 g02513(n12648, n4970, new_n2890);
and_5  g02514(n11296, n7388, new_n2891);
and_5  g02515(n9241, n6126, new_n2892);
xor_4  g02516(new_n2892, new_n2891, new_n2893);
xor_4  g02517(new_n2893, new_n2890, new_n2894);
xor_4  g02518(new_n2894, new_n2889, new_n2895);
xor_4  g02519(new_n2895, new_n2885, new_n2896);
and_5  g02520(new_n2686, new_n2685, new_n2897);
not_8  g02521(new_n2684, new_n2898);
nor_5  g02522(new_n2688, new_n2898, new_n2899);
or_5   g02523(new_n2899, new_n2897, new_n2900);
and_5  g02524(new_n2698, new_n2697, new_n2901);
nor_5  g02525(new_n2700, new_n2696, new_n2902_1);
nor_5  g02526(new_n2902_1, new_n2901, new_n2903);
xor_4  g02527(new_n2903, new_n2900, new_n2904);
nand_5 g02528(n11892, n6359, new_n2905);
and_5  g02529(n7546, n5331, new_n2906);
xor_4  g02530(new_n2906, new_n2905, new_n2907);
xor_4  g02531(new_n2907, new_n2904, new_n2908);
and_5  g02532(new_n2458, new_n2456, new_n2909);
and_5  g02533(new_n2464_1, new_n2459, new_n2910);
nor_5  g02534(new_n2910, new_n2909, new_n2911);
and_5  g02535(n8595, n8276, new_n2912);
and_5  g02536(n6611, n2393, new_n2913);
xor_4  g02537(new_n2913, new_n2912, new_n2914);
nand_5 g02538(n12925, n4499, new_n2915);
and_5  g02539(n11536, n5305, new_n2916);
xor_4  g02540(new_n2916, new_n2915, new_n2917);
xor_4  g02541(new_n2917, new_n2914, new_n2918);
xor_4  g02542(new_n2918, new_n2911, new_n2919);
xor_4  g02543(new_n2919, new_n2908, new_n2920);
and_5  g02544(new_n2682, new_n2680, new_n2921);
and_5  g02545(new_n2689, new_n2683, new_n2922);
nor_5  g02546(new_n2922, new_n2921, new_n2923);
and_5  g02547(new_n2575, new_n2574, new_n2924);
nor_5  g02548(new_n2577_1, new_n2573, new_n2925);
or_5   g02549(new_n2925, new_n2924, new_n2926);
nand_5 g02550(n4086, n3986, new_n2927);
and_5  g02551(n7733, n3616, new_n2928);
xor_4  g02552(new_n2928, new_n2927, new_n2929);
xor_4  g02553(new_n2929, new_n2926, new_n2930);
xor_4  g02554(new_n2930, new_n2923, new_n2931);
xor_4  g02555(new_n2931, new_n2920, new_n2932);
xor_4  g02556(new_n2932, new_n2896, new_n2933);
nor_5  g02557(new_n2705, new_n2670, new_n2934);
nor_5  g02558(new_n2727, new_n2707, new_n2935);
or_5   g02559(new_n2935, new_n2934, new_n2936);
and_5  g02560(n5860, n217, new_n2937);
xor_4  g02561(new_n2937, new_n2936, new_n2938);
nor_5  g02562(new_n2476, new_n2442, new_n2939);
nor_5  g02563(new_n2478, new_n2441, new_n2940);
or_5   g02564(new_n2940, new_n2939, new_n2941);
nor_5  g02565(new_n2578, new_n2571, new_n2942);
and_5  g02566(new_n2579, new_n2567, new_n2943);
or_5   g02567(new_n2943, new_n2942, new_n2944);
and_5  g02568(n12299, n8065, new_n2945);
and_5  g02569(n10510, n3602, new_n2946);
xor_4  g02570(new_n2946, new_n2945, new_n2947);
nand_5 g02571(n10644, n3719, new_n2948);
and_5  g02572(n7965, n1357, new_n2949);
xor_4  g02573(new_n2949, new_n2948, new_n2950);
and_5  g02574(n10439, n7436, new_n2951);
and_5  g02575(n8759, n4190, new_n2952);
xor_4  g02576(new_n2952, new_n2951, new_n2953);
xor_4  g02577(new_n2953, new_n2950, new_n2954);
xor_4  g02578(new_n2954, new_n2947, new_n2955);
and_5  g02579(new_n2308, new_n2307, new_n2956);
nor_5  g02580(new_n2310, new_n2306, new_n2957);
nor_5  g02581(new_n2957, new_n2956, new_n2958);
and_5  g02582(n9637, n1097, new_n2959);
xor_4  g02583(new_n2959, new_n2958, new_n2960);
xor_4  g02584(new_n2960, new_n2955, new_n2961);
xor_4  g02585(new_n2961, new_n2944, new_n2962);
or_5   g02586(new_n2453, new_n2445, new_n2963);
not_8  g02587(new_n2465, new_n2964);
nand_5 g02588(new_n2964, new_n2454, new_n2965);
nand_5 g02589(new_n2965, new_n2963, new_n2966);
nor_5  g02590(new_n2328, new_n2315, new_n2967);
nor_5  g02591(new_n2967, new_n2313, new_n2968);
xor_4  g02592(new_n2968, new_n2966, new_n2969);
xor_4  g02593(new_n2969, new_n2962, new_n2970);
and_5  g02594(new_n2472, new_n2470, new_n2971);
nor_5  g02595(new_n2474, new_n2467, new_n2972);
nor_5  g02596(new_n2972, new_n2971, new_n2973);
and_5  g02597(new_n2449, new_n2448, new_n2974);
nor_5  g02598(new_n2451, new_n2447, new_n2975);
nor_5  g02599(new_n2975, new_n2974, new_n2976);
and_5  g02600(n4312, n2577, new_n2977);
xor_4  g02601(new_n2977, new_n2976, new_n2978);
nor_5  g02602(new_n2462, new_n2461, new_n2979);
nand_5 g02603(n9241, n3602, new_n2980);
and_5  g02604(new_n2462, new_n2461, new_n2981);
nor_5  g02605(new_n2981, new_n2980, new_n2982);
or_5   g02606(new_n2982, new_n2979, new_n2983);
and_5  g02607(n11257, n4921, new_n2984);
and_5  g02608(n12705, n3842, new_n2985);
xor_4  g02609(new_n2985, new_n2984, new_n2986);
xor_4  g02610(new_n2986, new_n2983, new_n2987);
xor_4  g02611(new_n2987, new_n2978, new_n2988);
and_5  g02612(n8433, n45, new_n2989);
and_5  g02613(n12025, n11917, new_n2990);
xor_4  g02614(new_n2990, new_n2989, new_n2991);
and_5  g02615(new_n2323, new_n2322, new_n2992);
nor_5  g02616(new_n2325, new_n2321, new_n2993);
nor_5  g02617(new_n2993, new_n2992, new_n2994);
nand_5 g02618(n5964, n1835, new_n2995);
and_5  g02619(n5857, n405, new_n2996);
xor_4  g02620(new_n2996, new_n2995, new_n2997);
xor_4  g02621(new_n2997, new_n2994, new_n2998);
xor_4  g02622(new_n2998, new_n2991, new_n2999);
nor_5  g02623(new_n2318, new_n2317, new_n3000);
and_5  g02624(new_n2326, new_n2319, new_n3001);
nor_5  g02625(new_n3001, new_n3000, new_n3002);
and_5  g02626(n10391, n6776, new_n3003);
xor_4  g02627(new_n3003, new_n3002, new_n3004);
xor_4  g02628(new_n3004, new_n2999, new_n3005);
xor_4  g02629(new_n3005, new_n2988, new_n3006);
xor_4  g02630(new_n3006, new_n2973, new_n3007);
xor_4  g02631(new_n3007, new_n2970, new_n3008);
xor_4  g02632(new_n3008, new_n2941, new_n3009);
xor_4  g02633(new_n3009, new_n2938, new_n3010);
xor_4  g02634(new_n3010, new_n2933, new_n3011);
and_5  g02635(new_n2729, new_n2606, new_n3012);
nor_5  g02636(new_n2775, new_n2730, new_n3013);
nor_5  g02637(new_n3013, new_n3012, new_n3014);
and_5  g02638(new_n2676, new_n2674, new_n3015);
and_5  g02639(new_n2703, new_n2678, new_n3016);
or_5   g02640(new_n3016, new_n3015, new_n3017);
and_5  g02641(new_n2334, new_n2332, new_n3018);
nor_5  g02642(new_n2336, new_n2329, new_n3019);
nor_5  g02643(new_n3019, new_n3018, new_n3020);
xor_4  g02644(new_n3020, new_n3017, new_n3021);
xor_4  g02645(new_n3021, new_n3014, new_n3022_1);
xor_4  g02646(new_n3022_1, new_n3011, new_n3023);
xor_4  g02647(new_n3023, new_n2882, new_n3024);
nor_5  g02648(new_n2582, new_n2548, new_n3025);
nor_5  g02649(new_n2604, new_n2584, new_n3026);
or_5   g02650(new_n3026, new_n3025, new_n3027);
nor_5  g02651(new_n2338, new_n2300, new_n3028);
nor_5  g02652(new_n2358, new_n2340, new_n3029);
nor_5  g02653(new_n3029, new_n3028, new_n3030);
xor_4  g02654(new_n3030, new_n3027, new_n3031);
and_5  g02655(new_n2553, new_n2551_1, new_n3032);
and_5  g02656(new_n2580, new_n2555, new_n3033);
or_5   g02657(new_n3033, new_n3032, new_n3034);
and_5  g02658(new_n2701, new_n2694, new_n3035);
not_8  g02659(new_n2690, new_n3036);
and_5  g02660(new_n2702, new_n3036, new_n3037);
nor_5  g02661(new_n3037, new_n3035, new_n3038);
nand_5 g02662(n10547, n9956, new_n3039);
nand_5 g02663(n10965, n8476, new_n3040);
and_5  g02664(n7690, n4826, new_n3041);
xor_4  g02665(new_n3041, new_n3040, new_n3042);
and_5  g02666(n10545, n7610, new_n3043);
and_5  g02667(n2530, n503, new_n3044);
xor_4  g02668(new_n3044, new_n3043, new_n3045);
xor_4  g02669(new_n3045, new_n3042, new_n3046);
xor_4  g02670(new_n3046, new_n3039, new_n3047);
xor_4  g02671(new_n3047, new_n3038, new_n3048);
xor_4  g02672(new_n3048, new_n3034, new_n3049);
xor_4  g02673(new_n3049, new_n3031, new_n3050);
xor_4  g02674(new_n3050, new_n3024, new_n3051);
xor_4  g02675(new_n3051, new_n2879_1, n837);
nand_5 g02676(n11917, n11757, new_n3053);
not_8  g02677(new_n3053, new_n3054);
nand_5 g02678(n9956, n5240, new_n3055);
nand_5 g02679(n11757, n4921, new_n3056);
and_5  g02680(n11917, n3172, new_n3057);
xor_4  g02681(new_n3057, new_n3055, new_n3058);
not_8  g02682(new_n3058, new_n3059);
and_5  g02683(new_n3059, new_n3056, new_n3060);
nor_5  g02684(new_n3060, new_n3055, new_n3061);
nor_5  g02685(new_n3061, new_n3054, new_n3062);
nand_5 g02686(n4921, n3172, new_n3063);
not_8  g02687(new_n3063, new_n3064);
nor_5  g02688(new_n3064, new_n3061, new_n3065);
nor_5  g02689(new_n3065, new_n3053, new_n3066);
or_5   g02690(new_n3066, new_n3062, new_n3067);
not_8  g02691(new_n3067, new_n3068);
nand_5 g02692(n5240, n4921, new_n3069);
nand_5 g02693(n11821, n9956, new_n3070);
xor_4  g02694(new_n3070, new_n3069, new_n3071_1);
nor_5  g02695(new_n3071_1, new_n3068, new_n3072);
and_5  g02696(new_n3071_1, new_n3068, new_n3073);
or_5   g02697(new_n3073, new_n3072, new_n3074);
nand_5 g02698(n2577, n1333, new_n3075);
nand_5 g02699(n3842, n3172, new_n3076);
xor_4  g02700(new_n3076, new_n3075, new_n3077);
not_8  g02701(new_n3077, new_n3078);
xor_4  g02702(new_n3078, new_n3074, new_n3079);
nand_5 g02703(n3842, n1333, new_n3080);
not_8  g02704(new_n3080, new_n3081);
nand_5 g02705(n11757, n9956, new_n3082);
nand_5 g02706(n11917, n1333, new_n3083);
and_5  g02707(new_n3083, new_n3082, new_n3084);
nor_5  g02708(new_n3083, new_n3082, new_n3085);
nor_5  g02709(new_n3085, new_n3064, new_n3086);
or_5   g02710(new_n3086, new_n3084, new_n3087);
not_8  g02711(new_n3087, new_n3088);
and_5  g02712(new_n3088, new_n3081, new_n3089);
xor_4  g02713(new_n3059, new_n3056, new_n3090);
nor_5  g02714(new_n3088, new_n3081, new_n3091);
or_5   g02715(new_n3091, new_n3089, new_n3092);
nor_5  g02716(new_n3092, new_n3090, new_n3093);
or_5   g02717(new_n3093, new_n3089, new_n3094);
xor_4  g02718(new_n3094, new_n3079, new_n3095);
not_8  g02719(new_n3095, new_n3096);
nand_5 g02720(n7862, n2577, new_n3097);
not_8  g02721(new_n3097, new_n3098);
xor_4  g02722(new_n3092, new_n3090, new_n3099);
and_5  g02723(new_n3099, new_n3098, new_n3100);
nand_5 g02724(n7862, n3842, new_n3101);
nand_5 g02725(n9956, n3172, new_n3102);
nand_5 g02726(n11917, n7862, new_n3103);
nor_5  g02727(new_n3103, new_n3102, new_n3104);
and_5  g02728(new_n3103, new_n3102, new_n3105);
nand_5 g02729(n4921, n1333, new_n3106);
nor_5  g02730(new_n3106, new_n3105, new_n3107);
nor_5  g02731(new_n3107, new_n3104, new_n3108);
nor_5  g02732(new_n3108, new_n3101, new_n3109);
xor_4  g02733(new_n3108, new_n3101, new_n3110);
not_8  g02734(new_n3110, new_n3111);
xor_4  g02735(new_n3083, new_n3082, new_n3112);
xor_4  g02736(new_n3112, new_n3063, new_n3113);
nor_5  g02737(new_n3113, new_n3111, new_n3114);
or_5   g02738(new_n3114, new_n3109, new_n3115);
not_8  g02739(new_n3115, new_n3116);
xor_4  g02740(new_n3099, new_n3098, new_n3117);
not_8  g02741(new_n3117, new_n3118);
nor_5  g02742(new_n3118, new_n3116, new_n3119);
nor_5  g02743(new_n3119, new_n3100, new_n3120);
or_5   g02744(new_n3120, new_n3096, new_n3121);
or_5   g02745(new_n3073, new_n3066, new_n3122);
nand_5 g02746(n9637, n1333, new_n3123);
nand_5 g02747(n3172, n2577, new_n3124_1);
nand_5 g02748(n7862, n1835, new_n3125);
xor_4  g02749(new_n3125, new_n3124_1, new_n3126);
xor_4  g02750(new_n3126, new_n3123, new_n3127);
not_8  g02751(new_n3127, new_n3128);
xor_4  g02752(new_n3128, new_n3122, new_n3129);
or_5   g02753(new_n3070, new_n3069, new_n3130);
not_8  g02754(new_n3130, new_n3131);
nand_5 g02755(n11757, n3842, new_n3132);
not_8  g02756(new_n3132, new_n3133);
xor_4  g02757(new_n3133, new_n3131, new_n3134);
nand_5 g02758(n11821, n4921, new_n3135);
nand_5 g02759(n9956, n9080, new_n3136);
nand_5 g02760(n11917, n5240, new_n3137);
xor_4  g02761(new_n3137, new_n3136, new_n3138);
not_8  g02762(new_n3138, new_n3139);
xor_4  g02763(new_n3139, new_n3135, new_n3140);
xor_4  g02764(new_n3140, new_n3134, new_n3141);
xor_4  g02765(new_n3141, new_n3129, new_n3142);
not_8  g02766(new_n3142, new_n3143);
nor_5  g02767(new_n3078, new_n3074, new_n3144);
or_5   g02768(new_n3076, new_n3075, new_n3145);
nand_5 g02769(new_n3094, new_n3079, new_n3146_1);
xor_4  g02770(new_n3146_1, new_n3145, new_n3147);
nor_5  g02771(new_n3147, new_n3144, new_n3148);
xor_4  g02772(new_n3148, new_n3143, new_n3149);
not_8  g02773(new_n3149, new_n3150);
xor_4  g02774(new_n3150, new_n3121, new_n3151);
not_8  g02775(new_n3151, new_n3152);
nand_5 g02776(n9637, n7862, new_n3153);
xor_4  g02777(new_n3120, new_n3096, new_n3154);
not_8  g02778(new_n3154, new_n3155);
nor_5  g02779(new_n3155, new_n3153, new_n3156);
and_5  g02780(new_n3113, new_n3111, new_n3157);
or_5   g02781(new_n3157, new_n3114, new_n3158);
xor_4  g02782(new_n3103, new_n3102, new_n3159);
nand_5 g02783(n9956, n1333, new_n3160);
nand_5 g02784(n7862, n4921, new_n3161);
or_5   g02785(new_n3161, new_n3160, new_n3162);
or_5   g02786(new_n3162, new_n3159, new_n3163);
or_5   g02787(new_n3163, new_n3158, new_n3164);
xor_4  g02788(new_n3118, new_n3115, new_n3165);
or_5   g02789(new_n3165, new_n3164, new_n3166);
not_8  g02790(new_n3166, new_n3167);
xor_4  g02791(new_n3155, new_n3153, new_n3168);
and_5  g02792(new_n3168, new_n3167, new_n3169);
nor_5  g02793(new_n3169, new_n3156, new_n3170);
xor_4  g02794(new_n3170, new_n3152, new_n3171);
xor_4  g02795(new_n3168, new_n3167, new_n3172_1);
not_8  g02796(new_n3172_1, new_n3173);
nand_5 g02797(n8595, n6877, new_n3174);
and_5  g02798(n6877, n6126, new_n3175);
and_5  g02799(n3719, n2464, new_n3176);
nor_5  g02800(new_n3176, new_n3175, new_n3177);
nand_5 g02801(n6877, n3719, new_n3178);
nand_5 g02802(n6126, n2464, new_n3179);
nor_5  g02803(new_n3179, new_n3178, new_n3180);
nand_5 g02804(n9400, n3602, new_n3181);
not_8  g02805(new_n3181, new_n3182);
nor_5  g02806(new_n3182, new_n3180, new_n3183);
nor_5  g02807(new_n3183, new_n3177, new_n3184);
not_8  g02808(new_n3184, new_n3185);
xor_4  g02809(new_n3185, new_n3174, new_n3186);
nand_5 g02810(n3602, n2464, new_n3187);
not_8  g02811(new_n3187, new_n3188);
nand_5 g02812(n9400, n6126, new_n3189);
nand_5 g02813(n11311, n3719, new_n3190);
xor_4  g02814(new_n3190, new_n3189, new_n3191);
xor_4  g02815(new_n3191, new_n3188, new_n3192);
xor_4  g02816(new_n3192, new_n3186, new_n3193);
not_8  g02817(new_n3178, new_n3194);
or_5   g02818(new_n3181, new_n3194, new_n3195);
not_8  g02819(new_n3195, new_n3196);
nor_5  g02820(new_n3180, new_n3177, new_n3197);
nor_5  g02821(new_n3197, new_n3196, new_n3198);
not_8  g02822(new_n3198, new_n3199);
or_5   g02823(new_n3199, new_n3181, new_n3200);
not_8  g02824(new_n3200, new_n3201);
nand_5 g02825(new_n3201, new_n3193, new_n3202);
not_8  g02826(new_n3202, new_n3203);
nand_5 g02827(n10439, n6877, new_n3204);
not_8  g02828(new_n3204, new_n3205);
nand_5 g02829(n9400, n8595, new_n3206);
not_8  g02830(new_n3206, new_n3207);
and_5  g02831(new_n3190, new_n3189, new_n3208);
nor_5  g02832(new_n3190, new_n3189, new_n3209);
nor_5  g02833(new_n3209, new_n3188, new_n3210);
or_5   g02834(new_n3210, new_n3208, new_n3211);
not_8  g02835(new_n3211, new_n3212);
and_5  g02836(new_n3212, new_n3207, new_n3213);
nor_5  g02837(new_n3212, new_n3207, new_n3214_1);
or_5   g02838(new_n3214_1, new_n3213, new_n3215);
nand_5 g02839(n11311, n3602, new_n3216);
not_8  g02840(new_n3216, new_n3217);
nand_5 g02841(n4187, n3719, new_n3218);
xor_4  g02842(new_n3218, new_n3179, new_n3219);
not_8  g02843(new_n3219, new_n3220);
xor_4  g02844(new_n3220, new_n3217, new_n3221);
xor_4  g02845(new_n3221, new_n3215, new_n3222);
xor_4  g02846(new_n3222, new_n3205, new_n3223);
not_8  g02847(new_n3223, new_n3224);
nor_5  g02848(new_n3185, new_n3174, new_n3225);
and_5  g02849(new_n3192, new_n3186, new_n3226);
nor_5  g02850(new_n3226, new_n3225, new_n3227);
xor_4  g02851(new_n3227, new_n3224, new_n3228);
nand_5 g02852(new_n3228, new_n3203, new_n3229);
not_8  g02853(new_n3229, new_n3230_1);
nand_5 g02854(n8065, n6877, new_n3231);
not_8  g02855(new_n3231, new_n3232);
nand_5 g02856(n11311, n6126, new_n3233);
nand_5 g02857(n4203, n3719, new_n3234);
nand_5 g02858(n4187, n3602, new_n3235);
xor_4  g02859(new_n3235, new_n3234, new_n3236);
not_8  g02860(new_n3236, new_n3237);
xor_4  g02861(new_n3237, new_n3233, new_n3238);
and_5  g02862(new_n3218, new_n3179, new_n3239);
nor_5  g02863(new_n3220, new_n3217, new_n3240);
or_5   g02864(new_n3240, new_n3239, new_n3241);
not_8  g02865(new_n3241, new_n3242);
xor_4  g02866(new_n3242, new_n3238, new_n3243);
nand_5 g02867(n10439, n9400, new_n3244);
nand_5 g02868(n8595, n2464, new_n3245);
xor_4  g02869(new_n3245, new_n3244, new_n3246);
xor_4  g02870(new_n3246, new_n3243, new_n3247);
nor_5  g02871(new_n3221, new_n3215, new_n3248);
nor_5  g02872(new_n3248, new_n3213, new_n3249);
xor_4  g02873(new_n3249, new_n3247, new_n3250);
and_5  g02874(new_n3222, new_n3205, new_n3251);
nor_5  g02875(new_n3227, new_n3224, new_n3252);
nor_5  g02876(new_n3252, new_n3251, new_n3253);
xor_4  g02877(new_n3253, new_n3250, new_n3254);
xor_4  g02878(new_n3254, new_n3232, new_n3255);
not_8  g02879(new_n3255, new_n3256);
xor_4  g02880(new_n3256, new_n3230_1, new_n3257);
not_8  g02881(new_n3257, new_n3258);
xor_4  g02882(new_n3228, new_n3203, new_n3259);
xor_4  g02883(new_n3200, new_n3193, new_n3260);
not_8  g02884(new_n3260, new_n3261);
or_5   g02885(new_n3195, new_n3177, new_n3262);
nand_5 g02886(new_n3262, new_n3199, new_n3263);
and_5  g02887(n8433, n7236, new_n3264);
not_8  g02888(new_n3264, new_n3265);
nand_5 g02889(n12925, n4805, new_n3266);
or_5   g02890(new_n3266, new_n3265, new_n3267);
and_5  g02891(n7733, n4805, new_n3268);
and_5  g02892(n12925, n11478, new_n3269);
xnor_4 g02893(new_n3269, new_n3268, new_n3270);
and_5  g02894(new_n3270, new_n3267, new_n3271);
xor_4  g02895(new_n3269, new_n3268, new_n3272_1);
xor_4  g02896(new_n3272_1, new_n3267, new_n3273);
not_8  g02897(new_n3273, new_n3274);
nand_5 g02898(n7236, n405, new_n3275);
and_5  g02899(n8433, n3992, new_n3276);
xor_4  g02900(new_n3276, new_n3275, new_n3277);
and_5  g02901(new_n3277, new_n3274, new_n3278);
or_5   g02902(new_n3278, new_n3271, new_n3279);
not_8  g02903(new_n3279, new_n3280);
nand_5 g02904(n3992, n405, new_n3281);
nor_5  g02905(new_n3281, new_n3264, new_n3282);
not_8  g02906(new_n3282, new_n3283);
and_5  g02907(n8433, n8384, new_n3284);
and_5  g02908(n7236, n4086, new_n3285);
or_5   g02909(new_n3285, new_n3284, new_n3286);
not_8  g02910(new_n3286, new_n3287_1);
and_5  g02911(new_n3287_1, new_n3283, new_n3288);
and_5  g02912(new_n3285, new_n3284, new_n3289);
or_5   g02913(new_n3289, new_n3288, new_n3290);
nor_5  g02914(new_n3287_1, new_n3283, new_n3291);
nor_5  g02915(new_n3291, new_n3290, new_n3292);
xor_4  g02916(new_n3292, new_n3280, new_n3293);
and_5  g02917(n11478, n7733, new_n3294);
and_5  g02918(new_n3294, new_n3266, new_n3295);
not_8  g02919(new_n3295, new_n3296);
nand_5 g02920(n12925, n5283, new_n3297);
nand_5 g02921(n4826, n4805, new_n3298);
nand_5 g02922(new_n3298, new_n3297, new_n3299);
nor_5  g02923(new_n3299, new_n3296, new_n3300);
xnor_4 g02924(new_n3298, new_n3297, new_n3301);
not_8  g02925(new_n3301, new_n3302);
and_5  g02926(new_n3302, new_n3296, new_n3303);
nor_5  g02927(new_n3303, new_n3300, new_n3304);
xor_4  g02928(new_n3304, new_n3293, new_n3305);
nor_5  g02929(new_n3305, new_n3263, new_n3306);
xor_4  g02930(new_n3305, new_n3263, new_n3307);
not_8  g02931(new_n3307, new_n3308);
xor_4  g02932(new_n3277, new_n3274, new_n3309);
and_5  g02933(n9400, n3719, new_n3310);
and_5  g02934(n6877, n3602, new_n3311);
xor_4  g02935(new_n3311, new_n3310, new_n3312);
not_8  g02936(new_n3312, new_n3313);
nor_5  g02937(new_n3313, new_n3309, new_n3314);
xor_4  g02938(new_n3266, new_n3264, new_n3315);
not_8  g02939(new_n3315, new_n3316);
nand_5 g02940(new_n3316, new_n3194, new_n3317);
xor_4  g02941(new_n3312, new_n3309, new_n3318);
nor_5  g02942(new_n3318, new_n3317, new_n3319);
nor_5  g02943(new_n3319, new_n3314, new_n3320);
nor_5  g02944(new_n3320, new_n3308, new_n3321);
or_5   g02945(new_n3321, new_n3306, new_n3322);
nor_5  g02946(new_n3322, new_n3261, new_n3323);
nand_5 g02947(n7610, n4805, new_n3324);
nor_5  g02948(new_n3298, new_n3297, new_n3325);
nand_5 g02949(n11478, n7733, new_n3326);
not_8  g02950(new_n3299, new_n3327);
nor_5  g02951(new_n3327, new_n3326, new_n3328);
nor_5  g02952(new_n3328, new_n3325, new_n3329);
xor_4  g02953(new_n3329, new_n3324, new_n3330);
not_8  g02954(new_n3330, new_n3331);
nand_5 g02955(n7733, n5283, new_n3332);
nand_5 g02956(n12925, n137, new_n3333);
nand_5 g02957(n11478, n4826, new_n3334);
xnor_4 g02958(new_n3334, new_n3333, new_n3335);
not_8  g02959(new_n3335, new_n3336);
xor_4  g02960(new_n3336, new_n3332, new_n3337);
xor_4  g02961(new_n3337, new_n3331, new_n3338);
nand_5 g02962(new_n3269, new_n3268, new_n3339_1);
or_5   g02963(new_n3302, new_n3339_1, new_n3340);
not_8  g02964(new_n3340, new_n3341);
xor_4  g02965(new_n3341, new_n3338, new_n3342_1);
nand_5 g02966(n7236, n217, new_n3343);
not_8  g02967(new_n3343, new_n3344);
not_8  g02968(new_n3281, new_n3345);
nor_5  g02969(new_n3289, new_n3345, new_n3346);
nor_5  g02970(new_n3346, new_n3287_1, new_n3347);
not_8  g02971(new_n3347, new_n3348);
xor_4  g02972(new_n3348, new_n3344, new_n3349);
nand_5 g02973(n8384, n405, new_n3350);
nand_5 g02974(n8433, n6358, new_n3351);
nand_5 g02975(n4086, n3992, new_n3352);
xnor_4 g02976(new_n3352, new_n3351, new_n3353);
not_8  g02977(new_n3353, new_n3354);
xor_4  g02978(new_n3354, new_n3350, new_n3355);
xor_4  g02979(new_n3355, new_n3349, new_n3356);
and_5  g02980(new_n3290, new_n3345, new_n3357);
not_8  g02981(new_n3357, new_n3358);
xnor_4 g02982(new_n3358, new_n3356, new_n3359);
xor_4  g02983(new_n3359, new_n3342_1, new_n3360);
nor_5  g02984(new_n3292, new_n3280, new_n3361);
and_5  g02985(new_n3304, new_n3293, new_n3362);
nor_5  g02986(new_n3362, new_n3361, new_n3363);
xor_4  g02987(new_n3363, new_n3360, new_n3364);
xor_4  g02988(new_n3322, new_n3261, new_n3365);
not_8  g02989(new_n3365, new_n3366);
nor_5  g02990(new_n3366, new_n3364, new_n3367);
or_5   g02991(new_n3367, new_n3323, new_n3368);
not_8  g02992(new_n3368, new_n3369);
nor_5  g02993(new_n3369, new_n3259, new_n3370);
and_5  g02994(new_n3369, new_n3259, new_n3371);
nand_5 g02995(new_n3357, new_n3356, new_n3372);
nand_5 g02996(n7236, n6611, new_n3373);
nand_5 g02997(n3992, n217, new_n3374);
not_8  g02998(new_n3374, new_n3375);
and_5  g02999(new_n3352, new_n3351, new_n3376);
and_5  g03000(new_n3354, new_n3350, new_n3377);
or_5   g03001(new_n3377, new_n3376, new_n3378);
not_8  g03002(new_n3378, new_n3379);
xor_4  g03003(new_n3379, new_n3375, new_n3380);
nand_5 g03004(n6358, n405, new_n3381);
nand_5 g03005(n8384, n4086, new_n3382);
nand_5 g03006(n8433, n5198, new_n3383);
xor_4  g03007(new_n3383, new_n3382, new_n3384);
not_8  g03008(new_n3384, new_n3385);
xor_4  g03009(new_n3385, new_n3381, new_n3386);
xor_4  g03010(new_n3386, new_n3380, new_n3387);
not_8  g03011(new_n3387, new_n3388);
xor_4  g03012(new_n3388, new_n3373, new_n3389);
nor_5  g03013(new_n3348, new_n3343, new_n3390);
nor_5  g03014(new_n3355, new_n3349, new_n3391);
or_5   g03015(new_n3391, new_n3390, new_n3392);
xor_4  g03016(new_n3392, new_n3389, new_n3393);
not_8  g03017(new_n3393, new_n3394);
xor_4  g03018(new_n3394, new_n3372, new_n3395);
nand_5 g03019(new_n3341, new_n3338, new_n3396);
nand_5 g03020(n4970, n4805, new_n3397);
nand_5 g03021(n11478, n7610, new_n3398);
not_8  g03022(new_n3398, new_n3399);
and_5  g03023(new_n3334, new_n3333, new_n3400);
and_5  g03024(new_n3336, new_n3332, new_n3401);
or_5   g03025(new_n3401, new_n3400, new_n3402);
not_8  g03026(new_n3402, new_n3403);
xor_4  g03027(new_n3403, new_n3399, new_n3404);
nand_5 g03028(n7733, n137, new_n3405);
nand_5 g03029(n5283, n4826, new_n3406);
nand_5 g03030(n12925, n6294, new_n3407);
xor_4  g03031(new_n3407, new_n3406, new_n3408);
not_8  g03032(new_n3408, new_n3409);
xor_4  g03033(new_n3409, new_n3405, new_n3410);
xor_4  g03034(new_n3410, new_n3404, new_n3411);
not_8  g03035(new_n3411, new_n3412);
xor_4  g03036(new_n3412, new_n3397, new_n3413);
nor_5  g03037(new_n3329, new_n3324, new_n3414);
nor_5  g03038(new_n3337, new_n3331, new_n3415);
or_5   g03039(new_n3415, new_n3414, new_n3416);
xor_4  g03040(new_n3416, new_n3413, new_n3417);
not_8  g03041(new_n3417, new_n3418);
xor_4  g03042(new_n3418, new_n3396, new_n3419);
nor_5  g03043(new_n3359, new_n3342_1, new_n3420);
not_8  g03044(new_n3360, new_n3421);
nor_5  g03045(new_n3363, new_n3421, new_n3422);
nor_5  g03046(new_n3422, new_n3420, new_n3423);
xor_4  g03047(new_n3423, new_n3419, new_n3424);
not_8  g03048(new_n3424, new_n3425);
xor_4  g03049(new_n3425, new_n3395, new_n3426);
not_8  g03050(new_n3426, new_n3427);
nor_5  g03051(new_n3427, new_n3371, new_n3428);
or_5   g03052(new_n3428, new_n3370, new_n3429);
not_8  g03053(new_n3429, new_n3430);
xor_4  g03054(new_n3430, new_n3258, new_n3431);
or_5   g03055(new_n3394, new_n3372, new_n3432);
nand_5 g03056(n7236, n6359, new_n3433);
not_8  g03057(new_n3433, new_n3434);
nand_5 g03058(n6358, n4086, new_n3435);
not_8  g03059(new_n3435, new_n3436);
and_5  g03060(new_n3383, new_n3382, new_n3437);
not_8  g03061(new_n3381, new_n3438);
nor_5  g03062(new_n3385, new_n3438, new_n3439);
or_5   g03063(new_n3439, new_n3437, new_n3440);
not_8  g03064(new_n3440, new_n3441);
xor_4  g03065(new_n3441, new_n3436, new_n3442);
nand_5 g03066(n5198, n405, new_n3443);
nand_5 g03067(n8433, n1471, new_n3444);
xor_4  g03068(new_n3444, new_n3443, new_n3445);
xor_4  g03069(new_n3445, new_n3442, new_n3446);
not_8  g03070(new_n3446, new_n3447);
nand_5 g03071(n8384, n217, new_n3448);
nand_5 g03072(n6611, n3992, new_n3449);
xor_4  g03073(new_n3449, new_n3448, new_n3450);
not_8  g03074(new_n3450, new_n3451);
xor_4  g03075(new_n3451, new_n3447, new_n3452);
and_5  g03076(new_n3379, new_n3375, new_n3453);
and_5  g03077(new_n3386, new_n3380, new_n3454);
or_5   g03078(new_n3454, new_n3453, new_n3455);
not_8  g03079(new_n3455, new_n3456_1);
xor_4  g03080(new_n3456_1, new_n3452, new_n3457);
nor_5  g03081(new_n3388, new_n3373, new_n3458);
and_5  g03082(new_n3392, new_n3389, new_n3459);
nor_5  g03083(new_n3459, new_n3458, new_n3460);
xor_4  g03084(new_n3460, new_n3457, new_n3461);
xor_4  g03085(new_n3461, new_n3434, new_n3462);
not_8  g03086(new_n3462, new_n3463);
xor_4  g03087(new_n3463, new_n3432, new_n3464);
or_5   g03088(new_n3418, new_n3396, new_n3465);
not_8  g03089(new_n3465, new_n3466);
nand_5 g03090(n4805, n503, new_n3467);
not_8  g03091(new_n3467, new_n3468);
nand_5 g03092(n4826, n137, new_n3469);
nand_5 g03093(n7733, n6294, new_n3470);
nand_5 g03094(n12925, n6797, new_n3471);
xor_4  g03095(new_n3471, new_n3470, new_n3472);
not_8  g03096(new_n3472, new_n3473);
xor_4  g03097(new_n3473, new_n3469, new_n3474);
and_5  g03098(new_n3407, new_n3406, new_n3475);
not_8  g03099(new_n3405, new_n3476);
nor_5  g03100(new_n3409, new_n3476, new_n3477);
or_5   g03101(new_n3477, new_n3475, new_n3478);
not_8  g03102(new_n3478, new_n3479);
xor_4  g03103(new_n3479, new_n3474, new_n3480);
nand_5 g03104(n11478, n4970, new_n3481);
nand_5 g03105(n7610, n5283, new_n3482);
xor_4  g03106(new_n3482, new_n3481, new_n3483);
xor_4  g03107(new_n3483, new_n3480, new_n3484);
and_5  g03108(new_n3403, new_n3399, new_n3485);
and_5  g03109(new_n3410, new_n3404, new_n3486);
nor_5  g03110(new_n3486, new_n3485, new_n3487);
xor_4  g03111(new_n3487, new_n3484, new_n3488);
nor_5  g03112(new_n3412, new_n3397, new_n3489);
and_5  g03113(new_n3416, new_n3413, new_n3490);
nor_5  g03114(new_n3490, new_n3489, new_n3491);
xor_4  g03115(new_n3491, new_n3488, new_n3492);
xor_4  g03116(new_n3492, new_n3468, new_n3493);
not_8  g03117(new_n3493, new_n3494);
nand_5 g03118(new_n3494, new_n3466, new_n3495);
or_5   g03119(new_n3494, new_n3466, new_n3496);
and_5  g03120(new_n3496, new_n3495, new_n3497);
xor_4  g03121(new_n3497, new_n3464, new_n3498);
nor_5  g03122(new_n3423, new_n3419, new_n3499);
nor_5  g03123(new_n3425, new_n3395, new_n3500);
nor_5  g03124(new_n3500, new_n3499, new_n3501);
xor_4  g03125(new_n3501, new_n3498, new_n3502);
xor_4  g03126(new_n3502, new_n3431, new_n3503);
and_5  g03127(new_n3503, new_n3173, new_n3504);
nor_5  g03128(new_n3503, new_n3173, new_n3505);
xor_4  g03129(new_n3165, new_n3164, new_n3506);
not_8  g03130(new_n3506, new_n3507);
xor_4  g03131(new_n3369, new_n3259, new_n3508);
xor_4  g03132(new_n3508, new_n3426, new_n3509);
or_5   g03133(new_n3509, new_n3507, new_n3510);
xor_4  g03134(new_n3163, new_n3158, new_n3511);
not_8  g03135(new_n3511, new_n3512);
xor_4  g03136(new_n3366, new_n3364, new_n3513);
nor_5  g03137(new_n3513, new_n3512, new_n3514);
or_5   g03138(new_n3319, new_n3314, new_n3515);
xor_4  g03139(new_n3515, new_n3308, new_n3516);
not_8  g03140(new_n3106, new_n3517);
nand_5 g03141(n9956, n7862, new_n3518);
and_5  g03142(new_n3518, new_n3517, new_n3519);
nor_5  g03143(new_n3519, new_n3159, new_n3520);
nand_5 g03144(new_n3103, new_n3102, new_n3521);
and_5  g03145(new_n3519, new_n3521, new_n3522);
or_5   g03146(new_n3522, new_n3520, new_n3523);
and_5  g03147(new_n3523, new_n3516, new_n3524);
nor_5  g03148(new_n3522, new_n3520, new_n3525);
xor_4  g03149(new_n3525, new_n3516, new_n3526);
not_8  g03150(new_n3518, new_n3527);
xor_4  g03151(new_n3316, new_n3194, new_n3528);
nand_5 g03152(new_n3528, new_n3527, new_n3529);
xnor_4 g03153(new_n3161, new_n3160, new_n3530);
and_5  g03154(new_n3530, new_n3529, new_n3531);
xor_4  g03155(new_n3318, new_n3317, new_n3532);
xor_4  g03156(new_n3530, new_n3529, new_n3533);
not_8  g03157(new_n3533, new_n3534);
nor_5  g03158(new_n3534, new_n3532, new_n3535);
or_5   g03159(new_n3535, new_n3531, new_n3536);
not_8  g03160(new_n3536, new_n3537);
nor_5  g03161(new_n3537, new_n3526, new_n3538);
or_5   g03162(new_n3538, new_n3524, new_n3539);
xor_4  g03163(new_n3513, new_n3511, new_n3540);
or_5   g03164(new_n3540, new_n3539, new_n3541);
not_8  g03165(new_n3541, new_n3542);
nor_5  g03166(new_n3542, new_n3514, new_n3543);
not_8  g03167(new_n3543, new_n3544);
xor_4  g03168(new_n3509, new_n3506, new_n3545);
not_8  g03169(new_n3545, new_n3546);
nand_5 g03170(new_n3546, new_n3544, new_n3547);
nand_5 g03171(new_n3547, new_n3510, new_n3548);
nor_5  g03172(new_n3548, new_n3505, new_n3549);
or_5   g03173(new_n3549, new_n3504, new_n3550);
not_8  g03174(new_n3550, new_n3551);
or_5   g03175(new_n3551, new_n3171, new_n3552);
nand_5 g03176(new_n3551, new_n3171, new_n3553);
and_5  g03177(new_n3553, new_n3552, new_n3554);
or_5   g03178(new_n3253, new_n3250, new_n3555);
nand_5 g03179(n9400, n8065, new_n3556);
nand_5 g03180(n10439, n2464, new_n3557);
and_5  g03181(n10391, n6877, new_n3558);
xor_4  g03182(new_n3558, new_n3557, new_n3559);
not_8  g03183(new_n3559, new_n3560);
xor_4  g03184(new_n3560, new_n3556, new_n3561);
nor_5  g03185(new_n3237, new_n3233, new_n3562);
and_5  g03186(new_n3242, new_n3238, new_n3563);
or_5   g03187(new_n3563, new_n3562, new_n3564);
not_8  g03188(new_n3564, new_n3565);
xor_4  g03189(new_n3565, new_n3561, new_n3566);
or_5   g03190(new_n3235, new_n3234, new_n3567);
not_8  g03191(new_n3567, new_n3568);
nand_5 g03192(n11311, n8595, new_n3569);
not_8  g03193(new_n3569, new_n3570);
xor_4  g03194(new_n3570, new_n3568, new_n3571);
nand_5 g03195(n4203, n3602, new_n3572);
nand_5 g03196(n6126, n4187, new_n3573);
nand_5 g03197(n12753, n3719, new_n3574);
xor_4  g03198(new_n3574, new_n3573, new_n3575);
not_8  g03199(new_n3575, new_n3576);
xor_4  g03200(new_n3576, new_n3572, new_n3577);
xor_4  g03201(new_n3577, new_n3571, new_n3578);
xor_4  g03202(new_n3578, new_n3566, new_n3579);
not_8  g03203(new_n3579, new_n3580);
and_5  g03204(new_n3246, new_n3243, new_n3581);
or_5   g03205(new_n3245, new_n3244, new_n3582);
not_8  g03206(new_n3582, new_n3583);
not_8  g03207(new_n3247, new_n3584);
or_5   g03208(new_n3249, new_n3584, new_n3585);
not_8  g03209(new_n3585, new_n3586);
xor_4  g03210(new_n3586, new_n3583, new_n3587);
nor_5  g03211(new_n3587, new_n3581, new_n3588);
xor_4  g03212(new_n3588, new_n3580, new_n3589);
not_8  g03213(new_n3589, new_n3590);
xor_4  g03214(new_n3590, new_n3555, new_n3591);
nor_5  g03215(new_n3254, new_n3232, new_n3592);
nor_5  g03216(new_n3256, new_n3230_1, new_n3593);
or_5   g03217(new_n3593, new_n3592, new_n3594);
xor_4  g03218(new_n3594, new_n3591, new_n3595);
not_8  g03219(new_n3595, new_n3596);
or_5   g03220(new_n3491, new_n3488, new_n3597);
not_8  g03221(new_n3597, new_n3598);
nand_5 g03222(n10965, n4805, new_n3599);
not_8  g03223(new_n3599, new_n3600);
nand_5 g03224(n5283, n4970, new_n3601);
nand_5 g03225(n11478, n503, new_n3602_1);
xor_4  g03226(new_n3602_1, new_n3601, new_n3603);
not_8  g03227(new_n3603, new_n3604);
xor_4  g03228(new_n3604, new_n3600, new_n3605);
nor_5  g03229(new_n3473, new_n3469, new_n3606);
and_5  g03230(new_n3479, new_n3474, new_n3607);
or_5   g03231(new_n3607, new_n3606, new_n3608);
not_8  g03232(new_n3608, new_n3609);
xor_4  g03233(new_n3609, new_n3605, new_n3610);
or_5   g03234(new_n3471, new_n3470, new_n3611);
not_8  g03235(new_n3611, new_n3612);
nand_5 g03236(n7610, n137, new_n3613);
not_8  g03237(new_n3613, new_n3614);
xor_4  g03238(new_n3614, new_n3612, new_n3615);
and_5  g03239(n7733, n6797, new_n3616_1);
nand_5 g03240(n6294, n4826, new_n3617);
nand_5 g03241(n12925, n3146, new_n3618);
xor_4  g03242(new_n3618, new_n3617, new_n3619);
xor_4  g03243(new_n3619, new_n3616_1, new_n3620);
xor_4  g03244(new_n3620, new_n3615, new_n3621);
xor_4  g03245(new_n3621, new_n3610, new_n3622);
not_8  g03246(new_n3622, new_n3623);
and_5  g03247(new_n3483, new_n3480, new_n3624);
or_5   g03248(new_n3482, new_n3481, new_n3625);
not_8  g03249(new_n3625, new_n3626);
not_8  g03250(new_n3484, new_n3627_1);
or_5   g03251(new_n3487, new_n3627_1, new_n3628);
not_8  g03252(new_n3628, new_n3629);
xor_4  g03253(new_n3629, new_n3626, new_n3630);
nor_5  g03254(new_n3630, new_n3624, new_n3631);
xor_4  g03255(new_n3631, new_n3623, new_n3632);
not_8  g03256(new_n3632, new_n3633);
xnor_4 g03257(new_n3633, new_n3598, new_n3634);
not_8  g03258(new_n3634, new_n3635);
or_5   g03259(new_n3492, new_n3468, new_n3636);
nand_5 g03260(new_n3496, new_n3636, new_n3637);
xor_4  g03261(new_n3637, new_n3635, new_n3638);
not_8  g03262(new_n3638, new_n3639);
or_5   g03263(new_n3460, new_n3457, new_n3640);
not_8  g03264(new_n3640, new_n3641);
nand_5 g03265(n11296, n7236, new_n3642);
not_8  g03266(new_n3642, new_n3643);
nand_5 g03267(n8384, n6611, new_n3644);
nand_5 g03268(n6359, n3992, new_n3645);
xor_4  g03269(new_n3645, new_n3644, new_n3646);
not_8  g03270(new_n3646, new_n3647);
xor_4  g03271(new_n3647, new_n3643, new_n3648);
and_5  g03272(new_n3441, new_n3436, new_n3649);
and_5  g03273(new_n3445, new_n3442, new_n3650);
or_5   g03274(new_n3650, new_n3649, new_n3651);
not_8  g03275(new_n3651, new_n3652);
xor_4  g03276(new_n3652, new_n3648, new_n3653);
or_5   g03277(new_n3444, new_n3443, new_n3654_1);
not_8  g03278(new_n3654_1, new_n3655);
nand_5 g03279(n6358, n217, new_n3656);
not_8  g03280(new_n3656, new_n3657);
xor_4  g03281(new_n3657, new_n3655, new_n3658);
and_5  g03282(n1471, n405, new_n3659);
nand_5 g03283(n5198, n4086, new_n3660);
nand_5 g03284(n8433, n7646, new_n3661_1);
xor_4  g03285(new_n3661_1, new_n3660, new_n3662);
xor_4  g03286(new_n3662, new_n3659, new_n3663);
xor_4  g03287(new_n3663, new_n3658, new_n3664);
xor_4  g03288(new_n3664, new_n3653, new_n3665);
not_8  g03289(new_n3665, new_n3666);
nor_5  g03290(new_n3451, new_n3447, new_n3667);
or_5   g03291(new_n3449, new_n3448, new_n3668);
not_8  g03292(new_n3668, new_n3669);
nand_5 g03293(new_n3455, new_n3452, new_n3670);
not_8  g03294(new_n3670, new_n3671);
xor_4  g03295(new_n3671, new_n3669, new_n3672);
nor_5  g03296(new_n3672, new_n3667, new_n3673);
xor_4  g03297(new_n3673, new_n3666, new_n3674);
not_8  g03298(new_n3674, new_n3675);
xnor_4 g03299(new_n3675, new_n3641, new_n3676);
or_5   g03300(new_n3461, new_n3434, new_n3677_1);
nor_5  g03301(new_n3394, new_n3372, new_n3678);
or_5   g03302(new_n3463, new_n3678, new_n3679);
nand_5 g03303(new_n3679, new_n3677_1, new_n3680);
xor_4  g03304(new_n3680, new_n3676, new_n3681);
not_8  g03305(new_n3681, new_n3682);
xnor_4 g03306(new_n3682, new_n3639, new_n3683);
not_8  g03307(new_n3497, new_n3684);
nor_5  g03308(new_n3684, new_n3464, new_n3685);
nor_5  g03309(new_n3501, new_n3498, new_n3686);
or_5   g03310(new_n3686, new_n3685, new_n3687);
not_8  g03311(new_n3687, new_n3688);
xor_4  g03312(new_n3688, new_n3683, new_n3689);
xor_4  g03313(new_n3689, new_n3596, new_n3690);
and_5  g03314(new_n3430, new_n3258, new_n3691);
not_8  g03315(new_n3431, new_n3692);
nor_5  g03316(new_n3502, new_n3692, new_n3693);
or_5   g03317(new_n3693, new_n3691, new_n3694);
not_8  g03318(new_n3694, new_n3695);
and_5  g03319(new_n3695, new_n3690, new_n3696);
nor_5  g03320(new_n3695, new_n3690, new_n3697);
or_5   g03321(new_n3697, new_n3696, new_n3698);
xor_4  g03322(new_n3698, new_n3554, n844);
nand_5 g03323(n7456, n6687, new_n3700);
not_8  g03324(new_n3700, new_n3701);
and_5  g03325(n12591, n6687, new_n3702);
and_5  g03326(n4189, n1798, new_n3703);
nor_5  g03327(new_n3703, new_n3702, new_n3704);
nand_5 g03328(n6687, n1798, new_n3705);
nand_5 g03329(n12591, n4189, new_n3706);
nor_5  g03330(new_n3706, new_n3705, new_n3707);
and_5  g03331(n3932, n2564, new_n3708);
nor_5  g03332(new_n3708, new_n3707, new_n3709);
or_5   g03333(new_n3709, new_n3704, new_n3710);
not_8  g03334(new_n3710, new_n3711);
and_5  g03335(new_n3711, new_n3701, new_n3712);
nor_5  g03336(new_n3711, new_n3701, new_n3713);
or_5   g03337(new_n3713, new_n3712, new_n3714);
nand_5 g03338(n4189, n3932, new_n3715);
not_8  g03339(new_n3715, new_n3716);
nand_5 g03340(n12591, n2564, new_n3717);
nand_5 g03341(n6770, n1798, new_n3718);
xor_4  g03342(new_n3718, new_n3717, new_n3719_1);
xor_4  g03343(new_n3719_1, new_n3716, new_n3720);
xor_4  g03344(new_n3720, new_n3714, new_n3721);
nand_5 g03345(new_n3708, new_n3705, new_n3722);
not_8  g03346(new_n3722, new_n3723);
nor_5  g03347(new_n3707, new_n3704, new_n3724);
or_5   g03348(new_n3724, new_n3723, new_n3725);
not_8  g03349(new_n3725, new_n3726);
nand_5 g03350(new_n3726, new_n3708, new_n3727);
xor_4  g03351(new_n3727, new_n3721, new_n3728);
not_8  g03352(new_n3728, new_n3729);
nor_5  g03353(new_n3722, new_n3704, new_n3730);
or_5   g03354(new_n3730, new_n3726, new_n3731);
nand_5 g03355(n8336, n6703, new_n3732);
not_8  g03356(new_n3732, new_n3733);
nand_5 g03357(n11876, n11222, new_n3734);
nand_5 g03358(n12069, n5645, new_n3735);
xnor_4 g03359(new_n3735, new_n3734, new_n3736);
not_8  g03360(new_n3736, new_n3737);
nand_5 g03361(new_n3737, new_n3733, new_n3738);
nand_5 g03362(n9640, n8336, new_n3739);
and_5  g03363(n10928, n6703, new_n3740);
xor_4  g03364(new_n3740, new_n3739, new_n3741);
nor_5  g03365(new_n3741, new_n3738, new_n3742);
or_5   g03366(new_n3735, new_n3734, new_n3743);
and_5  g03367(n12391, n5645, new_n3744);
and_5  g03368(n12069, n1067, new_n3745);
xor_4  g03369(new_n3745, new_n3744, new_n3746);
xor_4  g03370(new_n3746, new_n3743, new_n3747);
not_8  g03371(new_n3747, new_n3748);
nand_5 g03372(n11222, n10898, new_n3749);
and_5  g03373(n11876, n11153, new_n3750);
xor_4  g03374(new_n3750, new_n3749, new_n3751);
xor_4  g03375(new_n3751, new_n3748, new_n3752);
xor_4  g03376(new_n3741, new_n3738, new_n3753);
not_8  g03377(new_n3753, new_n3754_1);
nor_5  g03378(new_n3754_1, new_n3752, new_n3755);
or_5   g03379(new_n3755, new_n3742, new_n3756);
not_8  g03380(new_n3756, new_n3757);
nand_5 g03381(n10928, n9640, new_n3758);
or_5   g03382(new_n3758, new_n3733, new_n3759);
not_8  g03383(new_n3759, new_n3760);
and_5  g03384(n6986, n6703, new_n3761);
and_5  g03385(n8336, n3022, new_n3762);
nor_5  g03386(new_n3762, new_n3761, new_n3763);
nand_5 g03387(n6986, n3022, new_n3764);
nor_5  g03388(new_n3764, new_n3732, new_n3765);
nor_5  g03389(new_n3765, new_n3763, new_n3766);
or_5   g03390(new_n3766, new_n3760, new_n3767);
not_8  g03391(new_n3767, new_n3768);
nor_5  g03392(new_n3763, new_n3759, new_n3769);
or_5   g03393(new_n3769, new_n3768, new_n3770);
xor_4  g03394(new_n3770, new_n3757, new_n3771);
nand_5 g03395(new_n3745, new_n3744, new_n3772);
and_5  g03396(n12069, n8665, new_n3773);
not_8  g03397(new_n3773, new_n3774);
nand_5 g03398(n12391, n1067, new_n3775);
and_5  g03399(n7891, n5645, new_n3776);
xor_4  g03400(new_n3776, new_n3775, new_n3777);
not_8  g03401(new_n3777, new_n3778);
xor_4  g03402(new_n3778, new_n3774, new_n3779);
xor_4  g03403(new_n3779, new_n3772, new_n3780);
not_8  g03404(new_n3743, new_n3781);
nor_5  g03405(new_n3746, new_n3781, new_n3782);
and_5  g03406(new_n3751, new_n3748, new_n3783);
or_5   g03407(new_n3783, new_n3782, new_n3784);
not_8  g03408(new_n3784, new_n3785);
not_8  g03409(new_n3734, new_n3786);
nand_5 g03410(n11153, n10898, new_n3787);
or_5   g03411(new_n3787, new_n3786, new_n3788);
and_5  g03412(n11876, n5314, new_n3789);
and_5  g03413(n11222, n3754, new_n3790);
or_5   g03414(new_n3790, new_n3789, new_n3791);
not_8  g03415(new_n3791, new_n3792);
and_5  g03416(new_n3792, new_n3788, new_n3793);
nand_5 g03417(n5314, n3754, new_n3794);
nor_5  g03418(new_n3794, new_n3734, new_n3795);
or_5   g03419(new_n3795, new_n3793, new_n3796);
not_8  g03420(new_n3796, new_n3797);
or_5   g03421(new_n3792, new_n3788, new_n3798);
and_5  g03422(new_n3798, new_n3797, new_n3799);
xor_4  g03423(new_n3799, new_n3785, new_n3800);
xor_4  g03424(new_n3800, new_n3780, new_n3801);
not_8  g03425(new_n3801, new_n3802);
xor_4  g03426(new_n3802, new_n3771, new_n3803);
nor_5  g03427(new_n3803, new_n3731, new_n3804);
not_8  g03428(new_n3705, new_n3805);
xor_4  g03429(new_n3737, new_n3733, new_n3806);
nand_5 g03430(new_n3806, new_n3805, new_n3807);
nand_5 g03431(n2564, n1798, new_n3808);
and_5  g03432(n6687, n3932, new_n3809);
xor_4  g03433(new_n3809, new_n3808, new_n3810);
and_5  g03434(new_n3810, new_n3807, new_n3811);
xnor_4 g03435(new_n3753, new_n3752, new_n3812);
xor_4  g03436(new_n3810, new_n3807, new_n3813);
not_8  g03437(new_n3813, new_n3814);
nor_5  g03438(new_n3814, new_n3812, new_n3815);
or_5   g03439(new_n3815, new_n3811, new_n3816);
not_8  g03440(new_n3816, new_n3817);
xor_4  g03441(new_n3803, new_n3731, new_n3818);
and_5  g03442(new_n3818, new_n3817, new_n3819);
nor_5  g03443(new_n3819, new_n3804, new_n3820);
xor_4  g03444(new_n3820, new_n3729, new_n3821);
not_8  g03445(new_n3821, new_n3822);
or_5   g03446(new_n3779, new_n3772, new_n3823);
not_8  g03447(new_n3823, new_n3824);
nand_5 g03448(n12069, n11922, new_n3825);
not_8  g03449(new_n3825, new_n3826);
nand_5 g03450(n7891, n5645, new_n3827);
and_5  g03451(new_n3827, new_n3775, new_n3828);
and_5  g03452(new_n3778, new_n3774, new_n3829);
nor_5  g03453(new_n3829, new_n3828, new_n3830);
not_8  g03454(new_n3830, new_n3831);
xor_4  g03455(new_n3831, new_n3826, new_n3832);
and_5  g03456(n7160, n5645, new_n3833);
not_8  g03457(new_n3833, new_n3834);
nand_5 g03458(n7891, n1067, new_n3835);
and_5  g03459(n12391, n8665, new_n3836);
xor_4  g03460(new_n3836, new_n3835, new_n3837);
not_8  g03461(new_n3837, new_n3838);
xor_4  g03462(new_n3838, new_n3834, new_n3839);
xor_4  g03463(new_n3839, new_n3832, new_n3840);
not_8  g03464(new_n3840, new_n3841);
xor_4  g03465(new_n3841, new_n3824, new_n3842_1);
nand_5 g03466(n11222, n2749, new_n3843);
not_8  g03467(new_n3787, new_n3844);
nor_5  g03468(new_n3795, new_n3844, new_n3845);
or_5   g03469(new_n3845, new_n3792, new_n3846);
not_8  g03470(new_n3846, new_n3847);
xor_4  g03471(new_n3847, new_n3843, new_n3848);
and_5  g03472(n10898, n5314, new_n3849_1);
not_8  g03473(new_n3849_1, new_n3850);
nand_5 g03474(n11153, n3754, new_n3851);
and_5  g03475(n11876, n996, new_n3852);
xor_4  g03476(new_n3852, new_n3851, new_n3853);
not_8  g03477(new_n3853, new_n3854);
xor_4  g03478(new_n3854, new_n3850, new_n3855);
xor_4  g03479(new_n3855, new_n3848, new_n3856);
nor_5  g03480(new_n3797, new_n3787, new_n3857);
xnor_4 g03481(new_n3857, new_n3856, new_n3858);
xor_4  g03482(new_n3858, new_n3842_1, new_n3859);
not_8  g03483(new_n3859, new_n3860);
nor_5  g03484(new_n3799, new_n3785, new_n3861);
not_8  g03485(new_n3780, new_n3862);
and_5  g03486(new_n3800, new_n3862, new_n3863);
nor_5  g03487(new_n3863, new_n3861, new_n3864);
xor_4  g03488(new_n3864, new_n3860, new_n3865_1);
not_8  g03489(new_n3865_1, new_n3866);
nand_5 g03490(n11023, n8336, new_n3867);
not_8  g03491(new_n3867, new_n3868);
not_8  g03492(new_n3758, new_n3869);
nor_5  g03493(new_n3765, new_n3869, new_n3870);
nor_5  g03494(new_n3870, new_n3763, new_n3871);
not_8  g03495(new_n3871, new_n3872);
xor_4  g03496(new_n3872, new_n3868, new_n3873);
nand_5 g03497(n9640, n6986, new_n3874);
not_8  g03498(new_n3874, new_n3875);
nand_5 g03499(n10928, n3022, new_n3876);
nand_5 g03500(n6703, n2226, new_n3877);
xor_4  g03501(new_n3877, new_n3876, new_n3878);
xor_4  g03502(new_n3878, new_n3875, new_n3879);
not_8  g03503(new_n3879, new_n3880);
xor_4  g03504(new_n3880, new_n3873, new_n3881);
nand_5 g03505(new_n3768, new_n3869, new_n3882);
xor_4  g03506(new_n3882, new_n3881, new_n3883);
not_8  g03507(new_n3883, new_n3884);
and_5  g03508(new_n3770, new_n3757, new_n3885);
and_5  g03509(new_n3802, new_n3771, new_n3886);
or_5   g03510(new_n3886, new_n3885, new_n3887);
not_8  g03511(new_n3887, new_n3888);
xor_4  g03512(new_n3888, new_n3884, new_n3889);
xor_4  g03513(new_n3889, new_n3866, new_n3890);
xnor_4 g03514(new_n3890, new_n3822, n911);
nand_5 g03515(n6687, n3842, new_n3892);
not_8  g03516(new_n3892, new_n3893);
and_5  g03517(n11917, n6687, new_n3894);
and_5  g03518(n9956, n4189, new_n3895);
nor_5  g03519(new_n3895, new_n3894, new_n3896);
nand_5 g03520(n9956, n6687, new_n3897);
nand_5 g03521(n11917, n4189, new_n3898);
nor_5  g03522(new_n3898, new_n3897, new_n3899);
nand_5 g03523(n4921, n2564, new_n3900);
not_8  g03524(new_n3900, new_n3901);
nor_5  g03525(new_n3901, new_n3899, new_n3902);
nor_5  g03526(new_n3902, new_n3896, new_n3903);
not_8  g03527(new_n3903, new_n3904);
xor_4  g03528(new_n3904, new_n3893, new_n3905);
nand_5 g03529(n4921, n4189, new_n3906);
not_8  g03530(new_n3906, new_n3907);
nand_5 g03531(n11917, n2564, new_n3908);
nand_5 g03532(n9956, n6770, new_n3909);
xor_4  g03533(new_n3909, new_n3908, new_n3910);
xor_4  g03534(new_n3910, new_n3907, new_n3911);
not_8  g03535(new_n3911, new_n3912);
xor_4  g03536(new_n3912, new_n3905, new_n3913);
nor_5  g03537(new_n3899, new_n3896, new_n3914);
nand_5 g03538(n9956, n2564, new_n3915);
nand_5 g03539(n6687, n4921, new_n3916);
or_5   g03540(new_n3916, new_n3915, new_n3917);
or_5   g03541(new_n3917, new_n3914, new_n3918);
not_8  g03542(new_n3918, new_n3919);
nand_5 g03543(new_n3919, new_n3913, new_n3920);
not_8  g03544(new_n3920, new_n3921);
nand_5 g03545(n6687, n2577, new_n3922);
nor_5  g03546(new_n3904, new_n3892, new_n3923);
nor_5  g03547(new_n3912, new_n3905, new_n3924);
nor_5  g03548(new_n3924, new_n3923, new_n3925);
xor_4  g03549(new_n3925, new_n3922, new_n3926);
not_8  g03550(new_n3926, new_n3927);
nand_5 g03551(n3842, n2564, new_n3928);
not_8  g03552(new_n3928, new_n3929);
and_5  g03553(new_n3909, new_n3908, new_n3930);
nor_5  g03554(new_n3909, new_n3908, new_n3931);
nor_5  g03555(new_n3931, new_n3907, new_n3932_1);
or_5   g03556(new_n3932_1, new_n3930, new_n3933);
not_8  g03557(new_n3933, new_n3934);
and_5  g03558(new_n3934, new_n3929, new_n3935);
nor_5  g03559(new_n3934, new_n3929, new_n3936);
or_5   g03560(new_n3936, new_n3935, new_n3937);
nand_5 g03561(n6770, n4921, new_n3938);
not_8  g03562(new_n3938, new_n3939);
nand_5 g03563(n9956, n9920, new_n3940);
xor_4  g03564(new_n3940, new_n3898, new_n3941);
not_8  g03565(new_n3941, new_n3942);
xor_4  g03566(new_n3942, new_n3939, new_n3943);
xor_4  g03567(new_n3943, new_n3937, new_n3944);
not_8  g03568(new_n3944, new_n3945);
xor_4  g03569(new_n3945, new_n3927, new_n3946);
xor_4  g03570(new_n3946, new_n3921, new_n3947);
not_8  g03571(new_n3947, new_n3948);
xor_4  g03572(new_n3919, new_n3913, new_n3949);
nand_5 g03573(n8595, n8336, new_n3950);
not_8  g03574(new_n3950, new_n3951);
and_5  g03575(n8336, n6126, new_n3952);
and_5  g03576(n6986, n3719, new_n3953);
nor_5  g03577(new_n3953, new_n3952, new_n3954);
nand_5 g03578(n8336, n3719, new_n3955);
nand_5 g03579(n6986, n6126, new_n3956);
nor_5  g03580(new_n3956, new_n3955, new_n3957);
nand_5 g03581(n10928, n3602, new_n3958);
not_8  g03582(new_n3958, new_n3959);
nor_5  g03583(new_n3959, new_n3957, new_n3960);
nor_5  g03584(new_n3960, new_n3954, new_n3961);
not_8  g03585(new_n3961, new_n3962);
xor_4  g03586(new_n3962, new_n3951, new_n3963);
nand_5 g03587(n6986, n3602, new_n3964);
not_8  g03588(new_n3964, new_n3965);
nand_5 g03589(n10928, n6126, new_n3966);
nand_5 g03590(n3719, n2226, new_n3967);
xor_4  g03591(new_n3967, new_n3966, new_n3968);
xor_4  g03592(new_n3968, new_n3965, new_n3969);
not_8  g03593(new_n3969, new_n3970);
xor_4  g03594(new_n3970, new_n3963, new_n3971);
not_8  g03595(new_n3955, new_n3972);
or_5   g03596(new_n3958, new_n3972, new_n3973);
not_8  g03597(new_n3973, new_n3974);
nor_5  g03598(new_n3957, new_n3954, new_n3975);
or_5   g03599(new_n3975, new_n3974, new_n3976);
not_8  g03600(new_n3976, new_n3977);
nand_5 g03601(new_n3977, new_n3959, new_n3978);
xor_4  g03602(new_n3978, new_n3971, new_n3979);
not_8  g03603(new_n3979, new_n3980);
nand_5 g03604(n12069, n7610, new_n3981);
not_8  g03605(new_n3981, new_n3982);
and_5  g03606(n12069, n4826, new_n3983);
and_5  g03607(n12925, n7891, new_n3984);
nor_5  g03608(new_n3984, new_n3983, new_n3985);
nand_5 g03609(n12925, n12069, new_n3986_1);
nand_5 g03610(n7891, n4826, new_n3987);
nor_5  g03611(new_n3987, new_n3986_1, new_n3988);
and_5  g03612(n12391, n7733, new_n3989);
nor_5  g03613(new_n3989, new_n3988, new_n3990);
nor_5  g03614(new_n3990, new_n3985, new_n3991);
not_8  g03615(new_n3991, new_n3992_1);
xor_4  g03616(new_n3992_1, new_n3982, new_n3993);
nand_5 g03617(n7891, n7733, new_n3994);
nand_5 g03618(n12925, n7160, new_n3995);
nand_5 g03619(n12391, n4826, new_n3996);
xnor_4 g03620(new_n3996, new_n3995, new_n3997);
not_8  g03621(new_n3997, new_n3998);
xor_4  g03622(new_n3998, new_n3994, new_n3999);
nor_5  g03623(new_n3999, new_n3993, new_n4000);
and_5  g03624(new_n3999, new_n3993, new_n4001);
or_5   g03625(new_n4001, new_n4000, new_n4002);
nor_5  g03626(new_n3988, new_n3985, new_n4003);
and_5  g03627(n12925, n12391, new_n4004);
and_5  g03628(n12069, n7733, new_n4005_1);
nand_5 g03629(new_n4005_1, new_n4004, new_n4006);
or_5   g03630(new_n4006, new_n4003, new_n4007);
xor_4  g03631(new_n4007, new_n4002, new_n4008);
nand_5 g03632(n11222, n217, new_n4009);
nand_5 g03633(n8433, n5314, new_n4010);
nand_5 g03634(n11222, n4086, new_n4011);
nand_5 g03635(new_n4011, new_n4010, new_n4012);
not_8  g03636(new_n4012, new_n4013);
nor_5  g03637(new_n4011, new_n4010, new_n4014);
nand_5 g03638(n11153, n405, new_n4015);
not_8  g03639(new_n4015, new_n4016);
nor_5  g03640(new_n4016, new_n4014, new_n4017);
nor_5  g03641(new_n4017, new_n4013, new_n4018);
not_8  g03642(new_n4018, new_n4019);
xor_4  g03643(new_n4019, new_n4009, new_n4020);
nand_5 g03644(n5314, n405, new_n4021);
not_8  g03645(new_n4021, new_n4022);
nand_5 g03646(n8433, n996, new_n4023);
nand_5 g03647(n11153, n4086, new_n4024);
xor_4  g03648(new_n4024, new_n4023, new_n4025);
xor_4  g03649(new_n4025, new_n4022, new_n4026);
xor_4  g03650(new_n4026, new_n4020, new_n4027);
nand_5 g03651(n11222, n8433, new_n4028);
not_8  g03652(new_n4028, new_n4029);
or_5   g03653(new_n4029, new_n4015, new_n4030);
and_5  g03654(new_n4030, new_n4013, new_n4031);
or_5   g03655(new_n4031, new_n4014, new_n4032);
not_8  g03656(new_n4032, new_n4033);
nor_5  g03657(new_n4033, new_n4015, new_n4034);
xor_4  g03658(new_n4034, new_n4027, new_n4035);
not_8  g03659(new_n4035, new_n4036);
xor_4  g03660(new_n4036, new_n4008, new_n4037);
or_5   g03661(new_n4028, new_n3986_1, new_n4038);
not_8  g03662(new_n4038, new_n4039);
and_5  g03663(n11153, n8433, new_n4040);
and_5  g03664(n11222, n405, new_n4041);
xor_4  g03665(new_n4041, new_n4040, new_n4042);
nor_5  g03666(new_n4042, new_n4039, new_n4043);
xor_4  g03667(new_n4042, new_n4038, new_n4044);
not_8  g03668(new_n4044, new_n4045);
xnor_4 g03669(new_n4005_1, new_n4004, new_n4046);
and_5  g03670(new_n4046, new_n4045, new_n4047);
or_5   g03671(new_n4047, new_n4043, new_n4048);
not_8  g03672(new_n4048, new_n4049);
or_5   g03673(new_n4030, new_n4013, new_n4050);
and_5  g03674(new_n4050, new_n4033, new_n4051);
nor_5  g03675(new_n4051, new_n4049, new_n4052);
xor_4  g03676(new_n4051, new_n4048, new_n4053);
nand_5 g03677(new_n3989, new_n3986_1, new_n4054);
not_8  g03678(new_n4054, new_n4055);
nor_5  g03679(new_n4055, new_n4003, new_n4056);
nor_5  g03680(new_n4054, new_n3985, new_n4057);
nor_5  g03681(new_n4057, new_n4056, new_n4058);
nor_5  g03682(new_n4058, new_n4053, new_n4059);
nor_5  g03683(new_n4059, new_n4052, new_n4060);
xor_4  g03684(new_n4060, new_n4037, new_n4061);
xor_4  g03685(new_n4061, new_n3980, new_n4062);
nor_5  g03686(new_n3973, new_n3954, new_n4063);
or_5   g03687(new_n4063, new_n3977, new_n4064);
xor_4  g03688(new_n4058, new_n4053, new_n4065);
nor_5  g03689(new_n4065, new_n4064, new_n4066);
xor_4  g03690(new_n4065, new_n4064, new_n4067);
not_8  g03691(new_n4067, new_n4068);
xor_4  g03692(new_n4046, new_n4045, new_n4069);
nand_5 g03693(n10928, n3719, new_n4070);
and_5  g03694(n8336, n3602, new_n4071);
xor_4  g03695(new_n4071, new_n4070, new_n4072);
nor_5  g03696(new_n4072, new_n4069, new_n4073);
xor_4  g03697(new_n4028, new_n3986_1, new_n4074);
not_8  g03698(new_n4074, new_n4075);
or_5   g03699(new_n4075, new_n3955, new_n4076);
not_8  g03700(new_n4076, new_n4077);
xor_4  g03701(new_n4072, new_n4069, new_n4078);
and_5  g03702(new_n4078, new_n4077, new_n4079);
nor_5  g03703(new_n4079, new_n4073, new_n4080);
nor_5  g03704(new_n4080, new_n4068, new_n4081);
nor_5  g03705(new_n4081, new_n4066, new_n4082);
xor_4  g03706(new_n4082, new_n4062, new_n4083);
nor_5  g03707(new_n4083, new_n3949, new_n4084);
xor_4  g03708(new_n4080, new_n4068, new_n4085);
not_8  g03709(new_n3897, new_n4086_1);
or_5   g03710(new_n3900, new_n4086_1, new_n4087);
not_8  g03711(new_n4087, new_n4088_1);
nor_5  g03712(new_n4088_1, new_n3914, new_n4089);
nor_5  g03713(new_n4087, new_n3896, new_n4090);
nor_5  g03714(new_n4090, new_n4089, new_n4091);
nor_5  g03715(new_n4091, new_n4085, new_n4092);
or_5   g03716(new_n4090, new_n4089, new_n4093);
xor_4  g03717(new_n4093, new_n4085, new_n4094_1);
xor_4  g03718(new_n4075, new_n3955, new_n4095);
nand_5 g03719(new_n4095, new_n4086_1, new_n4096);
xnor_4 g03720(new_n3916, new_n3915, new_n4097);
and_5  g03721(new_n4097, new_n4096, new_n4098);
xor_4  g03722(new_n4078, new_n4077, new_n4099);
xor_4  g03723(new_n4097, new_n4096, new_n4100);
not_8  g03724(new_n4100, new_n4101);
nor_5  g03725(new_n4101, new_n4099, new_n4102);
nor_5  g03726(new_n4102, new_n4098, new_n4103);
nor_5  g03727(new_n4103, new_n4094_1, new_n4104);
or_5   g03728(new_n4104, new_n4092, new_n4105);
not_8  g03729(new_n3949, new_n4106);
xor_4  g03730(new_n4083, new_n4106, new_n4107);
not_8  g03731(new_n4107, new_n4108);
and_5  g03732(new_n4108, new_n4105, new_n4109);
nor_5  g03733(new_n4109, new_n4084, new_n4110);
xor_4  g03734(new_n4110, new_n3948, new_n4111);
not_8  g03735(new_n4111, new_n4112);
not_8  g03736(new_n3978, new_n4113);
nand_5 g03737(new_n4113, new_n3971, new_n4114);
not_8  g03738(new_n4114, new_n4115);
nand_5 g03739(n10439, n8336, new_n4116);
nor_5  g03740(new_n3962, new_n3950, new_n4117);
nor_5  g03741(new_n3970, new_n3963, new_n4118);
nor_5  g03742(new_n4118, new_n4117, new_n4119);
xor_4  g03743(new_n4119, new_n4116, new_n4120);
not_8  g03744(new_n4120, new_n4121);
nand_5 g03745(n10928, n8595, new_n4122);
not_8  g03746(new_n4122, new_n4123);
and_5  g03747(new_n3967, new_n3966, new_n4124);
nor_5  g03748(new_n3967, new_n3966, new_n4125);
nor_5  g03749(new_n4125, new_n3965, new_n4126);
or_5   g03750(new_n4126, new_n4124, new_n4127);
not_8  g03751(new_n4127, new_n4128);
and_5  g03752(new_n4128, new_n4123, new_n4129);
nor_5  g03753(new_n4128, new_n4123, new_n4130);
or_5   g03754(new_n4130, new_n4129, new_n4131);
nand_5 g03755(n3602, n2226, new_n4132);
not_8  g03756(new_n4132, new_n4133);
nand_5 g03757(n3719, n1094, new_n4134);
xor_4  g03758(new_n4134, new_n3956, new_n4135);
not_8  g03759(new_n4135, new_n4136);
xor_4  g03760(new_n4136, new_n4133, new_n4137);
xor_4  g03761(new_n4137, new_n4131, new_n4138);
not_8  g03762(new_n4138, new_n4139);
xor_4  g03763(new_n4139, new_n4121, new_n4140);
xor_4  g03764(new_n4140, new_n4115, new_n4141_1);
not_8  g03765(new_n4141_1, new_n4142);
nand_5 g03766(new_n4034, new_n4027, new_n4143);
not_8  g03767(new_n4143, new_n4144);
nand_5 g03768(n11222, n6611, new_n4145);
not_8  g03769(new_n4145, new_n4146);
nand_5 g03770(n11153, n217, new_n4147);
nand_5 g03771(n996, n405, new_n4148);
not_8  g03772(new_n4148, new_n4149);
nand_5 g03773(n5314, n4086, new_n4150);
nand_5 g03774(n8433, n5767, new_n4151);
xor_4  g03775(new_n4151, new_n4150, new_n4152);
xor_4  g03776(new_n4152, new_n4149, new_n4153);
not_8  g03777(new_n4153, new_n4154);
xor_4  g03778(new_n4154, new_n4147, new_n4155_1);
and_5  g03779(new_n4024, new_n4023, new_n4156);
nor_5  g03780(new_n4024, new_n4023, new_n4157);
nor_5  g03781(new_n4157, new_n4022, new_n4158);
or_5   g03782(new_n4158, new_n4156, new_n4159_1);
not_8  g03783(new_n4159_1, new_n4160);
xor_4  g03784(new_n4160, new_n4155_1, new_n4161);
xor_4  g03785(new_n4161, new_n4146, new_n4162);
or_5   g03786(new_n4019, new_n4009, new_n4163);
not_8  g03787(new_n4163, new_n4164);
and_5  g03788(new_n4026, new_n4020, new_n4165);
or_5   g03789(new_n4165, new_n4164, new_n4166);
xor_4  g03790(new_n4166, new_n4162, new_n4167);
not_8  g03791(new_n4167, new_n4168);
xor_4  g03792(new_n4168, new_n4144, new_n4169);
not_8  g03793(new_n4169, new_n4170);
or_5   g03794(new_n4007, new_n4002, new_n4171);
nand_5 g03795(n12069, n4970, new_n4172);
nand_5 g03796(n12391, n7610, new_n4173);
not_8  g03797(new_n4173, new_n4174);
and_5  g03798(new_n3996, new_n3995, new_n4175);
and_5  g03799(new_n3998, new_n3994, new_n4176);
or_5   g03800(new_n4176, new_n4175, new_n4177);
not_8  g03801(new_n4177, new_n4178);
xor_4  g03802(new_n4178, new_n4174, new_n4179);
nand_5 g03803(n7733, n7160, new_n4180);
nand_5 g03804(n12925, n4828, new_n4181);
xor_4  g03805(new_n4181, new_n3987, new_n4182);
not_8  g03806(new_n4182, new_n4183);
xor_4  g03807(new_n4183, new_n4180, new_n4184);
xor_4  g03808(new_n4184, new_n4179, new_n4185);
not_8  g03809(new_n4185, new_n4186);
xor_4  g03810(new_n4186, new_n4172, new_n4187_1);
or_5   g03811(new_n3992_1, new_n3981, new_n4188);
or_5   g03812(new_n3999, new_n3993, new_n4189_1);
nand_5 g03813(new_n4189_1, new_n4188, new_n4190_1);
xor_4  g03814(new_n4190_1, new_n4187_1, new_n4191);
not_8  g03815(new_n4191, new_n4192);
xor_4  g03816(new_n4192, new_n4171, new_n4193);
not_8  g03817(new_n4008, new_n4194);
and_5  g03818(new_n4036, new_n4194, new_n4195);
nor_5  g03819(new_n4060, new_n4037, new_n4196);
nor_5  g03820(new_n4196, new_n4195, new_n4197);
xor_4  g03821(new_n4197, new_n4193, new_n4198);
not_8  g03822(new_n4198, new_n4199);
nand_5 g03823(new_n4199, new_n4170, new_n4200);
or_5   g03824(new_n4199, new_n4170, new_n4201);
and_5  g03825(new_n4201, new_n4200, new_n4202);
xor_4  g03826(new_n4202, new_n4142, new_n4203_1);
nor_5  g03827(new_n4061, new_n3979, new_n4204);
nor_5  g03828(new_n4082, new_n4062, new_n4205);
nor_5  g03829(new_n4205, new_n4204, new_n4206);
xor_4  g03830(new_n4206, new_n4203_1, new_n4207);
not_8  g03831(new_n4207, new_n4208);
xor_4  g03832(new_n4208, new_n4112, n992);
nand_5 g03833(n7265, n6687, new_n4210);
not_8  g03834(new_n4210, new_n4211);
nand_5 g03835(n8336, n7946, new_n4212);
nand_5 g03836(n11222, n9763, new_n4213);
nand_5 g03837(n12069, n2558, new_n4214);
xor_4  g03838(new_n4214, new_n4213, new_n4215);
not_8  g03839(new_n4215, new_n4216);
xor_4  g03840(new_n4216, new_n4212, new_n4217);
xor_4  g03841(new_n4217, new_n4211, n1020);
xor_4  g03842(new_n2056, new_n2054, n1136);
not_8  g03843(new_n4105, new_n4220);
xor_4  g03844(new_n4108, new_n4220, n1138);
nand_5 g03845(n12591, n11757, new_n4222);
nand_5 g03846(n5240, n3932, new_n4223);
nand_5 g03847(n11821, n1798, new_n4224);
xor_4  g03848(new_n4224, new_n4223, new_n4225);
not_8  g03849(new_n4225, new_n4226_1);
xor_4  g03850(new_n4226_1, new_n4222, new_n4227);
nand_5 g03851(n5240, n1798, new_n4228);
nand_5 g03852(n12591, n3172, new_n4229);
and_5  g03853(new_n4229, new_n4228, new_n4230_1);
nor_5  g03854(new_n4229, new_n4228, new_n4231);
nand_5 g03855(n11757, n3932, new_n4232);
not_8  g03856(new_n4232, new_n4233);
nor_5  g03857(new_n4233, new_n4231, new_n4234);
or_5   g03858(new_n4234, new_n4230_1, new_n4235);
not_8  g03859(new_n4235, new_n4236);
xor_4  g03860(new_n4236, new_n4227, new_n4237);
and_5  g03861(n7456, n1333, new_n4238);
nand_5 g03862(n11757, n1798, new_n4239);
nand_5 g03863(n12591, n1333, new_n4240);
and_5  g03864(new_n4240, new_n4239, new_n4241);
nor_5  g03865(new_n4240, new_n4239, new_n4242);
nand_5 g03866(n3932, n3172, new_n4243);
not_8  g03867(new_n4243, new_n4244);
nor_5  g03868(new_n4244, new_n4242, new_n4245);
or_5   g03869(new_n4245, new_n4241, new_n4246);
not_8  g03870(new_n4246, new_n4247);
and_5  g03871(new_n4247, new_n4238, new_n4248);
nor_5  g03872(new_n4247, new_n4238, new_n4249);
or_5   g03873(new_n4249, new_n4248, new_n4250);
xor_4  g03874(new_n4229, new_n4228, new_n4251);
xor_4  g03875(new_n4251, new_n4232, new_n4252);
nor_5  g03876(new_n4252, new_n4250, new_n4253);
or_5   g03877(new_n4253, new_n4248, new_n4254);
not_8  g03878(new_n4254, new_n4255);
nand_5 g03879(n11662, n1333, new_n4256);
nand_5 g03880(n7456, n3172, new_n4257);
xor_4  g03881(new_n4257, new_n4256, new_n4258);
not_8  g03882(new_n4258, new_n4259);
xor_4  g03883(new_n4259, new_n4255, new_n4260);
xor_4  g03884(new_n4260, new_n4237, new_n4261);
nand_5 g03885(n11662, n7862, new_n4262);
not_8  g03886(new_n4262, new_n4263);
xor_4  g03887(new_n4252, new_n4250, new_n4264);
nor_5  g03888(new_n4264, new_n4263, new_n4265);
xor_4  g03889(new_n4264, new_n4263, new_n4266);
not_8  g03890(new_n4266, new_n4267);
nand_5 g03891(n7862, n7456, new_n4268);
nand_5 g03892(n3172, n1798, new_n4269);
nand_5 g03893(n12591, n7862, new_n4270);
nor_5  g03894(new_n4270, new_n4269, new_n4271);
and_5  g03895(new_n4270, new_n4269, new_n4272);
nand_5 g03896(n3932, n1333, new_n4273);
nor_5  g03897(new_n4273, new_n4272, new_n4274);
nor_5  g03898(new_n4274, new_n4271, new_n4275);
nor_5  g03899(new_n4275, new_n4268, new_n4276);
xor_4  g03900(new_n4275, new_n4268, new_n4277);
not_8  g03901(new_n4277, new_n4278);
xor_4  g03902(new_n4240, new_n4239, new_n4279);
xor_4  g03903(new_n4279, new_n4243, new_n4280);
nor_5  g03904(new_n4280, new_n4278, new_n4281);
or_5   g03905(new_n4281, new_n4276, new_n4282);
nor_5  g03906(new_n4282, new_n4267, new_n4283);
or_5   g03907(new_n4283, new_n4265, new_n4284);
not_8  g03908(new_n4284, new_n4285);
nand_5 g03909(new_n4285, new_n4261, new_n4286);
nor_5  g03910(new_n4226_1, new_n4222, new_n4287);
and_5  g03911(new_n4236, new_n4227, new_n4288);
or_5   g03912(new_n4288, new_n4287, new_n4289);
nand_5 g03913(n10327, n1333, new_n4290);
not_8  g03914(new_n4290, new_n4291);
nand_5 g03915(n11662, n3172, new_n4292);
nand_5 g03916(n9583, n7862, new_n4293);
xor_4  g03917(new_n4293, new_n4292, new_n4294);
not_8  g03918(new_n4294, new_n4295);
xor_4  g03919(new_n4295, new_n4291, new_n4296);
not_8  g03920(new_n4296, new_n4297);
xor_4  g03921(new_n4297, new_n4289, new_n4298);
or_5   g03922(new_n4224, new_n4223, new_n4299);
nand_5 g03923(n11757, n7456, new_n4300_1);
not_8  g03924(new_n4300_1, new_n4301);
xor_4  g03925(new_n4301, new_n4299, new_n4302);
nand_5 g03926(n11821, n3932, new_n4303);
nand_5 g03927(n12591, n5240, new_n4304);
nand_5 g03928(n9080, n1798, new_n4305);
xor_4  g03929(new_n4305, new_n4304, new_n4306);
xor_4  g03930(new_n4306, new_n4303, new_n4307);
xor_4  g03931(new_n4307, new_n4302, new_n4308);
xor_4  g03932(new_n4308, new_n4298, new_n4309);
not_8  g03933(new_n4309, new_n4310);
nor_5  g03934(new_n4259, new_n4255, new_n4311);
or_5   g03935(new_n4257, new_n4256, new_n4312_1);
nand_5 g03936(new_n4260, new_n4237, new_n4313);
xor_4  g03937(new_n4313, new_n4312_1, new_n4314);
nor_5  g03938(new_n4314, new_n4311, new_n4315);
xor_4  g03939(new_n4315, new_n4310, new_n4316);
not_8  g03940(new_n4316, new_n4317);
nor_5  g03941(new_n4317, new_n4286, new_n4318);
and_5  g03942(new_n4317, new_n4286, new_n4319);
or_5   g03943(new_n4319, new_n4318, new_n4320);
nand_5 g03944(n10327, n7862, new_n4321);
not_8  g03945(new_n4321, new_n4322);
xor_4  g03946(new_n4285, new_n4261, new_n4323);
and_5  g03947(new_n4323, new_n4322, new_n4324);
and_5  g03948(new_n4280, new_n4278, new_n4325);
or_5   g03949(new_n4325, new_n4281, new_n4326_1);
xor_4  g03950(new_n4270, new_n4269, new_n4327);
nand_5 g03951(n1798, n1333, new_n4328);
nand_5 g03952(n7862, n3932, new_n4329);
or_5   g03953(new_n4329, new_n4328, new_n4330);
or_5   g03954(new_n4330, new_n4327, new_n4331);
or_5   g03955(new_n4331, new_n4326_1, new_n4332);
xor_4  g03956(new_n4282, new_n4267, new_n4333_1);
or_5   g03957(new_n4333_1, new_n4332, new_n4334);
xor_4  g03958(new_n4323, new_n4322, new_n4335);
not_8  g03959(new_n4335, new_n4336);
nor_5  g03960(new_n4336, new_n4334, new_n4337);
nor_5  g03961(new_n4337, new_n4324, new_n4338);
xor_4  g03962(new_n4338, new_n4320, new_n4339);
not_8  g03963(new_n4339, new_n4340);
nand_5 g03964(n11311, n3022, new_n4341);
nand_5 g03965(n9640, n4187, new_n4342);
nand_5 g03966(n6703, n4203, new_n4343);
xor_4  g03967(new_n4343, new_n4342, new_n4344);
not_8  g03968(new_n4344, new_n4345);
xor_4  g03969(new_n4345, new_n4341, new_n4346);
nand_5 g03970(n6703, n4187, new_n4347);
nand_5 g03971(n3022, n2464, new_n4348);
and_5  g03972(new_n4348, new_n4347, new_n4349);
nor_5  g03973(new_n4348, new_n4347, new_n4350);
nand_5 g03974(n11311, n9640, new_n4351);
not_8  g03975(new_n4351, new_n4352);
nor_5  g03976(new_n4352, new_n4350, new_n4353);
or_5   g03977(new_n4353, new_n4349, new_n4354);
not_8  g03978(new_n4354, new_n4355);
xor_4  g03979(new_n4355, new_n4346, new_n4356);
nand_5 g03980(n10451, n9400, new_n4357);
nand_5 g03981(n11023, n2464, new_n4358);
xor_4  g03982(new_n4358, new_n4357, new_n4359);
xor_4  g03983(new_n4359, new_n4356, new_n4360);
not_8  g03984(new_n4360, new_n4361);
nand_5 g03985(n11023, n9400, new_n4362);
not_8  g03986(new_n4362, new_n4363);
nand_5 g03987(n11311, n6703, new_n4364);
nand_5 g03988(n9400, n3022, new_n4365);
and_5  g03989(new_n4365, new_n4364, new_n4366);
nor_5  g03990(new_n4365, new_n4364, new_n4367);
nand_5 g03991(n9640, n2464, new_n4368);
not_8  g03992(new_n4368, new_n4369);
nor_5  g03993(new_n4369, new_n4367, new_n4370_1);
or_5   g03994(new_n4370_1, new_n4366, new_n4371);
not_8  g03995(new_n4371, new_n4372);
and_5  g03996(new_n4372, new_n4363, new_n4373);
nor_5  g03997(new_n4372, new_n4363, new_n4374);
or_5   g03998(new_n4374, new_n4373, new_n4375);
xor_4  g03999(new_n4348, new_n4347, new_n4376);
xor_4  g04000(new_n4376, new_n4351, new_n4377);
nor_5  g04001(new_n4377, new_n4375, new_n4378_1);
nor_5  g04002(new_n4378_1, new_n4373, new_n4379);
xor_4  g04003(new_n4379, new_n4361, new_n4380);
not_8  g04004(new_n4380, new_n4381);
nand_5 g04005(n10451, n6877, new_n4382);
not_8  g04006(new_n4382, new_n4383);
xor_4  g04007(new_n4377, new_n4375, new_n4384);
and_5  g04008(new_n4384, new_n4383, new_n4385);
nand_5 g04009(n11023, n6877, new_n4386);
not_8  g04010(new_n4386, new_n4387);
nand_5 g04011(n6703, n2464, new_n4388);
nand_5 g04012(n6877, n3022, new_n4389);
and_5  g04013(new_n4389, new_n4388, new_n4390);
nor_5  g04014(new_n4389, new_n4388, new_n4391);
nand_5 g04015(n9640, n9400, new_n4392);
not_8  g04016(new_n4392, new_n4393);
nor_5  g04017(new_n4393, new_n4391, new_n4394);
or_5   g04018(new_n4394, new_n4390, new_n4395);
not_8  g04019(new_n4395, new_n4396);
and_5  g04020(new_n4396, new_n4387, new_n4397_1);
nor_5  g04021(new_n4396, new_n4387, new_n4398);
or_5   g04022(new_n4398, new_n4397_1, new_n4399);
xor_4  g04023(new_n4365, new_n4364, new_n4400);
xor_4  g04024(new_n4400, new_n4368, new_n4401);
nor_5  g04025(new_n4401, new_n4399, new_n4402);
or_5   g04026(new_n4402, new_n4397_1, new_n4403);
not_8  g04027(new_n4403, new_n4404);
xor_4  g04028(new_n4384, new_n4383, new_n4405);
not_8  g04029(new_n4405, new_n4406);
nor_5  g04030(new_n4406, new_n4404, new_n4407);
nor_5  g04031(new_n4407, new_n4385, new_n4408);
or_5   g04032(new_n4408, new_n4381, new_n4409);
not_8  g04033(new_n4409, new_n4410);
nor_5  g04034(new_n4345, new_n4341, new_n4411);
and_5  g04035(new_n4355, new_n4346, new_n4412);
or_5   g04036(new_n4412, new_n4411, new_n4413);
nand_5 g04037(n10278, n9400, new_n4414);
nand_5 g04038(n10451, n2464, new_n4415);
nand_5 g04039(n11423, n6877, new_n4416);
xor_4  g04040(new_n4416, new_n4415, new_n4417);
xor_4  g04041(new_n4417, new_n4414, new_n4418);
not_8  g04042(new_n4418, new_n4419);
xor_4  g04043(new_n4419, new_n4413, new_n4420);
or_5   g04044(new_n4343, new_n4342, new_n4421);
not_8  g04045(new_n4421, new_n4422);
nand_5 g04046(n11311, n11023, new_n4423);
not_8  g04047(new_n4423, new_n4424);
xor_4  g04048(new_n4424, new_n4422, new_n4425);
and_5  g04049(n9640, n4203, new_n4426);
nand_5 g04050(n4187, n3022, new_n4427);
nand_5 g04051(n12753, n6703, new_n4428);
xor_4  g04052(new_n4428, new_n4427, new_n4429);
xor_4  g04053(new_n4429, new_n4426, new_n4430);
xor_4  g04054(new_n4430, new_n4425, new_n4431);
xor_4  g04055(new_n4431, new_n4420, new_n4432);
not_8  g04056(new_n4432, new_n4433);
nand_5 g04057(new_n4359, new_n4356, new_n4434);
or_5   g04058(new_n4358, new_n4357, new_n4435);
or_5   g04059(new_n4379, new_n4361, new_n4436_1);
not_8  g04060(new_n4436_1, new_n4437);
xor_4  g04061(new_n4437, new_n4435, new_n4438);
and_5  g04062(new_n4438, new_n4434, new_n4439);
xor_4  g04063(new_n4439, new_n4433, new_n4440);
xnor_4 g04064(new_n4440, new_n4410, new_n4441);
nand_5 g04065(n10278, n6877, new_n4442);
xor_4  g04066(new_n4408, new_n4381, new_n4443);
not_8  g04067(new_n4443, new_n4444);
nor_5  g04068(new_n4444, new_n4442, new_n4445);
xor_4  g04069(new_n4401, new_n4399, new_n4446);
nand_5 g04070(n6877, n6703, new_n4447);
not_8  g04071(new_n4447, new_n4448);
or_5   g04072(new_n4448, new_n4392, new_n4449);
xnor_4 g04073(new_n4389, new_n4388, new_n4450);
and_5  g04074(new_n4450, new_n4449, new_n4451);
not_8  g04075(new_n4451, new_n4452);
or_5   g04076(new_n4452, new_n4392, new_n4453);
not_8  g04077(new_n4453, new_n4454);
nand_5 g04078(new_n4454, new_n4446, new_n4455);
not_8  g04079(new_n4455, new_n4456);
xor_4  g04080(new_n4406, new_n4404, new_n4457);
nand_5 g04081(new_n4457, new_n4456, new_n4458);
not_8  g04082(new_n4458, new_n4459);
xor_4  g04083(new_n4444, new_n4442, new_n4460);
and_5  g04084(new_n4460, new_n4459, new_n4461);
nor_5  g04085(new_n4461, new_n4445, new_n4462);
xor_4  g04086(new_n4462, new_n4441, new_n4463);
nand_5 g04087(n12826, n4805, new_n4464);
not_8  g04088(new_n4464, new_n4465);
nand_5 g04089(n8665, n137, new_n4466);
nand_5 g04090(n6294, n1067, new_n4467);
nand_5 g04091(n6797, n5645, new_n4468);
xor_4  g04092(new_n4468, new_n4467, new_n4469);
not_8  g04093(new_n4469, new_n4470);
xor_4  g04094(new_n4470, new_n4466, new_n4471);
nand_5 g04095(n6294, n5645, new_n4472);
nand_5 g04096(n8665, n5283, new_n4473);
and_5  g04097(new_n4473, new_n4472, new_n4474);
nand_5 g04098(n1067, n137, new_n4475);
not_8  g04099(new_n4475, new_n4476);
xor_4  g04100(new_n4473, new_n4472, new_n4477);
not_8  g04101(new_n4477, new_n4478);
nor_5  g04102(new_n4478, new_n4476, new_n4479);
or_5   g04103(new_n4479, new_n4474, new_n4480);
not_8  g04104(new_n4480, new_n4481);
xor_4  g04105(new_n4481, new_n4471, new_n4482);
nand_5 g04106(n11922, n11478, new_n4483);
not_8  g04107(new_n4483, new_n4484);
nand_5 g04108(n5283, n1067, new_n4485);
nand_5 g04109(n11478, n8665, new_n4486);
and_5  g04110(new_n4486, new_n4485, new_n4487);
and_5  g04111(n5645, n137, new_n4488);
xor_4  g04112(new_n4486, new_n4485, new_n4489);
not_8  g04113(new_n4489, new_n4490);
nor_5  g04114(new_n4490, new_n4488, new_n4491);
or_5   g04115(new_n4491, new_n4487, new_n4492);
not_8  g04116(new_n4492, new_n4493);
and_5  g04117(new_n4493, new_n4484, new_n4494);
xor_4  g04118(new_n4478, new_n4476, new_n4495);
not_8  g04119(new_n4495, new_n4496);
xor_4  g04120(new_n4493, new_n4484, new_n4497);
and_5  g04121(new_n4497, new_n4496, new_n4498);
or_5   g04122(new_n4498, new_n4494, new_n4499_1);
not_8  g04123(new_n4499_1, new_n4500);
nand_5 g04124(n11478, n2551, new_n4501);
nand_5 g04125(n11922, n5283, new_n4502);
xor_4  g04126(new_n4502, new_n4501, new_n4503);
not_8  g04127(new_n4503, new_n4504);
xor_4  g04128(new_n4504, new_n4500, new_n4505);
xor_4  g04129(new_n4505, new_n4482, new_n4506);
nand_5 g04130(n4805, n2551, new_n4507);
nand_5 g04131(n11922, n4805, new_n4508);
nand_5 g04132(n5645, n5283, new_n4509);
nand_5 g04133(n8665, n4805, new_n4510);
nor_5  g04134(new_n4510, new_n4509, new_n4511);
nand_5 g04135(new_n4510, new_n4509, new_n4512);
not_8  g04136(new_n4512, new_n4513);
nand_5 g04137(n11478, n1067, new_n4514);
nor_5  g04138(new_n4514, new_n4513, new_n4515);
nor_5  g04139(new_n4515, new_n4511, new_n4516_1);
nor_5  g04140(new_n4516_1, new_n4508, new_n4517);
xor_4  g04141(new_n4516_1, new_n4508, new_n4518);
not_8  g04142(new_n4518, new_n4519);
xor_4  g04143(new_n4490, new_n4488, new_n4520);
nor_5  g04144(new_n4520, new_n4519, new_n4521);
or_5   g04145(new_n4521, new_n4517, new_n4522);
not_8  g04146(new_n4522, new_n4523);
and_5  g04147(new_n4523, new_n4507, new_n4524);
xor_4  g04148(new_n4497, new_n4496, new_n4525);
not_8  g04149(new_n4525, new_n4526);
xor_4  g04150(new_n4523, new_n4507, new_n4527);
and_5  g04151(new_n4527, new_n4526, new_n4528);
or_5   g04152(new_n4528, new_n4524, new_n4529);
not_8  g04153(new_n4529, new_n4530);
xor_4  g04154(new_n4530, new_n4506, new_n4531);
and_5  g04155(new_n4531, new_n4465, new_n4532);
xor_4  g04156(new_n4520, new_n4519, new_n4533);
xnor_4 g04157(new_n4510, new_n4509, new_n4534);
not_8  g04158(new_n4534, new_n4535);
and_5  g04159(n4805, n1067, new_n4536);
and_5  g04160(n11478, n5645, new_n4537);
nand_5 g04161(new_n4537, new_n4536, new_n4538);
or_5   g04162(new_n4538, new_n4535, new_n4539);
not_8  g04163(new_n4539, new_n4540);
nand_5 g04164(new_n4540, new_n4533, new_n4541);
xor_4  g04165(new_n4527, new_n4526, new_n4542);
or_5   g04166(new_n4542, new_n4541, new_n4543);
not_8  g04167(new_n4543, new_n4544);
xor_4  g04168(new_n4531, new_n4465, new_n4545);
and_5  g04169(new_n4545, new_n4544, new_n4546);
or_5   g04170(new_n4546, new_n4532, new_n4547);
not_8  g04171(new_n4547, new_n4548);
and_5  g04172(new_n4530, new_n4506, new_n4549);
nand_5 g04173(n12826, n11478, new_n4550);
nand_5 g04174(n5283, n2551, new_n4551);
and_5  g04175(n4805, n4094, new_n4552);
xor_4  g04176(new_n4552, new_n4551, new_n4553_1);
not_8  g04177(new_n4553_1, new_n4554);
xor_4  g04178(new_n4554, new_n4550, new_n4555);
nor_5  g04179(new_n4470, new_n4466, new_n4556);
and_5  g04180(new_n4481, new_n4471, new_n4557);
or_5   g04181(new_n4557, new_n4556, new_n4558);
not_8  g04182(new_n4558, new_n4559);
xor_4  g04183(new_n4559, new_n4555, new_n4560);
or_5   g04184(new_n4468, new_n4467, new_n4561);
not_8  g04185(new_n4561, new_n4562);
nand_5 g04186(n11922, n137, new_n4563);
not_8  g04187(new_n4563, new_n4564);
xor_4  g04188(new_n4564, new_n4562, new_n4565);
nand_5 g04189(n6797, n1067, new_n4566);
nand_5 g04190(n8665, n6294, new_n4567);
nand_5 g04191(n5645, n3146, new_n4568);
xor_4  g04192(new_n4568, new_n4567, new_n4569);
not_8  g04193(new_n4569, new_n4570);
xor_4  g04194(new_n4570, new_n4566, new_n4571);
xor_4  g04195(new_n4571, new_n4565, new_n4572);
xor_4  g04196(new_n4572, new_n4560, new_n4573);
not_8  g04197(new_n4573, new_n4574);
or_5   g04198(new_n4504, new_n4500, new_n4575);
or_5   g04199(new_n4502, new_n4501, new_n4576);
and_5  g04200(new_n4505, new_n4482, new_n4577);
xor_4  g04201(new_n4577, new_n4576, new_n4578);
and_5  g04202(new_n4578, new_n4575, new_n4579);
xor_4  g04203(new_n4579, new_n4574, new_n4580);
not_8  g04204(new_n4580, new_n4581);
xnor_4 g04205(new_n4581, new_n4549, new_n4582);
xnor_4 g04206(new_n4582, new_n4548, new_n4583);
nand_5 g04207(n3992, n2749, new_n4584);
not_8  g04208(new_n4584, new_n4585);
nand_5 g04209(n11876, n6358, new_n4586);
nand_5 g04210(n3992, n3754, new_n4587);
and_5  g04211(new_n4587, new_n4586, new_n4588);
and_5  g04212(n10898, n8384, new_n4589);
xor_4  g04213(new_n4587, new_n4586, new_n4590);
not_8  g04214(new_n4590, new_n4591);
nor_5  g04215(new_n4591, new_n4589, new_n4592);
or_5   g04216(new_n4592, new_n4588, new_n4593);
not_8  g04217(new_n4593, new_n4594);
nand_5 g04218(new_n4594, new_n4585, new_n4595);
xor_4  g04219(new_n4594, new_n4584, new_n4596);
nand_5 g04220(n10898, n6358, new_n4597);
not_8  g04221(new_n4597, new_n4598);
nand_5 g04222(n11876, n5198, new_n4599);
nand_5 g04223(n8384, n3754, new_n4600);
xor_4  g04224(new_n4600, new_n4599, new_n4601);
not_8  g04225(new_n4601, new_n4602);
xor_4  g04226(new_n4602, new_n4598, new_n4603);
nor_5  g04227(new_n4603, new_n4596, new_n4604);
not_8  g04228(new_n4604, new_n4605);
and_5  g04229(new_n4605, new_n4595, new_n4606);
nand_5 g04230(n8384, n2749, new_n4607);
nand_5 g04231(n3992, n159, new_n4608);
xor_4  g04232(new_n4608, new_n4607, new_n4609);
xor_4  g04233(new_n4609, new_n4606, new_n4610);
not_8  g04234(new_n4610, new_n4611);
nand_5 g04235(n6358, n3754, new_n4612);
not_8  g04236(new_n4612, new_n4613);
nand_5 g04237(n10898, n5198, new_n4614);
nand_5 g04238(n11876, n1471, new_n4615);
xor_4  g04239(new_n4615, new_n4614, new_n4616);
xor_4  g04240(new_n4616, new_n4613, new_n4617);
and_5  g04241(new_n4600, new_n4599, new_n4618);
nor_5  g04242(new_n4602, new_n4598, new_n4619);
nor_5  g04243(new_n4619, new_n4618, new_n4620);
xor_4  g04244(new_n4620, new_n4617, new_n4621);
xor_4  g04245(new_n4621, new_n4611, new_n4622);
nand_5 g04246(n7236, n159, new_n4623);
not_8  g04247(new_n4623, new_n4624);
nand_5 g04248(n7236, n2749, new_n4625);
not_8  g04249(new_n4625, new_n4626);
and_5  g04250(n11876, n8384, new_n4627);
and_5  g04251(n7236, n3754, new_n4628);
nor_5  g04252(new_n4628, new_n4627, new_n4629);
nand_5 g04253(n11876, n7236, new_n4630);
nor_5  g04254(new_n4630, new_n4600, new_n4631);
and_5  g04255(n10898, n3992, new_n4632);
nor_5  g04256(new_n4632, new_n4631, new_n4633);
or_5   g04257(new_n4633, new_n4629, new_n4634_1);
not_8  g04258(new_n4634_1, new_n4635);
and_5  g04259(new_n4635, new_n4626, new_n4636);
nor_5  g04260(new_n4635, new_n4626, new_n4637);
or_5   g04261(new_n4637, new_n4636, new_n4638);
xor_4  g04262(new_n4591, new_n4589, new_n4639);
nor_5  g04263(new_n4639, new_n4638, new_n4640);
or_5   g04264(new_n4640, new_n4636, new_n4641);
nor_5  g04265(new_n4641, new_n4624, new_n4642);
xor_4  g04266(new_n4603, new_n4596, new_n4643);
xor_4  g04267(new_n4641, new_n4624, new_n4644);
not_8  g04268(new_n4644, new_n4645);
nor_5  g04269(new_n4645, new_n4643, new_n4646);
nor_5  g04270(new_n4646, new_n4642, new_n4647);
nand_5 g04271(new_n4647, new_n4622, new_n4648);
or_5   g04272(new_n4615, new_n4614, new_n4649);
not_8  g04273(new_n4649, new_n4650);
nand_5 g04274(n6358, n2749, new_n4651);
not_8  g04275(new_n4651, new_n4652);
xor_4  g04276(new_n4652, new_n4650, new_n4653);
nand_5 g04277(n10898, n1471, new_n4654);
nand_5 g04278(n5198, n3754, new_n4655);
nand_5 g04279(n11876, n7646, new_n4656);
xor_4  g04280(new_n4656, new_n4655, new_n4657);
not_8  g04281(new_n4657, new_n4658);
xor_4  g04282(new_n4658, new_n4654, new_n4659);
xor_4  g04283(new_n4659, new_n4653, new_n4660);
nor_5  g04284(new_n4616, new_n4613, new_n4661);
not_8  g04285(new_n4617, new_n4662);
nor_5  g04286(new_n4620, new_n4662, new_n4663);
or_5   g04287(new_n4663, new_n4661, new_n4664);
not_8  g04288(new_n4664, new_n4665);
nand_5 g04289(n3992, n1510, new_n4666);
not_8  g04290(new_n4666, new_n4667);
nand_5 g04291(n8384, n159, new_n4668);
nand_5 g04292(n12247, n7236, new_n4669);
xor_4  g04293(new_n4669, new_n4668, new_n4670);
not_8  g04294(new_n4670, new_n4671);
xor_4  g04295(new_n4671, new_n4667, new_n4672);
xor_4  g04296(new_n4672, new_n4665, new_n4673);
xor_4  g04297(new_n4673, new_n4660, new_n4674);
not_8  g04298(new_n4609, new_n4675);
nor_5  g04299(new_n4675, new_n4606, new_n4676);
or_5   g04300(new_n4608, new_n4607, new_n4677);
not_8  g04301(new_n4677, new_n4678);
and_5  g04302(new_n4621, new_n4611, new_n4679);
xor_4  g04303(new_n4679, new_n4678, new_n4680);
nor_5  g04304(new_n4680, new_n4676, new_n4681);
xor_4  g04305(new_n4681, new_n4674, new_n4682);
not_8  g04306(new_n4682, new_n4683);
nor_5  g04307(new_n4683, new_n4648, new_n4684);
and_5  g04308(new_n4683, new_n4648, new_n4685);
or_5   g04309(new_n4685, new_n4684, new_n4686_1);
nand_5 g04310(n7236, n1510, new_n4687);
xnor_4 g04311(new_n4647, new_n4622, new_n4688);
nor_5  g04312(new_n4688, new_n4687, new_n4689_1);
xor_4  g04313(new_n4639, new_n4638, new_n4690);
nor_5  g04314(new_n4631, new_n4629, new_n4691);
nand_5 g04315(n11876, n3992, new_n4692);
and_5  g04316(n10898, n7236, new_n4693);
not_8  g04317(new_n4693, new_n4694);
or_5   g04318(new_n4694, new_n4692, new_n4695);
or_5   g04319(new_n4695, new_n4691, new_n4696);
not_8  g04320(new_n4696, new_n4697);
nand_5 g04321(new_n4697, new_n4690, new_n4698);
xor_4  g04322(new_n4645, new_n4643, new_n4699);
or_5   g04323(new_n4699, new_n4698, new_n4700);
xor_4  g04324(new_n4688, new_n4687, new_n4701);
not_8  g04325(new_n4701, new_n4702);
nor_5  g04326(new_n4702, new_n4700, new_n4703);
nor_5  g04327(new_n4703, new_n4689_1, new_n4704);
xor_4  g04328(new_n4704, new_n4686_1, new_n4705);
xor_4  g04329(new_n4705, new_n4583, new_n4706);
not_8  g04330(new_n4706, new_n4707);
xor_4  g04331(new_n4545, new_n4544, new_n4708);
xor_4  g04332(new_n4702, new_n4700, new_n4709);
nor_5  g04333(new_n4709, new_n4708, new_n4710);
xor_4  g04334(new_n4709, new_n4708, new_n4711);
not_8  g04335(new_n4698, new_n4712);
xor_4  g04336(new_n4699, new_n4712, new_n4713);
not_8  g04337(new_n4713, new_n4714);
xor_4  g04338(new_n4540, new_n4533, new_n4715);
xor_4  g04339(new_n4697, new_n4690, new_n4716);
nor_5  g04340(new_n4716, new_n4715, new_n4717);
xor_4  g04341(new_n4693, new_n4692, new_n4718);
not_8  g04342(new_n4718, new_n4719);
xor_4  g04343(new_n4537, new_n4536, new_n4720);
nor_5  g04344(new_n4720, new_n4719, new_n4721);
nand_5 g04345(n5645, n4805, new_n4722_1);
nor_5  g04346(new_n4722_1, new_n4630, new_n4723);
not_8  g04347(new_n4723, new_n4724);
xor_4  g04348(new_n4720, new_n4719, new_n4725);
and_5  g04349(new_n4725, new_n4724, new_n4726);
or_5   g04350(new_n4726, new_n4721, new_n4727);
not_8  g04351(new_n4727, new_n4728);
and_5  g04352(n11478, n1067, new_n4729);
and_5  g04353(new_n4722_1, new_n4729, new_n4730);
not_8  g04354(new_n4730, new_n4731);
nor_5  g04355(new_n4731, new_n4512, new_n4732);
and_5  g04356(new_n4731, new_n4535, new_n4733_1);
nor_5  g04357(new_n4733_1, new_n4732, new_n4734);
not_8  g04358(new_n4734, new_n4735);
nor_5  g04359(new_n4735, new_n4728, new_n4736);
xor_4  g04360(new_n4735, new_n4728, new_n4737);
nand_5 g04361(new_n4632, new_n4630, new_n4738);
not_8  g04362(new_n4738, new_n4739);
nor_5  g04363(new_n4739, new_n4691, new_n4740);
nor_5  g04364(new_n4738, new_n4629, new_n4741);
or_5   g04365(new_n4741, new_n4740, new_n4742);
and_5  g04366(new_n4742, new_n4737, new_n4743);
or_5   g04367(new_n4743, new_n4736, new_n4744);
not_8  g04368(new_n4744, new_n4745);
xor_4  g04369(new_n4716, new_n4715, new_n4746);
not_8  g04370(new_n4746, new_n4747);
nor_5  g04371(new_n4747, new_n4745, new_n4748);
nor_5  g04372(new_n4748, new_n4717, new_n4749);
nor_5  g04373(new_n4749, new_n4714, new_n4750);
xor_4  g04374(new_n4542, new_n4541, new_n4751);
xor_4  g04375(new_n4749, new_n4714, new_n4752);
not_8  g04376(new_n4752, new_n4753);
nor_5  g04377(new_n4753, new_n4751, new_n4754);
or_5   g04378(new_n4754, new_n4750, new_n4755);
and_5  g04379(new_n4755, new_n4711, new_n4756);
nor_5  g04380(new_n4756, new_n4710, new_n4757_1);
xor_4  g04381(new_n4757_1, new_n4707, new_n4758);
xor_4  g04382(new_n4758, new_n4463, new_n4759);
xor_4  g04383(new_n4460, new_n4459, new_n4760);
xor_4  g04384(new_n4755, new_n4711, new_n4761);
not_8  g04385(new_n4761, new_n4762);
nor_5  g04386(new_n4762, new_n4760, new_n4763);
xor_4  g04387(new_n4457, new_n4456, new_n4764);
not_8  g04388(new_n4764, new_n4765);
xor_4  g04389(new_n4454, new_n4446, new_n4766);
not_8  g04390(new_n4766, new_n4767);
xor_4  g04391(new_n4747, new_n4745, new_n4768);
nor_5  g04392(new_n4768, new_n4767, new_n4769);
xor_4  g04393(new_n4768, new_n4766, new_n4770);
xor_4  g04394(new_n4742, new_n4737, new_n4771);
nor_5  g04395(new_n4449, new_n4390, new_n4772);
or_5   g04396(new_n4772, new_n4451, new_n4773);
nor_5  g04397(new_n4773, new_n4771, new_n4774);
xor_4  g04398(new_n4773, new_n4771, new_n4775);
not_8  g04399(new_n4775, new_n4776);
xor_4  g04400(new_n4725, new_n4724, new_n4777);
not_8  g04401(new_n4777, new_n4778);
nand_5 g04402(n9400, n6703, new_n4779);
and_5  g04403(n9640, n6877, new_n4780);
xor_4  g04404(new_n4780, new_n4779, new_n4781);
not_8  g04405(new_n4781, new_n4782);
and_5  g04406(new_n4782, new_n4778, new_n4783);
xor_4  g04407(new_n4722_1, new_n4630, new_n4784);
not_8  g04408(new_n4784, new_n4785);
or_5   g04409(new_n4785, new_n4447, new_n4786);
xor_4  g04410(new_n4781, new_n4778, new_n4787);
nor_5  g04411(new_n4787, new_n4786, new_n4788);
nor_5  g04412(new_n4788, new_n4783, new_n4789);
nor_5  g04413(new_n4789, new_n4776, new_n4790);
nor_5  g04414(new_n4790, new_n4774, new_n4791);
nor_5  g04415(new_n4791, new_n4770, new_n4792);
or_5   g04416(new_n4792, new_n4769, new_n4793);
not_8  g04417(new_n4793, new_n4794);
and_5  g04418(new_n4794, new_n4765, new_n4795);
xor_4  g04419(new_n4753, new_n4751, new_n4796);
not_8  g04420(new_n4796, new_n4797);
nor_5  g04421(new_n4794, new_n4765, new_n4798);
or_5   g04422(new_n4798, new_n4795, new_n4799);
nor_5  g04423(new_n4799, new_n4797, new_n4800);
or_5   g04424(new_n4800, new_n4795, new_n4801);
xor_4  g04425(new_n4762, new_n4760, new_n4802);
and_5  g04426(new_n4802, new_n4801, new_n4803);
nor_5  g04427(new_n4803, new_n4763, new_n4804);
xor_4  g04428(new_n4804, new_n4759, new_n4805_1);
nor_5  g04429(new_n4805_1, new_n4340, new_n4806);
xor_4  g04430(new_n4805_1, new_n4339, new_n4807);
xor_4  g04431(new_n4336, new_n4334, new_n4808);
not_8  g04432(new_n4808, new_n4809);
not_8  g04433(new_n4801, new_n4810);
xnor_4 g04434(new_n4802, new_n4810, new_n4811);
or_5   g04435(new_n4811, new_n4809, new_n4812);
xor_4  g04436(new_n4333_1, new_n4332, new_n4813);
xor_4  g04437(new_n4799, new_n4796, new_n4814);
nor_5  g04438(new_n4814, new_n4813, new_n4815);
not_8  g04439(new_n4813, new_n4816);
xor_4  g04440(new_n4814, new_n4816, new_n4817_1);
not_8  g04441(new_n4817_1, new_n4818);
xor_4  g04442(new_n4331, new_n4326_1, new_n4819);
xor_4  g04443(new_n4791, new_n4770, new_n4820);
nor_5  g04444(new_n4820, new_n4819, new_n4821);
or_5   g04445(new_n4788, new_n4783, new_n4822);
xor_4  g04446(new_n4822, new_n4776, new_n4823);
not_8  g04447(new_n4273, new_n4824);
nand_5 g04448(n7862, n1798, new_n4825);
and_5  g04449(new_n4825, new_n4824, new_n4826_1);
nor_5  g04450(new_n4826_1, new_n4327, new_n4827);
nand_5 g04451(new_n4270, new_n4269, new_n4828_1);
and_5  g04452(new_n4826_1, new_n4828_1, new_n4829);
or_5   g04453(new_n4829, new_n4827, new_n4830);
and_5  g04454(new_n4830, new_n4823, new_n4831);
nor_5  g04455(new_n4829, new_n4827, new_n4832);
xor_4  g04456(new_n4832, new_n4823, new_n4833);
not_8  g04457(new_n4833, new_n4834);
not_8  g04458(new_n4825, new_n4835);
xor_4  g04459(new_n4785, new_n4447, new_n4836);
nand_5 g04460(new_n4836, new_n4835, new_n4837);
xnor_4 g04461(new_n4329, new_n4328, new_n4838);
and_5  g04462(new_n4838, new_n4837, new_n4839);
xor_4  g04463(new_n4787, new_n4786, new_n4840);
xor_4  g04464(new_n4838, new_n4837, new_n4841);
not_8  g04465(new_n4841, new_n4842);
nor_5  g04466(new_n4842, new_n4840, new_n4843);
or_5   g04467(new_n4843, new_n4839, new_n4844);
and_5  g04468(new_n4844, new_n4834, new_n4845);
or_5   g04469(new_n4845, new_n4831, new_n4846);
not_8  g04470(new_n4819, new_n4847);
xor_4  g04471(new_n4820, new_n4847, new_n4848);
not_8  g04472(new_n4848, new_n4849);
and_5  g04473(new_n4849, new_n4846, new_n4850);
or_5   g04474(new_n4850, new_n4821, new_n4851);
and_5  g04475(new_n4851, new_n4818, new_n4852);
or_5   g04476(new_n4852, new_n4815, new_n4853);
not_8  g04477(new_n4853, new_n4854);
xor_4  g04478(new_n4811, new_n4808, new_n4855);
not_8  g04479(new_n4855, new_n4856);
nand_5 g04480(new_n4856, new_n4854, new_n4857);
and_5  g04481(new_n4857, new_n4812, new_n4858);
nor_5  g04482(new_n4858, new_n4807, new_n4859);
or_5   g04483(new_n4859, new_n4806, new_n4860);
and_5  g04484(new_n4440, new_n4410, new_n4861);
nor_5  g04485(new_n4462, new_n4441, new_n4862);
nor_5  g04486(new_n4862, new_n4861, new_n4863);
and_5  g04487(n7862, n753, new_n4864);
nand_5 g04488(new_n4559, new_n4555, new_n4865);
not_8  g04489(new_n4572, new_n4866);
nand_5 g04490(new_n4866, new_n4560, new_n4867);
and_5  g04491(new_n4867, new_n4865, new_n4868);
xor_4  g04492(new_n4868, new_n4864, new_n4869);
and_5  g04493(new_n4564, new_n4562, new_n4870);
and_5  g04494(new_n4571, new_n4565, new_n4871);
or_5   g04495(new_n4871, new_n4870, new_n4872);
and_5  g04496(n3146, n1067, new_n4873);
and_5  g04497(n2551, n137, new_n4874);
xor_4  g04498(new_n4874, new_n4873, new_n4875);
and_5  g04499(n12826, n5283, new_n4876);
and_5  g04500(n8665, n6797, new_n4877);
xor_4  g04501(new_n4877, new_n4876, new_n4878);
xor_4  g04502(new_n4878, new_n4875, new_n4879);
xor_4  g04503(new_n4879, new_n4872, new_n4880);
and_5  g04504(new_n4652, new_n4650, new_n4881);
and_5  g04505(new_n4659, new_n4653, new_n4882);
or_5   g04506(new_n4882, new_n4881, new_n4883);
and_5  g04507(new_n4669, new_n4668, new_n4884);
nor_5  g04508(new_n4671, new_n4667, new_n4885);
nor_5  g04509(new_n4885, new_n4884, new_n4886);
nand_5 g04510(n8384, n1510, new_n4887);
and_5  g04511(n5198, n2749, new_n4888);
xor_4  g04512(new_n4888, new_n4887, new_n4889);
xor_4  g04513(new_n4889, new_n4886, new_n4890);
xor_4  g04514(new_n4890, new_n4883, new_n4891);
xor_4  g04515(new_n4891, new_n4880, new_n4892);
xor_4  g04516(new_n4892, new_n4869, new_n4893);
xor_4  g04517(new_n4893, new_n4863, new_n4894);
nor_5  g04518(new_n4313, new_n4312_1, new_n4895);
nor_5  g04519(new_n4315, new_n4310, new_n4896);
nor_5  g04520(new_n4896, new_n4895, new_n4897);
not_8  g04521(new_n4576, new_n4898);
and_5  g04522(new_n4577, new_n4898, new_n4899);
nor_5  g04523(new_n4579, new_n4574, new_n4900);
nor_5  g04524(new_n4900, new_n4899, new_n4901);
xor_4  g04525(new_n4901, new_n4897, new_n4902);
nand_5 g04526(n12511, n7236, new_n4903_1);
and_5  g04527(n6826, n1798, new_n4904);
xor_4  g04528(new_n4904, new_n4903_1, new_n4905);
and_5  g04529(new_n4568, new_n4567, new_n4906);
not_8  g04530(new_n4566, new_n4907);
nor_5  g04531(new_n4570, new_n4907, new_n4908);
or_5   g04532(new_n4908, new_n4906, new_n4909);
and_5  g04533(new_n4656, new_n4655, new_n4910);
not_8  g04534(new_n4654, new_n4911);
nor_5  g04535(new_n4658, new_n4911, new_n4912);
nor_5  g04536(new_n4912, new_n4910, new_n4913);
xor_4  g04537(new_n4913, new_n4909, new_n4914);
xor_4  g04538(new_n4914, new_n4905, new_n4915);
and_5  g04539(n6358, n159, new_n4916);
and_5  g04540(new_n4554, new_n4550, new_n4917);
or_5   g04541(new_n4917, new_n4551, new_n4918);
not_8  g04542(new_n4918, new_n4919);
and_5  g04543(n11478, n4094, new_n4920);
and_5  g04544(new_n4920, new_n4919, new_n4921_1);
and_5  g04545(new_n4920, new_n4464, new_n4922);
nor_5  g04546(new_n4922, new_n4919, new_n4923);
nor_5  g04547(new_n4923, new_n4921_1, new_n4924);
xor_4  g04548(new_n4924, new_n4916, new_n4925);
xor_4  g04549(new_n4925, new_n4915, new_n4926);
xor_4  g04550(new_n4926, new_n4902, new_n4927);
xor_4  g04551(new_n4927, new_n4894, new_n4928_1);
and_5  g04552(new_n4679, new_n4678, new_n4929);
nor_5  g04553(new_n4681, new_n4674, new_n4930);
nor_5  g04554(new_n4930, new_n4929, new_n4931);
nand_5 g04555(n5645, n4938, new_n4932);
and_5  g04556(n10898, n7646, new_n4933);
xor_4  g04557(new_n4933, new_n4932, new_n4934);
xor_4  g04558(new_n4934, new_n4931, new_n4935);
xor_4  g04559(new_n4935, new_n4928_1, new_n4936);
nor_5  g04560(new_n4705, new_n4583, new_n4937);
nor_5  g04561(new_n4757_1, new_n4707, new_n4938_1);
nor_5  g04562(new_n4938_1, new_n4937, new_n4939);
and_5  g04563(n11922, n6294, new_n4940);
not_8  g04564(new_n4549, new_n4941);
nor_5  g04565(new_n4581, new_n4941, new_n4942);
and_5  g04566(new_n4582, new_n4547, new_n4943);
nor_5  g04567(new_n4943, new_n4942, new_n4944);
xor_4  g04568(new_n4944, new_n4940, new_n4945);
nor_5  g04569(new_n4338, new_n4320, new_n4946);
or_5   g04570(new_n4946, new_n4318, new_n4947);
not_8  g04571(new_n4435, new_n4948);
nand_5 g04572(new_n4437, new_n4948, new_n4949);
not_8  g04573(new_n4949, new_n4950);
nor_5  g04574(new_n4439, new_n4433, new_n4951);
nor_5  g04575(new_n4951, new_n4950, new_n4952);
or_5   g04576(new_n4419, new_n4413, new_n4953);
not_8  g04577(new_n4431, new_n4954);
nand_5 g04578(new_n4954, new_n4420, new_n4955);
nand_5 g04579(new_n4955, new_n4953, new_n4956);
nor_5  g04580(new_n4428, new_n4427, new_n4957);
nand_5 g04581(n9640, n4203, new_n4958);
and_5  g04582(new_n4428, new_n4427, new_n4959);
nor_5  g04583(new_n4959, new_n4958, new_n4960);
nor_5  g04584(new_n4960, new_n4957, new_n4961);
nand_5 g04585(n4203, n3022, new_n4962);
and_5  g04586(n11023, n4187, new_n4963);
xor_4  g04587(new_n4963, new_n4962, new_n4964);
xor_4  g04588(new_n4964, new_n4961, new_n4965);
nand_5 g04589(n7456, n5240, new_n4966);
and_5  g04590(n12753, n9640, new_n4967);
xor_4  g04591(new_n4967, new_n4966, new_n4968);
nand_5 g04592(n9583, n1333, new_n4969);
and_5  g04593(n12591, n11821, new_n4970_1);
xor_4  g04594(new_n4970_1, new_n4969, new_n4971_1);
xor_4  g04595(new_n4971_1, new_n4968, new_n4972);
xor_4  g04596(new_n4972, new_n4965, new_n4973);
xor_4  g04597(new_n4973, new_n4956, new_n4974);
nor_5  g04598(new_n4297, new_n4289, new_n4975);
nor_5  g04599(new_n4224, new_n4223, new_n4976);
xor_4  g04600(new_n4301, new_n4976, new_n4977);
xor_4  g04601(new_n4307, new_n4977, new_n4978);
and_5  g04602(new_n4978, new_n4298, new_n4979);
or_5   g04603(new_n4979, new_n4975, new_n4980);
nand_5 g04604(n9080, n3932, new_n4981);
nand_5 g04605(n10174, n6703, new_n4982);
and_5  g04606(n6877, n2278, new_n4983);
xor_4  g04607(new_n4983, new_n4982, new_n4984);
xor_4  g04608(new_n4984, new_n4981, new_n4985);
xor_4  g04609(new_n4985, new_n4980, new_n4986);
xor_4  g04610(new_n4986, new_n4974, new_n4987);
xor_4  g04611(new_n4987, new_n4952, new_n4988);
xor_4  g04612(new_n4988, new_n4947, new_n4989);
xor_4  g04613(new_n4989, new_n4945, new_n4990);
xor_4  g04614(new_n4990, new_n4939, new_n4991);
xor_4  g04615(new_n4991, new_n4936, new_n4992);
xor_4  g04616(new_n4992, new_n4860, new_n4993);
not_8  g04617(new_n4672, new_n4994);
nor_5  g04618(new_n4994, new_n4665, new_n4995);
nor_5  g04619(new_n4673, new_n4660, new_n4996);
or_5   g04620(new_n4996, new_n4995, new_n4997);
nor_5  g04621(new_n4300_1, new_n4299, new_n4998);
nor_5  g04622(new_n4307, new_n4302, new_n4999);
or_5   g04623(new_n4999, new_n4998, new_n5000);
nor_5  g04624(new_n4416, new_n4415, new_n5001);
and_5  g04625(new_n4416, new_n4415, new_n5002);
nor_5  g04626(new_n5002, new_n4414, new_n5003);
nor_5  g04627(new_n5003, new_n5001, new_n5004);
xor_4  g04628(new_n5004, new_n5000, new_n5005);
and_5  g04629(new_n4293, new_n4292, new_n5006);
nor_5  g04630(new_n4295, new_n4291, new_n5007);
or_5   g04631(new_n5007, new_n5006, new_n5008);
nor_5  g04632(new_n4305, new_n4304, new_n5009);
and_5  g04633(new_n4305, new_n4304, new_n5010);
nor_5  g04634(new_n5010, new_n4303, new_n5011);
or_5   g04635(new_n5011, new_n5009, new_n5012);
nand_5 g04636(n10278, n2464, new_n5013);
and_5  g04637(n11757, n11662, new_n5014);
xor_4  g04638(new_n5014, new_n5013, new_n5015);
nand_5 g04639(n10327, n3172, new_n5016);
and_5  g04640(n11423, n9400, new_n5017);
xor_4  g04641(new_n5017, new_n5016, new_n5018);
xor_4  g04642(new_n5018, new_n5015, new_n5019);
xor_4  g04643(new_n5019, new_n5012, new_n5020);
xor_4  g04644(new_n5020, new_n5008, new_n5021);
xor_4  g04645(new_n5021, new_n5005, new_n5022);
xor_4  g04646(new_n5022, new_n4997, new_n5023);
and_5  g04647(n3754, n1471, new_n5024);
and_5  g04648(n11311, n10451, new_n5025);
xor_4  g04649(new_n5025, new_n5024, new_n5026);
and_5  g04650(new_n4424, new_n4422, new_n5027);
and_5  g04651(new_n4430, new_n4425, new_n5028);
nor_5  g04652(new_n5028, new_n5027, new_n5029);
and_5  g04653(n11876, n4722, new_n5030_1);
nand_5 g04654(n10685, n4805, new_n5031);
and_5  g04655(n12247, n3992, new_n5032);
xor_4  g04656(new_n5032, new_n5031, new_n5033);
xor_4  g04657(new_n5033, new_n5030_1, new_n5034_1);
xor_4  g04658(new_n5034_1, new_n5029, new_n5035);
xor_4  g04659(new_n5035, new_n5026, new_n5036);
xor_4  g04660(new_n5036, new_n5023, new_n5037);
nor_5  g04661(new_n4704, new_n4686_1, new_n5038);
nor_5  g04662(new_n5038, new_n4684, new_n5039);
not_8  g04663(new_n4758, new_n5040);
nor_5  g04664(new_n5040, new_n4463, new_n5041);
nor_5  g04665(new_n4804, new_n4759, new_n5042);
nor_5  g04666(new_n5042, new_n5041, new_n5043);
xor_4  g04667(new_n5043, new_n5039, new_n5044);
xor_4  g04668(new_n5044, new_n5037, new_n5045);
xor_4  g04669(new_n5045, new_n4993, n1269);
nand_5 g04670(n10223, n4312, new_n5047);
not_8  g04671(new_n5047, new_n5048);
nand_5 g04672(n12705, n7265, new_n5049);
nand_5 g04673(n4312, n2879, new_n5050);
not_8  g04674(new_n5050, new_n5051);
xor_4  g04675(new_n5049, new_n1034, new_n5052);
not_8  g04676(new_n5052, new_n5053);
nor_5  g04677(new_n5053, new_n5051, new_n5054);
nor_5  g04678(new_n5054, new_n5049, new_n5055);
nor_5  g04679(new_n5055, new_n5048, new_n5056);
nor_5  g04680(new_n5055, new_n1045, new_n5057);
nor_5  g04681(new_n5057, new_n5047, new_n5058);
or_5   g04682(new_n5058, new_n5056, new_n5059);
not_8  g04683(new_n5059, new_n5060);
nand_5 g04684(n12025, n7265, new_n5061);
nand_5 g04685(n12705, n2879, new_n5062);
xor_4  g04686(new_n5062, new_n5061, new_n5063);
nor_5  g04687(new_n5063, new_n5060, new_n5064);
and_5  g04688(new_n5063, new_n5060, new_n5065);
or_5   g04689(new_n5065, new_n5064, new_n5066);
nand_5 g04690(n9195, n5964, new_n5067);
nand_5 g04691(n4634, n1097, new_n5068);
xor_4  g04692(new_n5068, new_n5067, new_n5069_1);
not_8  g04693(new_n5069_1, new_n5070);
xor_4  g04694(new_n5070, new_n5066, new_n5071);
nand_5 g04695(n5964, n4634, new_n5072);
not_8  g04696(new_n5072, new_n5073);
and_5  g04697(new_n1047, new_n1046, new_n5074);
nor_5  g04698(new_n1047, new_n1046, new_n5075);
nor_5  g04699(new_n5075, new_n1045, new_n5076);
or_5   g04700(new_n5076, new_n5074, new_n5077);
not_8  g04701(new_n5077, new_n5078);
and_5  g04702(new_n5078, new_n5073, new_n5079);
xor_4  g04703(new_n5053, new_n5051, new_n5080);
nor_5  g04704(new_n5078, new_n5073, new_n5081);
or_5   g04705(new_n5081, new_n5079, new_n5082);
nor_5  g04706(new_n5082, new_n5080, new_n5083);
or_5   g04707(new_n5083, new_n5079, new_n5084);
xor_4  g04708(new_n5084, new_n5071, new_n5085);
nand_5 g04709(n9195, n5305, new_n5086);
nor_5  g04710(new_n1050, new_n1043, new_n5087);
or_5   g04711(new_n5087, new_n1041, new_n5088);
not_8  g04712(new_n5088, new_n5089);
and_5  g04713(new_n5089, new_n5086, new_n5090);
xor_4  g04714(new_n5082, new_n5080, new_n5091);
not_8  g04715(new_n5091, new_n5092);
xor_4  g04716(new_n5089, new_n5086, new_n5093);
and_5  g04717(new_n5093, new_n5092, new_n5094_1);
or_5   g04718(new_n5094_1, new_n5090, new_n5095);
not_8  g04719(new_n5095, new_n5096);
nand_5 g04720(new_n5096, new_n5085, new_n5097);
or_5   g04721(new_n5065, new_n5058, new_n5098);
nand_5 g04722(n5964, n2253, new_n5099);
not_8  g04723(new_n5099, new_n5100);
nand_5 g04724(n9195, n1097, new_n5101);
nand_5 g04725(n5305, n3865, new_n5102);
xor_4  g04726(new_n5102, new_n5101, new_n5103);
not_8  g04727(new_n5103, new_n5104);
xor_4  g04728(new_n5104, new_n5100, new_n5105_1);
not_8  g04729(new_n5105_1, new_n5106);
xor_4  g04730(new_n5106, new_n5098, new_n5107);
or_5   g04731(new_n5062, new_n5061, new_n5108);
not_8  g04732(new_n5108, new_n5109);
nand_5 g04733(n4634, n4312, new_n5110);
not_8  g04734(new_n5110, new_n5111);
xor_4  g04735(new_n5111, new_n5109, new_n5112);
nand_5 g04736(n12025, n2879, new_n5113);
nand_5 g04737(n11257, n7265, new_n5114);
nand_5 g04738(n12705, n10223, new_n5115);
xor_4  g04739(new_n5115, new_n5114, new_n5116);
not_8  g04740(new_n5116, new_n5117);
xor_4  g04741(new_n5117, new_n5113, new_n5118);
xor_4  g04742(new_n5118, new_n5112, new_n5119);
xor_4  g04743(new_n5119, new_n5107, new_n5120);
not_8  g04744(new_n5120, new_n5121);
nor_5  g04745(new_n5070, new_n5066, new_n5122);
or_5   g04746(new_n5068, new_n5067, new_n5123);
nand_5 g04747(new_n5084, new_n5071, new_n5124);
xor_4  g04748(new_n5124, new_n5123, new_n5125);
nor_5  g04749(new_n5125, new_n5122, new_n5126);
xor_4  g04750(new_n5126, new_n5121, new_n5127);
not_8  g04751(new_n5127, new_n5128);
xor_4  g04752(new_n5128, new_n5097, new_n5129);
nand_5 g04753(n5305, n2253, new_n5130);
not_8  g04754(new_n5130, new_n5131);
xor_4  g04755(new_n5096, new_n5085, new_n5132_1);
and_5  g04756(new_n5132_1, new_n5131, new_n5133);
nand_5 g04757(new_n1059, new_n1051, new_n5134);
xor_4  g04758(new_n5093, new_n5092, new_n5135);
or_5   g04759(new_n5135, new_n5134, new_n5136);
not_8  g04760(new_n5136, new_n5137);
xor_4  g04761(new_n5132_1, new_n5131, new_n5138);
and_5  g04762(new_n5138, new_n5137, new_n5139);
or_5   g04763(new_n5139, new_n5133, new_n5140);
xor_4  g04764(new_n5140, new_n5129, new_n5141);
not_8  g04765(new_n5141, new_n5142);
xor_4  g04766(new_n5138, new_n5137, new_n5143);
nand_5 g04767(new_n1173, new_n1170, new_n5144);
not_8  g04768(new_n5144, new_n5145);
nand_5 g04769(n12145, n8759, new_n5146);
nor_5  g04770(new_n1161, new_n1155, new_n5147);
nor_5  g04771(new_n1169, new_n1162, new_n5148);
nor_5  g04772(new_n5148, new_n5147, new_n5149);
xor_4  g04773(new_n5149, new_n5146, new_n5150);
not_8  g04774(new_n5150, new_n5151);
nand_5 g04775(n6776, n2522, new_n5152);
not_8  g04776(new_n5152, new_n5153_1);
and_5  g04777(new_n1166, new_n1165, new_n5154);
nor_5  g04778(new_n1166, new_n1165, new_n5155);
nor_5  g04779(new_n5155, new_n1164, new_n5156);
or_5   g04780(new_n5156, new_n5154, new_n5157);
not_8  g04781(new_n5157, new_n5158);
and_5  g04782(new_n5158, new_n5153_1, new_n5159);
nor_5  g04783(new_n5158, new_n5153_1, new_n5160);
or_5   g04784(new_n5160, new_n5159, new_n5161);
nand_5 g04785(n7436, n2024, new_n5162);
not_8  g04786(new_n5162, new_n5163);
nand_5 g04787(n12299, n9189, new_n5164);
nand_5 g04788(n8276, n7946, new_n5165);
xor_4  g04789(new_n5165, new_n5164, new_n5166);
not_8  g04790(new_n5166, new_n5167);
xor_4  g04791(new_n5167, new_n5163, new_n5168);
xor_4  g04792(new_n5168, new_n5161, new_n5169);
not_8  g04793(new_n5169, new_n5170);
xor_4  g04794(new_n5170, new_n5151, new_n5171);
nand_5 g04795(new_n5171, new_n5145, new_n5172);
not_8  g04796(new_n5172, new_n5173);
nand_5 g04797(n12221, n8759, new_n5174);
nor_5  g04798(new_n5168, new_n5161, new_n5175);
or_5   g04799(new_n5175, new_n5159, new_n5176);
not_8  g04800(new_n5176, new_n5177);
nand_5 g04801(n12145, n6776, new_n5178);
nand_5 g04802(n12299, n2522, new_n5179);
xor_4  g04803(new_n5179, new_n5178, new_n5180);
not_8  g04804(new_n5180, new_n5181);
xor_4  g04805(new_n5181, new_n5177, new_n5182);
nand_5 g04806(n9189, n7436, new_n5183);
not_8  g04807(new_n5183, new_n5184);
nor_5  g04808(new_n5167, new_n5163, new_n5185);
nor_5  g04809(new_n5185, new_n5165, new_n5186);
nor_5  g04810(new_n5186, new_n5184, new_n5187);
nor_5  g04811(new_n5186, new_n1164, new_n5188);
nor_5  g04812(new_n5188, new_n5183, new_n5189);
or_5   g04813(new_n5189, new_n5187, new_n5190);
not_8  g04814(new_n5190, new_n5191_1);
nand_5 g04815(n8276, n2024, new_n5192);
nand_5 g04816(n9241, n7946, new_n5193);
xor_4  g04817(new_n5193, new_n5192, new_n5194);
nor_5  g04818(new_n5194, new_n5191_1, new_n5195);
and_5  g04819(new_n5194, new_n5191_1, new_n5196);
or_5   g04820(new_n5196, new_n5195, new_n5197);
xor_4  g04821(new_n5197, new_n5182, new_n5198_1);
nor_5  g04822(new_n5149, new_n5146, new_n5199);
nor_5  g04823(new_n5170, new_n5151, new_n5200);
nor_5  g04824(new_n5200, new_n5199, new_n5201);
xor_4  g04825(new_n5201, new_n5198_1, new_n5202);
not_8  g04826(new_n5202, new_n5203);
xor_4  g04827(new_n5203, new_n5174, new_n5204);
xor_4  g04828(new_n5204, new_n5173, new_n5205);
xor_4  g04829(new_n5171, new_n5145, new_n5206);
not_8  g04830(new_n5206, new_n5207);
nand_5 g04831(new_n1200, new_n1197, new_n5208);
not_8  g04832(new_n5208, new_n5209);
nand_5 g04833(n6016, n5331, new_n5210);
not_8  g04834(new_n5210, new_n5211);
nand_5 g04835(n8476, n521, new_n5212_1);
nand_5 g04836(n8476, n5579, new_n5213);
and_5  g04837(new_n5213, new_n1192, new_n5214);
and_5  g04838(new_n1195, new_n1191, new_n5215);
nor_5  g04839(new_n5215, new_n5214, new_n5216);
not_8  g04840(new_n5216, new_n5217);
xor_4  g04841(new_n5217, new_n5212_1, new_n5218);
nand_5 g04842(n12648, n2498, new_n5219);
not_8  g04843(new_n5219, new_n5220);
nand_5 g04844(n10545, n2558, new_n5221);
xor_4  g04845(new_n5221, new_n1125, new_n5222);
xor_4  g04846(new_n5222, new_n5220, new_n5223);
xor_4  g04847(new_n5223, new_n5218, new_n5224);
not_8  g04848(new_n5224, new_n5225);
xor_4  g04849(new_n5225, new_n5211, new_n5226);
nor_5  g04850(new_n1196, new_n1189, new_n5227);
nor_5  g04851(new_n5227, new_n1187, new_n5228);
xor_4  g04852(new_n5228, new_n5226, new_n5229);
not_8  g04853(new_n5229, new_n5230);
xor_4  g04854(new_n5230, new_n5209, new_n5231);
not_8  g04855(new_n1218, new_n5232);
nor_5  g04856(new_n5232, new_n1217, new_n5233);
not_8  g04857(new_n5233, new_n5234);
nand_5 g04858(n7965, n7270, new_n5235);
not_8  g04859(new_n5235, new_n5236);
nand_5 g04860(n7388, n806, new_n5237);
nand_5 g04861(n7388, n3342, new_n5238);
and_5  g04862(new_n5238, new_n1210, new_n5239);
and_5  g04863(new_n1213, new_n1209_1, new_n5240_1);
nor_5  g04864(new_n5240_1, new_n5239, new_n5241);
not_8  g04865(new_n5241, new_n5242);
xor_4  g04866(new_n5242, new_n5237, new_n5243);
nand_5 g04867(n9111, n2393, new_n5244);
not_8  g04868(new_n5244, new_n5245);
nand_5 g04869(n9763, n5860, new_n5246);
xor_4  g04870(new_n5246, new_n1106, new_n5247);
xor_4  g04871(new_n5247, new_n5245, new_n5248);
xor_4  g04872(new_n5248, new_n5243, new_n5249);
not_8  g04873(new_n5249, new_n5250);
xor_4  g04874(new_n5250, new_n5236, new_n5251);
nor_5  g04875(new_n1205, new_n1202, new_n5252);
nor_5  g04876(new_n1215, new_n5252, new_n5253);
xor_4  g04877(new_n5253, new_n5251, new_n5254);
not_8  g04878(new_n5254, new_n5255);
xor_4  g04879(new_n5255, new_n5234, new_n5256);
xor_4  g04880(new_n5256, new_n5231, new_n5257_1);
nor_5  g04881(new_n1219, new_n1201, new_n5258);
nor_5  g04882(new_n1224, new_n1221, new_n5259);
nor_5  g04883(new_n5259, new_n5258, new_n5260);
xor_4  g04884(new_n5260, new_n5257_1, new_n5261);
nor_5  g04885(new_n5261, new_n5207, new_n5262);
and_5  g04886(new_n1180, new_n1174, new_n5263);
nor_5  g04887(new_n1225, new_n1181, new_n5264);
nor_5  g04888(new_n5264, new_n5263, new_n5265);
xor_4  g04889(new_n5261, new_n5207, new_n5266);
not_8  g04890(new_n5266, new_n5267);
nor_5  g04891(new_n5267, new_n5265, new_n5268);
nor_5  g04892(new_n5268, new_n5262, new_n5269);
xor_4  g04893(new_n5269, new_n5205, new_n5270);
or_5   g04894(new_n5230, new_n5208, new_n5271);
not_8  g04895(new_n5271, new_n5272);
nand_5 g04896(n5798, n5331, new_n5273);
nand_5 g04897(n12648, n5579, new_n5274);
nand_5 g04898(n10545, n2498, new_n5275);
nand_5 g04899(n7690, n2558, new_n5276);
xor_4  g04900(new_n5276, new_n5275, new_n5277);
not_8  g04901(new_n5277, new_n5278);
xor_4  g04902(new_n5278, new_n5274, new_n5279);
and_5  g04903(new_n5221, new_n1125, new_n5280);
nor_5  g04904(new_n5221, new_n1125, new_n5281);
nor_5  g04905(new_n5281, new_n5220, new_n5282);
or_5   g04906(new_n5282, new_n5280, new_n5283_1);
not_8  g04907(new_n5283_1, new_n5284);
xor_4  g04908(new_n5284, new_n5279, new_n5285);
nand_5 g04909(n8476, n6016, new_n5286);
nand_5 g04910(n2530, n521, new_n5287);
xor_4  g04911(new_n5287, new_n5286, new_n5288);
xor_4  g04912(new_n5288, new_n5285, new_n5289);
not_8  g04913(new_n5289, new_n5290);
nor_5  g04914(new_n5217, new_n5212_1, new_n5291);
and_5  g04915(new_n5223, new_n5218, new_n5292);
nor_5  g04916(new_n5292, new_n5291, new_n5293);
xor_4  g04917(new_n5293, new_n5290, new_n5294);
not_8  g04918(new_n5294, new_n5295);
nor_5  g04919(new_n5225, new_n5210, new_n5296);
nor_5  g04920(new_n5228, new_n5226, new_n5297);
nor_5  g04921(new_n5297, new_n5296, new_n5298);
xor_4  g04922(new_n5298, new_n5295, new_n5299);
not_8  g04923(new_n5299, new_n5300);
xor_4  g04924(new_n5300, new_n5273, new_n5301);
xor_4  g04925(new_n5301, new_n5272, new_n5302);
not_8  g04926(new_n5302, new_n5303);
or_5   g04927(new_n5255, new_n5234, new_n5304);
not_8  g04928(new_n5304, new_n5305_1);
nand_5 g04929(n7965, n5153, new_n5306);
not_8  g04930(new_n5306, new_n5307);
nand_5 g04931(n3342, n2393, new_n5308);
nand_5 g04932(n9763, n3986, new_n5309);
nand_5 g04933(n9111, n5860, new_n5310);
xor_4  g04934(new_n5310, new_n5309, new_n5311);
not_8  g04935(new_n5311, new_n5312);
xor_4  g04936(new_n5312, new_n5308, new_n5313);
and_5  g04937(new_n5246, new_n1106, new_n5314_1);
nor_5  g04938(new_n5246, new_n1106, new_n5315);
nor_5  g04939(new_n5315, new_n5245, new_n5316);
or_5   g04940(new_n5316, new_n5314_1, new_n5317);
not_8  g04941(new_n5317, new_n5318);
xor_4  g04942(new_n5318, new_n5313, new_n5319_1);
nand_5 g04943(n7388, n7270, new_n5320_1);
nand_5 g04944(n11892, n806, new_n5321);
xor_4  g04945(new_n5321, new_n5320_1, new_n5322);
xor_4  g04946(new_n5322, new_n5319_1, new_n5323);
nor_5  g04947(new_n5242, new_n5237, new_n5324);
and_5  g04948(new_n5248, new_n5243, new_n5325);
nor_5  g04949(new_n5325, new_n5324, new_n5326);
xor_4  g04950(new_n5326, new_n5323, new_n5327);
nor_5  g04951(new_n5250, new_n5235, new_n5328);
nor_5  g04952(new_n5253, new_n5251, new_n5329);
nor_5  g04953(new_n5329, new_n5328, new_n5330);
xor_4  g04954(new_n5330, new_n5327, new_n5331_1);
xor_4  g04955(new_n5331_1, new_n5307, new_n5332);
not_8  g04956(new_n5332, new_n5333);
nand_5 g04957(new_n5333, new_n5305_1, new_n5334);
or_5   g04958(new_n5333, new_n5305_1, new_n5335);
and_5  g04959(new_n5335, new_n5334, new_n5336);
xnor_4 g04960(new_n5336, new_n5303, new_n5337);
not_8  g04961(new_n5231, new_n5338);
nor_5  g04962(new_n5256, new_n5338, new_n5339);
nor_5  g04963(new_n5260, new_n5257_1, new_n5340);
nor_5  g04964(new_n5340, new_n5339, new_n5341);
xor_4  g04965(new_n5341, new_n5337, new_n5342);
xor_4  g04966(new_n5342, new_n5270, new_n5343);
nor_5  g04967(new_n5343, new_n5143, new_n5344);
not_8  g04968(new_n5143, new_n5345);
xor_4  g04969(new_n5343, new_n5345, new_n5346);
not_8  g04970(new_n5346, new_n5347);
xor_4  g04971(new_n5135, new_n5134, new_n5348);
not_8  g04972(new_n5348, new_n5349);
not_8  g04973(new_n5265, new_n5350);
xor_4  g04974(new_n5267, new_n5350, new_n5351);
and_5  g04975(new_n5351, new_n5349, new_n5352);
nor_5  g04976(new_n1152, new_n1061, new_n5353);
not_8  g04977(new_n1226, new_n5354);
nor_5  g04978(new_n5354, new_n1154, new_n5355);
or_5   g04979(new_n5355, new_n5353, new_n5356);
xor_4  g04980(new_n5351, new_n5348, new_n5357);
nor_5  g04981(new_n5357, new_n5356, new_n5358);
or_5   g04982(new_n5358, new_n5352, new_n5359);
and_5  g04983(new_n5359, new_n5347, new_n5360);
nor_5  g04984(new_n5360, new_n5344, new_n5361);
xor_4  g04985(new_n5361, new_n5142, new_n5362);
not_8  g04986(new_n5362, new_n5363);
nor_5  g04987(new_n5203, new_n5174, new_n5364);
and_5  g04988(new_n5204, new_n5173, new_n5365);
or_5   g04989(new_n5365, new_n5364, new_n5366);
or_5   g04990(new_n5201, new_n5198_1, new_n5367);
or_5   g04991(new_n5196, new_n5189, new_n5368);
nand_5 g04992(n12221, n6776, new_n5369);
not_8  g04993(new_n5369, new_n5370);
nand_5 g04994(n12299, n12145, new_n5371);
nand_5 g04995(n10217, n8759, new_n5372);
xor_4  g04996(new_n5372, new_n5371, new_n5373);
not_8  g04997(new_n5373, new_n5374);
xor_4  g04998(new_n5374, new_n5370, new_n5375);
not_8  g04999(new_n5375, new_n5376);
xor_4  g05000(new_n5376, new_n5368, new_n5377);
or_5   g05001(new_n5193, new_n5192, new_n5378);
not_8  g05002(new_n5378, new_n5379);
nand_5 g05003(n7436, n2522, new_n5380);
not_8  g05004(new_n5380, new_n5381);
xor_4  g05005(new_n5381, new_n5379, new_n5382);
and_5  g05006(n9241, n2024, new_n5383);
nand_5 g05007(n10510, n7946, new_n5384);
nand_5 g05008(n9189, n8276, new_n5385);
xor_4  g05009(new_n5385, new_n5384, new_n5386);
xor_4  g05010(new_n5386, new_n5383, new_n5387);
xor_4  g05011(new_n5387, new_n5382, new_n5388);
xor_4  g05012(new_n5388, new_n5377, new_n5389);
not_8  g05013(new_n5389, new_n5390);
nor_5  g05014(new_n5181, new_n5177, new_n5391);
or_5   g05015(new_n5179, new_n5178, new_n5392);
not_8  g05016(new_n5392, new_n5393);
not_8  g05017(new_n5182, new_n5394);
or_5   g05018(new_n5197, new_n5394, new_n5395);
not_8  g05019(new_n5395, new_n5396);
xor_4  g05020(new_n5396, new_n5393, new_n5397);
nor_5  g05021(new_n5397, new_n5391, new_n5398);
xor_4  g05022(new_n5398, new_n5390, new_n5399);
not_8  g05023(new_n5399, new_n5400);
xor_4  g05024(new_n5400, new_n5367, new_n5401);
xor_4  g05025(new_n5401, new_n5366, new_n5402);
not_8  g05026(new_n5205, new_n5403);
nor_5  g05027(new_n5269, new_n5403, new_n5404);
nor_5  g05028(new_n5342, new_n5270, new_n5405);
nor_5  g05029(new_n5405, new_n5404, new_n5406);
xor_4  g05030(new_n5406, new_n5402, new_n5407);
or_5   g05031(new_n5298, new_n5295, new_n5408);
not_8  g05032(new_n5408, new_n5409);
nand_5 g05033(n8476, n5798, new_n5410);
nand_5 g05034(n6016, n2530, new_n5411_1);
and_5  g05035(n5331, n2347, new_n5412);
xor_4  g05036(new_n5412, new_n5411_1, new_n5413);
not_8  g05037(new_n5413, new_n5414);
xor_4  g05038(new_n5414, new_n5410, new_n5415);
not_8  g05039(new_n5415, new_n5416);
nor_5  g05040(new_n5278, new_n5274, new_n5417);
and_5  g05041(new_n5284, new_n5279, new_n5418);
or_5   g05042(new_n5418, new_n5417, new_n5419);
xor_4  g05043(new_n5419, new_n5416, new_n5420);
or_5   g05044(new_n5276, new_n5275, new_n5421);
not_8  g05045(new_n5421, new_n5422);
nand_5 g05046(n12648, n521, new_n5423);
not_8  g05047(new_n5423, new_n5424);
xor_4  g05048(new_n5424, new_n5422, new_n5425);
nand_5 g05049(n7690, n2498, new_n5426);
nand_5 g05050(n10545, n5579, new_n5427);
nand_5 g05051(n3616, n2558, new_n5428);
xor_4  g05052(new_n5428, new_n5427, new_n5429);
not_8  g05053(new_n5429, new_n5430);
xor_4  g05054(new_n5430, new_n5426, new_n5431);
xor_4  g05055(new_n5431, new_n5425, new_n5432);
xor_4  g05056(new_n5432, new_n5420, new_n5433);
not_8  g05057(new_n5433, new_n5434);
nand_5 g05058(new_n5288, new_n5285, new_n5435_1);
or_5   g05059(new_n5287, new_n5286, new_n5436);
or_5   g05060(new_n5293, new_n5290, new_n5437);
not_8  g05061(new_n5437, new_n5438);
xor_4  g05062(new_n5438, new_n5436, new_n5439);
and_5  g05063(new_n5439, new_n5435_1, new_n5440);
xor_4  g05064(new_n5440, new_n5434, new_n5441);
xor_4  g05065(new_n5441, new_n5409, new_n5442);
not_8  g05066(new_n5442, new_n5443);
nor_5  g05067(new_n5300, new_n5273, new_n5444);
and_5  g05068(new_n5301, new_n5272, new_n5445);
nor_5  g05069(new_n5445, new_n5444, new_n5446);
xor_4  g05070(new_n5446, new_n5443, new_n5447);
not_8  g05071(new_n5447, new_n5448);
or_5   g05072(new_n5330, new_n5327, new_n5449);
not_8  g05073(new_n5449, new_n5450);
nor_5  g05074(new_n5312, new_n5308, new_n5451);
and_5  g05075(new_n5318, new_n5313, new_n5452);
or_5   g05076(new_n5452, new_n5451, new_n5453);
nand_5 g05077(n7388, n5153, new_n5454);
not_8  g05078(new_n5454, new_n5455);
nand_5 g05079(n11892, n7270, new_n5456);
nand_5 g05080(n7965, n2507, new_n5457);
xor_4  g05081(new_n5457, new_n5456, new_n5458);
not_8  g05082(new_n5458, new_n5459);
xor_4  g05083(new_n5459, new_n5455, new_n5460);
not_8  g05084(new_n5460, new_n5461);
xor_4  g05085(new_n5461, new_n5453, new_n5462);
or_5   g05086(new_n5310, new_n5309, new_n5463);
not_8  g05087(new_n5463, new_n5464);
nand_5 g05088(n2393, n806, new_n5465);
not_8  g05089(new_n5465, new_n5466);
xor_4  g05090(new_n5466, new_n5464, new_n5467);
nand_5 g05091(n9111, n3986, new_n5468);
nand_5 g05092(n5860, n3342, new_n5469);
nand_5 g05093(n9763, n5857, new_n5470);
xor_4  g05094(new_n5470, new_n5469, new_n5471);
not_8  g05095(new_n5471, new_n5472);
xor_4  g05096(new_n5472, new_n5468, new_n5473);
xor_4  g05097(new_n5473, new_n5467, new_n5474);
xor_4  g05098(new_n5474, new_n5462, new_n5475);
not_8  g05099(new_n5475, new_n5476);
nand_5 g05100(new_n5322, new_n5319_1, new_n5477);
or_5   g05101(new_n5321, new_n5320_1, new_n5478);
not_8  g05102(new_n5323, new_n5479);
or_5   g05103(new_n5326, new_n5479, new_n5480);
not_8  g05104(new_n5480, new_n5481);
xor_4  g05105(new_n5481, new_n5478, new_n5482);
and_5  g05106(new_n5482, new_n5477, new_n5483);
xor_4  g05107(new_n5483, new_n5476, new_n5484);
xor_4  g05108(new_n5484, new_n5450, new_n5485);
not_8  g05109(new_n5485, new_n5486);
or_5   g05110(new_n5331_1, new_n5307, new_n5487);
nand_5 g05111(new_n5335, new_n5487, new_n5488);
xor_4  g05112(new_n5488, new_n5486, new_n5489);
xor_4  g05113(new_n5489, new_n5448, new_n5490);
and_5  g05114(new_n5336, new_n5303, new_n5491);
nor_5  g05115(new_n5341, new_n5337, new_n5492);
nor_5  g05116(new_n5492, new_n5491, new_n5493);
xor_4  g05117(new_n5493, new_n5490, new_n5494);
xor_4  g05118(new_n5494, new_n5407, new_n5495);
xor_4  g05119(new_n5495, new_n5363, n1523);
nand_5 g05120(n6687, n4634, new_n5497);
nand_5 g05121(n10223, n4189, new_n5498);
nor_5  g05122(new_n5498, new_n4210, new_n5499);
and_5  g05123(n10223, n6687, new_n5500);
and_5  g05124(n7265, n4189, new_n5501);
nor_5  g05125(new_n5501, new_n5500, new_n5502);
nand_5 g05126(n2879, n2564, new_n5503);
nor_5  g05127(new_n5503, new_n5502, new_n5504);
nor_5  g05128(new_n5504, new_n5499, new_n5505);
xor_4  g05129(new_n5505, new_n5497, new_n5506);
not_8  g05130(new_n5506, new_n5507);
nand_5 g05131(n4189, n2879, new_n5508);
not_8  g05132(new_n5508, new_n5509);
nand_5 g05133(n10223, n2564, new_n5510);
nand_5 g05134(n7265, n6770, new_n5511);
xor_4  g05135(new_n5511, new_n5510, new_n5512);
not_8  g05136(new_n5512, new_n5513);
xor_4  g05137(new_n5513, new_n5509, new_n5514);
nor_5  g05138(new_n5514, new_n5507, new_n5515);
and_5  g05139(new_n5514, new_n5507, new_n5516);
or_5   g05140(new_n5516, new_n5515, new_n5517);
nor_5  g05141(new_n5502, new_n5499, new_n5518);
nand_5 g05142(n7265, n2564, new_n5519);
nand_5 g05143(n6687, n2879, new_n5520);
or_5   g05144(new_n5520, new_n5519, new_n5521);
or_5   g05145(new_n5521, new_n5518, new_n5522);
or_5   g05146(new_n5522, new_n5517, new_n5523);
nand_5 g05147(n9195, n6687, new_n5524);
not_8  g05148(new_n5524, new_n5525);
nand_5 g05149(n4634, n2564, new_n5526);
nand_5 g05150(n6770, n2879, new_n5527);
not_8  g05151(new_n5527, new_n5528);
nand_5 g05152(n9920, n7265, new_n5529);
xor_4  g05153(new_n5529, new_n5498, new_n5530);
not_8  g05154(new_n5530, new_n5531);
xor_4  g05155(new_n5531, new_n5528, new_n5532);
xor_4  g05156(new_n5532, new_n5526, new_n5533);
and_5  g05157(new_n5511, new_n5510, new_n5534);
nor_5  g05158(new_n5513, new_n5509, new_n5535);
or_5   g05159(new_n5535, new_n5534, new_n5536);
not_8  g05160(new_n5536, new_n5537);
xor_4  g05161(new_n5537, new_n5533, new_n5538);
xor_4  g05162(new_n5538, new_n5525, new_n5539);
not_8  g05163(new_n5539, new_n5540);
nor_5  g05164(new_n5505, new_n5497, new_n5541);
nor_5  g05165(new_n5515, new_n5541, new_n5542);
xor_4  g05166(new_n5542, new_n5540, new_n5543);
not_8  g05167(new_n5543, new_n5544);
xor_4  g05168(new_n5544, new_n5523, new_n5545);
not_8  g05169(new_n5545, new_n5546);
nand_5 g05170(n8336, n2522, new_n5547);
not_8  g05171(new_n5547, new_n5548);
and_5  g05172(n9189, n8336, new_n5549);
and_5  g05173(n7946, n6986, new_n5550);
nor_5  g05174(new_n5550, new_n5549, new_n5551);
nand_5 g05175(n9189, n6986, new_n5552);
nor_5  g05176(new_n5552, new_n4212, new_n5553);
nand_5 g05177(n10928, n2024, new_n5554);
not_8  g05178(new_n5554, new_n5555);
nor_5  g05179(new_n5555, new_n5553, new_n5556);
nor_5  g05180(new_n5556, new_n5551, new_n5557);
not_8  g05181(new_n5557, new_n5558);
xor_4  g05182(new_n5558, new_n5548, new_n5559);
nand_5 g05183(n6986, n2024, new_n5560);
not_8  g05184(new_n5560, new_n5561);
nand_5 g05185(n10928, n9189, new_n5562);
nand_5 g05186(n7946, n2226, new_n5563);
xor_4  g05187(new_n5563, new_n5562, new_n5564);
xor_4  g05188(new_n5564, new_n5561, new_n5565);
not_8  g05189(new_n5565, new_n5566);
xor_4  g05190(new_n5566, new_n5559, new_n5567);
not_8  g05191(new_n4212, new_n5568);
or_5   g05192(new_n5554, new_n5568, new_n5569);
not_8  g05193(new_n5569, new_n5570);
nor_5  g05194(new_n5553, new_n5551, new_n5571);
or_5   g05195(new_n5571, new_n5570, new_n5572);
not_8  g05196(new_n5572, new_n5573);
nand_5 g05197(new_n5573, new_n5555, new_n5574);
not_8  g05198(new_n5574, new_n5575);
nand_5 g05199(new_n5575, new_n5567, new_n5576);
not_8  g05200(new_n5576, new_n5577);
nand_5 g05201(n12145, n8336, new_n5578);
not_8  g05202(new_n5578, new_n5579_1);
nand_5 g05203(n10928, n2522, new_n5580);
not_8  g05204(new_n5580, new_n5581);
and_5  g05205(new_n5563, new_n5562, new_n5582);
nor_5  g05206(new_n5563, new_n5562, new_n5583);
nor_5  g05207(new_n5583, new_n5561, new_n5584);
nor_5  g05208(new_n5584, new_n5582, new_n5585);
not_8  g05209(new_n5585, new_n5586);
xor_4  g05210(new_n5586, new_n5581, new_n5587);
nand_5 g05211(n2226, n2024, new_n5588);
not_8  g05212(new_n5588, new_n5589);
nand_5 g05213(n7946, n1094, new_n5590);
xor_4  g05214(new_n5590, new_n5552, new_n5591);
not_8  g05215(new_n5591, new_n5592);
xor_4  g05216(new_n5592, new_n5589, new_n5593);
xor_4  g05217(new_n5593, new_n5587, new_n5594);
xor_4  g05218(new_n5594, new_n5579_1, new_n5595);
nor_5  g05219(new_n5558, new_n5547, new_n5596);
nor_5  g05220(new_n5566, new_n5559, new_n5597);
or_5   g05221(new_n5597, new_n5596, new_n5598);
xor_4  g05222(new_n5598, new_n5595, new_n5599);
not_8  g05223(new_n5599, new_n5600);
xor_4  g05224(new_n5600, new_n5577, new_n5601);
not_8  g05225(new_n5601, new_n5602);
xor_4  g05226(new_n5574, new_n5567, new_n5603);
nand_5 g05227(n12069, n521, new_n5604);
not_8  g05228(new_n5604, new_n5605);
nand_5 g05229(n7891, n5579, new_n5606);
nor_5  g05230(new_n5606, new_n4214, new_n5607);
and_5  g05231(n12069, n5579, new_n5608);
and_5  g05232(n7891, n2558, new_n5609);
nor_5  g05233(new_n5609, new_n5608, new_n5610);
nand_5 g05234(n12391, n2498, new_n5611);
nor_5  g05235(new_n5611, new_n5610, new_n5612);
nor_5  g05236(new_n5612, new_n5607, new_n5613);
xor_4  g05237(new_n5613, new_n5605, new_n5614);
not_8  g05238(new_n5614, new_n5615);
nand_5 g05239(n7891, n2498, new_n5616);
not_8  g05240(new_n5616, new_n5617);
nand_5 g05241(n12391, n5579, new_n5618);
nand_5 g05242(n7160, n2558, new_n5619);
xor_4  g05243(new_n5619, new_n5618, new_n5620);
xor_4  g05244(new_n5620, new_n5617, new_n5621);
and_5  g05245(new_n5621, new_n5615, new_n5622);
nor_5  g05246(new_n5621, new_n5615, new_n5623);
or_5   g05247(new_n5623, new_n5622, new_n5624);
nor_5  g05248(new_n5610, new_n5607, new_n5625);
and_5  g05249(n12391, n2558, new_n5626);
and_5  g05250(n12069, n2498, new_n5627);
nand_5 g05251(new_n5627, new_n5626, new_n5628);
or_5   g05252(new_n5628, new_n5625, new_n5629);
not_8  g05253(new_n5629, new_n5630);
xor_4  g05254(new_n5630, new_n5624, new_n5631);
nand_5 g05255(n11222, n806, new_n5632);
and_5  g05256(n11222, n3342, new_n5633);
and_5  g05257(n9763, n5314, new_n5634);
or_5   g05258(new_n5634, new_n5633, new_n5635);
not_8  g05259(new_n5635, new_n5636);
nand_5 g05260(n5314, n3342, new_n5637);
nor_5  g05261(new_n5637, new_n4213, new_n5638);
nand_5 g05262(n11153, n9111, new_n5639);
not_8  g05263(new_n5639, new_n5640);
nor_5  g05264(new_n5640, new_n5638, new_n5641_1);
nor_5  g05265(new_n5641_1, new_n5636, new_n5642);
not_8  g05266(new_n5642, new_n5643);
xor_4  g05267(new_n5643, new_n5632, new_n5644);
nand_5 g05268(n9111, n5314, new_n5645_1);
not_8  g05269(new_n5645_1, new_n5646);
nand_5 g05270(n11153, n3342, new_n5647);
nand_5 g05271(n9763, n996, new_n5648);
xor_4  g05272(new_n5648, new_n5647, new_n5649);
xor_4  g05273(new_n5649, new_n5646, new_n5650);
xor_4  g05274(new_n5650, new_n5644, new_n5651);
not_8  g05275(new_n4213, new_n5652);
or_5   g05276(new_n5639, new_n5652, new_n5653);
and_5  g05277(new_n5653, new_n5636, new_n5654);
or_5   g05278(new_n5654, new_n5638, new_n5655);
not_8  g05279(new_n5655, new_n5656);
nor_5  g05280(new_n5656, new_n5639, new_n5657);
xor_4  g05281(new_n5657, new_n5651, new_n5658);
not_8  g05282(new_n5658, new_n5659);
xnor_4 g05283(new_n5659, new_n5631, new_n5660);
or_5   g05284(new_n5653, new_n5636, new_n5661);
nand_5 g05285(new_n5661, new_n5656, new_n5662);
or_5   g05286(new_n4214, new_n4213, new_n5663);
not_8  g05287(new_n5663, new_n5664);
xor_4  g05288(new_n5627, new_n5626, new_n5665);
nor_5  g05289(new_n5665, new_n5664, new_n5666);
xor_4  g05290(new_n5665, new_n5663, new_n5667);
not_8  g05291(new_n5667, new_n5668);
nand_5 g05292(n11153, n9763, new_n5669);
and_5  g05293(n11222, n9111, new_n5670_1);
xor_4  g05294(new_n5670_1, new_n5669, new_n5671);
and_5  g05295(new_n5671, new_n5668, new_n5672);
or_5   g05296(new_n5672, new_n5666, new_n5673);
and_5  g05297(new_n5673, new_n5662, new_n5674);
nor_5  g05298(new_n5672, new_n5666, new_n5675);
xor_4  g05299(new_n5675, new_n5662, new_n5676);
not_8  g05300(new_n5611, new_n5677);
and_5  g05301(new_n5677, new_n4214, new_n5678);
nor_5  g05302(new_n5678, new_n5625, new_n5679);
or_5   g05303(new_n5609, new_n5608, new_n5680);
and_5  g05304(new_n5678, new_n5680, new_n5681);
nor_5  g05305(new_n5681, new_n5679, new_n5682);
nor_5  g05306(new_n5682, new_n5676, new_n5683);
nor_5  g05307(new_n5683, new_n5674, new_n5684);
xor_4  g05308(new_n5684, new_n5660, new_n5685);
nor_5  g05309(new_n5685, new_n5603, new_n5686);
not_8  g05310(new_n5603, new_n5687);
xor_4  g05311(new_n5685, new_n5687, new_n5688);
nor_5  g05312(new_n5569, new_n5551, new_n5689);
or_5   g05313(new_n5689, new_n5573, new_n5690);
xor_4  g05314(new_n5682, new_n5676, new_n5691);
nor_5  g05315(new_n5691, new_n5690, new_n5692);
xor_4  g05316(new_n5691, new_n5690, new_n5693_1);
not_8  g05317(new_n5693_1, new_n5694_1);
xor_4  g05318(new_n5671, new_n5668, new_n5695);
nand_5 g05319(n10928, n7946, new_n5696);
and_5  g05320(n8336, n2024, new_n5697);
xor_4  g05321(new_n5697, new_n5696, new_n5698);
nor_5  g05322(new_n5698, new_n5695, new_n5699);
or_5   g05323(new_n4216, new_n4212, new_n5700);
not_8  g05324(new_n5700, new_n5701);
xor_4  g05325(new_n5698, new_n5695, new_n5702);
and_5  g05326(new_n5702, new_n5701, new_n5703);
nor_5  g05327(new_n5703, new_n5699, new_n5704);
nor_5  g05328(new_n5704, new_n5694_1, new_n5705);
nor_5  g05329(new_n5705, new_n5692, new_n5706);
nor_5  g05330(new_n5706, new_n5688, new_n5707);
nor_5  g05331(new_n5707, new_n5686, new_n5708);
xor_4  g05332(new_n5708, new_n5602, new_n5709);
or_5   g05333(new_n5629, new_n5624, new_n5710);
nand_5 g05334(n12069, n6016, new_n5711);
not_8  g05335(new_n5711, new_n5712);
nand_5 g05336(n12391, n521, new_n5713);
not_8  g05337(new_n5713, new_n5714);
and_5  g05338(new_n5619, new_n5618, new_n5715);
nor_5  g05339(new_n5619, new_n5618, new_n5716);
nor_5  g05340(new_n5716, new_n5617, new_n5717);
nor_5  g05341(new_n5717, new_n5715, new_n5718);
not_8  g05342(new_n5718, new_n5719);
xor_4  g05343(new_n5719, new_n5714, new_n5720);
and_5  g05344(n7160, n2498, new_n5721);
not_8  g05345(new_n5721, new_n5722);
and_5  g05346(n4828, n2558, new_n5723);
xor_4  g05347(new_n5723, new_n5606, new_n5724);
not_8  g05348(new_n5724, new_n5725);
xor_4  g05349(new_n5725, new_n5722, new_n5726);
xor_4  g05350(new_n5726, new_n5720, new_n5727);
xor_4  g05351(new_n5727, new_n5712, new_n5728);
not_8  g05352(new_n5728, new_n5729);
nor_5  g05353(new_n5613, new_n5604, new_n5730);
nor_5  g05354(new_n5622, new_n5730, new_n5731);
xor_4  g05355(new_n5731, new_n5729, new_n5732);
not_8  g05356(new_n5732, new_n5733);
xor_4  g05357(new_n5733, new_n5710, new_n5734);
nand_5 g05358(new_n5657, new_n5651, new_n5735);
not_8  g05359(new_n5735, new_n5736);
nand_5 g05360(n11222, n7270, new_n5737);
not_8  g05361(new_n5737, new_n5738);
nand_5 g05362(n11153, n806, new_n5739);
and_5  g05363(new_n5648, new_n5647, new_n5740);
nor_5  g05364(new_n5648, new_n5647, new_n5741);
nor_5  g05365(new_n5741, new_n5646, new_n5742);
nor_5  g05366(new_n5742, new_n5740, new_n5743);
not_8  g05367(new_n5743, new_n5744);
xor_4  g05368(new_n5744, new_n5739, new_n5745);
nand_5 g05369(n9111, n996, new_n5746);
not_8  g05370(new_n5746, new_n5747);
nand_5 g05371(n9763, n5767, new_n5748);
xor_4  g05372(new_n5748, new_n5637, new_n5749);
xor_4  g05373(new_n5749, new_n5747, new_n5750);
xor_4  g05374(new_n5750, new_n5745, new_n5751);
xor_4  g05375(new_n5751, new_n5738, new_n5752);
or_5   g05376(new_n5643, new_n5632, new_n5753);
not_8  g05377(new_n5753, new_n5754);
and_5  g05378(new_n5650, new_n5644, new_n5755);
or_5   g05379(new_n5755, new_n5754, new_n5756);
xor_4  g05380(new_n5756, new_n5752, new_n5757);
not_8  g05381(new_n5757, new_n5758);
xor_4  g05382(new_n5758, new_n5736, new_n5759);
xor_4  g05383(new_n5759, new_n5734, new_n5760_1);
and_5  g05384(new_n5659, new_n5631, new_n5761);
nor_5  g05385(new_n5684, new_n5660, new_n5762);
nor_5  g05386(new_n5762, new_n5761, new_n5763);
xor_4  g05387(new_n5763, new_n5760_1, new_n5764);
xor_4  g05388(new_n5764, new_n5709, new_n5765);
xor_4  g05389(new_n5765, new_n5546, new_n5766);
not_8  g05390(new_n5766, new_n5767_1);
xor_4  g05391(new_n5522, new_n5517, new_n5768);
xor_4  g05392(new_n5706, new_n5688, new_n5769);
nor_5  g05393(new_n5769, new_n5768, new_n5770);
or_5   g05394(new_n5703, new_n5699, new_n5771);
xor_4  g05395(new_n5771, new_n5694_1, new_n5772);
not_8  g05396(new_n5503, new_n5773);
and_5  g05397(new_n5773, new_n4210, new_n5774);
nor_5  g05398(new_n5774, new_n5518, new_n5775);
or_5   g05399(new_n5501, new_n5500, new_n5776);
and_5  g05400(new_n5774, new_n5776, new_n5777);
or_5   g05401(new_n5777, new_n5775, new_n5778);
and_5  g05402(new_n5778, new_n5772, new_n5779);
nor_5  g05403(new_n5777, new_n5775, new_n5780);
xor_4  g05404(new_n5780, new_n5772, new_n5781);
nand_5 g05405(new_n4217, new_n4211, new_n5782);
xnor_4 g05406(new_n5520, new_n5519, new_n5783);
and_5  g05407(new_n5783, new_n5782, new_n5784);
xor_4  g05408(new_n5702, new_n5701, new_n5785);
xor_4  g05409(new_n5783, new_n5782, new_n5786);
not_8  g05410(new_n5786, new_n5787);
nor_5  g05411(new_n5787, new_n5785, new_n5788);
or_5   g05412(new_n5788, new_n5784, new_n5789);
not_8  g05413(new_n5789, new_n5790);
nor_5  g05414(new_n5790, new_n5781, new_n5791);
or_5   g05415(new_n5791, new_n5779, new_n5792);
not_8  g05416(new_n5768, new_n5793);
xor_4  g05417(new_n5769, new_n5793, new_n5794);
not_8  g05418(new_n5794, new_n5795);
and_5  g05419(new_n5795, new_n5792, new_n5796);
or_5   g05420(new_n5796, new_n5770, new_n5797);
nor_5  g05421(new_n5797, new_n5767_1, new_n5798_1);
and_5  g05422(new_n5797, new_n5767_1, new_n5799);
or_5   g05423(new_n5799, new_n5798_1, n1658);
nand_5 g05424(n7862, n4634, new_n5801);
not_8  g05425(new_n5801, new_n5802);
and_5  g05426(n10223, n7862, new_n5803);
and_5  g05427(n7265, n3172, new_n5804);
or_5   g05428(new_n5804, new_n5803, new_n5805);
not_8  g05429(new_n5805, new_n5806);
nand_5 g05430(n7862, n7265, new_n5807);
nand_5 g05431(n10223, n3172, new_n5808);
nor_5  g05432(new_n5808, new_n5807, new_n5809);
nand_5 g05433(n2879, n1333, new_n5810);
not_8  g05434(new_n5810, new_n5811);
nor_5  g05435(new_n5811, new_n5809, new_n5812);
or_5   g05436(new_n5812, new_n5806, new_n5813);
not_8  g05437(new_n5813, new_n5814_1);
xor_4  g05438(new_n5814_1, new_n5802, new_n5815);
nand_5 g05439(n3172, n2879, new_n5816);
not_8  g05440(new_n5816, new_n5817);
nand_5 g05441(n10223, n1333, new_n5818);
nand_5 g05442(n11757, n7265, new_n5819);
xor_4  g05443(new_n5819, new_n5818, new_n5820);
xor_4  g05444(new_n5820, new_n5817, new_n5821);
xor_4  g05445(new_n5821, new_n5815, new_n5822);
not_8  g05446(new_n5807, new_n5823);
or_5   g05447(new_n5810, new_n5823, new_n5824);
and_5  g05448(new_n5824, new_n5806, new_n5825);
or_5   g05449(new_n5825, new_n5809, new_n5826);
not_8  g05450(new_n5826, new_n5827);
or_5   g05451(new_n5827, new_n5810, new_n5828);
xor_4  g05452(new_n5828, new_n5822, new_n5829);
not_8  g05453(new_n5829, new_n5830);
nand_5 g05454(n6877, n2522, new_n5831);
nand_5 g05455(n2464, n2024, new_n5832);
not_8  g05456(new_n5832, new_n5833);
nand_5 g05457(n9400, n9189, new_n5834);
nand_5 g05458(n11311, n7946, new_n5835);
xor_4  g05459(new_n5835, new_n5834, new_n5836);
not_8  g05460(new_n5836, new_n5837);
xor_4  g05461(new_n5837, new_n5833, new_n5838);
xor_4  g05462(new_n5838, new_n5831, new_n5839);
and_5  g05463(n9189, n6877, new_n5840);
and_5  g05464(n7946, n2464, new_n5841);
nor_5  g05465(new_n5841, new_n5840, new_n5842);
nand_5 g05466(n7946, n6877, new_n5843);
nand_5 g05467(n9189, n2464, new_n5844);
nor_5  g05468(new_n5844, new_n5843, new_n5845);
nand_5 g05469(n9400, n2024, new_n5846);
not_8  g05470(new_n5846, new_n5847);
nor_5  g05471(new_n5847, new_n5845, new_n5848);
or_5   g05472(new_n5848, new_n5842, new_n5849);
not_8  g05473(new_n5849, new_n5850);
xor_4  g05474(new_n5850, new_n5839, new_n5851);
not_8  g05475(new_n5843, new_n5852);
or_5   g05476(new_n5846, new_n5852, new_n5853);
not_8  g05477(new_n5853, new_n5854);
nor_5  g05478(new_n5845, new_n5842, new_n5855);
nor_5  g05479(new_n5855, new_n5854, new_n5856);
not_8  g05480(new_n5856, new_n5857_1);
or_5   g05481(new_n5857_1, new_n5846, new_n5858);
xor_4  g05482(new_n5858, new_n5851, new_n5859);
not_8  g05483(new_n5859, new_n5860_1);
or_5   g05484(new_n5853, new_n5842, new_n5861);
and_5  g05485(new_n5861, new_n5857_1, new_n5862);
not_8  g05486(new_n5862, new_n5863);
nand_5 g05487(n4805, n2558, new_n5864);
nand_5 g05488(n9763, n7236, new_n5865);
xnor_4 g05489(new_n5865, new_n5864, new_n5866);
not_8  g05490(new_n5866, new_n5867);
nand_5 g05491(new_n5867, new_n5852, new_n5868);
nand_5 g05492(n9400, n7946, new_n5869);
and_5  g05493(n6877, n2024, new_n5870);
xor_4  g05494(new_n5870, new_n5869, new_n5871);
nor_5  g05495(new_n5871, new_n5868, new_n5872);
or_5   g05496(new_n5865, new_n5864, new_n5873);
and_5  g05497(n9111, n7236, new_n5874);
and_5  g05498(n9763, n3992, new_n5875);
xor_4  g05499(new_n5875, new_n5874, new_n5876);
xor_4  g05500(new_n5876, new_n5873, new_n5877);
not_8  g05501(new_n5877, new_n5878);
nand_5 g05502(n4805, n2498, new_n5879);
and_5  g05503(n11478, n2558, new_n5880);
xor_4  g05504(new_n5880, new_n5879, new_n5881);
xor_4  g05505(new_n5881, new_n5878, new_n5882);
not_8  g05506(new_n5871, new_n5883);
xor_4  g05507(new_n5883, new_n5868, new_n5884);
nor_5  g05508(new_n5884, new_n5882, new_n5885);
or_5   g05509(new_n5885, new_n5872, new_n5886);
not_8  g05510(new_n5886, new_n5887);
and_5  g05511(new_n5887, new_n5863, new_n5888);
not_8  g05512(new_n5873, new_n5889);
nor_5  g05513(new_n5876, new_n5889, new_n5890);
and_5  g05514(new_n5881, new_n5878, new_n5891);
or_5   g05515(new_n5891, new_n5890, new_n5892);
not_8  g05516(new_n5864, new_n5893);
nand_5 g05517(n11478, n2498, new_n5894);
or_5   g05518(new_n5894, new_n5893, new_n5895);
nand_5 g05519(n5283, n2558, new_n5896);
nand_5 g05520(n5579, n4805, new_n5897);
xnor_4 g05521(new_n5897, new_n5896, new_n5898);
and_5  g05522(new_n5898, new_n5895, new_n5899);
and_5  g05523(new_n5897, new_n5896, new_n5900);
nor_5  g05524(new_n5900, new_n5895, new_n5901);
or_5   g05525(new_n5901, new_n5899, new_n5902);
not_8  g05526(new_n5902, new_n5903);
xor_4  g05527(new_n5903, new_n5892, new_n5904);
and_5  g05528(n9111, n3992, new_n5905);
and_5  g05529(new_n5905, new_n5865, new_n5906);
not_8  g05530(new_n5906, new_n5907);
nand_5 g05531(n9763, n8384, new_n5908);
nand_5 g05532(n7236, n3342, new_n5909);
nand_5 g05533(new_n5909, new_n5908, new_n5910);
nor_5  g05534(new_n5910, new_n5907, new_n5911);
xnor_4 g05535(new_n5909, new_n5908, new_n5912);
not_8  g05536(new_n5912, new_n5913);
and_5  g05537(new_n5913, new_n5907, new_n5914);
nor_5  g05538(new_n5914, new_n5911, new_n5915);
xor_4  g05539(new_n5915, new_n5904, new_n5916);
xor_4  g05540(new_n5887, new_n5862, new_n5917);
nor_5  g05541(new_n5917, new_n5916, new_n5918);
or_5   g05542(new_n5918, new_n5888, new_n5919);
not_8  g05543(new_n5919, new_n5920);
xor_4  g05544(new_n5920, new_n5860_1, new_n5921);
nand_5 g05545(n4805, n521, new_n5922);
not_8  g05546(new_n5922, new_n5923);
not_8  g05547(new_n5894, new_n5924);
nor_5  g05548(new_n5897, new_n5896, new_n5925);
nor_5  g05549(new_n5925, new_n5924, new_n5926);
or_5   g05550(new_n5926, new_n5900, new_n5927);
not_8  g05551(new_n5927, new_n5928);
and_5  g05552(new_n5928, new_n5923, new_n5929);
nor_5  g05553(new_n5928, new_n5923, new_n5930);
or_5   g05554(new_n5930, new_n5929, new_n5931);
nand_5 g05555(n5283, n2498, new_n5932);
not_8  g05556(new_n5932, new_n5933);
nand_5 g05557(n2558, n137, new_n5934_1);
nand_5 g05558(n11478, n5579, new_n5935);
xor_4  g05559(new_n5935, new_n5934_1, new_n5936);
xor_4  g05560(new_n5936, new_n5933, new_n5937);
xor_4  g05561(new_n5937, new_n5931, new_n5938);
not_8  g05562(new_n5899, new_n5939);
or_5   g05563(new_n5939, new_n5894, new_n5940);
not_8  g05564(new_n5940, new_n5941);
xor_4  g05565(new_n5941, new_n5938, new_n5942);
not_8  g05566(new_n5942, new_n5943);
nand_5 g05567(n7236, n806, new_n5944);
nor_5  g05568(new_n5909, new_n5908, new_n5945);
nand_5 g05569(n9111, n3992, new_n5946);
not_8  g05570(new_n5910, new_n5947);
nor_5  g05571(new_n5947, new_n5946, new_n5948);
nor_5  g05572(new_n5948, new_n5945, new_n5949);
xor_4  g05573(new_n5949, new_n5944, new_n5950);
not_8  g05574(new_n5950, new_n5951);
nand_5 g05575(n9111, n8384, new_n5952);
not_8  g05576(new_n5952, new_n5953);
nand_5 g05577(n9763, n6358, new_n5954);
nand_5 g05578(n3992, n3342, new_n5955);
xor_4  g05579(new_n5955, new_n5954, new_n5956);
xor_4  g05580(new_n5956, new_n5953, new_n5957);
not_8  g05581(new_n5957, new_n5958);
xor_4  g05582(new_n5958, new_n5951, new_n5959);
nand_5 g05583(new_n5875, new_n5874, new_n5960);
or_5   g05584(new_n5913, new_n5960, new_n5961);
not_8  g05585(new_n5961, new_n5962);
xor_4  g05586(new_n5962, new_n5959, new_n5963);
xnor_4 g05587(new_n5963, new_n5943, new_n5964_1);
and_5  g05588(new_n5902, new_n5892, new_n5965);
not_8  g05589(new_n5915, new_n5966);
nor_5  g05590(new_n5966, new_n5904, new_n5967);
nor_5  g05591(new_n5967, new_n5965, new_n5968);
xor_4  g05592(new_n5968, new_n5964_1, new_n5969);
xor_4  g05593(new_n5969, new_n5921, new_n5970);
xor_4  g05594(new_n5970, new_n5830, new_n5971);
or_5   g05595(new_n5824, new_n5806, new_n5972);
nand_5 g05596(new_n5972, new_n5827, new_n5973);
not_8  g05597(new_n5916, new_n5974);
xnor_4 g05598(new_n5917, new_n5974, new_n5975);
nor_5  g05599(new_n5975, new_n5973, new_n5976);
xor_4  g05600(new_n5867, new_n5852, new_n5977);
nand_5 g05601(new_n5977, new_n5823, new_n5978);
nand_5 g05602(n7265, n1333, new_n5979);
and_5  g05603(n7862, n2879, new_n5980);
xor_4  g05604(new_n5980, new_n5979, new_n5981);
and_5  g05605(new_n5981, new_n5978, new_n5982);
xor_4  g05606(new_n5884, new_n5882, new_n5983);
xor_4  g05607(new_n5981, new_n5978, new_n5984);
not_8  g05608(new_n5984, new_n5985);
nor_5  g05609(new_n5985, new_n5983, new_n5986);
or_5   g05610(new_n5986, new_n5982, new_n5987);
xor_4  g05611(new_n5975, new_n5973, new_n5988);
not_8  g05612(new_n5988, new_n5989);
nor_5  g05613(new_n5989, new_n5987, new_n5990);
or_5   g05614(new_n5990, new_n5976, new_n5991);
not_8  g05615(new_n5991, new_n5992);
xor_4  g05616(new_n5992, new_n5971, n1847);
nand_5 g05617(n5305, n1798, new_n5994);
not_8  g05618(new_n5994, new_n5995);
nand_5 g05619(n8759, n6703, new_n5996);
nand_5 g05620(n5645, n5331, new_n5997);
nand_5 g05621(n11876, n7965, new_n5998);
xor_4  g05622(new_n5998, new_n5997, new_n5999);
not_8  g05623(new_n5999, new_n6000);
xor_4  g05624(new_n6000, new_n5996, new_n6001);
nand_5 g05625(new_n6001, new_n5995, new_n6002);
nand_5 g05626(n5305, n3932, new_n6003);
nand_5 g05627(n5964, n1798, new_n6004);
xor_4  g05628(new_n6004, new_n6003, new_n6005);
not_8  g05629(new_n6005, new_n6006);
xor_4  g05630(new_n6006, new_n6002, new_n6007);
not_8  g05631(new_n6007, new_n6008);
or_5   g05632(new_n6000, new_n5996, new_n6009);
nand_5 g05633(n9640, n8759, new_n6010);
and_5  g05634(n6776, n6703, new_n6011);
xor_4  g05635(new_n6011, new_n6010, new_n6012);
xor_4  g05636(new_n6012, new_n6009, new_n6013);
or_5   g05637(new_n5998, new_n5997, new_n6014);
not_8  g05638(new_n6014, new_n6015);
and_5  g05639(n10898, n7965, new_n6016_1);
and_5  g05640(n11876, n7388, new_n6017);
xor_4  g05641(new_n6017, new_n6016_1, new_n6018);
not_8  g05642(new_n6018, new_n6019);
xor_4  g05643(new_n6019, new_n6015, new_n6020);
nand_5 g05644(n5331, n1067, new_n6021);
nand_5 g05645(n8476, n5645, new_n6022);
xor_4  g05646(new_n6022, new_n6021, new_n6023);
not_8  g05647(new_n6023, new_n6024);
xor_4  g05648(new_n6024, new_n6020, new_n6025);
xor_4  g05649(new_n6025, new_n6013, new_n6026);
not_8  g05650(new_n6026, new_n6027);
xor_4  g05651(new_n6027, new_n6008, n2096);
xnor_4 g05652(new_n3546, new_n3543, n2131);
nand_5 g05653(n7456, n2564, new_n6030);
and_5  g05654(new_n3718, new_n3717, new_n6031);
nor_5  g05655(new_n3718, new_n3717, new_n6032);
nor_5  g05656(new_n6032, new_n3716, new_n6033);
nor_5  g05657(new_n6033, new_n6031, new_n6034);
not_8  g05658(new_n6034, new_n6035);
nor_5  g05659(new_n6035, new_n6030, new_n6036);
not_8  g05660(new_n6030, new_n6037);
xor_4  g05661(new_n6035, new_n6037, new_n6038_1);
nand_5 g05662(n6770, n3932, new_n6039);
not_8  g05663(new_n6039, new_n6040);
nand_5 g05664(n9920, n1798, new_n6041);
xor_4  g05665(new_n6041, new_n3706, new_n6042);
xor_4  g05666(new_n6042, new_n6040, new_n6043);
not_8  g05667(new_n6043, new_n6044);
nor_5  g05668(new_n6044, new_n6038_1, new_n6045);
or_5   g05669(new_n6045, new_n6036, new_n6046);
nand_5 g05670(n11662, n2564, new_n6047);
nand_5 g05671(n7456, n4189, new_n6048);
xor_4  g05672(new_n6048, new_n6047, new_n6049);
xor_4  g05673(new_n6049, new_n6046, new_n6050);
not_8  g05674(new_n6050, new_n6051);
nand_5 g05675(n12591, n6770, new_n6052);
nand_5 g05676(n3627, n1798, new_n6053);
nand_5 g05677(n9920, n3932, new_n6054);
xor_4  g05678(new_n6054, new_n6053, new_n6055);
not_8  g05679(new_n6055, new_n6056);
xor_4  g05680(new_n6056, new_n6052, new_n6057);
and_5  g05681(new_n6041, new_n3706, new_n6058);
nor_5  g05682(new_n6041, new_n3706, new_n6059);
nor_5  g05683(new_n6059, new_n6040, new_n6060);
or_5   g05684(new_n6060, new_n6058, new_n6061);
not_8  g05685(new_n6061, new_n6062);
xor_4  g05686(new_n6062, new_n6057, new_n6063);
not_8  g05687(new_n6063, new_n6064);
xor_4  g05688(new_n6064, new_n6051, new_n6065);
nand_5 g05689(n11662, n6687, new_n6066);
not_8  g05690(new_n3720, new_n6067);
nor_5  g05691(new_n6067, new_n3714, new_n6068);
nor_5  g05692(new_n6068, new_n3712, new_n6069);
and_5  g05693(new_n6069, new_n6066, new_n6070);
xor_4  g05694(new_n6044, new_n6038_1, new_n6071);
not_8  g05695(new_n6071, new_n6072);
not_8  g05696(new_n6066, new_n6073);
xor_4  g05697(new_n6069, new_n6073, new_n6074);
not_8  g05698(new_n6074, new_n6075);
and_5  g05699(new_n6075, new_n6072, new_n6076);
or_5   g05700(new_n6076, new_n6070, new_n6077);
not_8  g05701(new_n6077, new_n6078);
nand_5 g05702(new_n6078, new_n6065, new_n6079);
nor_5  g05703(new_n6056, new_n6052, new_n6080);
and_5  g05704(new_n6062, new_n6057, new_n6081);
or_5   g05705(new_n6081, new_n6080, new_n6082);
nand_5 g05706(n10327, n2564, new_n6083);
not_8  g05707(new_n6083, new_n6084);
nand_5 g05708(n11662, n4189, new_n6085);
nand_5 g05709(n9583, n6687, new_n6086);
xor_4  g05710(new_n6086, new_n6085, new_n6087);
not_8  g05711(new_n6087, new_n6088);
xor_4  g05712(new_n6088, new_n6084, new_n6089_1);
not_8  g05713(new_n6089_1, new_n6090);
xor_4  g05714(new_n6090, new_n6082, new_n6091);
or_5   g05715(new_n6054, new_n6053, new_n6092);
nand_5 g05716(n7456, n6770, new_n6093);
not_8  g05717(new_n6093, new_n6094);
xor_4  g05718(new_n6094, new_n6092, new_n6095);
nand_5 g05719(n3932, n3627, new_n6096);
nand_5 g05720(n12591, n9920, new_n6097);
nand_5 g05721(n4516, n1798, new_n6098);
xor_4  g05722(new_n6098, new_n6097, new_n6099);
xor_4  g05723(new_n6099, new_n6096, new_n6100);
xor_4  g05724(new_n6100, new_n6095, new_n6101);
xor_4  g05725(new_n6101, new_n6091, new_n6102);
not_8  g05726(new_n6102, new_n6103);
and_5  g05727(new_n6049, new_n6046, new_n6104);
or_5   g05728(new_n6048, new_n6047, new_n6105);
or_5   g05729(new_n6064, new_n6051, new_n6106);
xor_4  g05730(new_n6106, new_n6105, new_n6107);
nor_5  g05731(new_n6107, new_n6104, new_n6108);
xor_4  g05732(new_n6108, new_n6103, new_n6109);
not_8  g05733(new_n6109, new_n6110);
xor_4  g05734(new_n6110, new_n6079, new_n6111);
not_8  g05735(new_n6111, new_n6112);
nand_5 g05736(n10327, n6687, new_n6113);
not_8  g05737(new_n6113, new_n6114);
xor_4  g05738(new_n6078, new_n6065, new_n6115);
and_5  g05739(new_n6115, new_n6114, new_n6116);
or_5   g05740(new_n3727, new_n3721, new_n6117);
xor_4  g05741(new_n6075, new_n6072, new_n6118);
or_5   g05742(new_n6118, new_n6117, new_n6119);
xor_4  g05743(new_n6115, new_n6114, new_n6120);
not_8  g05744(new_n6120, new_n6121);
nor_5  g05745(new_n6121, new_n6119, new_n6122);
nor_5  g05746(new_n6122, new_n6116, new_n6123);
xor_4  g05747(new_n6123, new_n6112, new_n6124);
nand_5 g05748(n3022, n2226, new_n6125);
nand_5 g05749(n9640, n1094, new_n6126_1);
nand_5 g05750(n10678, n6703, new_n6127);
xor_4  g05751(new_n6127, new_n6126_1, new_n6128);
not_8  g05752(new_n6128, new_n6129);
xor_4  g05753(new_n6129, new_n6125, new_n6130);
nand_5 g05754(n6703, n1094, new_n6131);
and_5  g05755(new_n6131, new_n3764, new_n6132);
nor_5  g05756(new_n6131, new_n3764, new_n6133);
nand_5 g05757(n9640, n2226, new_n6134);
not_8  g05758(new_n6134, new_n6135);
nor_5  g05759(new_n6135, new_n6133, new_n6136);
or_5   g05760(new_n6136, new_n6132, new_n6137);
not_8  g05761(new_n6137, new_n6138);
xor_4  g05762(new_n6138, new_n6130, new_n6139);
nand_5 g05763(n10928, n10451, new_n6140);
nand_5 g05764(n11023, n6986, new_n6141);
xor_4  g05765(new_n6141, new_n6140, new_n6142);
xor_4  g05766(new_n6142, new_n6139, new_n6143);
nand_5 g05767(n11023, n10928, new_n6144);
and_5  g05768(new_n3877, new_n3876, new_n6145);
nor_5  g05769(new_n3877, new_n3876, new_n6146);
nor_5  g05770(new_n6146, new_n3875, new_n6147);
nor_5  g05771(new_n6147, new_n6145, new_n6148);
not_8  g05772(new_n6148, new_n6149);
nor_5  g05773(new_n6149, new_n6144, new_n6150);
not_8  g05774(new_n6144, new_n6151);
xor_4  g05775(new_n6149, new_n6151, new_n6152);
xor_4  g05776(new_n6131, new_n3764, new_n6153);
xor_4  g05777(new_n6153, new_n6134, new_n6154);
nor_5  g05778(new_n6154, new_n6152, new_n6155);
or_5   g05779(new_n6155, new_n6150, new_n6156);
xnor_4 g05780(new_n6156, new_n6143, new_n6157);
nand_5 g05781(n10451, n8336, new_n6158);
not_8  g05782(new_n6158, new_n6159);
xor_4  g05783(new_n6154, new_n6152, new_n6160);
and_5  g05784(new_n6160, new_n6159, new_n6161);
nor_5  g05785(new_n3872, new_n3867, new_n6162);
nor_5  g05786(new_n3880, new_n3873, new_n6163);
or_5   g05787(new_n6163, new_n6162, new_n6164);
xor_4  g05788(new_n6160, new_n6159, new_n6165);
and_5  g05789(new_n6165, new_n6164, new_n6166);
nor_5  g05790(new_n6166, new_n6161, new_n6167);
or_5   g05791(new_n6167, new_n6157, new_n6168);
not_8  g05792(new_n6168, new_n6169);
nor_5  g05793(new_n6129, new_n6125, new_n6170);
and_5  g05794(new_n6138, new_n6130, new_n6171);
or_5   g05795(new_n6171, new_n6170, new_n6172);
nand_5 g05796(n10928, n10278, new_n6173);
not_8  g05797(new_n6173, new_n6174);
nand_5 g05798(n10451, n6986, new_n6175);
nand_5 g05799(n11423, n8336, new_n6176);
xor_4  g05800(new_n6176, new_n6175, new_n6177);
not_8  g05801(new_n6177, new_n6178);
xor_4  g05802(new_n6178, new_n6174, new_n6179);
not_8  g05803(new_n6179, new_n6180);
xor_4  g05804(new_n6180, new_n6172, new_n6181);
or_5   g05805(new_n6127, new_n6126_1, new_n6182);
not_8  g05806(new_n6182, new_n6183);
nand_5 g05807(n11023, n2226, new_n6184);
not_8  g05808(new_n6184, new_n6185);
xor_4  g05809(new_n6185, new_n6183, new_n6186);
nand_5 g05810(n10678, n9640, new_n6187);
nand_5 g05811(n3022, n1094, new_n6188);
nand_5 g05812(n7320, n6703, new_n6189);
xor_4  g05813(new_n6189, new_n6188, new_n6190);
not_8  g05814(new_n6190, new_n6191);
xor_4  g05815(new_n6191, new_n6187, new_n6192_1);
xor_4  g05816(new_n6192_1, new_n6186, new_n6193);
xor_4  g05817(new_n6193, new_n6181, new_n6194);
not_8  g05818(new_n6194, new_n6195);
and_5  g05819(new_n6142, new_n6139, new_n6196);
or_5   g05820(new_n6141, new_n6140, new_n6197);
not_8  g05821(new_n6197, new_n6198);
nand_5 g05822(new_n6156, new_n6143, new_n6199);
not_8  g05823(new_n6199, new_n6200);
xor_4  g05824(new_n6200, new_n6198, new_n6201);
nor_5  g05825(new_n6201, new_n6196, new_n6202);
xor_4  g05826(new_n6202, new_n6195, new_n6203);
not_8  g05827(new_n6203, new_n6204);
xor_4  g05828(new_n6204, new_n6169, new_n6205);
nand_5 g05829(n10278, n8336, new_n6206);
not_8  g05830(new_n6206, new_n6207);
xor_4  g05831(new_n6167, new_n6157, new_n6208);
nor_5  g05832(new_n6208, new_n6207, new_n6209);
not_8  g05833(new_n3882, new_n6210);
nand_5 g05834(new_n6210, new_n3881, new_n6211);
xor_4  g05835(new_n6165, new_n6164, new_n6212);
not_8  g05836(new_n6212, new_n6213);
or_5   g05837(new_n6213, new_n6211, new_n6214);
not_8  g05838(new_n6214, new_n6215);
xor_4  g05839(new_n6208, new_n6207, new_n6216);
not_8  g05840(new_n6216, new_n6217);
nor_5  g05841(new_n6217, new_n6215, new_n6218);
or_5   g05842(new_n6218, new_n6209, new_n6219);
xor_4  g05843(new_n6219, new_n6205, new_n6220);
not_8  g05844(new_n6220, new_n6221);
nand_5 g05845(n8665, n7160, new_n6222);
nand_5 g05846(n4828, n1067, new_n6223);
nand_5 g05847(n5645, n2515, new_n6224);
xor_4  g05848(new_n6224, new_n6223, new_n6225);
not_8  g05849(new_n6225, new_n6226);
xor_4  g05850(new_n6226, new_n6222, new_n6227);
nand_5 g05851(n5645, n4828, new_n6228);
nand_5 g05852(n8665, n7891, new_n6229);
and_5  g05853(new_n6229, new_n6228, new_n6230);
nand_5 g05854(n7160, n1067, new_n6231);
not_8  g05855(new_n6231, new_n6232);
xor_4  g05856(new_n6229, new_n6228, new_n6233);
not_8  g05857(new_n6233, new_n6234);
nor_5  g05858(new_n6234, new_n6232, new_n6235);
or_5   g05859(new_n6235, new_n6230, new_n6236);
not_8  g05860(new_n6236, new_n6237);
xor_4  g05861(new_n6237, new_n6227, new_n6238);
nand_5 g05862(n12391, n2551, new_n6239);
nand_5 g05863(n11922, n7891, new_n6240);
xor_4  g05864(new_n6240, new_n6239, new_n6241);
xor_4  g05865(new_n6241, new_n6238, new_n6242);
nand_5 g05866(n12391, n11922, new_n6243);
nand_5 g05867(n12391, n8665, new_n6244);
and_5  g05868(new_n6244, new_n3835, new_n6245);
and_5  g05869(new_n3838, new_n3834, new_n6246);
nor_5  g05870(new_n6246, new_n6245, new_n6247);
not_8  g05871(new_n6247, new_n6248);
nor_5  g05872(new_n6248, new_n6243, new_n6249);
xor_4  g05873(new_n6234, new_n6232, new_n6250);
not_8  g05874(new_n6250, new_n6251);
xor_4  g05875(new_n6248, new_n6243, new_n6252);
and_5  g05876(new_n6252, new_n6251, new_n6253);
nor_5  g05877(new_n6253, new_n6249, new_n6254_1);
xor_4  g05878(new_n6254_1, new_n6242, new_n6255);
nand_5 g05879(n12069, n2551, new_n6256);
xor_4  g05880(new_n6252, new_n6251, new_n6257);
not_8  g05881(new_n6257, new_n6258);
nor_5  g05882(new_n6258, new_n6256, new_n6259);
and_5  g05883(new_n6258, new_n6256, new_n6260);
nor_5  g05884(new_n3831, new_n3825, new_n6261);
nor_5  g05885(new_n3839, new_n3832, new_n6262);
nor_5  g05886(new_n6262, new_n6261, new_n6263);
nor_5  g05887(new_n6263, new_n6260, new_n6264);
nor_5  g05888(new_n6264, new_n6259, new_n6265);
or_5   g05889(new_n6265, new_n6255, new_n6266);
not_8  g05890(new_n6266, new_n6267);
nor_5  g05891(new_n6226, new_n6222, new_n6268);
and_5  g05892(new_n6237, new_n6227, new_n6269);
or_5   g05893(new_n6269, new_n6268, new_n6270);
not_8  g05894(new_n6270, new_n6271);
nand_5 g05895(n12826, n12391, new_n6272);
not_8  g05896(new_n6272, new_n6273_1);
nand_5 g05897(n7891, n2551, new_n6274);
nand_5 g05898(n12069, n4094, new_n6275);
xor_4  g05899(new_n6275, new_n6274, new_n6276);
not_8  g05900(new_n6276, new_n6277);
xor_4  g05901(new_n6277, new_n6273_1, new_n6278);
xor_4  g05902(new_n6278, new_n6271, new_n6279);
or_5   g05903(new_n6224, new_n6223, new_n6280);
not_8  g05904(new_n6280, new_n6281);
nand_5 g05905(n11922, n7160, new_n6282);
not_8  g05906(new_n6282, new_n6283);
xor_4  g05907(new_n6283, new_n6281, new_n6284);
and_5  g05908(n2515, n1067, new_n6285);
nand_5 g05909(n8665, n4828, new_n6286);
nand_5 g05910(n5645, n1199, new_n6287);
xor_4  g05911(new_n6287, new_n6286, new_n6288);
xor_4  g05912(new_n6288, new_n6285, new_n6289);
xor_4  g05913(new_n6289, new_n6284, new_n6290);
xor_4  g05914(new_n6290, new_n6279, new_n6291);
not_8  g05915(new_n6291, new_n6292);
and_5  g05916(new_n6241, new_n6238, new_n6293);
or_5   g05917(new_n6240, new_n6239, new_n6294_1);
not_8  g05918(new_n6294_1, new_n6295);
not_8  g05919(new_n6242, new_n6296);
or_5   g05920(new_n6254_1, new_n6296, new_n6297);
not_8  g05921(new_n6297, new_n6298);
xor_4  g05922(new_n6298, new_n6295, new_n6299);
nor_5  g05923(new_n6299, new_n6293, new_n6300);
xor_4  g05924(new_n6300, new_n6292, new_n6301);
not_8  g05925(new_n6301, new_n6302);
xor_4  g05926(new_n6302, new_n6267, new_n6303);
nand_5 g05927(n12826, n12069, new_n6304);
not_8  g05928(new_n6304, new_n6305);
xor_4  g05929(new_n6265, new_n6255, new_n6306);
nor_5  g05930(new_n6306, new_n6305, new_n6307);
or_5   g05931(new_n3841, new_n3823, new_n6308);
xor_4  g05932(new_n6258, new_n6256, new_n6309);
xor_4  g05933(new_n6309, new_n6263, new_n6310);
or_5   g05934(new_n6310, new_n6308, new_n6311);
not_8  g05935(new_n6311, new_n6312);
xor_4  g05936(new_n6306, new_n6305, new_n6313);
not_8  g05937(new_n6313, new_n6314);
nor_5  g05938(new_n6314, new_n6312, new_n6315);
or_5   g05939(new_n6315, new_n6307, new_n6316);
xor_4  g05940(new_n6316, new_n6303, new_n6317);
not_8  g05941(new_n6317, new_n6318);
nand_5 g05942(n3754, n996, new_n6319);
nand_5 g05943(n10898, n5767, new_n6320);
nand_5 g05944(n11876, n5319, new_n6321);
xor_4  g05945(new_n6321, new_n6320, new_n6322);
not_8  g05946(new_n6322, new_n6323);
xor_4  g05947(new_n6323, new_n6319, new_n6324);
nand_5 g05948(n10898, n996, new_n6325);
and_5  g05949(new_n6325, new_n3794, new_n6326);
nand_5 g05950(n11876, n5767, new_n6327);
not_8  g05951(new_n6327, new_n6328);
xor_4  g05952(new_n6325, new_n3794, new_n6329);
not_8  g05953(new_n6329, new_n6330);
nor_5  g05954(new_n6330, new_n6328, new_n6331);
or_5   g05955(new_n6331, new_n6326, new_n6332);
not_8  g05956(new_n6332, new_n6333);
xor_4  g05957(new_n6333, new_n6324, new_n6334);
nand_5 g05958(n11153, n159, new_n6335);
nand_5 g05959(n5314, n2749, new_n6336);
xor_4  g05960(new_n6336, new_n6335, new_n6337);
xor_4  g05961(new_n6337, new_n6334, new_n6338);
nand_5 g05962(n11153, n2749, new_n6339);
nand_5 g05963(n11876, n996, new_n6340);
and_5  g05964(new_n6340, new_n3851, new_n6341);
and_5  g05965(new_n3854, new_n3850, new_n6342);
nor_5  g05966(new_n6342, new_n6341, new_n6343);
not_8  g05967(new_n6343, new_n6344);
nor_5  g05968(new_n6344, new_n6339, new_n6345);
not_8  g05969(new_n6339, new_n6346);
xor_4  g05970(new_n6344, new_n6346, new_n6347);
xor_4  g05971(new_n6330, new_n6328, new_n6348);
nor_5  g05972(new_n6348, new_n6347, new_n6349);
nor_5  g05973(new_n6349, new_n6345, new_n6350);
xor_4  g05974(new_n6350, new_n6338, new_n6351);
nand_5 g05975(n11222, n159, new_n6352);
xor_4  g05976(new_n6348, new_n6347, new_n6353);
not_8  g05977(new_n6353, new_n6354);
nor_5  g05978(new_n6354, new_n6352, new_n6355);
nand_5 g05979(new_n6354, new_n6352, new_n6356);
not_8  g05980(new_n3843, new_n6357);
and_5  g05981(new_n3847, new_n6357, new_n6358_1);
nor_5  g05982(new_n3855, new_n3848, new_n6359_1);
nor_5  g05983(new_n6359_1, new_n6358_1, new_n6360);
not_8  g05984(new_n6360, new_n6361);
and_5  g05985(new_n6361, new_n6356, new_n6362);
nor_5  g05986(new_n6362, new_n6355, new_n6363);
or_5   g05987(new_n6363, new_n6351, new_n6364);
not_8  g05988(new_n6364, new_n6365);
and_5  g05989(new_n6337, new_n6334, new_n6366);
or_5   g05990(new_n6336, new_n6335, new_n6367);
not_8  g05991(new_n6367, new_n6368);
not_8  g05992(new_n6338, new_n6369);
or_5   g05993(new_n6350, new_n6369, new_n6370);
not_8  g05994(new_n6370, new_n6371);
xor_4  g05995(new_n6371, new_n6368, new_n6372);
or_5   g05996(new_n6372, new_n6366, new_n6373);
nor_5  g05997(new_n6323, new_n6319, new_n6374);
and_5  g05998(new_n6333, new_n6324, new_n6375);
or_5   g05999(new_n6375, new_n6374, new_n6376);
not_8  g06000(new_n6376, new_n6377);
nand_5 g06001(n11153, n1510, new_n6378);
not_8  g06002(new_n6378, new_n6379);
nand_5 g06003(n5314, n159, new_n6380);
nand_5 g06004(n12247, n11222, new_n6381);
xor_4  g06005(new_n6381, new_n6380, new_n6382);
not_8  g06006(new_n6382, new_n6383);
xor_4  g06007(new_n6383, new_n6379, new_n6384);
xor_4  g06008(new_n6384, new_n6377, new_n6385);
or_5   g06009(new_n6321, new_n6320, new_n6386);
not_8  g06010(new_n6386, new_n6387);
nand_5 g06011(n2749, n996, new_n6388);
not_8  g06012(new_n6388, new_n6389);
xor_4  g06013(new_n6389, new_n6387, new_n6390);
nand_5 g06014(n10898, n5319, new_n6391);
nand_5 g06015(n11876, n9457, new_n6392);
nand_5 g06016(n5767, n3754, new_n6393);
xor_4  g06017(new_n6393, new_n6392, new_n6394);
not_8  g06018(new_n6394, new_n6395);
xor_4  g06019(new_n6395, new_n6391, new_n6396);
xor_4  g06020(new_n6396, new_n6390, new_n6397);
xor_4  g06021(new_n6397, new_n6385, new_n6398);
xor_4  g06022(new_n6398, new_n6373, new_n6399);
not_8  g06023(new_n6399, new_n6400);
xor_4  g06024(new_n6400, new_n6365, new_n6401);
nand_5 g06025(n11222, n1510, new_n6402);
not_8  g06026(new_n6402, new_n6403);
xor_4  g06027(new_n6363, new_n6351, new_n6404);
nor_5  g06028(new_n6404, new_n6403, new_n6405);
nand_5 g06029(new_n3857, new_n3856, new_n6406);
not_8  g06030(new_n6352, new_n6407);
xor_4  g06031(new_n6354, new_n6407, new_n6408);
xor_4  g06032(new_n6408, new_n6361, new_n6409);
or_5   g06033(new_n6409, new_n6406, new_n6410);
not_8  g06034(new_n6410, new_n6411);
xor_4  g06035(new_n6404, new_n6403, new_n6412);
not_8  g06036(new_n6412, new_n6413);
nor_5  g06037(new_n6413, new_n6411, new_n6414);
or_5   g06038(new_n6414, new_n6405, new_n6415);
xor_4  g06039(new_n6415, new_n6401, new_n6416);
and_5  g06040(new_n6413, new_n6411, new_n6417);
or_5   g06041(new_n6417, new_n6414, new_n6418);
and_5  g06042(new_n6314, new_n6312, new_n6419);
or_5   g06043(new_n6419, new_n6315, new_n6420);
and_5  g06044(new_n6420, new_n6418, new_n6421);
nor_5  g06045(new_n6420, new_n6418, new_n6422);
xor_4  g06046(new_n6310, new_n6308, new_n6423);
and_5  g06047(new_n3858, new_n3842_1, new_n6424);
nor_5  g06048(new_n3864, new_n3860, new_n6425);
nor_5  g06049(new_n6425, new_n6424, new_n6426);
nor_5  g06050(new_n6426, new_n6423, new_n6427);
xor_4  g06051(new_n6409, new_n6406, new_n6428);
xor_4  g06052(new_n6426, new_n6423, new_n6429_1);
not_8  g06053(new_n6429_1, new_n6430);
nor_5  g06054(new_n6430, new_n6428, new_n6431_1);
or_5   g06055(new_n6431_1, new_n6427, new_n6432);
nor_5  g06056(new_n6432, new_n6422, new_n6433);
nor_5  g06057(new_n6433, new_n6421, new_n6434);
not_8  g06058(new_n6434, new_n6435);
xor_4  g06059(new_n6435, new_n6416, new_n6436);
xor_4  g06060(new_n6436, new_n6318, new_n6437);
xor_4  g06061(new_n6437, new_n6221, new_n6438);
and_5  g06062(new_n6217, new_n6215, new_n6439);
or_5   g06063(new_n6439, new_n6218, new_n6440);
not_8  g06064(new_n6440, new_n6441_1);
not_8  g06065(new_n6211, new_n6442);
xor_4  g06066(new_n6213, new_n6442, new_n6443);
xor_4  g06067(new_n6430, new_n6428, new_n6444);
nor_5  g06068(new_n6444, new_n6443, new_n6445_1);
and_5  g06069(new_n3888, new_n3884, new_n6446);
and_5  g06070(new_n3889, new_n3866, new_n6447);
or_5   g06071(new_n6447, new_n6446, new_n6448);
xor_4  g06072(new_n6444, new_n6443, new_n6449);
and_5  g06073(new_n6449, new_n6448, new_n6450);
nor_5  g06074(new_n6450, new_n6445_1, new_n6451);
nor_5  g06075(new_n6451, new_n6441_1, new_n6452);
xor_4  g06076(new_n6451, new_n6441_1, new_n6453);
not_8  g06077(new_n6453, new_n6454);
xnor_4 g06078(new_n6420, new_n6418, new_n6455);
xor_4  g06079(new_n6455, new_n6432, new_n6456);
not_8  g06080(new_n6456, new_n6457);
nor_5  g06081(new_n6457, new_n6454, new_n6458);
or_5   g06082(new_n6458, new_n6452, new_n6459);
xor_4  g06083(new_n6459, new_n6438, new_n6460);
not_8  g06084(new_n6460, new_n6461);
xor_4  g06085(new_n6461, new_n6124, new_n6462);
xor_4  g06086(new_n6121, new_n6119, new_n6463);
xor_4  g06087(new_n6457, new_n6454, new_n6464);
and_5  g06088(new_n6464, new_n6463, new_n6465);
or_5   g06089(new_n6464, new_n6463, new_n6466);
xor_4  g06090(new_n6118, new_n6117, new_n6467);
xor_4  g06091(new_n6449, new_n6448, new_n6468);
nor_5  g06092(new_n6468, new_n6467, new_n6469);
nor_5  g06093(new_n3820, new_n3729, new_n6470);
not_8  g06094(new_n3890, new_n6471);
nor_5  g06095(new_n6471, new_n3822, new_n6472);
nor_5  g06096(new_n6472, new_n6470, new_n6473);
not_8  g06097(new_n6467, new_n6474);
xor_4  g06098(new_n6468, new_n6474, new_n6475);
not_8  g06099(new_n6475, new_n6476);
and_5  g06100(new_n6476, new_n6473, new_n6477);
or_5   g06101(new_n6477, new_n6469, new_n6478);
not_8  g06102(new_n6478, new_n6479);
and_5  g06103(new_n6479, new_n6466, new_n6480);
nor_5  g06104(new_n6480, new_n6465, new_n6481);
xor_4  g06105(new_n6481, new_n6462, n2301);
xor_4  g06106(new_n3818, new_n3817, n2316);
nand_5 g06107(n4634, n1333, new_n6484);
not_8  g06108(new_n6484, new_n6485);
and_5  g06109(new_n5819, new_n5818, new_n6486);
nor_5  g06110(new_n5819, new_n5818, new_n6487);
nor_5  g06111(new_n6487, new_n5817, new_n6488);
or_5   g06112(new_n6488, new_n6486, new_n6489);
not_8  g06113(new_n6489, new_n6490);
and_5  g06114(new_n6490, new_n6485, new_n6491);
nor_5  g06115(new_n6490, new_n6485, new_n6492);
or_5   g06116(new_n6492, new_n6491, new_n6493);
nand_5 g06117(n11757, n2879, new_n6494);
not_8  g06118(new_n6494, new_n6495);
nand_5 g06119(n7265, n5240, new_n6496);
xor_4  g06120(new_n6496, new_n5808, new_n6497);
xor_4  g06121(new_n6497, new_n6495, new_n6498);
not_8  g06122(new_n6498, new_n6499);
nor_5  g06123(new_n6499, new_n6493, new_n6500);
or_5   g06124(new_n6500, new_n6491, new_n6501);
not_8  g06125(new_n6501, new_n6502);
nand_5 g06126(n4634, n3172, new_n6503);
nand_5 g06127(n9195, n1333, new_n6504);
xor_4  g06128(new_n6504, new_n6503, new_n6505);
not_8  g06129(new_n6505, new_n6506);
xor_4  g06130(new_n6506, new_n6502, new_n6507);
nand_5 g06131(n11757, n10223, new_n6508);
not_8  g06132(new_n6508, new_n6509);
nand_5 g06133(n5240, n2879, new_n6510);
nand_5 g06134(n11821, n7265, new_n6511);
xor_4  g06135(new_n6511, new_n6510, new_n6512);
xor_4  g06136(new_n6512, new_n6509, new_n6513);
and_5  g06137(new_n6496, new_n5808, new_n6514);
nor_5  g06138(new_n6496, new_n5808, new_n6515);
nor_5  g06139(new_n6515, new_n6495, new_n6516);
nor_5  g06140(new_n6516, new_n6514, new_n6517);
xor_4  g06141(new_n6517, new_n6513, new_n6518);
xor_4  g06142(new_n6518, new_n6507, new_n6519);
nand_5 g06143(n9195, n7862, new_n6520);
not_8  g06144(new_n6520, new_n6521);
xor_4  g06145(new_n6499, new_n6493, new_n6522);
and_5  g06146(new_n6522, new_n6521, new_n6523);
and_5  g06147(new_n5814_1, new_n5802, new_n6524);
and_5  g06148(new_n5821, new_n5815, new_n6525);
or_5   g06149(new_n6525, new_n6524, new_n6526);
not_8  g06150(new_n6526, new_n6527);
xor_4  g06151(new_n6522, new_n6521, new_n6528);
not_8  g06152(new_n6528, new_n6529);
nor_5  g06153(new_n6529, new_n6527, new_n6530);
or_5   g06154(new_n6530, new_n6523, new_n6531);
nand_5 g06155(new_n6531, new_n6519, new_n6532);
nor_5  g06156(new_n6512, new_n6509, new_n6533);
not_8  g06157(new_n6513, new_n6534);
nor_5  g06158(new_n6517, new_n6534, new_n6535);
or_5   g06159(new_n6535, new_n6533, new_n6536);
not_8  g06160(new_n6536, new_n6537);
nand_5 g06161(n2253, n1333, new_n6538);
nand_5 g06162(n9195, n3172, new_n6539);
nand_5 g06163(n7862, n3865, new_n6540);
xor_4  g06164(new_n6540, new_n6539, new_n6541);
xor_4  g06165(new_n6541, new_n6538, new_n6542);
not_8  g06166(new_n6542, new_n6543);
nor_5  g06167(new_n6543, new_n6537, new_n6544);
and_5  g06168(new_n6543, new_n6537, new_n6545);
or_5   g06169(new_n6545, new_n6544, new_n6546);
or_5   g06170(new_n6511, new_n6510, new_n6547);
not_8  g06171(new_n6547, new_n6548);
and_5  g06172(n11757, n4634, new_n6549);
xor_4  g06173(new_n6549, new_n6548, new_n6550);
nand_5 g06174(n11821, n2879, new_n6551);
not_8  g06175(new_n6551, new_n6552);
nand_5 g06176(n10223, n5240, new_n6553);
nand_5 g06177(n9080, n7265, new_n6554);
xor_4  g06178(new_n6554, new_n6553, new_n6555);
not_8  g06179(new_n6555, new_n6556);
xor_4  g06180(new_n6556, new_n6552, new_n6557);
xor_4  g06181(new_n6557, new_n6550, new_n6558);
not_8  g06182(new_n6558, new_n6559);
xor_4  g06183(new_n6559, new_n6546, new_n6560);
nor_5  g06184(new_n6506, new_n6502, new_n6561);
or_5   g06185(new_n6504, new_n6503, new_n6562);
not_8  g06186(new_n6562, new_n6563);
and_5  g06187(new_n6518, new_n6507, new_n6564);
xor_4  g06188(new_n6564, new_n6563, new_n6565);
nor_5  g06189(new_n6565, new_n6561, new_n6566);
xor_4  g06190(new_n6566, new_n6560, new_n6567);
not_8  g06191(new_n6567, new_n6568);
nor_5  g06192(new_n6568, new_n6532, new_n6569);
and_5  g06193(new_n6568, new_n6532, new_n6570);
or_5   g06194(new_n6570, new_n6569, new_n6571);
nand_5 g06195(n7862, n2253, new_n6572);
xor_4  g06196(new_n6531, new_n6519, new_n6573);
not_8  g06197(new_n6573, new_n6574);
nor_5  g06198(new_n6574, new_n6572, new_n6575);
not_8  g06199(new_n5828, new_n6576);
nand_5 g06200(new_n6576, new_n5822, new_n6577);
not_8  g06201(new_n6577, new_n6578_1);
xor_4  g06202(new_n6529, new_n6527, new_n6579);
nand_5 g06203(new_n6579, new_n6578_1, new_n6580);
not_8  g06204(new_n6580, new_n6581);
xor_4  g06205(new_n6574, new_n6572, new_n6582);
and_5  g06206(new_n6582, new_n6581, new_n6583);
nor_5  g06207(new_n6583, new_n6575, new_n6584);
xor_4  g06208(new_n6584, new_n6571, new_n6585);
xor_4  g06209(new_n6582, new_n6581, new_n6586);
xor_4  g06210(new_n6579, new_n6578_1, new_n6587);
not_8  g06211(new_n5858, new_n6588);
nand_5 g06212(new_n6588, new_n5851, new_n6589);
not_8  g06213(new_n6589, new_n6590);
nand_5 g06214(n12145, n6877, new_n6591);
nand_5 g06215(n9400, n2522, new_n6592);
and_5  g06216(n11311, n2024, new_n6593);
nand_5 g06217(n7946, n4187, new_n6594);
xor_4  g06218(new_n6594, new_n5844, new_n6595);
xor_4  g06219(new_n6595, new_n6593, new_n6596);
xor_4  g06220(new_n6596, new_n6592, new_n6597);
and_5  g06221(new_n5835, new_n5834, new_n6598);
nor_5  g06222(new_n5837, new_n5833, new_n6599);
nor_5  g06223(new_n6599, new_n6598, new_n6600);
xor_4  g06224(new_n6600, new_n6597, new_n6601);
xor_4  g06225(new_n6601, new_n6591, new_n6602);
not_8  g06226(new_n6602, new_n6603);
nor_5  g06227(new_n5838, new_n5831, new_n6604_1);
and_5  g06228(new_n5850, new_n5839, new_n6605);
nor_5  g06229(new_n6605, new_n6604_1, new_n6606);
xor_4  g06230(new_n6606, new_n6603, new_n6607);
xor_4  g06231(new_n6607, new_n6590, new_n6608);
and_5  g06232(new_n5920, new_n5860_1, new_n6609);
xor_4  g06233(new_n5963, new_n5943, new_n6610);
xor_4  g06234(new_n5968, new_n6610, new_n6611_1);
and_5  g06235(new_n6611_1, new_n5921, new_n6612);
nor_5  g06236(new_n6612, new_n6609, new_n6613);
not_8  g06237(new_n6613, new_n6614);
xor_4  g06238(new_n6614, new_n6608, new_n6615);
or_5   g06239(new_n5940, new_n5938, new_n6616);
not_8  g06240(new_n6616, new_n6617);
nand_5 g06241(n11478, n521, new_n6618);
not_8  g06242(new_n6618, new_n6619);
and_5  g06243(new_n5935, new_n5934_1, new_n6620);
nor_5  g06244(new_n5935, new_n5934_1, new_n6621);
nor_5  g06245(new_n6621, new_n5933, new_n6622);
or_5   g06246(new_n6622, new_n6620, new_n6623);
not_8  g06247(new_n6623, new_n6624);
and_5  g06248(new_n6624, new_n6619, new_n6625);
nor_5  g06249(new_n6624, new_n6619, new_n6626);
or_5   g06250(new_n6626, new_n6625, new_n6627);
nand_5 g06251(n2498, n137, new_n6628);
not_8  g06252(new_n6628, new_n6629);
nand_5 g06253(n5579, n5283, new_n6630);
nand_5 g06254(n6294, n2558, new_n6631);
xor_4  g06255(new_n6631, new_n6630, new_n6632);
xor_4  g06256(new_n6632, new_n6629, new_n6633);
not_8  g06257(new_n6633, new_n6634);
xor_4  g06258(new_n6634, new_n6627, new_n6635);
not_8  g06259(new_n6635, new_n6636);
nand_5 g06260(n6016, n4805, new_n6637);
not_8  g06261(new_n6637, new_n6638);
not_8  g06262(new_n5937, new_n6639);
nor_5  g06263(new_n6639, new_n5931, new_n6640);
nor_5  g06264(new_n6640, new_n5929, new_n6641);
not_8  g06265(new_n6641, new_n6642);
xor_4  g06266(new_n6642, new_n6638, new_n6643);
xor_4  g06267(new_n6643, new_n6636, new_n6644);
xor_4  g06268(new_n6644, new_n6617, new_n6645_1);
not_8  g06269(new_n6645_1, new_n6646);
and_5  g06270(new_n5962, new_n5959, new_n6647);
not_8  g06271(new_n6647, new_n6648);
and_5  g06272(n7270, n7236, new_n6649);
nor_5  g06273(new_n5949, new_n5944, new_n6650);
nor_5  g06274(new_n5958, new_n5951, new_n6651);
or_5   g06275(new_n6651, new_n6650, new_n6652);
not_8  g06276(new_n6652, new_n6653);
xor_4  g06277(new_n6653, new_n6649, new_n6654);
and_5  g06278(n3992, n806, new_n6655);
and_5  g06279(new_n5955, new_n5954, new_n6656);
nor_5  g06280(new_n5955, new_n5954, new_n6657);
nor_5  g06281(new_n6657, new_n5953, new_n6658);
or_5   g06282(new_n6658, new_n6656, new_n6659);
not_8  g06283(new_n6659, new_n6660);
and_5  g06284(new_n6660, new_n6655, new_n6661);
nor_5  g06285(new_n6660, new_n6655, new_n6662);
or_5   g06286(new_n6662, new_n6661, new_n6663);
nand_5 g06287(n9111, n6358, new_n6664);
not_8  g06288(new_n6664, new_n6665);
nand_5 g06289(n8384, n3342, new_n6666);
nand_5 g06290(n9763, n5198, new_n6667);
xor_4  g06291(new_n6667, new_n6666, new_n6668);
not_8  g06292(new_n6668, new_n6669);
xor_4  g06293(new_n6669, new_n6665, new_n6670);
xor_4  g06294(new_n6670, new_n6663, new_n6671);
xor_4  g06295(new_n6671, new_n6654, new_n6672);
xor_4  g06296(new_n6672, new_n6648, new_n6673);
xor_4  g06297(new_n6673, new_n6646, new_n6674);
nor_5  g06298(new_n5963, new_n5943, new_n6675);
nor_5  g06299(new_n5968, new_n5964_1, new_n6676);
or_5   g06300(new_n6676, new_n6675, new_n6677);
xor_4  g06301(new_n6677, new_n6674, new_n6678);
xor_4  g06302(new_n6678, new_n6615, new_n6679);
not_8  g06303(new_n6679, new_n6680);
nor_5  g06304(new_n6680, new_n6587, new_n6681);
xor_4  g06305(new_n6679, new_n6587, new_n6682);
not_8  g06306(new_n6682, new_n6683);
and_5  g06307(new_n5970, new_n5829, new_n6684);
nor_5  g06308(new_n5970, new_n5829, new_n6685);
nor_5  g06309(new_n5991, new_n6685, new_n6686);
or_5   g06310(new_n6686, new_n6684, new_n6687_1);
and_5  g06311(new_n6687_1, new_n6683, new_n6688);
nor_5  g06312(new_n6688, new_n6681, new_n6689_1);
or_5   g06313(new_n6689_1, new_n6586, new_n6690);
or_5   g06314(new_n6614, new_n6608, new_n6691);
not_8  g06315(new_n6691, new_n6692);
and_5  g06316(new_n6678, new_n6615, new_n6693);
nor_5  g06317(new_n6693, new_n6692, new_n6694);
nand_5 g06318(new_n6607, new_n6590, new_n6695);
nand_5 g06319(n12221, n6877, new_n6696);
nor_5  g06320(new_n6601, new_n6591, new_n6697);
nor_5  g06321(new_n6606, new_n6603, new_n6698);
or_5   g06322(new_n6698, new_n6697, new_n6699);
not_8  g06323(new_n6699, new_n6700);
not_8  g06324(new_n6592, new_n6701);
nor_5  g06325(new_n6596, new_n6701, new_n6702);
nor_5  g06326(new_n6600, new_n6597, new_n6703_1);
or_5   g06327(new_n6703_1, new_n6702, new_n6704);
not_8  g06328(new_n6704, new_n6705);
nand_5 g06329(n11311, n9189, new_n6706);
not_8  g06330(new_n6706, new_n6707);
nand_5 g06331(n7946, n4203, new_n6708);
nand_5 g06332(n4187, n2024, new_n6709);
xor_4  g06333(new_n6709, new_n6708, new_n6710);
xor_4  g06334(new_n6710, new_n6707, new_n6711);
not_8  g06335(new_n6711, new_n6712);
and_5  g06336(new_n6594, new_n5844, new_n6713);
nor_5  g06337(new_n6594, new_n5844, new_n6714);
nor_5  g06338(new_n6714, new_n6593, new_n6715);
nor_5  g06339(new_n6715, new_n6713, new_n6716);
xor_4  g06340(new_n6716, new_n6712, new_n6717);
not_8  g06341(new_n6717, new_n6718);
nand_5 g06342(n12145, n9400, new_n6719);
nand_5 g06343(n2522, n2464, new_n6720);
xor_4  g06344(new_n6720, new_n6719, new_n6721);
xor_4  g06345(new_n6721, new_n6718, new_n6722);
xor_4  g06346(new_n6722, new_n6705, new_n6723);
xor_4  g06347(new_n6723, new_n6700, new_n6724);
xor_4  g06348(new_n6724, new_n6696, new_n6725);
not_8  g06349(new_n6725, new_n6726);
xor_4  g06350(new_n6726, new_n6695, new_n6727);
xor_4  g06351(new_n6727, new_n6694, new_n6728);
or_5   g06352(new_n6672, new_n6648, new_n6729);
nand_5 g06353(n7236, n5153, new_n6730);
not_8  g06354(new_n6730, new_n6731);
nand_5 g06355(n6358, n3342, new_n6732);
nand_5 g06356(n9111, n5198, new_n6733);
nand_5 g06357(n9763, n1471, new_n6734);
xor_4  g06358(new_n6734, new_n6733, new_n6735);
not_8  g06359(new_n6735, new_n6736);
xor_4  g06360(new_n6736, new_n6732, new_n6737);
and_5  g06361(new_n6667, new_n6666, new_n6738);
nor_5  g06362(new_n6669, new_n6665, new_n6739);
or_5   g06363(new_n6739, new_n6738, new_n6740);
not_8  g06364(new_n6740, new_n6741);
xor_4  g06365(new_n6741, new_n6737, new_n6742_1);
nand_5 g06366(n7270, n3992, new_n6743);
nand_5 g06367(n8384, n806, new_n6744);
xor_4  g06368(new_n6744, new_n6743, new_n6745);
xor_4  g06369(new_n6745, new_n6742_1, new_n6746);
not_8  g06370(new_n6746, new_n6747);
nor_5  g06371(new_n6670, new_n6663, new_n6748);
nor_5  g06372(new_n6748, new_n6661, new_n6749);
xor_4  g06373(new_n6749, new_n6747, new_n6750);
not_8  g06374(new_n6750, new_n6751);
nand_5 g06375(n7270, n7236, new_n6752);
and_5  g06376(new_n6653, new_n6752, new_n6753);
nor_5  g06377(new_n6671, new_n6654, new_n6754);
nor_5  g06378(new_n6754, new_n6753, new_n6755);
not_8  g06379(new_n6755, new_n6756);
xor_4  g06380(new_n6756, new_n6751, new_n6757);
xor_4  g06381(new_n6757, new_n6731, new_n6758);
xor_4  g06382(new_n6758, new_n6729, new_n6759);
or_5   g06383(new_n6644, new_n6616, new_n6760);
nand_5 g06384(n5798, n4805, new_n6761);
not_8  g06385(new_n6761, new_n6762);
nand_5 g06386(n5579, n137, new_n6763);
nand_5 g06387(n6797, n2558, new_n6764);
nand_5 g06388(n6294, n2498, new_n6765);
xor_4  g06389(new_n6765, new_n6764, new_n6766);
not_8  g06390(new_n6766, new_n6767);
xor_4  g06391(new_n6767, new_n6763, new_n6768);
and_5  g06392(new_n6631, new_n6630, new_n6769);
nor_5  g06393(new_n6631, new_n6630, new_n6770_1);
nor_5  g06394(new_n6770_1, new_n6629, new_n6771);
or_5   g06395(new_n6771, new_n6769, new_n6772);
not_8  g06396(new_n6772, new_n6773);
xor_4  g06397(new_n6773, new_n6768, new_n6774);
nand_5 g06398(n11478, n6016, new_n6775);
nand_5 g06399(n5283, n521, new_n6776_1);
xor_4  g06400(new_n6776_1, new_n6775, new_n6777);
xor_4  g06401(new_n6777, new_n6774, new_n6778);
not_8  g06402(new_n6778, new_n6779);
nor_5  g06403(new_n6634, new_n6627, new_n6780);
nor_5  g06404(new_n6780, new_n6625, new_n6781);
xor_4  g06405(new_n6781, new_n6779, new_n6782);
not_8  g06406(new_n6782, new_n6783);
nor_5  g06407(new_n6642, new_n6638, new_n6784);
and_5  g06408(new_n6643, new_n6636, new_n6785);
nor_5  g06409(new_n6785, new_n6784, new_n6786);
not_8  g06410(new_n6786, new_n6787);
xor_4  g06411(new_n6787, new_n6783, new_n6788);
xor_4  g06412(new_n6788, new_n6762, new_n6789);
xor_4  g06413(new_n6789, new_n6760, new_n6790);
not_8  g06414(new_n6790, new_n6791);
xor_4  g06415(new_n6791, new_n6759, new_n6792);
nor_5  g06416(new_n6673, new_n6646, new_n6793);
and_5  g06417(new_n6677, new_n6674, new_n6794);
nor_5  g06418(new_n6794, new_n6793, new_n6795);
xor_4  g06419(new_n6795, new_n6792, new_n6796);
xor_4  g06420(new_n6796, new_n6728, new_n6797_1);
not_8  g06421(new_n6586, new_n6798);
xor_4  g06422(new_n6689_1, new_n6798, new_n6799);
not_8  g06423(new_n6799, new_n6800);
nand_5 g06424(new_n6800, new_n6797_1, new_n6801);
and_5  g06425(new_n6801, new_n6690, new_n6802);
nor_5  g06426(new_n6802, new_n6585, new_n6803);
not_8  g06427(new_n6585, new_n6804);
xor_4  g06428(new_n6802, new_n6804, new_n6805);
not_8  g06429(new_n6805, new_n6806_1);
not_8  g06430(new_n6723, new_n6807);
or_5   g06431(new_n6807, new_n6700, new_n6808);
nor_5  g06432(new_n6710, new_n6707, new_n6809_1);
nor_5  g06433(new_n6716, new_n6712, new_n6810);
or_5   g06434(new_n6810, new_n6809_1, new_n6811);
not_8  g06435(new_n6811, new_n6812);
nand_5 g06436(n12221, n9400, new_n6813);
not_8  g06437(new_n6813, new_n6814);
nand_5 g06438(n12145, n2464, new_n6815);
nand_5 g06439(n10217, n6877, new_n6816);
xor_4  g06440(new_n6816, new_n6815, new_n6817);
not_8  g06441(new_n6817, new_n6818);
xor_4  g06442(new_n6818, new_n6814, new_n6819);
not_8  g06443(new_n6819, new_n6820);
nor_5  g06444(new_n6820, new_n6812, new_n6821);
and_5  g06445(new_n6820, new_n6812, new_n6822_1);
or_5   g06446(new_n6822_1, new_n6821, new_n6823);
or_5   g06447(new_n6709, new_n6708, new_n6824);
nand_5 g06448(n11311, n2522, new_n6825);
not_8  g06449(new_n6825, new_n6826_1);
xor_4  g06450(new_n6826_1, new_n6824, new_n6827);
nand_5 g06451(n4203, n2024, new_n6828);
nand_5 g06452(n9189, n4187, new_n6829);
nand_5 g06453(n12753, n7946, new_n6830);
xor_4  g06454(new_n6830, new_n6829, new_n6831);
xor_4  g06455(new_n6831, new_n6828, new_n6832);
xor_4  g06456(new_n6832, new_n6827, new_n6833);
xor_4  g06457(new_n6833, new_n6823, new_n6834);
and_5  g06458(new_n6721, new_n6718, new_n6835);
or_5   g06459(new_n6720, new_n6719, new_n6836);
or_5   g06460(new_n6721, new_n6718, new_n6837);
nand_5 g06461(new_n6837, new_n6705, new_n6838);
xor_4  g06462(new_n6838, new_n6836, new_n6839);
nor_5  g06463(new_n6839, new_n6835, new_n6840);
xor_4  g06464(new_n6840, new_n6834, new_n6841);
not_8  g06465(new_n6841, new_n6842);
xor_4  g06466(new_n6842, new_n6808, new_n6843);
not_8  g06467(new_n6843, new_n6844);
nor_5  g06468(new_n6724, new_n6696, new_n6845);
nor_5  g06469(new_n6726, new_n6695, new_n6846);
nor_5  g06470(new_n6846, new_n6845, new_n6847);
xor_4  g06471(new_n6847, new_n6844, new_n6848);
not_8  g06472(new_n6848, new_n6849);
or_5   g06473(new_n6787, new_n6783, new_n6850);
nand_5 g06474(n4805, n2347, new_n6851);
not_8  g06475(new_n6851, new_n6852);
nand_5 g06476(n6016, n5283, new_n6853);
nand_5 g06477(n11478, n5798, new_n6854);
xor_4  g06478(new_n6854, new_n6853, new_n6855);
not_8  g06479(new_n6855, new_n6856);
xor_4  g06480(new_n6856, new_n6852, new_n6857);
not_8  g06481(new_n6857, new_n6858);
nor_5  g06482(new_n6767, new_n6763, new_n6859);
and_5  g06483(new_n6773, new_n6768, new_n6860_1);
or_5   g06484(new_n6860_1, new_n6859, new_n6861);
xor_4  g06485(new_n6861, new_n6858, new_n6862);
or_5   g06486(new_n6765, new_n6764, new_n6863);
not_8  g06487(new_n6863, new_n6864);
nand_5 g06488(n521, n137, new_n6865);
not_8  g06489(new_n6865, new_n6866);
xor_4  g06490(new_n6866, new_n6864, new_n6867);
nand_5 g06491(n6797, n2498, new_n6868);
nand_5 g06492(n6294, n5579, new_n6869);
nand_5 g06493(n3146, n2558, new_n6870);
xor_4  g06494(new_n6870, new_n6869, new_n6871);
not_8  g06495(new_n6871, new_n6872);
xor_4  g06496(new_n6872, new_n6868, new_n6873);
xor_4  g06497(new_n6873, new_n6867, new_n6874);
xor_4  g06498(new_n6874, new_n6862, new_n6875);
not_8  g06499(new_n6875, new_n6876);
nand_5 g06500(new_n6777, new_n6774, new_n6877_1);
or_5   g06501(new_n6776_1, new_n6775, new_n6878);
or_5   g06502(new_n6781, new_n6779, new_n6879);
not_8  g06503(new_n6879, new_n6880);
xor_4  g06504(new_n6880, new_n6878, new_n6881);
and_5  g06505(new_n6881, new_n6877_1, new_n6882);
xor_4  g06506(new_n6882, new_n6876, new_n6883);
xnor_4 g06507(new_n6883, new_n6850, new_n6884);
not_8  g06508(new_n6884, new_n6885);
and_5  g06509(new_n6788, new_n6762, new_n6886);
nor_5  g06510(new_n6788, new_n6762, new_n6887);
nor_5  g06511(new_n6887, new_n6760, new_n6888);
nor_5  g06512(new_n6888, new_n6886, new_n6889);
xor_4  g06513(new_n6889, new_n6885, new_n6890);
not_8  g06514(new_n6890, new_n6891);
or_5   g06515(new_n6756, new_n6751, new_n6892);
and_5  g06516(new_n6745, new_n6742_1, new_n6893);
or_5   g06517(new_n6744, new_n6743, new_n6894);
not_8  g06518(new_n6894, new_n6895);
or_5   g06519(new_n6749, new_n6747, new_n6896);
not_8  g06520(new_n6896, new_n6897);
xor_4  g06521(new_n6897, new_n6895, new_n6898);
or_5   g06522(new_n6898, new_n6893, new_n6899);
or_5   g06523(new_n6734, new_n6733, new_n6900);
not_8  g06524(new_n6900, new_n6901);
nand_5 g06525(n6358, n806, new_n6902);
not_8  g06526(new_n6902, new_n6903);
xor_4  g06527(new_n6903, new_n6901, new_n6904);
nand_5 g06528(n9111, n1471, new_n6905);
not_8  g06529(new_n6905, new_n6906);
nand_5 g06530(n5198, n3342, new_n6907);
nand_5 g06531(n9763, n7646, new_n6908);
xor_4  g06532(new_n6908, new_n6907, new_n6909);
xor_4  g06533(new_n6909, new_n6906, new_n6910);
xor_4  g06534(new_n6910, new_n6904, new_n6911);
nor_5  g06535(new_n6736, new_n6732, new_n6912);
and_5  g06536(new_n6741, new_n6737, new_n6913);
or_5   g06537(new_n6913, new_n6912, new_n6914);
not_8  g06538(new_n6914, new_n6915);
nand_5 g06539(n5153, n3992, new_n6916);
not_8  g06540(new_n6916, new_n6917);
nand_5 g06541(n8384, n7270, new_n6918);
nand_5 g06542(n7236, n2507, new_n6919);
xor_4  g06543(new_n6919, new_n6918, new_n6920);
not_8  g06544(new_n6920, new_n6921);
xor_4  g06545(new_n6921, new_n6917, new_n6922);
xor_4  g06546(new_n6922, new_n6915, new_n6923);
xor_4  g06547(new_n6923, new_n6911, new_n6924);
xor_4  g06548(new_n6924, new_n6899, new_n6925);
not_8  g06549(new_n6925, new_n6926);
xor_4  g06550(new_n6926, new_n6892, new_n6927);
nor_5  g06551(new_n6757, new_n6731, new_n6928);
nor_5  g06552(new_n6672, new_n6648, new_n6929);
and_5  g06553(new_n6757, new_n6731, new_n6930);
nor_5  g06554(new_n6930, new_n6929, new_n6931);
or_5   g06555(new_n6931, new_n6928, new_n6932);
not_8  g06556(new_n6932, new_n6933);
xor_4  g06557(new_n6933, new_n6927, new_n6934);
xor_4  g06558(new_n6934, new_n6891, new_n6935);
xor_4  g06559(new_n6758, new_n6929, new_n6936);
nor_5  g06560(new_n6791, new_n6936, new_n6937);
nor_5  g06561(new_n6795, new_n6792, new_n6938);
nor_5  g06562(new_n6938, new_n6937, new_n6939);
xor_4  g06563(new_n6939, new_n6935, new_n6940);
xor_4  g06564(new_n6940, new_n6849, new_n6941);
not_8  g06565(new_n6941, new_n6942);
or_5   g06566(new_n6693, new_n6692, new_n6943);
not_8  g06567(new_n6727, new_n6944);
nor_5  g06568(new_n6944, new_n6943, new_n6945);
xor_4  g06569(new_n6727, new_n6943, new_n6946);
nor_5  g06570(new_n6796, new_n6946, new_n6947);
nor_5  g06571(new_n6947, new_n6945, new_n6948);
xor_4  g06572(new_n6948, new_n6942, new_n6949);
not_8  g06573(new_n6949, new_n6950);
and_5  g06574(new_n6950, new_n6806_1, new_n6951);
or_5   g06575(new_n6951, new_n6803, new_n6952);
nor_5  g06576(new_n6940, new_n6849, new_n6953);
nor_5  g06577(new_n6948, new_n6942, new_n6954);
nor_5  g06578(new_n6954, new_n6953, new_n6955);
nand_5 g06579(n4805, n1576, new_n6956);
not_8  g06580(new_n6878, new_n6957);
nand_5 g06581(new_n6880, new_n6957, new_n6958);
not_8  g06582(new_n6958, new_n6959);
nor_5  g06583(new_n6882, new_n6876, new_n6960);
nor_5  g06584(new_n6960, new_n6959, new_n6961);
xor_4  g06585(new_n6961, new_n6956, new_n6962);
xor_4  g06586(new_n6962, new_n6955, new_n6963);
nor_5  g06587(new_n6842, new_n6808, new_n6964);
nor_5  g06588(new_n6847, new_n6844, new_n6965);
nor_5  g06589(new_n6965, new_n6964, new_n6966);
nor_5  g06590(new_n6926, new_n6892, new_n6967);
and_5  g06591(new_n6933, new_n6927, new_n6968);
nor_5  g06592(new_n6968, new_n6967, new_n6969);
nor_5  g06593(new_n6833, new_n6823, new_n6970);
or_5   g06594(new_n6970, new_n6821, new_n6971);
and_5  g06595(n9189, n4203, new_n6972);
and_5  g06596(n4187, n2522, new_n6973);
xor_4  g06597(new_n6973, new_n6972, new_n6974);
and_5  g06598(n9763, n4722, new_n6975);
and_5  g06599(n10217, n9400, new_n6976);
xor_4  g06600(new_n6976, new_n6975, new_n6977);
xor_4  g06601(new_n6977, new_n6974, new_n6978);
nand_5 g06602(n9111, n7646, new_n6979);
nand_5 g06603(n12221, n2464, new_n6980);
and_5  g06604(n12145, n11311, new_n6981);
xor_4  g06605(new_n6981, new_n6980, new_n6982);
xor_4  g06606(new_n6982, new_n6979, new_n6983);
xor_4  g06607(new_n6983, new_n6978, new_n6984);
xor_4  g06608(new_n6984, new_n6971, new_n6985);
xor_4  g06609(new_n6985, new_n6969, new_n6986_1);
xor_4  g06610(new_n6986_1, new_n6966, new_n6987);
nor_5  g06611(new_n6838, new_n6836, new_n6988);
nor_5  g06612(new_n6840, new_n6834, new_n6989);
nor_5  g06613(new_n6989, new_n6988, new_n6990);
and_5  g06614(new_n6897, new_n6895, new_n6991);
and_5  g06615(new_n6924, new_n6899, new_n6992);
nor_5  g06616(new_n6992, new_n6991, new_n6993);
xor_4  g06617(new_n6993, new_n6990, new_n6994);
nand_5 g06618(n11821, n10223, new_n6995);
and_5  g06619(n9080, n2879, new_n6996);
xor_4  g06620(new_n6996, new_n6995, new_n6997);
nand_5 g06621(n11757, n9195, new_n6998);
and_5  g06622(n7862, n2512, new_n6999);
xor_4  g06623(new_n6999, new_n6998, new_n7000);
xor_4  g06624(new_n7000, new_n6997, new_n7001);
nor_5  g06625(new_n6540, new_n6539, new_n7002);
and_5  g06626(new_n6540, new_n6539, new_n7003);
nor_5  g06627(new_n7003, new_n6538, new_n7004);
nor_5  g06628(new_n7004, new_n7002, new_n7005);
xor_4  g06629(new_n7005, new_n7001, new_n7006);
nand_5 g06630(n12753, n2024, new_n7007);
nand_5 g06631(n3865, n1333, new_n7008);
and_5  g06632(n5240, n4634, new_n7009);
xor_4  g06633(new_n7009, new_n7008, new_n7010);
xor_4  g06634(new_n7010, new_n7007, new_n7011);
xor_4  g06635(new_n7011, new_n7006, new_n7012);
xor_4  g06636(new_n7012, new_n6994, new_n7013);
and_5  g06637(new_n6564, new_n6563, new_n7014);
nor_5  g06638(new_n6566, new_n6560, new_n7015);
nor_5  g06639(new_n7015, new_n7014, new_n7016);
nor_5  g06640(new_n6559, new_n6546, new_n7017);
nor_5  g06641(new_n7017, new_n6544, new_n7018);
nor_5  g06642(new_n6825, new_n6824, new_n7019);
nor_5  g06643(new_n6832, new_n6827, new_n7020);
or_5   g06644(new_n7020, new_n7019, new_n7021);
and_5  g06645(n8384, n5153, new_n7022);
and_5  g06646(n7270, n6358, new_n7023);
xor_4  g06647(new_n7023, new_n7022, new_n7024);
nor_5  g06648(new_n6830, new_n6829, new_n7025);
and_5  g06649(new_n6830, new_n6829, new_n7026);
nor_5  g06650(new_n7026, new_n6828, new_n7027);
nor_5  g06651(new_n7027, new_n7025, new_n7028);
xor_4  g06652(new_n7028, new_n7024, new_n7029);
xor_4  g06653(new_n7029, new_n7021, new_n7030);
xor_4  g06654(new_n7030, new_n7018, new_n7031);
and_5  g06655(n5198, n806, new_n7032);
and_5  g06656(n3992, n2507, new_n7033);
xor_4  g06657(new_n7033, new_n7032, new_n7034);
nand_5 g06658(n7823, n6877, new_n7035);
and_5  g06659(n3342, n1471, new_n7036);
xor_4  g06660(new_n7036, new_n7035, new_n7037);
xor_4  g06661(new_n7037, new_n7034, new_n7038);
nor_5  g06662(new_n6908, new_n6907, new_n7039);
and_5  g06663(new_n6908, new_n6907, new_n7040);
nor_5  g06664(new_n7040, new_n6905, new_n7041);
nor_5  g06665(new_n7041, new_n7039, new_n7042);
xor_4  g06666(new_n7042, new_n7038, new_n7043);
xor_4  g06667(new_n7043, new_n7031, new_n7044);
and_5  g06668(new_n6922, new_n6915, new_n7045);
not_8  g06669(new_n6911, new_n7046);
and_5  g06670(new_n6923, new_n7046, new_n7047);
or_5   g06671(new_n7047, new_n7045, new_n7048);
and_5  g06672(new_n6816, new_n6815, new_n7049);
nor_5  g06673(new_n6818, new_n6814, new_n7050);
nor_5  g06674(new_n7050, new_n7049, new_n7051);
nand_5 g06675(n7236, n6431, new_n7052);
and_5  g06676(n10174, n7946, new_n7053);
xor_4  g06677(new_n7053, new_n7052, new_n7054);
xor_4  g06678(new_n7054, new_n7051, new_n7055);
xor_4  g06679(new_n7055, new_n7048, new_n7056);
xor_4  g06680(new_n7056, new_n7044, new_n7057);
xor_4  g06681(new_n7057, new_n7016, new_n7058);
xor_4  g06682(new_n7058, new_n7013, new_n7059);
xor_4  g06683(new_n7059, new_n6987, new_n7060);
not_8  g06684(new_n6934, new_n7061);
and_5  g06685(new_n7061, new_n6891, new_n7062);
nor_5  g06686(new_n6939, new_n6935, new_n7063);
nor_5  g06687(new_n7063, new_n7062, new_n7064);
nor_5  g06688(new_n6584, new_n6571, new_n7065);
nor_5  g06689(new_n7065, new_n6569, new_n7066);
not_8  g06690(new_n6883, new_n7067);
nor_5  g06691(new_n7067, new_n6850, new_n7068);
nor_5  g06692(new_n6889, new_n6885, new_n7069);
or_5   g06693(new_n7069, new_n7068, new_n7070);
and_5  g06694(new_n6903, new_n6901, new_n7071);
and_5  g06695(new_n6910, new_n6904, new_n7072);
nor_5  g06696(new_n7072, new_n7071, new_n7073);
and_5  g06697(new_n6866, new_n6864, new_n7074);
and_5  g06698(new_n6873, new_n6867, new_n7075);
nor_5  g06699(new_n7075, new_n7074, new_n7076);
xor_4  g06700(new_n7076, new_n7073, new_n7077);
nor_5  g06701(new_n6549, new_n6548, new_n7078);
and_5  g06702(new_n6557, new_n6550, new_n7079);
or_5   g06703(new_n7079, new_n7078, new_n7080);
nand_5 g06704(n3172, n2253, new_n7081);
and_5  g06705(n6797, n5579, new_n7082);
and_5  g06706(n5798, n5283, new_n7083);
xor_4  g06707(new_n7083, new_n7082, new_n7084);
xor_4  g06708(new_n7084, new_n7081, new_n7085);
xor_4  g06709(new_n7085, new_n7080, new_n7086);
and_5  g06710(new_n6854, new_n6853, new_n7087);
nor_5  g06711(new_n6856, new_n6852, new_n7088);
nor_5  g06712(new_n7088, new_n7087, new_n7089);
and_5  g06713(new_n6870, new_n6869, new_n7090);
not_8  g06714(new_n6868, new_n7091);
nor_5  g06715(new_n6872, new_n7091, new_n7092);
nor_5  g06716(new_n7092, new_n7090, new_n7093);
xor_4  g06717(new_n7093, new_n7089, new_n7094);
nand_5 g06718(n11478, n2347, new_n7095);
and_5  g06719(n3146, n2498, new_n7096);
xor_4  g06720(new_n7096, new_n7095, new_n7097);
xor_4  g06721(new_n7097, new_n7094, new_n7098);
xor_4  g06722(new_n7098, new_n7086, new_n7099);
xor_4  g06723(new_n7099, new_n7077, new_n7100);
or_5   g06724(new_n6861, new_n6858, new_n7101);
not_8  g06725(new_n6874, new_n7102);
nand_5 g06726(new_n7102, new_n6862, new_n7103);
and_5  g06727(new_n7103, new_n7101, new_n7104);
and_5  g06728(new_n6554, new_n6553, new_n7105);
nor_5  g06729(new_n6556, new_n6552, new_n7106);
nor_5  g06730(new_n7106, new_n7105, new_n7107);
and_5  g06731(n6016, n137, new_n7108);
nand_5 g06732(n7265, n6826, new_n7109);
and_5  g06733(n6294, n521, new_n7110);
xor_4  g06734(new_n7110, new_n7109, new_n7111);
xor_4  g06735(new_n7111, new_n7108, new_n7112);
xor_4  g06736(new_n7112, new_n7107, new_n7113);
nand_5 g06737(n4938, n2558, new_n7114);
and_5  g06738(new_n6919, new_n6918, new_n7115);
nor_5  g06739(new_n6921, new_n6917, new_n7116);
nor_5  g06740(new_n7116, new_n7115, new_n7117);
xor_4  g06741(new_n7117, new_n7114, new_n7118);
xor_4  g06742(new_n7118, new_n7113, new_n7119);
xor_4  g06743(new_n7119, new_n7104, new_n7120);
xor_4  g06744(new_n7120, new_n7100, new_n7121);
xor_4  g06745(new_n7121, new_n7070, new_n7122);
xor_4  g06746(new_n7122, new_n7066, new_n7123);
xor_4  g06747(new_n7123, new_n7064, new_n7124);
xor_4  g06748(new_n7124, new_n7060, new_n7125);
xor_4  g06749(new_n7125, new_n6963, new_n7126);
xor_4  g06750(new_n7126, new_n6952, n2383);
xor_4  g06751(new_n5789, new_n5781, n2425);
xor_4  g06752(new_n2877, new_n2830, n2431);
xor_4  g06753(new_n2049, new_n2046, n2434);
xor_4  g06754(new_n4841, new_n4840, n2581);
xor_4  g06755(new_n6464, new_n6463, new_n7132);
xor_4  g06756(new_n7132, new_n6479, n2624);
nand_5 g06757(n11917, n6770, new_n7134);
not_8  g06758(new_n7134, new_n7135);
nand_5 g06759(n9920, n4921, new_n7136);
nand_5 g06760(n9956, n3627, new_n7137);
xor_4  g06761(new_n7137, new_n7136, new_n7138);
xor_4  g06762(new_n7138, new_n7135, new_n7139);
not_8  g06763(new_n7139, new_n7140);
and_5  g06764(new_n3940, new_n3898, new_n7141);
nor_5  g06765(new_n3942, new_n3939, new_n7142);
nor_5  g06766(new_n7142, new_n7141, new_n7143);
xor_4  g06767(new_n7143, new_n7140, new_n7144);
nand_5 g06768(n2577, n2564, new_n7145);
nand_5 g06769(n4189, n3842, new_n7146);
xor_4  g06770(new_n7146, new_n7145, new_n7147);
xor_4  g06771(new_n7147, new_n7144, new_n7148);
nor_5  g06772(new_n3943, new_n3937, new_n7149);
nor_5  g06773(new_n7149, new_n3935, new_n7150);
xor_4  g06774(new_n7150, new_n7148, new_n7151);
not_8  g06775(new_n7151, new_n7152);
nor_5  g06776(new_n3925, new_n3922, new_n7153);
nor_5  g06777(new_n3945, new_n3927, new_n7154);
nor_5  g06778(new_n7154, new_n7153, new_n7155);
or_5   g06779(new_n7155, new_n7152, new_n7156);
not_8  g06780(new_n7156, new_n7157);
or_5   g06781(new_n7137, new_n7136, new_n7158);
not_8  g06782(new_n7158, new_n7159_1);
and_5  g06783(n6770, n3842, new_n7160_1);
xor_4  g06784(new_n7160_1, new_n7159_1, new_n7161);
nand_5 g06785(n4921, n3627, new_n7162);
not_8  g06786(new_n7162, new_n7163);
nand_5 g06787(n11917, n9920, new_n7164);
nand_5 g06788(n9956, n4516, new_n7165);
xor_4  g06789(new_n7165, new_n7164, new_n7166);
not_8  g06790(new_n7166, new_n7167);
xor_4  g06791(new_n7167, new_n7163, new_n7168);
xor_4  g06792(new_n7168, new_n7161, new_n7169);
not_8  g06793(new_n7169, new_n7170);
nor_5  g06794(new_n7138, new_n7135, new_n7171);
nor_5  g06795(new_n7143, new_n7140, new_n7172);
or_5   g06796(new_n7172, new_n7171, new_n7173);
not_8  g06797(new_n7173, new_n7174);
nand_5 g06798(n9637, n2564, new_n7175);
nand_5 g06799(n4189, n2577, new_n7176);
nand_5 g06800(n6687, n1835, new_n7177);
xor_4  g06801(new_n7177, new_n7176, new_n7178);
not_8  g06802(new_n7178, new_n7179);
xor_4  g06803(new_n7179, new_n7175, new_n7180);
xor_4  g06804(new_n7180, new_n7174, new_n7181);
xor_4  g06805(new_n7181, new_n7170, new_n7182);
not_8  g06806(new_n7182, new_n7183);
not_8  g06807(new_n7147, new_n7184);
or_5   g06808(new_n7184, new_n7144, new_n7185);
or_5   g06809(new_n7146, new_n7145, new_n7186);
or_5   g06810(new_n7150, new_n7148, new_n7187);
not_8  g06811(new_n7187, new_n7188);
xor_4  g06812(new_n7188, new_n7186, new_n7189);
and_5  g06813(new_n7189, new_n7185, new_n7190);
xor_4  g06814(new_n7190, new_n7183, new_n7191);
xor_4  g06815(new_n7191, new_n7157, new_n7192);
not_8  g06816(new_n7192, new_n7193_1);
nand_5 g06817(n9637, n6687, new_n7194);
xor_4  g06818(new_n7155, new_n7152, new_n7195);
not_8  g06819(new_n7195, new_n7196);
nor_5  g06820(new_n7196, new_n7194, new_n7197);
nand_5 g06821(new_n3946, new_n3921, new_n7198);
not_8  g06822(new_n7198, new_n7199);
xor_4  g06823(new_n7196, new_n7194, new_n7200);
and_5  g06824(new_n7200, new_n7199, new_n7201);
nor_5  g06825(new_n7201, new_n7197, new_n7202);
xor_4  g06826(new_n7202, new_n7193_1, new_n7203);
not_8  g06827(new_n7203, new_n7204);
nand_5 g06828(n6126, n2226, new_n7205);
not_8  g06829(new_n7205, new_n7206);
nand_5 g06830(n3602, n1094, new_n7207);
nand_5 g06831(n10678, n3719, new_n7208);
xor_4  g06832(new_n7208, new_n7207, new_n7209);
xor_4  g06833(new_n7209, new_n7206, new_n7210);
not_8  g06834(new_n7210, new_n7211);
and_5  g06835(new_n4134, new_n3956, new_n7212);
nor_5  g06836(new_n4136, new_n4133, new_n7213);
nor_5  g06837(new_n7213, new_n7212, new_n7214);
xor_4  g06838(new_n7214, new_n7211, new_n7215);
nand_5 g06839(n10928, n10439, new_n7216);
nand_5 g06840(n8595, n6986, new_n7217);
xor_4  g06841(new_n7217, new_n7216, new_n7218);
xor_4  g06842(new_n7218, new_n7215, new_n7219);
not_8  g06843(new_n7219, new_n7220);
nor_5  g06844(new_n4137, new_n4131, new_n7221);
nor_5  g06845(new_n7221, new_n4129, new_n7222);
xor_4  g06846(new_n7222, new_n7220, new_n7223);
nor_5  g06847(new_n4119, new_n4116, new_n7224);
nor_5  g06848(new_n4139, new_n4121, new_n7225);
nor_5  g06849(new_n7225, new_n7224, new_n7226);
or_5   g06850(new_n7226, new_n7223, new_n7227);
not_8  g06851(new_n7227, new_n7228);
nor_5  g06852(new_n7209, new_n7206, new_n7229);
nor_5  g06853(new_n7214, new_n7211, new_n7230);
or_5   g06854(new_n7230, new_n7229, new_n7231);
not_8  g06855(new_n7231, new_n7232);
nand_5 g06856(n10928, n8065, new_n7233);
not_8  g06857(new_n7233, new_n7234);
nand_5 g06858(n10439, n6986, new_n7235);
nand_5 g06859(n10391, n8336, new_n7236_1);
xor_4  g06860(new_n7236_1, new_n7235, new_n7237);
not_8  g06861(new_n7237, new_n7238);
xor_4  g06862(new_n7238, new_n7234, new_n7239);
not_8  g06863(new_n7239, new_n7240);
xor_4  g06864(new_n7240, new_n7232, new_n7241);
or_5   g06865(new_n7208, new_n7207, new_n7242);
not_8  g06866(new_n7242, new_n7243);
nand_5 g06867(n8595, n2226, new_n7244);
not_8  g06868(new_n7244, new_n7245);
xor_4  g06869(new_n7245, new_n7243, new_n7246);
nand_5 g06870(n10678, n3602, new_n7247);
nand_5 g06871(n6126, n1094, new_n7248);
nand_5 g06872(n7320, n3719, new_n7249);
xor_4  g06873(new_n7249, new_n7248, new_n7250);
not_8  g06874(new_n7250, new_n7251);
xor_4  g06875(new_n7251, new_n7247, new_n7252);
xor_4  g06876(new_n7252, new_n7246, new_n7253);
xor_4  g06877(new_n7253, new_n7241, new_n7254);
not_8  g06878(new_n7254, new_n7255);
not_8  g06879(new_n7218, new_n7256);
or_5   g06880(new_n7256, new_n7215, new_n7257);
or_5   g06881(new_n7217, new_n7216, new_n7258);
or_5   g06882(new_n7222, new_n7219, new_n7259);
not_8  g06883(new_n7259, new_n7260);
xor_4  g06884(new_n7260, new_n7258, new_n7261);
and_5  g06885(new_n7261, new_n7257, new_n7262);
xor_4  g06886(new_n7262, new_n7255, new_n7263);
xor_4  g06887(new_n7263, new_n7228, new_n7264);
nand_5 g06888(n8336, n8065, new_n7265_1);
not_8  g06889(new_n7265_1, new_n7266);
xor_4  g06890(new_n7226, new_n7223, new_n7267);
nor_5  g06891(new_n7267, new_n7266, new_n7268);
nand_5 g06892(new_n4140, new_n4115, new_n7269);
not_8  g06893(new_n7269, new_n7270_1);
xor_4  g06894(new_n7267, new_n7266, new_n7271);
not_8  g06895(new_n7271, new_n7272);
nor_5  g06896(new_n7272, new_n7270_1, new_n7273);
or_5   g06897(new_n7273, new_n7268, new_n7274);
xor_4  g06898(new_n7274, new_n7264, new_n7275);
nand_5 g06899(n7160, n4826, new_n7276);
nand_5 g06900(n7733, n4828, new_n7277);
nand_5 g06901(n12925, n2515, new_n7278);
xor_4  g06902(new_n7278, new_n7277, new_n7279);
not_8  g06903(new_n7279, new_n7280);
xor_4  g06904(new_n7280, new_n7276, new_n7281);
and_5  g06905(new_n4181, new_n3987, new_n7282);
not_8  g06906(new_n4180, new_n7283);
nor_5  g06907(new_n4183, new_n7283, new_n7284);
or_5   g06908(new_n7284, new_n7282, new_n7285);
not_8  g06909(new_n7285, new_n7286);
xor_4  g06910(new_n7286, new_n7281, new_n7287);
nand_5 g06911(n12391, n4970, new_n7288);
nand_5 g06912(n7891, n7610, new_n7289);
xor_4  g06913(new_n7289, new_n7288, new_n7290);
xor_4  g06914(new_n7290, new_n7287, new_n7291);
not_8  g06915(new_n7291, new_n7292);
and_5  g06916(new_n4178, new_n4174, new_n7293);
and_5  g06917(new_n4184, new_n4179, new_n7294_1);
nor_5  g06918(new_n7294_1, new_n7293, new_n7295);
xor_4  g06919(new_n7295, new_n7292, new_n7296);
not_8  g06920(new_n7296, new_n7297);
nor_5  g06921(new_n4186, new_n4172, new_n7298);
and_5  g06922(new_n4190_1, new_n4187_1, new_n7299);
nor_5  g06923(new_n7299, new_n7298, new_n7300);
or_5   g06924(new_n7300, new_n7297, new_n7301);
nor_5  g06925(new_n7280, new_n7276, new_n7302);
and_5  g06926(new_n7286, new_n7281, new_n7303);
or_5   g06927(new_n7303, new_n7302, new_n7304);
not_8  g06928(new_n7304, new_n7305);
nand_5 g06929(n12391, n503, new_n7306);
not_8  g06930(new_n7306, new_n7307);
nand_5 g06931(n7891, n4970, new_n7308);
nand_5 g06932(n12069, n10965, new_n7309);
xor_4  g06933(new_n7309, new_n7308, new_n7310);
not_8  g06934(new_n7310, new_n7311);
xor_4  g06935(new_n7311, new_n7307, new_n7312);
xor_4  g06936(new_n7312, new_n7305, new_n7313);
or_5   g06937(new_n7278, new_n7277, new_n7314);
not_8  g06938(new_n7314, new_n7315);
nand_5 g06939(n7610, n7160, new_n7316);
not_8  g06940(new_n7316, new_n7317);
xor_4  g06941(new_n7317, new_n7315, new_n7318);
nand_5 g06942(n7733, n2515, new_n7319);
nand_5 g06943(n4828, n4826, new_n7320_1);
nand_5 g06944(n12925, n1199, new_n7321);
xor_4  g06945(new_n7321, new_n7320_1, new_n7322);
not_8  g06946(new_n7322, new_n7323);
xor_4  g06947(new_n7323, new_n7319, new_n7324);
xor_4  g06948(new_n7324, new_n7318, new_n7325);
xor_4  g06949(new_n7325, new_n7313, new_n7326);
not_8  g06950(new_n7326, new_n7327);
and_5  g06951(new_n7290, new_n7287, new_n7328);
or_5   g06952(new_n7289, new_n7288, new_n7329);
not_8  g06953(new_n7329, new_n7330);
or_5   g06954(new_n7295, new_n7292, new_n7331);
not_8  g06955(new_n7331, new_n7332);
xor_4  g06956(new_n7332, new_n7330, new_n7333);
nor_5  g06957(new_n7333, new_n7328, new_n7334);
xor_4  g06958(new_n7334, new_n7327, new_n7335);
not_8  g06959(new_n7335, new_n7336);
xor_4  g06960(new_n7336, new_n7301, new_n7337);
not_8  g06961(new_n7337, new_n7338);
nand_5 g06962(n12069, n503, new_n7339);
xor_4  g06963(new_n7300, new_n7297, new_n7340);
not_8  g06964(new_n7340, new_n7341);
nor_5  g06965(new_n7341, new_n7339, new_n7342);
or_5   g06966(new_n4192, new_n4171, new_n7343);
not_8  g06967(new_n7343, new_n7344);
xor_4  g06968(new_n7341, new_n7339, new_n7345);
and_5  g06969(new_n7345, new_n7344, new_n7346);
nor_5  g06970(new_n7346, new_n7342, new_n7347);
xor_4  g06971(new_n7347, new_n7338, new_n7348);
not_8  g06972(new_n7348, new_n7349);
nand_5 g06973(n11222, n6359, new_n7350);
nand_5 g06974(n4086, n996, new_n7351);
nand_5 g06975(n5767, n405, new_n7352);
nand_5 g06976(n8433, n5319, new_n7353);
xor_4  g06977(new_n7353, new_n7352, new_n7354_1);
not_8  g06978(new_n7354_1, new_n7355);
xor_4  g06979(new_n7355, new_n7351, new_n7356);
and_5  g06980(new_n4151, new_n4150, new_n7357);
nor_5  g06981(new_n4151, new_n4150, new_n7358);
nor_5  g06982(new_n7358, new_n4149, new_n7359);
or_5   g06983(new_n7359, new_n7357, new_n7360);
not_8  g06984(new_n7360, new_n7361);
xor_4  g06985(new_n7361, new_n7356, new_n7362);
nand_5 g06986(n11153, n6611, new_n7363);
nand_5 g06987(n5314, n217, new_n7364);
xor_4  g06988(new_n7364, new_n7363, new_n7365);
xor_4  g06989(new_n7365, new_n7362, new_n7366);
nor_5  g06990(new_n4154, new_n4147, new_n7367);
and_5  g06991(new_n4160, new_n4155_1, new_n7368);
or_5   g06992(new_n7368, new_n7367, new_n7369);
xor_4  g06993(new_n7369, new_n7366, new_n7370);
not_8  g06994(new_n7370, new_n7371);
and_5  g06995(new_n4161, new_n4146, new_n7372);
and_5  g06996(new_n4166, new_n4162, new_n7373);
nor_5  g06997(new_n7373, new_n7372, new_n7374);
xor_4  g06998(new_n7374, new_n7371, new_n7375);
not_8  g06999(new_n7375, new_n7376);
nor_5  g07000(new_n7376, new_n7350, new_n7377);
or_5   g07001(new_n4168, new_n4143, new_n7378);
not_8  g07002(new_n7378, new_n7379);
xor_4  g07003(new_n7376, new_n7350, new_n7380);
and_5  g07004(new_n7380, new_n7379, new_n7381);
or_5   g07005(new_n7381, new_n7377, new_n7382);
or_5   g07006(new_n7374, new_n7371, new_n7383);
not_8  g07007(new_n7383, new_n7384);
or_5   g07008(new_n7353, new_n7352, new_n7385);
not_8  g07009(new_n7385, new_n7386);
nand_5 g07010(n996, n217, new_n7387);
not_8  g07011(new_n7387, new_n7388_1);
xor_4  g07012(new_n7388_1, new_n7386, new_n7389);
nand_5 g07013(n5319, n405, new_n7390);
nand_5 g07014(n5767, n4086, new_n7391);
nand_5 g07015(n9457, n8433, new_n7392);
xor_4  g07016(new_n7392, new_n7391, new_n7393);
not_8  g07017(new_n7393, new_n7394);
xor_4  g07018(new_n7394, new_n7390, new_n7395);
xor_4  g07019(new_n7395, new_n7389, new_n7396);
not_8  g07020(new_n7396, new_n7397);
nand_5 g07021(n11153, n6359, new_n7398);
nand_5 g07022(n6611, n5314, new_n7399);
and_5  g07023(n11296, n11222, new_n7400);
xor_4  g07024(new_n7400, new_n7399, new_n7401);
not_8  g07025(new_n7401, new_n7402);
xor_4  g07026(new_n7402, new_n7398, new_n7403);
not_8  g07027(new_n7403, new_n7404);
nor_5  g07028(new_n7355, new_n7351, new_n7405);
and_5  g07029(new_n7361, new_n7356, new_n7406);
or_5   g07030(new_n7406, new_n7405, new_n7407);
xor_4  g07031(new_n7407, new_n7404, new_n7408);
xor_4  g07032(new_n7408, new_n7397, new_n7409);
and_5  g07033(new_n7365, new_n7362, new_n7410);
or_5   g07034(new_n7364, new_n7363, new_n7411);
not_8  g07035(new_n7411, new_n7412);
nand_5 g07036(new_n7369, new_n7366, new_n7413);
not_8  g07037(new_n7413, new_n7414);
xor_4  g07038(new_n7414, new_n7412, new_n7415);
nor_5  g07039(new_n7415, new_n7410, new_n7416);
xor_4  g07040(new_n7416, new_n7409, new_n7417);
not_8  g07041(new_n7417, new_n7418);
xor_4  g07042(new_n7418, new_n7384, new_n7419);
xor_4  g07043(new_n7419, new_n7382, new_n7420);
xor_4  g07044(new_n7420, new_n7349, new_n7421);
xor_4  g07045(new_n7345, new_n7344, new_n7422);
not_8  g07046(new_n7422, new_n7423);
xor_4  g07047(new_n7380, new_n7378, new_n7424);
and_5  g07048(new_n7424, new_n7423, new_n7425);
nor_5  g07049(new_n4197, new_n4193, new_n7426);
nor_5  g07050(new_n4199, new_n4170, new_n7427);
or_5   g07051(new_n7427, new_n7426, new_n7428);
xor_4  g07052(new_n7424, new_n7423, new_n7429);
and_5  g07053(new_n7429, new_n7428, new_n7430);
or_5   g07054(new_n7430, new_n7425, new_n7431);
xor_4  g07055(new_n7431, new_n7421, new_n7432);
not_8  g07056(new_n7432, new_n7433);
xor_4  g07057(new_n7433, new_n7275, new_n7434);
xor_4  g07058(new_n7272, new_n7269, new_n7435);
xor_4  g07059(new_n7429, new_n7428, new_n7436_1);
not_8  g07060(new_n7436_1, new_n7437);
or_5   g07061(new_n7437, new_n7435, new_n7438);
not_8  g07062(new_n7438, new_n7439);
xor_4  g07063(new_n7437, new_n7435, new_n7440);
nor_5  g07064(new_n4202, new_n4142, new_n7441);
or_5   g07065(new_n4205, new_n4204, new_n7442);
and_5  g07066(new_n7442, new_n4203_1, new_n7443);
or_5   g07067(new_n7443, new_n7441, new_n7444);
not_8  g07068(new_n7444, new_n7445);
and_5  g07069(new_n7445, new_n7440, new_n7446);
nor_5  g07070(new_n7446, new_n7439, new_n7447);
xor_4  g07071(new_n7447, new_n7434, new_n7448);
nor_5  g07072(new_n7448, new_n7204, new_n7449);
xor_4  g07073(new_n7200, new_n7199, new_n7450);
not_8  g07074(new_n7450, new_n7451);
and_5  g07075(new_n4110, new_n3947, new_n7452);
and_5  g07076(new_n4208, new_n4112, new_n7453);
or_5   g07077(new_n7453, new_n7452, new_n7454);
not_8  g07078(new_n7454, new_n7455);
and_5  g07079(new_n7455, new_n7451, new_n7456_1);
xor_4  g07080(new_n7445, new_n7440, new_n7457);
xor_4  g07081(new_n7455, new_n7451, new_n7458);
and_5  g07082(new_n7458, new_n7457, new_n7459);
or_5   g07083(new_n7459, new_n7456_1, new_n7460);
not_8  g07084(new_n7460, new_n7461);
xor_4  g07085(new_n7448, new_n7204, new_n7462);
and_5  g07086(new_n7462, new_n7461, new_n7463);
or_5   g07087(new_n7463, new_n7449, new_n7464);
and_5  g07088(new_n7332, new_n7330, new_n7465);
nor_5  g07089(new_n7334, new_n7327, new_n7466);
or_5   g07090(new_n7466, new_n7465, new_n7467);
and_5  g07091(new_n7317, new_n7315, new_n7468);
and_5  g07092(new_n7324, new_n7318, new_n7469);
nor_5  g07093(new_n7469, new_n7468, new_n7470);
and_5  g07094(new_n7177, new_n7176, new_n7471);
not_8  g07095(new_n7175, new_n7472);
nor_5  g07096(new_n7179, new_n7472, new_n7473);
or_5   g07097(new_n7473, new_n7471, new_n7474);
and_5  g07098(n6770, n2577, new_n7475);
xor_4  g07099(new_n7475, new_n7474, new_n7476);
nand_5 g07100(n9637, n4189, new_n7477);
and_5  g07101(n11917, n3627, new_n7478);
xor_4  g07102(new_n7478, new_n7477, new_n7479);
xor_4  g07103(new_n7479, new_n7476, new_n7480);
and_5  g07104(new_n7309, new_n7308, new_n7481);
nor_5  g07105(new_n7311, new_n7307, new_n7482);
nor_5  g07106(new_n7482, new_n7481, new_n7483);
nor_5  g07107(new_n7160_1, new_n7159_1, new_n7484);
and_5  g07108(new_n7168, new_n7161, new_n7485);
nor_5  g07109(new_n7485, new_n7484, new_n7486);
xor_4  g07110(new_n7486, new_n7483, new_n7487);
xor_4  g07111(new_n7487, new_n7480, new_n7488);
xor_4  g07112(new_n7488, new_n7470, new_n7489);
nand_5 g07113(new_n7312, new_n7305, new_n7490);
not_8  g07114(new_n7325, new_n7491);
nand_5 g07115(new_n7491, new_n7313, new_n7492);
nand_5 g07116(new_n7492, new_n7490, new_n7493);
and_5  g07117(new_n7249, new_n7248, new_n7494);
not_8  g07118(new_n7247, new_n7495);
nor_5  g07119(new_n7251, new_n7495, new_n7496);
or_5   g07120(new_n7496, new_n7494, new_n7497);
and_5  g07121(n7523, n3719, new_n7498);
and_5  g07122(n11222, n1357, new_n7499);
xor_4  g07123(new_n7499, new_n7498, new_n7500_1);
and_5  g07124(n8336, n4190, new_n7501);
and_5  g07125(n7320, n3602, new_n7502);
xor_4  g07126(new_n7502, new_n7501, new_n7503);
xor_4  g07127(new_n7503, new_n7500_1, new_n7504);
xor_4  g07128(new_n7504, new_n7497, new_n7505);
xor_4  g07129(new_n7505, new_n7493, new_n7506);
xor_4  g07130(new_n7506, new_n7489, new_n7507);
not_8  g07131(new_n7186, new_n7508);
nand_5 g07132(new_n7188, new_n7508, new_n7509);
not_8  g07133(new_n7509, new_n7510);
nor_5  g07134(new_n7190, new_n7183, new_n7511);
nor_5  g07135(new_n7511, new_n7510, new_n7512);
not_8  g07136(new_n7258, new_n7513);
nand_5 g07137(new_n7260, new_n7513, new_n7514);
not_8  g07138(new_n7514, new_n7515);
nor_5  g07139(new_n7262, new_n7255, new_n7516);
nor_5  g07140(new_n7516, new_n7515, new_n7517);
xor_4  g07141(new_n7517, new_n7512, new_n7518);
xor_4  g07142(new_n7518, new_n7507, new_n7519);
xor_4  g07143(new_n7519, new_n7467, new_n7520);
and_5  g07144(new_n7263, new_n7228, new_n7521);
not_8  g07145(new_n7264, new_n7522);
nor_5  g07146(new_n7274, new_n7522, new_n7523_1);
or_5   g07147(new_n7523_1, new_n7521, new_n7524);
and_5  g07148(new_n7236_1, new_n7235, new_n7525);
nor_5  g07149(new_n7238, new_n7234, new_n7526);
nor_5  g07150(new_n7526, new_n7525, new_n7527);
nand_5 g07151(n5319, n4086, new_n7528);
and_5  g07152(n10928, n10391, new_n7529);
xor_4  g07153(new_n7529, new_n7528, new_n7530);
xor_4  g07154(new_n7530, new_n7527, new_n7531);
xor_4  g07155(new_n7531, new_n7524, new_n7532);
xor_4  g07156(new_n7532, new_n7520, new_n7533);
nor_5  g07157(new_n7336, new_n7301, new_n7534);
nor_5  g07158(new_n7347, new_n7338, new_n7535);
nor_5  g07159(new_n7535, new_n7534, new_n7536);
and_5  g07160(new_n7417, new_n7384, new_n7537);
not_8  g07161(new_n7419, new_n7538);
and_5  g07162(new_n7538, new_n7382, new_n7539);
nor_5  g07163(new_n7539, new_n7537, new_n7540);
xor_4  g07164(new_n7540, new_n7536, new_n7541);
xor_4  g07165(new_n7541, new_n7533, new_n7542);
and_5  g07166(n4826, n2515, new_n7543);
and_5  g07167(n12925, n6578, new_n7544);
xor_4  g07168(new_n7544, new_n7543, new_n7545);
nand_5 g07169(n6359, n5314, new_n7546_1);
and_5  g07170(n12069, n7546, new_n7547);
xor_4  g07171(new_n7547, new_n7546_1, new_n7548);
xor_4  g07172(new_n7548, new_n7545, new_n7549);
and_5  g07173(new_n7392, new_n7391, new_n7550);
not_8  g07174(new_n7390, new_n7551);
nor_5  g07175(new_n7394, new_n7551, new_n7552);
nor_5  g07176(new_n7552, new_n7550, new_n7553);
and_5  g07177(new_n7402, new_n7398, new_n7554);
or_5   g07178(new_n7554, new_n7399, new_n7555);
not_8  g07179(new_n7555, new_n7556);
and_5  g07180(n11296, n11153, new_n7557);
and_5  g07181(new_n7557, new_n7556, new_n7558);
and_5  g07182(new_n7557, new_n7350, new_n7559);
nor_5  g07183(new_n7559, new_n7556, new_n7560);
nor_5  g07184(new_n7560, new_n7558, new_n7561);
xor_4  g07185(new_n7561, new_n7553, new_n7562);
xor_4  g07186(new_n7562, new_n7549, new_n7563);
xor_4  g07187(new_n7563, new_n7542, new_n7564);
xnor_4 g07188(new_n7274, new_n7264, new_n7565);
nor_5  g07189(new_n7433, new_n7565, new_n7566);
nor_5  g07190(new_n7447, new_n7434, new_n7567);
or_5   g07191(new_n7567, new_n7566, new_n7568_1);
and_5  g07192(new_n7420, new_n7349, new_n7569);
and_5  g07193(new_n7431, new_n7421, new_n7570);
nor_5  g07194(new_n7570, new_n7569, new_n7571);
and_5  g07195(new_n7191, new_n7157, new_n7572);
nor_5  g07196(new_n7202, new_n7193_1, new_n7573);
or_5   g07197(new_n7573, new_n7572, new_n7574);
and_5  g07198(new_n7414, new_n7412, new_n7575);
nor_5  g07199(new_n7416, new_n7409, new_n7576);
or_5   g07200(new_n7576, new_n7575, new_n7577);
and_5  g07201(new_n7180, new_n7174, new_n7578);
and_5  g07202(new_n7181, new_n7170, new_n7579);
nor_5  g07203(new_n7579, new_n7578, new_n7580);
or_5   g07204(new_n7240, new_n7232, new_n7581);
not_8  g07205(new_n7253, new_n7582);
nand_5 g07206(new_n7582, new_n7241, new_n7583);
and_5  g07207(new_n7583, new_n7581, new_n7584);
xor_4  g07208(new_n7584, new_n7580, new_n7585);
and_5  g07209(new_n7388_1, new_n7386, new_n7586);
and_5  g07210(new_n7395, new_n7389, new_n7587);
or_5   g07211(new_n7587, new_n7586, new_n7588);
nand_5 g07212(n8595, n1094, new_n7589);
and_5  g07213(n2564, n1835, new_n7590);
xor_4  g07214(new_n7590, new_n7589, new_n7591);
xor_4  g07215(new_n7591, new_n7588, new_n7592);
and_5  g07216(new_n7321, new_n7320_1, new_n7593);
not_8  g07217(new_n7319, new_n7594);
nor_5  g07218(new_n7323, new_n7594, new_n7595);
nor_5  g07219(new_n7595, new_n7593, new_n7596);
and_5  g07220(n12391, n10965, new_n7597);
nand_5 g07221(n7891, n503, new_n7598);
and_5  g07222(n9457, n405, new_n7599);
xor_4  g07223(new_n7599, new_n7598, new_n7600);
xor_4  g07224(new_n7600, new_n7597, new_n7601);
xor_4  g07225(new_n7601, new_n7596, new_n7602);
nand_5 g07226(n8065, n6986, new_n7603);
and_5  g07227(n10439, n2226, new_n7604);
xor_4  g07228(new_n7604, new_n7603, new_n7605);
xor_4  g07229(new_n7605, new_n7602, new_n7606);
xor_4  g07230(new_n7606, new_n7592, new_n7607);
and_5  g07231(new_n7165, new_n7164, new_n7608);
nor_5  g07232(new_n7167, new_n7163, new_n7609);
or_5   g07233(new_n7609, new_n7608, new_n7610_1);
and_5  g07234(n11536, n6687, new_n7611);
and_5  g07235(n6611, n996, new_n7612);
xor_4  g07236(new_n7612, new_n7611, new_n7613);
nand_5 g07237(n4921, n4516, new_n7614);
and_5  g07238(n9920, n3842, new_n7615);
xor_4  g07239(new_n7615, new_n7614, new_n7616);
xor_4  g07240(new_n7616, new_n7613, new_n7617);
xor_4  g07241(new_n7617, new_n7610_1, new_n7618);
nand_5 g07242(n9956, n2087, new_n7619);
and_5  g07243(n7733, n1199, new_n7620);
and_5  g07244(n5767, n217, new_n7621);
xor_4  g07245(new_n7621, new_n7620, new_n7622);
and_5  g07246(n7160, n4970, new_n7623);
and_5  g07247(n7610, n4828, new_n7624);
xor_4  g07248(new_n7624, new_n7623, new_n7625);
xor_4  g07249(new_n7625, new_n7622, new_n7626);
xor_4  g07250(new_n7626, new_n7619, new_n7627);
xor_4  g07251(new_n7627, new_n7618, new_n7628);
and_5  g07252(new_n7245, new_n7243, new_n7629);
and_5  g07253(new_n7252, new_n7246, new_n7630);
or_5   g07254(new_n7630, new_n7629, new_n7631);
nand_5 g07255(n8433, n4817, new_n7632);
and_5  g07256(n10678, n6126, new_n7633);
xor_4  g07257(new_n7633, new_n7632, new_n7634);
xor_4  g07258(new_n7634, new_n7631, new_n7635);
xor_4  g07259(new_n7635, new_n7628, new_n7636);
xor_4  g07260(new_n7636, new_n7607, new_n7637);
xor_4  g07261(new_n7637, new_n7585, new_n7638);
xor_4  g07262(new_n7638, new_n7577, new_n7639);
xor_4  g07263(new_n7639, new_n7574, new_n7640);
xor_4  g07264(new_n7640, new_n7571, new_n7641);
nor_5  g07265(new_n7407, new_n7404, new_n7642);
and_5  g07266(new_n7408, new_n7397, new_n7643);
nor_5  g07267(new_n7643, new_n7642, new_n7644);
xor_4  g07268(new_n7644, new_n7641, new_n7645);
xor_4  g07269(new_n7645, new_n7568_1, new_n7646_1);
xor_4  g07270(new_n7646_1, new_n7564, new_n7647);
xor_4  g07271(new_n7647, new_n7464, n2679);
or_5   g07272(new_n5544, new_n5523, new_n7649);
not_8  g07273(new_n7649, new_n7650);
nand_5 g07274(n6687, n2253, new_n7651);
not_8  g07275(new_n7651, new_n7652);
nand_5 g07276(n10223, n6770, new_n7653);
nand_5 g07277(n9920, n2879, new_n7654);
nand_5 g07278(n7265, n3627, new_n7655);
xor_4  g07279(new_n7655, new_n7654, new_n7656);
not_8  g07280(new_n7656, new_n7657);
xor_4  g07281(new_n7657, new_n7653, new_n7658);
and_5  g07282(new_n5529, new_n5498, new_n7659);
nor_5  g07283(new_n5531, new_n5528, new_n7660);
or_5   g07284(new_n7660, new_n7659, new_n7661);
not_8  g07285(new_n7661, new_n7662);
xor_4  g07286(new_n7662, new_n7658, new_n7663);
nand_5 g07287(n9195, n2564, new_n7664);
nand_5 g07288(n4634, n4189, new_n7665);
xor_4  g07289(new_n7665, new_n7664, new_n7666);
xor_4  g07290(new_n7666, new_n7663, new_n7667);
nor_5  g07291(new_n5532, new_n5526, new_n7668);
and_5  g07292(new_n5537, new_n5533, new_n7669);
nor_5  g07293(new_n7669, new_n7668, new_n7670);
xor_4  g07294(new_n7670, new_n7667, new_n7671);
and_5  g07295(new_n5538, new_n5525, new_n7672);
nor_5  g07296(new_n5542, new_n5540, new_n7673);
nor_5  g07297(new_n7673, new_n7672, new_n7674);
xor_4  g07298(new_n7674, new_n7671, new_n7675);
xor_4  g07299(new_n7675, new_n7652, new_n7676_1);
not_8  g07300(new_n7676_1, new_n7677);
and_5  g07301(new_n7677, new_n7650, new_n7678);
nor_5  g07302(new_n7677, new_n7650, new_n7679);
or_5   g07303(new_n7679, new_n7678, new_n7680);
not_8  g07304(new_n7680, new_n7681);
nor_5  g07305(new_n5765, new_n5545, new_n7682);
nor_5  g07306(new_n5799, new_n7682, new_n7683);
xor_4  g07307(new_n7683, new_n7681, new_n7684);
not_8  g07308(new_n7684, new_n7685);
or_5   g07309(new_n5600, new_n5576, new_n7686);
not_8  g07310(new_n7686, new_n7687);
nand_5 g07311(n12221, n8336, new_n7688);
nand_5 g07312(n9189, n2226, new_n7689);
nand_5 g07313(n2024, n1094, new_n7690_1);
nand_5 g07314(n10678, n7946, new_n7691);
xor_4  g07315(new_n7691, new_n7690_1, new_n7692);
not_8  g07316(new_n7692, new_n7693);
xor_4  g07317(new_n7693, new_n7689, new_n7694);
and_5  g07318(new_n5590, new_n5552, new_n7695);
nor_5  g07319(new_n5592, new_n5589, new_n7696);
or_5   g07320(new_n7696, new_n7695, new_n7697);
not_8  g07321(new_n7697, new_n7698);
xor_4  g07322(new_n7698, new_n7694, new_n7699);
nand_5 g07323(n12145, n10928, new_n7700);
nand_5 g07324(n6986, n2522, new_n7701);
xor_4  g07325(new_n7701, new_n7700, new_n7702);
xor_4  g07326(new_n7702, new_n7699, new_n7703);
not_8  g07327(new_n7703, new_n7704);
nor_5  g07328(new_n5586, new_n5580, new_n7705);
nor_5  g07329(new_n5593, new_n5587, new_n7706);
nor_5  g07330(new_n7706, new_n7705, new_n7707);
xor_4  g07331(new_n7707, new_n7704, new_n7708);
not_8  g07332(new_n7708, new_n7709);
and_5  g07333(new_n5594, new_n5579_1, new_n7710);
and_5  g07334(new_n5598, new_n5595, new_n7711);
nor_5  g07335(new_n7711, new_n7710, new_n7712);
xor_4  g07336(new_n7712, new_n7709, new_n7713);
not_8  g07337(new_n7713, new_n7714);
xor_4  g07338(new_n7714, new_n7688, new_n7715);
xor_4  g07339(new_n7715, new_n7687, new_n7716);
nor_5  g07340(new_n5708, new_n5601, new_n7717);
nor_5  g07341(new_n5764, new_n5709, new_n7718);
nor_5  g07342(new_n7718, new_n7717, new_n7719);
xor_4  g07343(new_n7719, new_n7716, new_n7720);
not_8  g07344(new_n7720, new_n7721);
or_5   g07345(new_n5733, new_n5710, new_n7722);
not_8  g07346(new_n7722, new_n7723);
nand_5 g07347(n12069, n5798, new_n7724);
nand_5 g07348(n7160, n5579, new_n7725);
not_8  g07349(new_n7725, new_n7726);
not_8  g07350(new_n5723, new_n7727);
and_5  g07351(new_n5725, new_n5722, new_n7728);
nor_5  g07352(new_n7728, new_n7727, new_n7729);
nor_5  g07353(new_n7729, new_n7726, new_n7730_1);
nor_5  g07354(new_n7729, new_n5617, new_n7731);
nor_5  g07355(new_n7731, new_n7725, new_n7732);
or_5   g07356(new_n7732, new_n7730_1, new_n7733_1);
not_8  g07357(new_n7733_1, new_n7734);
nand_5 g07358(n4828, n2498, new_n7735);
nand_5 g07359(n2558, n2515, new_n7736);
xor_4  g07360(new_n7736, new_n7735, new_n7737);
nor_5  g07361(new_n7737, new_n7734, new_n7738);
and_5  g07362(new_n7737, new_n7734, new_n7739);
or_5   g07363(new_n7739, new_n7738, new_n7740);
nand_5 g07364(n12391, n6016, new_n7741);
nand_5 g07365(n7891, n521, new_n7742);
xor_4  g07366(new_n7742, new_n7741, new_n7743);
not_8  g07367(new_n7743, new_n7744);
xor_4  g07368(new_n7744, new_n7740, new_n7745);
nor_5  g07369(new_n5719, new_n5713, new_n7746);
nor_5  g07370(new_n5726, new_n5720, new_n7747);
nor_5  g07371(new_n7747, new_n7746, new_n7748);
xor_4  g07372(new_n7748, new_n7745, new_n7749);
not_8  g07373(new_n7749, new_n7750);
and_5  g07374(new_n5727, new_n5712, new_n7751);
nor_5  g07375(new_n5731, new_n5729, new_n7752);
or_5   g07376(new_n7752, new_n7751, new_n7753);
xor_4  g07377(new_n7753, new_n7750, new_n7754);
not_8  g07378(new_n7754, new_n7755);
xor_4  g07379(new_n7755, new_n7724, new_n7756);
xor_4  g07380(new_n7756, new_n7723, new_n7757);
not_8  g07381(new_n7757, new_n7758);
or_5   g07382(new_n5758, new_n5735, new_n7759);
not_8  g07383(new_n7759, new_n7760);
nand_5 g07384(n11222, n5153, new_n7761);
not_8  g07385(new_n7761, new_n7762);
nand_5 g07386(n3342, n996, new_n7763);
nand_5 g07387(n9111, n5767, new_n7764);
nand_5 g07388(n9763, n5319, new_n7765);
xor_4  g07389(new_n7765, new_n7764, new_n7766);
not_8  g07390(new_n7766, new_n7767);
xor_4  g07391(new_n7767, new_n7763, new_n7768);
and_5  g07392(new_n5748, new_n5637, new_n7769);
nor_5  g07393(new_n5748, new_n5637, new_n7770);
nor_5  g07394(new_n7770, new_n5747, new_n7771);
or_5   g07395(new_n7771, new_n7769, new_n7772);
not_8  g07396(new_n7772, new_n7773);
xor_4  g07397(new_n7773, new_n7768, new_n7774);
nand_5 g07398(n11153, n7270, new_n7775);
nand_5 g07399(n5314, n806, new_n7776);
xor_4  g07400(new_n7776, new_n7775, new_n7777);
xor_4  g07401(new_n7777, new_n7774, new_n7778);
nor_5  g07402(new_n5744, new_n5739, new_n7779);
and_5  g07403(new_n5750, new_n5745, new_n7780);
or_5   g07404(new_n7780, new_n7779, new_n7781);
xnor_4 g07405(new_n7781, new_n7778, new_n7782);
and_5  g07406(new_n5751, new_n5738, new_n7783);
and_5  g07407(new_n5756, new_n5752, new_n7784);
nor_5  g07408(new_n7784, new_n7783, new_n7785);
xor_4  g07409(new_n7785, new_n7782, new_n7786);
xor_4  g07410(new_n7786, new_n7762, new_n7787);
not_8  g07411(new_n7787, new_n7788);
nand_5 g07412(new_n7788, new_n7760, new_n7789);
or_5   g07413(new_n7788, new_n7760, new_n7790);
and_5  g07414(new_n7790, new_n7789, new_n7791);
xor_4  g07415(new_n7791, new_n7758, new_n7792);
not_8  g07416(new_n5734, new_n7793);
and_5  g07417(new_n5759, new_n7793, new_n7794);
nor_5  g07418(new_n5763, new_n5760_1, new_n7795);
or_5   g07419(new_n7795, new_n7794, new_n7796);
not_8  g07420(new_n7796, new_n7797);
xor_4  g07421(new_n7797, new_n7792, new_n7798);
and_5  g07422(new_n7798, new_n7721, new_n7799);
nor_5  g07423(new_n7798, new_n7721, new_n7800);
or_5   g07424(new_n7800, new_n7799, new_n7801);
xnor_4 g07425(new_n7801, new_n7685, n2708);
xor_4  g07426(new_n863, new_n862, n2818);
xor_4  g07427(new_n2051, new_n2024_1, n2902);
nand_5 g07428(n11407, n5305, new_n7805);
not_8  g07429(new_n7805, new_n7806);
nand_5 g07430(n12709, n8759, new_n7807);
nand_5 g07431(n12489, n5331, new_n7808);
nand_5 g07432(n10990, n7965, new_n7809);
xor_4  g07433(new_n7809, new_n7808, new_n7810);
not_8  g07434(new_n7810, new_n7811);
xor_4  g07435(new_n7811, new_n7807, new_n7812);
xor_4  g07436(new_n7812, new_n7806, n3071);
xnor_4 g07437(new_n2868, new_n2866, n3124);
nand_5 g07438(new_n7812, new_n7806, new_n7815);
nand_5 g07439(n11407, n5964, new_n7816);
and_5  g07440(n5305, n5212, new_n7817);
xor_4  g07441(new_n7817, new_n7816, new_n7818);
and_5  g07442(new_n7818, new_n7815, new_n7819);
or_5   g07443(new_n7811, new_n7807, new_n7820);
nand_5 g07444(n11728, n8759, new_n7821);
and_5  g07445(n12709, n6776, new_n7822);
xor_4  g07446(new_n7822, new_n7821, new_n7823_1);
not_8  g07447(new_n7823_1, new_n7824);
xor_4  g07448(new_n7824, new_n7820, new_n7825);
or_5   g07449(new_n7809, new_n7808, new_n7826);
and_5  g07450(n7159, n5331, new_n7827);
and_5  g07451(n12489, n8476, new_n7828);
xor_4  g07452(new_n7828, new_n7827, new_n7829);
xor_4  g07453(new_n7829, new_n7826, new_n7830);
and_5  g07454(n7965, n5760, new_n7831);
and_5  g07455(n10990, n7388, new_n7832);
xor_4  g07456(new_n7832, new_n7831, new_n7833);
xor_4  g07457(new_n7833, new_n7830, new_n7834);
xor_4  g07458(new_n7834, new_n7825, new_n7835);
xor_4  g07459(new_n7818, new_n7815, new_n7836);
not_8  g07460(new_n7836, new_n7837);
nor_5  g07461(new_n7837, new_n7835, new_n7838);
or_5   g07462(new_n7838, new_n7819, new_n7839);
not_8  g07463(new_n7839, new_n7840);
nand_5 g07464(n5964, n5212, new_n7841);
or_5   g07465(new_n7841, new_n7806, new_n7842);
nand_5 g07466(n11407, n1097, new_n7843);
nand_5 g07467(n11877, n5305, new_n7844);
xnor_4 g07468(new_n7844, new_n7843, new_n7845);
and_5  g07469(new_n7845, new_n7842, new_n7846);
and_5  g07470(new_n7844, new_n7843, new_n7847);
nor_5  g07471(new_n7847, new_n7842, new_n7848);
or_5   g07472(new_n7848, new_n7846, new_n7849);
not_8  g07473(new_n7849, new_n7850);
xor_4  g07474(new_n7850, new_n7840, new_n7851);
nor_5  g07475(new_n7823_1, new_n7820, new_n7852);
nor_5  g07476(new_n7834, new_n7825, new_n7853);
or_5   g07477(new_n7853, new_n7852, new_n7854);
not_8  g07478(new_n7854, new_n7855);
not_8  g07479(new_n7807, new_n7856);
nand_5 g07480(n11728, n6776, new_n7857);
or_5   g07481(new_n7857, new_n7856, new_n7858);
nand_5 g07482(n12709, n12299, new_n7859);
nand_5 g07483(n8759, n6429, new_n7860);
xnor_4 g07484(new_n7860, new_n7859, new_n7861);
and_5  g07485(new_n7861, new_n7858, new_n7862_1);
and_5  g07486(new_n7860, new_n7859, new_n7863);
nor_5  g07487(new_n7863, new_n7858, new_n7864);
or_5   g07488(new_n7864, new_n7862_1, new_n7865);
nor_5  g07489(new_n7865, new_n7855, new_n7866);
and_5  g07490(new_n7865, new_n7855, new_n7867);
or_5   g07491(new_n7867, new_n7866, new_n7868);
not_8  g07492(new_n7808, new_n7869);
nand_5 g07493(n8476, n7159, new_n7870);
or_5   g07494(new_n7870, new_n7869, new_n7871);
not_8  g07495(new_n7871, new_n7872);
and_5  g07496(n12489, n2530, new_n7873);
and_5  g07497(n12777, n5331, new_n7874);
nor_5  g07498(new_n7874, new_n7873, new_n7875);
nand_5 g07499(n12777, n2530, new_n7876);
nor_5  g07500(new_n7876, new_n7808, new_n7877);
nor_5  g07501(new_n7877, new_n7875, new_n7878);
or_5   g07502(new_n7878, new_n7872, new_n7879);
not_8  g07503(new_n7879, new_n7880);
nor_5  g07504(new_n7875, new_n7871, new_n7881);
or_5   g07505(new_n7881, new_n7880, new_n7882);
and_5  g07506(n7388, n5760, new_n7883);
nand_5 g07507(new_n7883, new_n7809, new_n7884);
not_8  g07508(new_n7884, new_n7885);
nand_5 g07509(n11892, n10990, new_n7886);
nand_5 g07510(n7965, n1478, new_n7887);
xor_4  g07511(new_n7887, new_n7886, new_n7888);
or_5   g07512(new_n7888, new_n7885, new_n7889);
and_5  g07513(new_n7887, new_n7886, new_n7890);
or_5   g07514(new_n7890, new_n7884, new_n7891_1);
nand_5 g07515(new_n7891_1, new_n7889, new_n7892);
xor_4  g07516(new_n7892, new_n7882, new_n7893);
not_8  g07517(new_n7826, new_n7894);
nor_5  g07518(new_n7829, new_n7894, new_n7895);
nor_5  g07519(new_n7833, new_n7830, new_n7896);
or_5   g07520(new_n7896, new_n7895, new_n7897);
not_8  g07521(new_n7897, new_n7898);
xor_4  g07522(new_n7898, new_n7893, new_n7899);
xor_4  g07523(new_n7899, new_n7868, new_n7900);
xnor_4 g07524(new_n7900, new_n7851, n3214);
xnor_4 g07525(new_n5357, new_n5356, n3230);
xor_4  g07526(new_n4858, new_n4807, n3272);
nand_5 g07527(n5964, n4370, new_n7904);
not_8  g07528(new_n7904, new_n7905);
nand_5 g07529(n11407, n4312, new_n7906);
nand_5 g07530(n11877, n5964, new_n7907);
and_5  g07531(new_n7907, new_n7906, new_n7908);
nor_5  g07532(new_n7907, new_n7906, new_n7909);
nand_5 g07533(n5212, n1097, new_n7910);
not_8  g07534(new_n7910, new_n7911);
nor_5  g07535(new_n7911, new_n7909, new_n7912);
or_5   g07536(new_n7912, new_n7908, new_n7913);
not_8  g07537(new_n7913, new_n7914);
and_5  g07538(new_n7914, new_n7905, new_n7915);
nor_5  g07539(new_n7914, new_n7905, new_n7916);
or_5   g07540(new_n7916, new_n7915, new_n7917);
nand_5 g07541(n5212, n4312, new_n7918);
not_8  g07542(new_n7918, new_n7919);
nand_5 g07543(n11877, n1097, new_n7920);
nand_5 g07544(n12705, n11407, new_n7921);
xor_4  g07545(new_n7921, new_n7920, new_n7922);
xor_4  g07546(new_n7922, new_n7919, new_n7923);
not_8  g07547(new_n7923, new_n7924);
nor_5  g07548(new_n7924, new_n7917, new_n7925);
or_5   g07549(new_n7925, new_n7915, new_n7926);
not_8  g07550(new_n7926, new_n7927);
nand_5 g07551(n5964, n5320, new_n7928);
nand_5 g07552(n4370, n1097, new_n7929);
xor_4  g07553(new_n7929, new_n7928, new_n7930);
not_8  g07554(new_n7930, new_n7931);
xor_4  g07555(new_n7931, new_n7927, new_n7932);
nand_5 g07556(n11877, n4312, new_n7933);
not_8  g07557(new_n7933, new_n7934);
nand_5 g07558(n12705, n5212, new_n7935);
nand_5 g07559(n12025, n11407, new_n7936);
xor_4  g07560(new_n7936, new_n7935, new_n7937);
xor_4  g07561(new_n7937, new_n7934, new_n7938);
and_5  g07562(new_n7921, new_n7920, new_n7939);
nor_5  g07563(new_n7921, new_n7920, new_n7940);
nor_5  g07564(new_n7940, new_n7919, new_n7941);
nor_5  g07565(new_n7941, new_n7939, new_n7942);
xor_4  g07566(new_n7942, new_n7938, new_n7943);
xor_4  g07567(new_n7943, new_n7932, new_n7944);
nand_5 g07568(n5320, n5305, new_n7945);
not_8  g07569(new_n7945, new_n7946_1);
xor_4  g07570(new_n7924, new_n7917, new_n7947);
nor_5  g07571(new_n7947, new_n7946_1, new_n7948);
xor_4  g07572(new_n7947, new_n7946_1, new_n7949);
not_8  g07573(new_n7949, new_n7950);
nand_5 g07574(n5305, n4370, new_n7951);
not_8  g07575(new_n7951, new_n7952);
not_8  g07576(new_n7841, new_n7953);
nor_5  g07577(new_n7844, new_n7843, new_n7954);
nor_5  g07578(new_n7954, new_n7953, new_n7955);
or_5   g07579(new_n7955, new_n7847, new_n7956);
not_8  g07580(new_n7956, new_n7957);
and_5  g07581(new_n7957, new_n7952, new_n7958);
nor_5  g07582(new_n7957, new_n7952, new_n7959);
or_5   g07583(new_n7959, new_n7958, new_n7960);
xor_4  g07584(new_n7907, new_n7906, new_n7961);
xor_4  g07585(new_n7961, new_n7910, new_n7962);
nor_5  g07586(new_n7962, new_n7960, new_n7963);
or_5   g07587(new_n7963, new_n7958, new_n7964);
nor_5  g07588(new_n7964, new_n7950, new_n7965_1);
or_5   g07589(new_n7965_1, new_n7948, new_n7966_1);
not_8  g07590(new_n7966_1, new_n7967);
nand_5 g07591(new_n7967, new_n7944, new_n7968);
nor_5  g07592(new_n7937, new_n7934, new_n7969);
not_8  g07593(new_n7938, new_n7970);
nor_5  g07594(new_n7942, new_n7970, new_n7971);
or_5   g07595(new_n7971, new_n7969, new_n7972);
not_8  g07596(new_n7972, new_n7973);
nand_5 g07597(n12000, n5964, new_n7974);
not_8  g07598(new_n7974, new_n7975);
nand_5 g07599(n5320, n1097, new_n7976);
nand_5 g07600(n9725, n5305, new_n7977);
xor_4  g07601(new_n7977, new_n7976, new_n7978);
not_8  g07602(new_n7978, new_n7979);
xor_4  g07603(new_n7979, new_n7975, new_n7980);
not_8  g07604(new_n7980, new_n7981_1);
nor_5  g07605(new_n7981_1, new_n7973, new_n7982);
and_5  g07606(new_n7981_1, new_n7973, new_n7983);
or_5   g07607(new_n7983, new_n7982, new_n7984);
or_5   g07608(new_n7936, new_n7935, new_n7985);
not_8  g07609(new_n7985, new_n7986);
and_5  g07610(n4370, n4312, new_n7987);
xor_4  g07611(new_n7987, new_n7986, new_n7988);
nand_5 g07612(n12025, n5212, new_n7989);
not_8  g07613(new_n7989, new_n7990);
nand_5 g07614(n12705, n11877, new_n7991);
nand_5 g07615(n11407, n11257, new_n7992);
xor_4  g07616(new_n7992, new_n7991, new_n7993);
not_8  g07617(new_n7993, new_n7994);
xor_4  g07618(new_n7994, new_n7990, new_n7995);
xor_4  g07619(new_n7995, new_n7988, new_n7996);
not_8  g07620(new_n7996, new_n7997);
xor_4  g07621(new_n7997, new_n7984, new_n7998);
nor_5  g07622(new_n7931, new_n7927, new_n7999);
or_5   g07623(new_n7929, new_n7928, new_n8000);
not_8  g07624(new_n8000, new_n8001);
and_5  g07625(new_n7943, new_n7932, new_n8002);
xor_4  g07626(new_n8002, new_n8001, new_n8003);
nor_5  g07627(new_n8003, new_n7999, new_n8004);
xor_4  g07628(new_n8004, new_n7998, new_n8005);
not_8  g07629(new_n8005, new_n8006);
nor_5  g07630(new_n8006, new_n7968, new_n8007);
and_5  g07631(new_n8006, new_n7968, new_n8008);
or_5   g07632(new_n8008, new_n8007, new_n8009);
nand_5 g07633(n12000, n5305, new_n8010);
not_8  g07634(new_n8010, new_n8011);
xor_4  g07635(new_n7967, new_n7944, new_n8012);
and_5  g07636(new_n8012, new_n8011, new_n8013);
xor_4  g07637(new_n7962, new_n7960, new_n8014);
not_8  g07638(new_n7846, new_n8015);
or_5   g07639(new_n8015, new_n7841, new_n8016);
not_8  g07640(new_n8016, new_n8017);
nand_5 g07641(new_n8017, new_n8014, new_n8018);
not_8  g07642(new_n7964, new_n8019);
xnor_4 g07643(new_n8019, new_n7950, new_n8020);
or_5   g07644(new_n8020, new_n8018, new_n8021);
not_8  g07645(new_n8021, new_n8022);
xor_4  g07646(new_n8012, new_n8011, new_n8023);
and_5  g07647(new_n8023, new_n8022, new_n8024);
nor_5  g07648(new_n8024, new_n8013, new_n8025);
xor_4  g07649(new_n8025, new_n8009, new_n8026);
not_8  g07650(new_n8026, new_n8027);
nand_5 g07651(n8759, n8717, new_n8028_1);
not_8  g07652(new_n8028_1, new_n8029);
nand_5 g07653(n7436, n6429, new_n8030);
not_8  g07654(new_n8030, new_n8031);
nand_5 g07655(n12709, n9241, new_n8032);
nand_5 g07656(n11728, n8276, new_n8033);
xor_4  g07657(new_n8033, new_n8032, new_n8034);
xor_4  g07658(new_n8034, new_n8031, new_n8035);
not_8  g07659(new_n8035, new_n8036);
nand_5 g07660(n12299, n6429, new_n8037);
nand_5 g07661(n12709, n8276, new_n8038);
and_5  g07662(new_n8038, new_n8037, new_n8039);
nor_5  g07663(new_n8038, new_n8037, new_n8040);
nand_5 g07664(n11728, n7436, new_n8041);
not_8  g07665(new_n8041, new_n8042);
nor_5  g07666(new_n8042, new_n8040, new_n8043);
nor_5  g07667(new_n8043, new_n8039, new_n8044);
xor_4  g07668(new_n8044, new_n8036, new_n8045);
not_8  g07669(new_n8045, new_n8046);
nand_5 g07670(n6776, n2433, new_n8047);
nand_5 g07671(n12299, n8819, new_n8048);
xor_4  g07672(new_n8048, new_n8047, new_n8049);
xor_4  g07673(new_n8049, new_n8046, new_n8050);
and_5  g07674(n8819, n6776, new_n8051);
nand_5 g07675(n12709, n7436, new_n8052);
nand_5 g07676(n6776, n6429, new_n8053);
and_5  g07677(new_n8053, new_n8052, new_n8054);
nor_5  g07678(new_n8053, new_n8052, new_n8055);
nand_5 g07679(n12299, n11728, new_n8056);
not_8  g07680(new_n8056, new_n8057);
nor_5  g07681(new_n8057, new_n8055, new_n8058);
or_5   g07682(new_n8058, new_n8054, new_n8059);
not_8  g07683(new_n8059, new_n8060);
and_5  g07684(new_n8060, new_n8051, new_n8061);
nor_5  g07685(new_n8060, new_n8051, new_n8062);
or_5   g07686(new_n8062, new_n8061, new_n8063);
xor_4  g07687(new_n8038, new_n8037, new_n8064);
xor_4  g07688(new_n8064, new_n8041, new_n8065_1);
nor_5  g07689(new_n8065_1, new_n8063, new_n8066);
or_5   g07690(new_n8066, new_n8061, new_n8067);
xor_4  g07691(new_n8067, new_n8050, new_n8068);
nand_5 g07692(n8759, n2433, new_n8069);
not_8  g07693(new_n8069, new_n8070);
xor_4  g07694(new_n8065_1, new_n8063, new_n8071);
nor_5  g07695(new_n8071, new_n8070, new_n8072);
xor_4  g07696(new_n8071, new_n8070, new_n8073);
not_8  g07697(new_n8073, new_n8074);
nand_5 g07698(n8819, n8759, new_n8075);
not_8  g07699(new_n8075, new_n8076);
not_8  g07700(new_n7857, new_n8077);
nor_5  g07701(new_n7860, new_n7859, new_n8078);
nor_5  g07702(new_n8078, new_n8077, new_n8079);
or_5   g07703(new_n8079, new_n7863, new_n8080);
not_8  g07704(new_n8080, new_n8081);
and_5  g07705(new_n8081, new_n8076, new_n8082);
nor_5  g07706(new_n8081, new_n8076, new_n8083);
or_5   g07707(new_n8083, new_n8082, new_n8084);
xor_4  g07708(new_n8053, new_n8052, new_n8085);
xor_4  g07709(new_n8085, new_n8056, new_n8086);
nor_5  g07710(new_n8086, new_n8084, new_n8087);
or_5   g07711(new_n8087, new_n8082, new_n8088);
nor_5  g07712(new_n8088, new_n8074, new_n8089);
or_5   g07713(new_n8089, new_n8072, new_n8090);
not_8  g07714(new_n8090, new_n8091);
xor_4  g07715(new_n8091, new_n8068, new_n8092);
and_5  g07716(new_n8092, new_n8029, new_n8093);
xor_4  g07717(new_n8086, new_n8084, new_n8094);
not_8  g07718(new_n7862_1, new_n8095);
or_5   g07719(new_n8095, new_n7857, new_n8096);
not_8  g07720(new_n8096, new_n8097);
nand_5 g07721(new_n8097, new_n8094, new_n8098);
not_8  g07722(new_n8088, new_n8099);
xnor_4 g07723(new_n8099, new_n8074, new_n8100_1);
or_5   g07724(new_n8100_1, new_n8098, new_n8101);
not_8  g07725(new_n8101, new_n8102);
xor_4  g07726(new_n8092, new_n8029, new_n8103);
and_5  g07727(new_n8103, new_n8102, new_n8104);
or_5   g07728(new_n8104, new_n8093, new_n8105);
not_8  g07729(new_n8105, new_n8106);
nand_5 g07730(new_n8091, new_n8068, new_n8107);
nor_5  g07731(new_n8034, new_n8031, new_n8108);
nor_5  g07732(new_n8044, new_n8036, new_n8109);
or_5   g07733(new_n8109, new_n8108, new_n8110);
not_8  g07734(new_n8110, new_n8111);
nand_5 g07735(n8717, n6776, new_n8112);
nand_5 g07736(n12299, n2433, new_n8113);
nand_5 g07737(n8759, n7730, new_n8114);
xor_4  g07738(new_n8114, new_n8113, new_n8115);
xor_4  g07739(new_n8115, new_n8112, new_n8116);
not_8  g07740(new_n8116, new_n8117);
nor_5  g07741(new_n8117, new_n8111, new_n8118);
and_5  g07742(new_n8117, new_n8111, new_n8119);
or_5   g07743(new_n8119, new_n8118, new_n8120);
or_5   g07744(new_n8033, new_n8032, new_n8121);
nand_5 g07745(n8819, n7436, new_n8122);
not_8  g07746(new_n8122, new_n8123);
xor_4  g07747(new_n8123, new_n8121, new_n8124);
nand_5 g07748(n11728, n9241, new_n8125);
not_8  g07749(new_n8125, new_n8126);
nand_5 g07750(n8276, n6429, new_n8127);
nand_5 g07751(n12709, n10510, new_n8128);
xor_4  g07752(new_n8128, new_n8127, new_n8129);
not_8  g07753(new_n8129, new_n8130);
xor_4  g07754(new_n8130, new_n8126, new_n8131);
xor_4  g07755(new_n8131, new_n8124, new_n8132);
xor_4  g07756(new_n8132, new_n8120, new_n8133);
and_5  g07757(new_n8049, new_n8046, new_n8134);
or_5   g07758(new_n8048, new_n8047, new_n8135);
not_8  g07759(new_n8135, new_n8136);
nand_5 g07760(new_n8067, new_n8050, new_n8137);
not_8  g07761(new_n8137, new_n8138_1);
xor_4  g07762(new_n8138_1, new_n8136, new_n8139);
nor_5  g07763(new_n8139, new_n8134, new_n8140);
xor_4  g07764(new_n8140, new_n8133, new_n8141);
not_8  g07765(new_n8141, new_n8142);
xor_4  g07766(new_n8142, new_n8107, new_n8143);
not_8  g07767(new_n8143, new_n8144);
xor_4  g07768(new_n8144, new_n8106, new_n8145);
nand_5 g07769(n2393, n1478, new_n8146);
nand_5 g07770(n5860, n5760, new_n8147);
nand_5 g07771(n10990, n3986, new_n8148);
xor_4  g07772(new_n8148, new_n8147, new_n8149);
not_8  g07773(new_n8149, new_n8150);
xor_4  g07774(new_n8150, new_n8146, new_n8151);
nand_5 g07775(n11892, n1478, new_n8152);
nand_5 g07776(n10990, n5860, new_n8153);
and_5  g07777(new_n8153, new_n8152, new_n8154);
nor_5  g07778(new_n8153, new_n8152, new_n8155);
nand_5 g07779(n5760, n2393, new_n8156);
not_8  g07780(new_n8156, new_n8157);
nor_5  g07781(new_n8157, new_n8155, new_n8158);
or_5   g07782(new_n8158, new_n8154, new_n8159);
not_8  g07783(new_n8159, new_n8160);
xor_4  g07784(new_n8160, new_n8151, new_n8161);
nand_5 g07785(n12947, n7388, new_n8162);
nand_5 g07786(n11892, n11791, new_n8163);
xor_4  g07787(new_n8163, new_n8162, new_n8164);
xor_4  g07788(new_n8164, new_n8161, new_n8165);
not_8  g07789(new_n8165, new_n8166);
nand_5 g07790(n11791, n7388, new_n8167);
not_8  g07791(new_n8167, new_n8168);
nand_5 g07792(n10990, n2393, new_n8169);
nand_5 g07793(n7388, n1478, new_n8170);
and_5  g07794(new_n8170, new_n8169, new_n8171);
nor_5  g07795(new_n8170, new_n8169, new_n8172);
nand_5 g07796(n11892, n5760, new_n8173);
not_8  g07797(new_n8173, new_n8174);
nor_5  g07798(new_n8174, new_n8172, new_n8175);
or_5   g07799(new_n8175, new_n8171, new_n8176);
not_8  g07800(new_n8176, new_n8177);
and_5  g07801(new_n8177, new_n8168, new_n8178);
nor_5  g07802(new_n8177, new_n8168, new_n8179);
or_5   g07803(new_n8179, new_n8178, new_n8180);
xor_4  g07804(new_n8153, new_n8152, new_n8181);
xor_4  g07805(new_n8181, new_n8156, new_n8182);
nor_5  g07806(new_n8182, new_n8180, new_n8183);
nor_5  g07807(new_n8183, new_n8178, new_n8184);
xor_4  g07808(new_n8184, new_n8166, new_n8185);
nand_5 g07809(n12947, n7965, new_n8186);
nand_5 g07810(n11791, n7965, new_n8187);
not_8  g07811(new_n8187, new_n8188);
nor_5  g07812(new_n7887, new_n7886, new_n8189);
nor_5  g07813(new_n8189, new_n7883, new_n8190);
or_5   g07814(new_n8190, new_n7890, new_n8191);
not_8  g07815(new_n8191, new_n8192);
and_5  g07816(new_n8192, new_n8188, new_n8193);
nor_5  g07817(new_n8192, new_n8188, new_n8194);
or_5   g07818(new_n8194, new_n8193, new_n8195);
xor_4  g07819(new_n8170, new_n8169, new_n8196);
xor_4  g07820(new_n8196, new_n8173, new_n8197);
nor_5  g07821(new_n8197, new_n8195, new_n8198);
nor_5  g07822(new_n8198, new_n8193, new_n8199);
and_5  g07823(new_n8199, new_n8186, new_n8200);
xor_4  g07824(new_n8182, new_n8180, new_n8201);
not_8  g07825(new_n8201, new_n8202_1);
not_8  g07826(new_n8186, new_n8203);
xor_4  g07827(new_n8199, new_n8203, new_n8204);
not_8  g07828(new_n8204, new_n8205);
and_5  g07829(new_n8205, new_n8202_1, new_n8206);
or_5   g07830(new_n8206, new_n8200, new_n8207);
not_8  g07831(new_n8207, new_n8208);
nand_5 g07832(new_n8208, new_n8185, new_n8209);
or_5   g07833(new_n8148, new_n8147, new_n8210);
not_8  g07834(new_n8210, new_n8211);
nand_5 g07835(n11791, n2393, new_n8212);
not_8  g07836(new_n8212, new_n8213);
xor_4  g07837(new_n8213, new_n8211, new_n8214);
nand_5 g07838(n5760, n3986, new_n8215);
not_8  g07839(new_n8215, new_n8216);
nand_5 g07840(n5860, n1478, new_n8217);
nand_5 g07841(n10990, n5857, new_n8218);
xor_4  g07842(new_n8218, new_n8217, new_n8219);
xor_4  g07843(new_n8219, new_n8216, new_n8220);
xor_4  g07844(new_n8220, new_n8214, new_n8221);
not_8  g07845(new_n8221, new_n8222);
nand_5 g07846(n7388, n6441, new_n8223);
nand_5 g07847(n12947, n11892, new_n8224);
and_5  g07848(n11999, n7965, new_n8225);
xor_4  g07849(new_n8225, new_n8224, new_n8226);
not_8  g07850(new_n8226, new_n8227);
xor_4  g07851(new_n8227, new_n8223, new_n8228);
not_8  g07852(new_n8228, new_n8229);
nor_5  g07853(new_n8150, new_n8146, new_n8230);
and_5  g07854(new_n8160, new_n8151, new_n8231);
or_5   g07855(new_n8231, new_n8230, new_n8232);
xor_4  g07856(new_n8232, new_n8229, new_n8233);
xor_4  g07857(new_n8233, new_n8222, new_n8234);
nand_5 g07858(new_n8164, new_n8161, new_n8235);
or_5   g07859(new_n8163, new_n8162, new_n8236_1);
or_5   g07860(new_n8184, new_n8166, new_n8237);
not_8  g07861(new_n8237, new_n8238);
xor_4  g07862(new_n8238, new_n8236_1, new_n8239);
and_5  g07863(new_n8239, new_n8235, new_n8240);
xor_4  g07864(new_n8240, new_n8234, new_n8241);
xnor_4 g07865(new_n8241, new_n8209, new_n8242);
not_8  g07866(new_n8242, new_n8243);
nand_5 g07867(n7965, n6441, new_n8244);
not_8  g07868(new_n8244, new_n8245);
xor_4  g07869(new_n8208, new_n8185, new_n8246);
and_5  g07870(new_n8246, new_n8245, new_n8247);
nor_5  g07871(new_n8246, new_n8245, new_n8248);
xor_4  g07872(new_n8196, new_n8174, new_n8249);
xor_4  g07873(new_n8249, new_n8195, new_n8250);
not_8  g07874(new_n7883, new_n8251);
or_5   g07875(new_n7889, new_n8251, new_n8252);
or_5   g07876(new_n8252, new_n8250, new_n8253);
xor_4  g07877(new_n8205, new_n8202_1, new_n8254);
or_5   g07878(new_n8254, new_n8253, new_n8255);
nor_5  g07879(new_n8255, new_n8248, new_n8256);
nor_5  g07880(new_n8256, new_n8247, new_n8257);
xor_4  g07881(new_n8257, new_n8243, new_n8258);
not_8  g07882(new_n8258, new_n8259);
nand_5 g07883(n12777, n12648, new_n8260);
nand_5 g07884(n10545, n7159, new_n8261);
nand_5 g07885(n12489, n7690, new_n8262);
xor_4  g07886(new_n8262, new_n8261, new_n8263);
not_8  g07887(new_n8263, new_n8264);
xor_4  g07888(new_n8264, new_n8260, new_n8265);
nand_5 g07889(n12489, n10545, new_n8266);
and_5  g07890(new_n8266, new_n7876, new_n8267);
nor_5  g07891(new_n8266, new_n7876, new_n8268);
nand_5 g07892(n12648, n7159, new_n8269);
not_8  g07893(new_n8269, new_n8270);
nor_5  g07894(new_n8270, new_n8268, new_n8271);
or_5   g07895(new_n8271, new_n8267, new_n8272);
not_8  g07896(new_n8272, new_n8273);
xor_4  g07897(new_n8273, new_n8265, new_n8274);
nand_5 g07898(n6254, n2530, new_n8275);
nand_5 g07899(n11967, n8476, new_n8276_1);
xor_4  g07900(new_n8276_1, new_n8275, new_n8277);
xor_4  g07901(new_n8277, new_n8274, new_n8278);
nand_5 g07902(n8476, n6254, new_n8279);
nand_5 g07903(n12648, n12489, new_n8280);
nand_5 g07904(n12777, n8476, new_n8281);
and_5  g07905(new_n8281, new_n8280, new_n8282);
nor_5  g07906(new_n8281, new_n8280, new_n8283);
nand_5 g07907(n7159, n2530, new_n8284);
not_8  g07908(new_n8284, new_n8285);
nor_5  g07909(new_n8285, new_n8283, new_n8286);
nor_5  g07910(new_n8286, new_n8282, new_n8287);
not_8  g07911(new_n8287, new_n8288);
nor_5  g07912(new_n8288, new_n8279, new_n8289);
xor_4  g07913(new_n8288, new_n8279, new_n8290);
xor_4  g07914(new_n8266, new_n7876, new_n8291);
xor_4  g07915(new_n8291, new_n8270, new_n8292);
and_5  g07916(new_n8292, new_n8290, new_n8293);
or_5   g07917(new_n8293, new_n8289, new_n8294);
xor_4  g07918(new_n8294, new_n8278, new_n8295);
nand_5 g07919(n11967, n5331, new_n8296);
not_8  g07920(new_n8296, new_n8297);
xor_4  g07921(new_n8292, new_n8290, new_n8298);
nor_5  g07922(new_n8298, new_n8297, new_n8299);
xor_4  g07923(new_n8298, new_n8297, new_n8300);
nand_5 g07924(n6254, n5331, new_n8301);
not_8  g07925(new_n7870, new_n8302);
nor_5  g07926(new_n7877, new_n8302, new_n8303_1);
nor_5  g07927(new_n8303_1, new_n7875, new_n8304);
not_8  g07928(new_n8304, new_n8305);
nor_5  g07929(new_n8305, new_n8301, new_n8306);
not_8  g07930(new_n8301, new_n8307);
xor_4  g07931(new_n8305, new_n8307, new_n8308);
xor_4  g07932(new_n8281, new_n8280, new_n8309);
xor_4  g07933(new_n8309, new_n8284, new_n8310);
nor_5  g07934(new_n8310, new_n8308, new_n8311);
or_5   g07935(new_n8311, new_n8306, new_n8312);
not_8  g07936(new_n8312, new_n8313);
and_5  g07937(new_n8313, new_n8300, new_n8314);
or_5   g07938(new_n8314, new_n8299, new_n8315);
not_8  g07939(new_n8315, new_n8316);
nand_5 g07940(new_n8316, new_n8295, new_n8317);
nand_5 g07941(n5331, n1353, new_n8318);
not_8  g07942(new_n8318, new_n8319);
nand_5 g07943(n11967, n2530, new_n8320);
nand_5 g07944(n8476, n447, new_n8321);
xor_4  g07945(new_n8321, new_n8320, new_n8322);
not_8  g07946(new_n8322, new_n8323);
xor_4  g07947(new_n8323, new_n8319, new_n8324);
not_8  g07948(new_n8324, new_n8325);
nor_5  g07949(new_n8264, new_n8260, new_n8326);
and_5  g07950(new_n8273, new_n8265, new_n8327);
or_5   g07951(new_n8327, new_n8326, new_n8328);
xor_4  g07952(new_n8328, new_n8325, new_n8329);
or_5   g07953(new_n8262, new_n8261, new_n8330);
not_8  g07954(new_n8330, new_n8331);
nand_5 g07955(n12648, n6254, new_n8332);
not_8  g07956(new_n8332, new_n8333);
xor_4  g07957(new_n8333, new_n8331, new_n8334);
nand_5 g07958(n7690, n7159, new_n8335);
nand_5 g07959(n12777, n10545, new_n8336_1);
nand_5 g07960(n12489, n3616, new_n8337);
xor_4  g07961(new_n8337, new_n8336_1, new_n8338);
not_8  g07962(new_n8338, new_n8339);
xor_4  g07963(new_n8339, new_n8335, new_n8340);
xor_4  g07964(new_n8340, new_n8334, new_n8341);
xor_4  g07965(new_n8341, new_n8329, new_n8342);
not_8  g07966(new_n8342, new_n8343);
and_5  g07967(new_n8277, new_n8274, new_n8344);
or_5   g07968(new_n8276_1, new_n8275, new_n8345);
not_8  g07969(new_n8345, new_n8346);
nand_5 g07970(new_n8294, new_n8278, new_n8347);
not_8  g07971(new_n8347, new_n8348);
xor_4  g07972(new_n8348, new_n8346, new_n8349);
nor_5  g07973(new_n8349, new_n8344, new_n8350);
xor_4  g07974(new_n8350, new_n8343, new_n8351);
not_8  g07975(new_n8351, new_n8352);
xor_4  g07976(new_n8352, new_n8317, new_n8353);
nand_5 g07977(n5331, n447, new_n8354);
not_8  g07978(new_n8354, new_n8355);
xor_4  g07979(new_n8316, new_n8295, new_n8356);
and_5  g07980(new_n8356, new_n8355, new_n8357);
nor_5  g07981(new_n8356, new_n8355, new_n8358);
xor_4  g07982(new_n8310, new_n8308, new_n8359);
nand_5 g07983(new_n7880, new_n8302, new_n8360);
not_8  g07984(new_n8360, new_n8361);
nand_5 g07985(new_n8361, new_n8359, new_n8362);
xnor_4 g07986(new_n8312, new_n8300, new_n8363);
or_5   g07987(new_n8363, new_n8362, new_n8364);
nor_5  g07988(new_n8364, new_n8358, new_n8365);
nor_5  g07989(new_n8365, new_n8357, new_n8366);
xor_4  g07990(new_n8366, new_n8353, new_n8367);
xor_4  g07991(new_n8367, new_n8259, new_n8368);
xor_4  g07992(new_n8246, new_n8245, new_n8369);
xor_4  g07993(new_n8369, new_n8255, new_n8370);
not_8  g07994(new_n8370, new_n8371);
not_8  g07995(new_n8364, new_n8372);
xor_4  g07996(new_n8356, new_n8355, new_n8373);
xor_4  g07997(new_n8373, new_n8372, new_n8374);
nor_5  g07998(new_n8374, new_n8371, new_n8375);
xor_4  g07999(new_n8363, new_n8362, new_n8376);
xor_4  g08000(new_n8254, new_n8253, new_n8377);
nor_5  g08001(new_n8377, new_n8376, new_n8378);
xor_4  g08002(new_n8377, new_n8376, new_n8379);
not_8  g08003(new_n8379, new_n8380);
xor_4  g08004(new_n8360, new_n8359, new_n8381);
xor_4  g08005(new_n8252, new_n8250, new_n8382);
not_8  g08006(new_n8382, new_n8383);
nor_5  g08007(new_n8383, new_n8381, new_n8384_1);
nor_5  g08008(new_n7892, new_n7882, new_n8385);
and_5  g08009(new_n7898, new_n7893, new_n8386);
or_5   g08010(new_n8386, new_n8385, new_n8387);
not_8  g08011(new_n8387, new_n8388);
xnor_4 g08012(new_n8382, new_n8381, new_n8389);
not_8  g08013(new_n8389, new_n8390);
nor_5  g08014(new_n8390, new_n8388, new_n8391);
or_5   g08015(new_n8391, new_n8384_1, new_n8392);
nor_5  g08016(new_n8392, new_n8380, new_n8393);
or_5   g08017(new_n8393, new_n8378, new_n8394);
xor_4  g08018(new_n8374, new_n8371, new_n8395);
and_5  g08019(new_n8395, new_n8394, new_n8396);
or_5   g08020(new_n8396, new_n8375, new_n8397);
xor_4  g08021(new_n8397, new_n8368, new_n8398_1);
xor_4  g08022(new_n8398_1, new_n8145, new_n8399);
xor_4  g08023(new_n8103, new_n8102, new_n8400);
not_8  g08024(new_n8400, new_n8401);
xor_4  g08025(new_n8395, new_n8394, new_n8402);
and_5  g08026(new_n8402, new_n8401, new_n8403);
xor_4  g08027(new_n8402, new_n8401, new_n8404);
not_8  g08028(new_n8404, new_n8405);
xor_4  g08029(new_n8100_1, new_n8098, new_n8406);
not_8  g08030(new_n8406, new_n8407);
xor_4  g08031(new_n8392, new_n8380, new_n8408);
nor_5  g08032(new_n8408, new_n8407, new_n8409);
xor_4  g08033(new_n8097, new_n8094, new_n8410);
xor_4  g08034(new_n8390, new_n8388, new_n8411);
and_5  g08035(new_n8411, new_n8410, new_n8412);
not_8  g08036(new_n8410, new_n8413);
xor_4  g08037(new_n8411, new_n8413, new_n8414);
not_8  g08038(new_n7899, new_n8415);
nor_5  g08039(new_n8415, new_n7868, new_n8416);
nor_5  g08040(new_n8416, new_n7866, new_n8417);
nor_5  g08041(new_n8417, new_n8414, new_n8418);
or_5   g08042(new_n8418, new_n8412, new_n8419);
not_8  g08043(new_n8419, new_n8420);
xor_4  g08044(new_n8408, new_n8407, new_n8421);
not_8  g08045(new_n8421, new_n8422);
nor_5  g08046(new_n8422, new_n8420, new_n8423);
or_5   g08047(new_n8423, new_n8409, new_n8424);
nor_5  g08048(new_n8424, new_n8405, new_n8425);
nor_5  g08049(new_n8425, new_n8403, new_n8426);
xor_4  g08050(new_n8426, new_n8399, new_n8427);
nor_5  g08051(new_n8427, new_n8027, new_n8428);
xor_4  g08052(new_n8427, new_n8027, new_n8429);
not_8  g08053(new_n8429, new_n8430);
xor_4  g08054(new_n8023, new_n8022, new_n8431);
not_8  g08055(new_n8431, new_n8432);
xor_4  g08056(new_n8424, new_n8405, new_n8433_1);
and_5  g08057(new_n8433_1, new_n8432, new_n8434);
xor_4  g08058(new_n8433_1, new_n8432, new_n8435);
not_8  g08059(new_n8435, new_n8436);
xor_4  g08060(new_n8020, new_n8018, new_n8437);
xor_4  g08061(new_n8422, new_n8420, new_n8438);
nor_5  g08062(new_n8438, new_n8437, new_n8439);
xor_4  g08063(new_n8438, new_n8437, new_n8440);
not_8  g08064(new_n8440, new_n8441);
xor_4  g08065(new_n8017, new_n8014, new_n8442);
xor_4  g08066(new_n8417, new_n8414, new_n8443);
nor_5  g08067(new_n8443, new_n8442, new_n8444);
and_5  g08068(new_n7850, new_n7840, new_n8445);
not_8  g08069(new_n7900, new_n8446);
and_5  g08070(new_n8446, new_n7851, new_n8447);
or_5   g08071(new_n8447, new_n8445, new_n8448);
xor_4  g08072(new_n8443, new_n8442, new_n8449);
not_8  g08073(new_n8449, new_n8450);
nor_5  g08074(new_n8450, new_n8448, new_n8451);
or_5   g08075(new_n8451, new_n8444, new_n8452);
not_8  g08076(new_n8452, new_n8453);
nor_5  g08077(new_n8453, new_n8441, new_n8454);
or_5   g08078(new_n8454, new_n8439, new_n8455);
not_8  g08079(new_n8455, new_n8456);
nor_5  g08080(new_n8456, new_n8436, new_n8457);
or_5   g08081(new_n8457, new_n8434, new_n8458);
nor_5  g08082(new_n8458, new_n8430, new_n8459);
nor_5  g08083(new_n8459, new_n8428, new_n8460);
not_8  g08084(new_n8145, new_n8461);
and_5  g08085(new_n8398_1, new_n8461, new_n8462);
nor_5  g08086(new_n8426, new_n8399, new_n8463);
nor_5  g08087(new_n8463, new_n8462, new_n8464);
nor_5  g08088(new_n8025, new_n8009, new_n8465);
or_5   g08089(new_n8465, new_n8007, new_n8466);
and_5  g08090(new_n7992, new_n7991, new_n8467);
nor_5  g08091(new_n7994, new_n7990, new_n8468);
nor_5  g08092(new_n8468, new_n8467, new_n8469);
and_5  g08093(new_n7977, new_n7976, new_n8470);
nor_5  g08094(new_n7979, new_n7975, new_n8471);
or_5   g08095(new_n8471, new_n8470, new_n8472);
and_5  g08096(n9725, n5964, new_n8473);
xor_4  g08097(new_n8473, new_n8472, new_n8474);
xor_4  g08098(new_n8474, new_n8469, new_n8475);
xor_4  g08099(new_n8475, new_n8466, new_n8476_1);
nor_5  g08100(new_n8142, new_n8107, new_n8477);
nor_5  g08101(new_n8144, new_n8106, new_n8478);
nor_5  g08102(new_n8478, new_n8477, new_n8479);
nor_5  g08103(new_n8352, new_n8317, new_n8480);
not_8  g08104(new_n8353, new_n8481);
nor_5  g08105(new_n8366, new_n8481, new_n8482);
nor_5  g08106(new_n8482, new_n8480, new_n8483);
xor_4  g08107(new_n8483, new_n8479, new_n8484);
not_8  g08108(new_n8241, new_n8485);
nor_5  g08109(new_n8485, new_n8209, new_n8486);
nor_5  g08110(new_n8257, new_n8243, new_n8487);
nor_5  g08111(new_n8487, new_n8486, new_n8488);
or_5   g08112(new_n8328, new_n8325, new_n8489);
not_8  g08113(new_n8341, new_n8490);
nand_5 g08114(new_n8490, new_n8329, new_n8491);
nand_5 g08115(new_n8491, new_n8489, new_n8492);
nor_5  g08116(new_n8114, new_n8113, new_n8493);
and_5  g08117(new_n8114, new_n8113, new_n8494);
nor_5  g08118(new_n8494, new_n8112, new_n8495);
or_5   g08119(new_n8495, new_n8493, new_n8496);
and_5  g08120(n3986, n1478, new_n8497);
nand_5 g08121(n9241, n6429, new_n8498);
and_5  g08122(n10022, n7965, new_n8499);
xor_4  g08123(new_n8499, new_n8498, new_n8500);
xor_4  g08124(new_n8500, new_n8497, new_n8501);
xor_4  g08125(new_n8501, new_n8496, new_n8502);
xor_4  g08126(new_n8502, new_n8492, new_n8503);
and_5  g08127(new_n8337, new_n8336_1, new_n8504);
not_8  g08128(new_n8335, new_n8505);
nor_5  g08129(new_n8339, new_n8505, new_n8506);
or_5   g08130(new_n8506, new_n8504, new_n8507);
and_5  g08131(new_n8227, new_n8223, new_n8508);
or_5   g08132(new_n8508, new_n8224, new_n8509);
not_8  g08133(new_n8509, new_n8510);
and_5  g08134(n11999, n7388, new_n8511);
and_5  g08135(new_n8511, new_n8510, new_n8512);
and_5  g08136(new_n8511, new_n8244, new_n8513);
nor_5  g08137(new_n8513, new_n8510, new_n8514);
nor_5  g08138(new_n8514, new_n8512, new_n8515);
xor_4  g08139(new_n8515, new_n8507, new_n8516);
and_5  g08140(new_n8333, new_n8331, new_n8517);
and_5  g08141(new_n8340, new_n8334, new_n8518);
or_5   g08142(new_n8518, new_n8517, new_n8519);
nor_5  g08143(new_n8218, new_n8217, new_n8520);
and_5  g08144(new_n8218, new_n8217, new_n8521);
nor_5  g08145(new_n8521, new_n8215, new_n8522);
or_5   g08146(new_n8522, new_n8520, new_n8523);
and_5  g08147(n2530, n447, new_n8524);
nand_5 g08148(n12777, n7690, new_n8525);
and_5  g08149(n8476, n1353, new_n8526);
xor_4  g08150(new_n8526, new_n8525, new_n8527);
xor_4  g08151(new_n8527, new_n8524, new_n8528);
xor_4  g08152(new_n8528, new_n8523, new_n8529);
xor_4  g08153(new_n8529, new_n8519, new_n8530);
xor_4  g08154(new_n8530, new_n8516, new_n8531);
and_5  g08155(n8759, n1198, new_n8532);
and_5  g08156(n11728, n10510, new_n8533);
xor_4  g08157(new_n8533, new_n8532, new_n8534);
nand_5 g08158(n12489, n4499, new_n8535);
and_5  g08159(n10545, n6254, new_n8536);
xor_4  g08160(new_n8536, new_n8535, new_n8537);
nand_5 g08161(n5331, n4436, new_n8538);
and_5  g08162(n12947, n2393, new_n8539);
xor_4  g08163(new_n8539, new_n8538, new_n8540);
xor_4  g08164(new_n8540, new_n8537, new_n8541);
xor_4  g08165(new_n8541, new_n8534, new_n8542);
and_5  g08166(n12648, n11967, new_n8543);
nand_5 g08167(n7159, n3616, new_n8544);
and_5  g08168(n12709, n10644, new_n8545);
xor_4  g08169(new_n8545, new_n8544, new_n8546);
xor_4  g08170(new_n8546, new_n8543, new_n8547);
nand_5 g08171(n8819, n8276, new_n8548);
and_5  g08172(n7730, n6776, new_n8549);
xor_4  g08173(new_n8549, new_n8548, new_n8550);
xor_4  g08174(new_n8550, new_n8547, new_n8551);
xor_4  g08175(new_n8551, new_n8542, new_n8552);
xor_4  g08176(new_n8552, new_n8531, new_n8553);
xor_4  g08177(new_n8553, new_n8503, new_n8554);
not_8  g08178(new_n8236_1, new_n8555);
nand_5 g08179(new_n8238, new_n8555, new_n8556);
not_8  g08180(new_n8556, new_n8557);
nor_5  g08181(new_n8240, new_n8234, new_n8558);
nor_5  g08182(new_n8558, new_n8557, new_n8559);
and_5  g08183(n12705, n4370, new_n8560);
nor_5  g08184(new_n7997, new_n7984, new_n8561);
or_5   g08185(new_n8561, new_n7982, new_n8562);
nor_5  g08186(new_n8232, new_n8229, new_n8563);
and_5  g08187(new_n8233, new_n8222, new_n8564);
nor_5  g08188(new_n8564, new_n8563, new_n8565);
xor_4  g08189(new_n8565, new_n8562, new_n8566);
xor_4  g08190(new_n8566, new_n8560, new_n8567);
xor_4  g08191(new_n8567, new_n8559, new_n8568);
xor_4  g08192(new_n8568, new_n8554, new_n8569);
xor_4  g08193(new_n8569, new_n8488, new_n8570);
xor_4  g08194(new_n8570, new_n8484, new_n8571);
xor_4  g08195(new_n8571, new_n8476_1, new_n8572);
and_5  g08196(new_n8367, new_n8259, new_n8573);
and_5  g08197(new_n8397, new_n8368, new_n8574);
nor_5  g08198(new_n8574, new_n8573, new_n8575);
and_5  g08199(new_n8138_1, new_n8136, new_n8576);
nor_5  g08200(new_n8140, new_n8133, new_n8577);
nor_5  g08201(new_n8577, new_n8576, new_n8578);
and_5  g08202(n11407, n10547, new_n8579);
and_5  g08203(n5320, n4312, new_n8580);
xor_4  g08204(new_n8580, new_n8579, new_n8581);
nand_5 g08205(n12299, n8717, new_n8582);
and_5  g08206(n5857, n5760, new_n8583);
xor_4  g08207(new_n8583, new_n8582, new_n8584);
nand_5 g08208(n12025, n11877, new_n8585);
and_5  g08209(n12000, n1097, new_n8586);
xor_4  g08210(new_n8586, new_n8585, new_n8587);
xor_4  g08211(new_n8587, new_n8584, new_n8588);
xor_4  g08212(new_n8588, new_n8581, new_n8589);
and_5  g08213(new_n8128, new_n8127, new_n8590);
nor_5  g08214(new_n8130, new_n8126, new_n8591);
nor_5  g08215(new_n8591, new_n8590, new_n8592);
and_5  g08216(n10990, n45, new_n8593);
xor_4  g08217(new_n8593, new_n8592, new_n8594);
xor_4  g08218(new_n8594, new_n8589, new_n8595_1);
nor_5  g08219(new_n8122, new_n8121, new_n8596);
nor_5  g08220(new_n8131, new_n8124, new_n8597);
nor_5  g08221(new_n8597, new_n8596, new_n8598);
and_5  g08222(n7436, n2433, new_n8599);
xor_4  g08223(new_n8599, new_n8598, new_n8600);
xor_4  g08224(new_n8600, new_n8595_1, new_n8601);
and_5  g08225(new_n8321, new_n8320, new_n8602);
nor_5  g08226(new_n8323, new_n8319, new_n8603);
nor_5  g08227(new_n8603, new_n8602, new_n8604);
nor_5  g08228(new_n8132, new_n8120, new_n8605);
nor_5  g08229(new_n8605, new_n8118, new_n8606);
xor_4  g08230(new_n8606, new_n8604, new_n8607);
xor_4  g08231(new_n8607, new_n8601, new_n8608);
xor_4  g08232(new_n8608, new_n8578, new_n8609);
and_5  g08233(new_n8348, new_n8346, new_n8610);
nor_5  g08234(new_n8350, new_n8343, new_n8611);
nor_5  g08235(new_n8611, new_n8610, new_n8612);
and_5  g08236(new_n8213, new_n8211, new_n8613);
and_5  g08237(new_n8220, new_n8214, new_n8614);
or_5   g08238(new_n8614, new_n8613, new_n8615);
nand_5 g08239(n11892, n6441, new_n8616);
and_5  g08240(n11791, n5860, new_n8617);
xor_4  g08241(new_n8617, new_n8616, new_n8618);
and_5  g08242(n11257, n5212, new_n8619);
and_5  g08243(n6604, n5305, new_n8620);
xor_4  g08244(new_n8620, new_n8619, new_n8621);
xor_4  g08245(new_n8621, new_n8618, new_n8622);
xor_4  g08246(new_n8622, new_n8615, new_n8623);
xor_4  g08247(new_n8623, new_n8612, new_n8624);
xor_4  g08248(new_n8624, new_n8609, new_n8625);
nor_5  g08249(new_n7987, new_n7986, new_n8626);
and_5  g08250(new_n7995, new_n7988, new_n8627);
nor_5  g08251(new_n8627, new_n8626, new_n8628);
and_5  g08252(new_n8002, new_n8001, new_n8629);
nor_5  g08253(new_n8004, new_n7998, new_n8630);
nor_5  g08254(new_n8630, new_n8629, new_n8631);
xor_4  g08255(new_n8631, new_n8628, new_n8632);
xor_4  g08256(new_n8632, new_n8625, new_n8633);
xor_4  g08257(new_n8633, new_n8575, new_n8634);
xor_4  g08258(new_n8634, new_n8572, new_n8635);
xor_4  g08259(new_n8635, new_n8464, new_n8636);
xor_4  g08260(new_n8636, new_n8460, n3287);
xor_4  g08261(new_n8455, new_n8436, n3339);
xor_4  g08262(new_n3813, new_n3812, n3456);
nand_5 g08263(n6687, n4005, new_n8640);
not_8  g08264(new_n8640, new_n8641);
nand_5 g08265(n12720, n6770, new_n8642);
not_8  g08266(new_n8642, new_n8643);
nand_5 g08267(n9920, n2509, new_n8644);
nand_5 g08268(n6038, n3627, new_n8645);
xor_4  g08269(new_n8645, new_n8644, new_n8646);
xor_4  g08270(new_n8646, new_n8643, new_n8647);
not_8  g08271(new_n8647, new_n8648);
nand_5 g08272(n9920, n6038, new_n8649);
nand_5 g08273(n12720, n4189, new_n8650);
and_5  g08274(new_n8650, new_n8649, new_n8651);
nand_5 g08275(n6770, n2509, new_n8652);
not_8  g08276(new_n8652, new_n8653);
xor_4  g08277(new_n8650, new_n8649, new_n8654);
not_8  g08278(new_n8654, new_n8655);
nor_5  g08279(new_n8655, new_n8653, new_n8656);
nor_5  g08280(new_n8656, new_n8651, new_n8657);
xor_4  g08281(new_n8657, new_n8648, new_n8658);
not_8  g08282(new_n8658, new_n8659);
nand_5 g08283(n2564, n2508, new_n8660);
not_8  g08284(new_n8660, new_n8661);
nand_5 g08285(n6770, n6038, new_n8662);
nand_5 g08286(n4189, n2509, new_n8663);
and_5  g08287(new_n8663, new_n8662, new_n8664);
nand_5 g08288(n12720, n2564, new_n8665_1);
xnor_4 g08289(new_n8663, new_n8662, new_n8666);
not_8  g08290(new_n8666, new_n8667);
and_5  g08291(new_n8667, new_n8665_1, new_n8668);
or_5   g08292(new_n8668, new_n8664, new_n8669);
not_8  g08293(new_n8669, new_n8670);
and_5  g08294(new_n8670, new_n8661, new_n8671);
xor_4  g08295(new_n8655, new_n8653, new_n8672);
not_8  g08296(new_n8672, new_n8673);
xor_4  g08297(new_n8670, new_n8661, new_n8674);
and_5  g08298(new_n8674, new_n8673, new_n8675);
or_5   g08299(new_n8675, new_n8671, new_n8676);
not_8  g08300(new_n8676, new_n8677);
nand_5 g08301(n2585, n2564, new_n8678);
nand_5 g08302(n4189, n2508, new_n8679);
xor_4  g08303(new_n8679, new_n8678, new_n8680);
not_8  g08304(new_n8680, new_n8681);
xor_4  g08305(new_n8681, new_n8677, new_n8682);
xor_4  g08306(new_n8682, new_n8659, new_n8683);
nand_5 g08307(n6687, n2585, new_n8684);
nand_5 g08308(n6687, n2508, new_n8685);
nor_5  g08309(new_n8650, new_n377, new_n8686);
and_5  g08310(n6038, n4189, new_n8687);
and_5  g08311(n12720, n6687, new_n8688);
nor_5  g08312(new_n8688, new_n8687, new_n8689);
nand_5 g08313(n2564, n2509, new_n8690);
nor_5  g08314(new_n8690, new_n8689, new_n8691);
nor_5  g08315(new_n8691, new_n8686, new_n8692);
nor_5  g08316(new_n8692, new_n8685, new_n8693);
not_8  g08317(new_n8685, new_n8694);
xor_4  g08318(new_n8692, new_n8694, new_n8695);
not_8  g08319(new_n8695, new_n8696);
not_8  g08320(new_n8665_1, new_n8697);
xor_4  g08321(new_n8667, new_n8697, new_n8698);
and_5  g08322(new_n8698, new_n8696, new_n8699);
nor_5  g08323(new_n8699, new_n8693, new_n8700);
and_5  g08324(new_n8700, new_n8684, new_n8701);
xor_4  g08325(new_n8674, new_n8673, new_n8702);
not_8  g08326(new_n8702, new_n8703);
not_8  g08327(new_n8684, new_n8704);
xor_4  g08328(new_n8700, new_n8704, new_n8705);
not_8  g08329(new_n8705, new_n8706);
and_5  g08330(new_n8706, new_n8703, new_n8707);
or_5   g08331(new_n8707, new_n8701, new_n8708);
not_8  g08332(new_n8708, new_n8709);
xor_4  g08333(new_n8709, new_n8683, new_n8710);
and_5  g08334(new_n8710, new_n8641, new_n8711);
nor_5  g08335(new_n8698, new_n8696, new_n8712);
or_5   g08336(new_n8712, new_n8699, new_n8713);
nor_5  g08337(new_n8689, new_n8686, new_n8714);
nand_5 g08338(n6687, n2509, new_n8715);
nand_5 g08339(n6038, n2564, new_n8716);
or_5   g08340(new_n8716, new_n8715, new_n8717_1);
or_5   g08341(new_n8717_1, new_n8714, new_n8718);
or_5   g08342(new_n8718, new_n8713, new_n8719);
xor_4  g08343(new_n8706, new_n8703, new_n8720);
or_5   g08344(new_n8720, new_n8719, new_n8721);
xor_4  g08345(new_n8710, new_n8641, new_n8722);
not_8  g08346(new_n8722, new_n8723);
nor_5  g08347(new_n8723, new_n8721, new_n8724);
or_5   g08348(new_n8724, new_n8711, new_n8725);
not_8  g08349(new_n8725, new_n8726);
nand_5 g08350(new_n8709, new_n8683, new_n8727);
nor_5  g08351(new_n8646, new_n8643, new_n8728);
nor_5  g08352(new_n8657, new_n8648, new_n8729);
or_5   g08353(new_n8729, new_n8728, new_n8730);
not_8  g08354(new_n8730, new_n8731);
nand_5 g08355(n4005, n2564, new_n8732);
not_8  g08356(new_n8732, new_n8733);
nand_5 g08357(n4189, n2585, new_n8734);
nand_5 g08358(n12706, n6687, new_n8735);
xor_4  g08359(new_n8735, new_n8734, new_n8736);
not_8  g08360(new_n8736, new_n8737);
xor_4  g08361(new_n8737, new_n8733, new_n8738);
not_8  g08362(new_n8738, new_n8739);
xor_4  g08363(new_n8739, new_n8731, new_n8740);
or_5   g08364(new_n8645, new_n8644, new_n8741);
not_8  g08365(new_n8741, new_n8742);
and_5  g08366(n6770, n2508, new_n8743);
xor_4  g08367(new_n8743, new_n8742, new_n8744);
nand_5 g08368(n3627, n2509, new_n8745);
nand_5 g08369(n12720, n9920, new_n8746);
nand_5 g08370(n6038, n4516, new_n8747);
xor_4  g08371(new_n8747, new_n8746, new_n8748);
xor_4  g08372(new_n8748, new_n8745, new_n8749);
not_8  g08373(new_n8749, new_n8750);
xnor_4 g08374(new_n8750, new_n8744, new_n8751);
xor_4  g08375(new_n8751, new_n8740, new_n8752);
nor_5  g08376(new_n8681, new_n8677, new_n8753);
or_5   g08377(new_n8679, new_n8678, new_n8754);
nand_5 g08378(new_n8682, new_n8659, new_n8755);
xor_4  g08379(new_n8755, new_n8754, new_n8756);
nor_5  g08380(new_n8756, new_n8753, new_n8757);
xor_4  g08381(new_n8757, new_n8752, new_n8758);
not_8  g08382(new_n8758, new_n8759_1);
xor_4  g08383(new_n8759_1, new_n8727, new_n8760);
not_8  g08384(new_n8760, new_n8761);
xor_4  g08385(new_n8761, new_n8726, new_n8762);
not_8  g08386(new_n8762, new_n8763);
nand_5 g08387(n8336, n5105, new_n8764);
nand_5 g08388(n10928, n7500, new_n8765);
nand_5 g08389(n8336, n1209, new_n8766);
nand_5 g08390(n7354, n6986, new_n8767);
nand_5 g08391(new_n8767, new_n8766, new_n8768);
not_8  g08392(new_n8768, new_n8769);
nor_5  g08393(new_n8769, new_n8765, new_n8770);
nor_5  g08394(new_n8767, new_n8766, new_n8771);
nor_5  g08395(new_n8771, new_n8770, new_n8772);
xor_4  g08396(new_n8772, new_n8764, new_n8773);
not_8  g08397(new_n8773, new_n8774);
nand_5 g08398(n7500, n6986, new_n8775);
not_8  g08399(new_n8775, new_n8776);
nand_5 g08400(n7354, n2226, new_n8777);
nand_5 g08401(n10928, n1209, new_n8778);
xor_4  g08402(new_n8778, new_n8777, new_n8779);
xor_4  g08403(new_n8779, new_n8776, new_n8780);
not_8  g08404(new_n8780, new_n8781);
xor_4  g08405(new_n8781, new_n8774, new_n8782);
xor_4  g08406(new_n8767, new_n8766, new_n8783);
nand_5 g08407(n10928, n7354, new_n8784);
nand_5 g08408(n8336, n7500, new_n8785);
or_5   g08409(new_n8785, new_n8784, new_n8786);
or_5   g08410(new_n8786, new_n8783, new_n8787);
not_8  g08411(new_n8787, new_n8788);
nand_5 g08412(new_n8788, new_n8782, new_n8789);
nand_5 g08413(n8336, n4141, new_n8790);
not_8  g08414(new_n8790, new_n8791);
nor_5  g08415(new_n8772, new_n8764, new_n8792);
nor_5  g08416(new_n8781, new_n8774, new_n8793);
or_5   g08417(new_n8793, new_n8792, new_n8794);
not_8  g08418(new_n8794, new_n8795);
xor_4  g08419(new_n8795, new_n8791, new_n8796);
and_5  g08420(n10928, n5105, new_n8797);
and_5  g08421(new_n8778, new_n8777, new_n8798);
nor_5  g08422(new_n8778, new_n8777, new_n8799);
nor_5  g08423(new_n8799, new_n8776, new_n8800);
or_5   g08424(new_n8800, new_n8798, new_n8801);
not_8  g08425(new_n8801, new_n8802);
and_5  g08426(new_n8802, new_n8797, new_n8803);
nor_5  g08427(new_n8802, new_n8797, new_n8804);
or_5   g08428(new_n8804, new_n8803, new_n8805);
nand_5 g08429(n6986, n1209, new_n8806);
not_8  g08430(new_n8806, new_n8807);
nand_5 g08431(n7354, n1094, new_n8808);
nand_5 g08432(n7500, n2226, new_n8809);
xor_4  g08433(new_n8809, new_n8808, new_n8810);
not_8  g08434(new_n8810, new_n8811);
xor_4  g08435(new_n8811, new_n8807, new_n8812);
xor_4  g08436(new_n8812, new_n8805, new_n8813);
xor_4  g08437(new_n8813, new_n8796, new_n8814);
or_5   g08438(new_n8814, new_n8789, new_n8815);
nand_5 g08439(n8336, n4928, new_n8816);
nand_5 g08440(n2226, n1209, new_n8817);
not_8  g08441(new_n8817, new_n8818);
and_5  g08442(new_n8809, new_n8808, new_n8819_1);
nor_5  g08443(new_n8811, new_n8807, new_n8820);
or_5   g08444(new_n8820, new_n8819_1, new_n8821);
not_8  g08445(new_n8821, new_n8822);
xor_4  g08446(new_n8822, new_n8818, new_n8823);
nand_5 g08447(n7500, n1094, new_n8824);
nand_5 g08448(n10678, n7354, new_n8825);
xor_4  g08449(new_n8825, new_n8824, new_n8826);
xor_4  g08450(new_n8826, new_n8823, new_n8827);
not_8  g08451(new_n8827, new_n8828);
nand_5 g08452(n10928, n4141, new_n8829);
nand_5 g08453(n6986, n5105, new_n8830);
xor_4  g08454(new_n8830, new_n8829, new_n8831);
not_8  g08455(new_n8831, new_n8832);
xor_4  g08456(new_n8832, new_n8828, new_n8833);
nor_5  g08457(new_n8812, new_n8805, new_n8834);
or_5   g08458(new_n8834, new_n8803, new_n8835);
xor_4  g08459(new_n8835, new_n8833, new_n8836);
not_8  g08460(new_n8836, new_n8837);
and_5  g08461(new_n8795, new_n8790, new_n8838);
nor_5  g08462(new_n8813, new_n8796, new_n8839);
or_5   g08463(new_n8839, new_n8838, new_n8840);
not_8  g08464(new_n8840, new_n8841);
xor_4  g08465(new_n8841, new_n8837, new_n8842);
xor_4  g08466(new_n8842, new_n8816, new_n8843);
xor_4  g08467(new_n8843, new_n8815, new_n8844);
nand_5 g08468(n11222, n7294, new_n8845);
nand_5 g08469(n11222, n1980, new_n8846);
nand_5 g08470(n8028, n5314, new_n8847);
nor_5  g08471(new_n8847, new_n8846, new_n8848);
and_5  g08472(new_n8847, new_n8846, new_n8849);
nand_5 g08473(n11153, n10848, new_n8850);
nor_5  g08474(new_n8850, new_n8849, new_n8851);
nor_5  g08475(new_n8851, new_n8848, new_n8852);
xor_4  g08476(new_n8852, new_n8845, new_n8853);
not_8  g08477(new_n8853, new_n8854);
and_5  g08478(n10848, n5314, new_n8855);
nand_5 g08479(n8028, n996, new_n8856);
nand_5 g08480(n11153, n1980, new_n8857);
xor_4  g08481(new_n8857, new_n8856, new_n8858);
xor_4  g08482(new_n8858, new_n8855, new_n8859);
not_8  g08483(new_n8859, new_n8860);
or_5   g08484(new_n8860, new_n8854, new_n8861);
nand_5 g08485(new_n8860, new_n8854, new_n8862);
and_5  g08486(new_n8862, new_n8861, new_n8863);
xor_4  g08487(new_n8847, new_n8846, new_n8864);
and_5  g08488(n11153, n8028, new_n8865);
and_5  g08489(n11222, n10848, new_n8866);
nand_5 g08490(new_n8866, new_n8865, new_n8867);
or_5   g08491(new_n8867, new_n8864, new_n8868);
not_8  g08492(new_n8868, new_n8869);
nand_5 g08493(new_n8869, new_n8863, new_n8870);
nor_5  g08494(new_n8852, new_n8845, new_n8871);
nor_5  g08495(new_n8860, new_n8854, new_n8872);
or_5   g08496(new_n8872, new_n8871, new_n8873);
nand_5 g08497(n12704, n11222, new_n8874);
not_8  g08498(new_n8874, new_n8875);
nand_5 g08499(n11153, n7294, new_n8876);
not_8  g08500(new_n8876, new_n8877);
and_5  g08501(new_n8857, new_n8856, new_n8878);
nor_5  g08502(new_n8857, new_n8856, new_n8879);
nor_5  g08503(new_n8879, new_n8855, new_n8880);
nor_5  g08504(new_n8880, new_n8878, new_n8881);
not_8  g08505(new_n8881, new_n8882);
xor_4  g08506(new_n8882, new_n8877, new_n8883);
nand_5 g08507(n10848, n996, new_n8884);
not_8  g08508(new_n8884, new_n8885);
nand_5 g08509(n5314, n1980, new_n8886);
nand_5 g08510(n8028, n5767, new_n8887);
xor_4  g08511(new_n8887, new_n8886, new_n8888);
xor_4  g08512(new_n8888, new_n8885, new_n8889);
not_8  g08513(new_n8889, new_n8890);
or_5   g08514(new_n8890, new_n8883, new_n8891);
nand_5 g08515(new_n8890, new_n8883, new_n8892);
and_5  g08516(new_n8892, new_n8891, new_n8893);
xor_4  g08517(new_n8893, new_n8875, new_n8894);
not_8  g08518(new_n8894, new_n8895);
xor_4  g08519(new_n8895, new_n8873, new_n8896);
or_5   g08520(new_n8896, new_n8870, new_n8897);
not_8  g08521(new_n8897, new_n8898);
nand_5 g08522(n11222, n5814, new_n8899);
not_8  g08523(new_n8899, new_n8900);
nand_5 g08524(n1980, n996, new_n8901);
nand_5 g08525(n8028, n5319, new_n8902);
nand_5 g08526(n10848, n5767, new_n8903);
xor_4  g08527(new_n8903, new_n8902, new_n8904);
not_8  g08528(new_n8904, new_n8905);
xor_4  g08529(new_n8905, new_n8901, new_n8906);
and_5  g08530(new_n8887, new_n8886, new_n8907);
nor_5  g08531(new_n8887, new_n8886, new_n8908);
nor_5  g08532(new_n8908, new_n8885, new_n8909);
or_5   g08533(new_n8909, new_n8907, new_n8910);
not_8  g08534(new_n8910, new_n8911);
xor_4  g08535(new_n8911, new_n8906, new_n8912);
nand_5 g08536(n12704, n11153, new_n8913);
nand_5 g08537(n7294, n5314, new_n8914);
xor_4  g08538(new_n8914, new_n8913, new_n8915);
xor_4  g08539(new_n8915, new_n8912, new_n8916);
or_5   g08540(new_n8882, new_n8876, new_n8917);
nand_5 g08541(new_n8891, new_n8917, new_n8918);
xor_4  g08542(new_n8918, new_n8916, new_n8919);
not_8  g08543(new_n8919, new_n8920);
nor_5  g08544(new_n8893, new_n8875, new_n8921);
nor_5  g08545(new_n8895, new_n8873, new_n8922);
nor_5  g08546(new_n8922, new_n8921, new_n8923);
not_8  g08547(new_n8923, new_n8924);
xor_4  g08548(new_n8924, new_n8920, new_n8925);
xor_4  g08549(new_n8925, new_n8900, new_n8926);
xor_4  g08550(new_n8926, new_n8898, new_n8927);
nand_5 g08551(n12069, n2802, new_n8928);
nand_5 g08552(n7891, n1564, new_n8929);
nand_5 g08553(n12069, n533, new_n8930);
and_5  g08554(new_n8930, new_n8929, new_n8931);
nand_5 g08555(n12391, n1512, new_n8932);
or_5   g08556(new_n8932, new_n8931, new_n8933);
not_8  g08557(new_n8933, new_n8934);
nor_5  g08558(new_n8930, new_n8929, new_n8935);
nor_5  g08559(new_n8935, new_n8934, new_n8936);
xor_4  g08560(new_n8936, new_n8928, new_n8937);
and_5  g08561(n7891, n1512, new_n8938);
nand_5 g08562(n7160, n1564, new_n8939);
and_5  g08563(n12391, n533, new_n8940);
xor_4  g08564(new_n8940, new_n8939, new_n8941);
not_8  g08565(new_n8941, new_n8942);
xor_4  g08566(new_n8942, new_n8938, new_n8943);
xor_4  g08567(new_n8943, new_n8937, new_n8944);
not_8  g08568(new_n8944, new_n8945);
xor_4  g08569(new_n8930, new_n8929, new_n8946);
nand_5 g08570(n12391, n1564, new_n8947);
nand_5 g08571(n12069, n1512, new_n8948);
or_5   g08572(new_n8948, new_n8947, new_n8949);
or_5   g08573(new_n8949, new_n8946, new_n8950);
or_5   g08574(new_n8950, new_n8945, new_n8951);
nand_5 g08575(n12069, n6806, new_n8952);
nand_5 g08576(n12391, n2802, new_n8953);
not_8  g08577(new_n8953, new_n8954);
nand_5 g08578(n12391, n533, new_n8955);
and_5  g08579(new_n8955, new_n8939, new_n8956);
not_8  g08580(new_n8938, new_n8957);
and_5  g08581(new_n8942, new_n8957, new_n8958);
nor_5  g08582(new_n8958, new_n8956, new_n8959);
not_8  g08583(new_n8959, new_n8960);
xor_4  g08584(new_n8960, new_n8954, new_n8961);
nand_5 g08585(n7891, n533, new_n8962);
not_8  g08586(new_n8962, new_n8963);
nand_5 g08587(n4828, n1564, new_n8964);
nand_5 g08588(n7160, n1512, new_n8965);
xor_4  g08589(new_n8965, new_n8964, new_n8966);
not_8  g08590(new_n8966, new_n8967);
xor_4  g08591(new_n8967, new_n8963, new_n8968);
xor_4  g08592(new_n8968, new_n8961, new_n8969);
xor_4  g08593(new_n8969, new_n8952, new_n8970);
not_8  g08594(new_n8970, new_n8971);
nor_5  g08595(new_n8936, new_n8928, new_n8972);
and_5  g08596(new_n8943, new_n8937, new_n8973);
or_5   g08597(new_n8973, new_n8972, new_n8974);
not_8  g08598(new_n8974, new_n8975);
xor_4  g08599(new_n8975, new_n8971, new_n8976);
nor_5  g08600(new_n8976, new_n8951, new_n8977);
not_8  g08601(new_n8977, new_n8978);
nand_5 g08602(n12069, n5069, new_n8979);
nand_5 g08603(n7160, n533, new_n8980);
nand_5 g08604(n2515, n1564, new_n8981);
nand_5 g08605(n4828, n1512, new_n8982);
xor_4  g08606(new_n8982, new_n8981, new_n8983);
not_8  g08607(new_n8983, new_n8984);
xor_4  g08608(new_n8984, new_n8980, new_n8985);
and_5  g08609(new_n8965, new_n8964, new_n8986);
nor_5  g08610(new_n8967, new_n8963, new_n8987);
or_5   g08611(new_n8987, new_n8986, new_n8988);
not_8  g08612(new_n8988, new_n8989);
xor_4  g08613(new_n8989, new_n8985, new_n8990);
nand_5 g08614(n7891, n2802, new_n8991);
nand_5 g08615(n12391, n6806, new_n8992);
xor_4  g08616(new_n8992, new_n8991, new_n8993);
xor_4  g08617(new_n8993, new_n8990, new_n8994);
not_8  g08618(new_n8994, new_n8995);
nor_5  g08619(new_n8960, new_n8953, new_n8996);
nor_5  g08620(new_n8968, new_n8961, new_n8997);
nor_5  g08621(new_n8997, new_n8996, new_n8998);
xor_4  g08622(new_n8998, new_n8995, new_n8999);
not_8  g08623(new_n8952, new_n9000);
nor_5  g08624(new_n8969, new_n9000, new_n9001);
and_5  g08625(new_n8975, new_n8971, new_n9002);
nor_5  g08626(new_n9002, new_n9001, new_n9003);
xor_4  g08627(new_n9003, new_n8999, new_n9004);
not_8  g08628(new_n9004, new_n9005);
xor_4  g08629(new_n9005, new_n8979, new_n9006);
xor_4  g08630(new_n9006, new_n8978, new_n9007);
xor_4  g08631(new_n9007, new_n8927, new_n9008);
xor_4  g08632(new_n8896, new_n8870, new_n9009);
xor_4  g08633(new_n8950, new_n8945, new_n9010);
xor_4  g08634(new_n8869, new_n8863, new_n9011);
nor_5  g08635(new_n9011, new_n9010, new_n9012);
and_5  g08636(n12391, n1512, new_n9013);
and_5  g08637(new_n9013, new_n381_1, new_n9014);
nor_5  g08638(new_n9014, new_n8946, new_n9015);
and_5  g08639(new_n8934, new_n381_1, new_n9016);
or_5   g08640(new_n9016, new_n9015, new_n9017);
and_5  g08641(n11153, n10848, new_n9018);
and_5  g08642(new_n9018, new_n380, new_n9019);
nor_5  g08643(new_n9019, new_n8864, new_n9020);
not_8  g08644(new_n9019, new_n9021);
nor_5  g08645(new_n9021, new_n8849, new_n9022);
nor_5  g08646(new_n9022, new_n9020, new_n9023);
not_8  g08647(new_n9023, new_n9024);
nor_5  g08648(new_n9024, new_n9017, new_n9025);
or_5   g08649(new_n381_1, new_n380, new_n9026);
not_8  g08650(new_n9026, new_n9027);
xor_4  g08651(new_n8866, new_n8865, new_n9028);
nor_5  g08652(new_n9028, new_n9027, new_n9029);
xor_4  g08653(new_n9028, new_n9026, new_n9030);
not_8  g08654(new_n9030, new_n9031);
xnor_4 g08655(new_n8948, new_n8947, new_n9032);
and_5  g08656(new_n9032, new_n9031, new_n9033);
or_5   g08657(new_n9033, new_n9029, new_n9034);
not_8  g08658(new_n9034, new_n9035);
xor_4  g08659(new_n9024, new_n9017, new_n9036);
and_5  g08660(new_n9036, new_n9035, new_n9037);
or_5   g08661(new_n9037, new_n9025, new_n9038);
not_8  g08662(new_n9038, new_n9039);
xor_4  g08663(new_n9011, new_n9010, new_n9040);
and_5  g08664(new_n9040, new_n9039, new_n9041);
nor_5  g08665(new_n9041, new_n9012, new_n9042);
nor_5  g08666(new_n9042, new_n9009, new_n9043);
xor_4  g08667(new_n8976, new_n8951, new_n9044);
xor_4  g08668(new_n9042, new_n9009, new_n9045);
not_8  g08669(new_n9045, new_n9046);
nor_5  g08670(new_n9046, new_n9044, new_n9047);
nor_5  g08671(new_n9047, new_n9043, new_n9048);
xor_4  g08672(new_n9048, new_n9008, new_n9049);
nor_5  g08673(new_n9049, new_n8844, new_n9050);
xor_4  g08674(new_n9049, new_n8844, new_n9051);
not_8  g08675(new_n9051, new_n9052);
xor_4  g08676(new_n8814, new_n8789, new_n9053);
not_8  g08677(new_n9053, new_n9054);
xor_4  g08678(new_n9046, new_n9044, new_n9055);
nor_5  g08679(new_n9055, new_n9054, new_n9056);
xor_4  g08680(new_n9055, new_n9053, new_n9057);
xor_4  g08681(new_n8788, new_n8782, new_n9058);
not_8  g08682(new_n9058, new_n9059);
xor_4  g08683(new_n9040, new_n9039, new_n9060);
nor_5  g08684(new_n9060, new_n9059, new_n9061);
xor_4  g08685(new_n9060, new_n9059, new_n9062);
not_8  g08686(new_n9062, new_n9063);
xor_4  g08687(new_n9036, new_n9035, new_n9064);
not_8  g08688(new_n9064, new_n9065);
not_8  g08689(new_n8765, new_n9066);
and_5  g08690(new_n9066, new_n379, new_n9067);
and_5  g08691(new_n9067, new_n8769, new_n9068);
not_8  g08692(new_n8783, new_n9069);
nor_5  g08693(new_n9067, new_n9069, new_n9070);
or_5   g08694(new_n9070, new_n9068, new_n9071);
not_8  g08695(new_n9071, new_n9072);
and_5  g08696(new_n9072, new_n9065, new_n9073);
xor_4  g08697(new_n9072, new_n9065, new_n9074);
xor_4  g08698(new_n9032, new_n9031, new_n9075);
xor_4  g08699(new_n8785, new_n8784, new_n9076);
not_8  g08700(new_n9076, new_n9077);
nor_5  g08701(new_n9077, new_n9075, new_n9078);
or_5   g08702(new_n383, new_n379, new_n9079);
not_8  g08703(new_n9079, new_n9080_1);
xor_4  g08704(new_n9077, new_n9075, new_n9081);
and_5  g08705(new_n9081, new_n9080_1, new_n9082);
or_5   g08706(new_n9082, new_n9078, new_n9083);
not_8  g08707(new_n9083, new_n9084);
and_5  g08708(new_n9084, new_n9074, new_n9085);
or_5   g08709(new_n9085, new_n9073, new_n9086);
nor_5  g08710(new_n9086, new_n9063, new_n9087);
nor_5  g08711(new_n9087, new_n9061, new_n9088);
nor_5  g08712(new_n9088, new_n9057, new_n9089);
nor_5  g08713(new_n9089, new_n9056, new_n9090);
nor_5  g08714(new_n9090, new_n9052, new_n9091);
or_5   g08715(new_n9091, new_n9050, new_n9092);
not_8  g08716(new_n9092, new_n9093);
nand_5 g08717(new_n8841, new_n8836, new_n9094);
and_5  g08718(new_n8822, new_n8818, new_n9095);
and_5  g08719(new_n8826, new_n8823, new_n9096);
or_5   g08720(new_n9096, new_n9095, new_n9097);
not_8  g08721(new_n9097, new_n9098);
nand_5 g08722(n10928, n4928, new_n9099);
not_8  g08723(new_n9099, new_n9100);
nand_5 g08724(n6986, n4141, new_n9101);
nand_5 g08725(n8336, n8236, new_n9102);
xor_4  g08726(new_n9102, new_n9101, new_n9103);
not_8  g08727(new_n9103, new_n9104);
xor_4  g08728(new_n9104, new_n9100, new_n9105);
xor_4  g08729(new_n9105, new_n9098, new_n9106);
or_5   g08730(new_n8825, new_n8824, new_n9107);
not_8  g08731(new_n9107, new_n9108);
nand_5 g08732(n5105, n2226, new_n9109);
not_8  g08733(new_n9109, new_n9110);
xor_4  g08734(new_n9110, new_n9108, new_n9111_1);
nand_5 g08735(n10678, n7500, new_n9112);
nand_5 g08736(n7354, n7320, new_n9113);
nand_5 g08737(n1209, n1094, new_n9114);
xor_4  g08738(new_n9114, new_n9113, new_n9115);
not_8  g08739(new_n9115, new_n9116);
xor_4  g08740(new_n9116, new_n9112, new_n9117);
xor_4  g08741(new_n9117, new_n9111_1, new_n9118);
xor_4  g08742(new_n9118, new_n9106, new_n9119);
not_8  g08743(new_n9119, new_n9120);
nor_5  g08744(new_n8832, new_n8828, new_n9121);
or_5   g08745(new_n8830, new_n8829, new_n9122);
not_8  g08746(new_n9122, new_n9123);
nand_5 g08747(new_n8835, new_n8833, new_n9124);
not_8  g08748(new_n9124, new_n9125);
xor_4  g08749(new_n9125, new_n9123, new_n9126);
nor_5  g08750(new_n9126, new_n9121, new_n9127);
xor_4  g08751(new_n9127, new_n9120, new_n9128);
not_8  g08752(new_n9128, new_n9129);
xor_4  g08753(new_n9129, new_n9094, new_n9130);
and_5  g08754(new_n8842, new_n8816, new_n9131);
and_5  g08755(new_n8843, new_n8815, new_n9132);
or_5   g08756(new_n9132, new_n9131, new_n9133);
not_8  g08757(new_n9133, new_n9134);
xor_4  g08758(new_n9134, new_n9130, new_n9135);
or_5   g08759(new_n8924, new_n8920, new_n9136);
nor_5  g08760(new_n8905, new_n8901, new_n9137_1);
and_5  g08761(new_n8911, new_n8906, new_n9138);
or_5   g08762(new_n9138, new_n9137_1, new_n9139);
nand_5 g08763(n11153, n5814, new_n9140);
not_8  g08764(new_n9140, new_n9141);
nand_5 g08765(n12704, n5314, new_n9142);
nand_5 g08766(n11222, n4903, new_n9143);
xor_4  g08767(new_n9143, new_n9142, new_n9144);
not_8  g08768(new_n9144, new_n9145);
xor_4  g08769(new_n9145, new_n9141, new_n9146);
not_8  g08770(new_n9146, new_n9147);
xor_4  g08771(new_n9147, new_n9139, new_n9148);
or_5   g08772(new_n8903, new_n8902, new_n9149);
not_8  g08773(new_n9149, new_n9150);
nand_5 g08774(n7294, n996, new_n9151);
not_8  g08775(new_n9151, new_n9152);
xor_4  g08776(new_n9152, new_n9150, new_n9153);
nand_5 g08777(n10848, n5319, new_n9154);
nand_5 g08778(n5767, n1980, new_n9155);
nand_5 g08779(n9457, n8028, new_n9156);
xor_4  g08780(new_n9156, new_n9155, new_n9157);
not_8  g08781(new_n9157, new_n9158);
xor_4  g08782(new_n9158, new_n9154, new_n9159);
xor_4  g08783(new_n9159, new_n9153, new_n9160);
xor_4  g08784(new_n9160, new_n9148, new_n9161);
not_8  g08785(new_n9161, new_n9162);
and_5  g08786(new_n8915, new_n8912, new_n9163);
or_5   g08787(new_n8914, new_n8913, new_n9164);
nand_5 g08788(new_n8918, new_n8916, new_n9165);
xor_4  g08789(new_n9165, new_n9164, new_n9166);
nor_5  g08790(new_n9166, new_n9163, new_n9167);
xor_4  g08791(new_n9167, new_n9162, new_n9168);
not_8  g08792(new_n9168, new_n9169);
xor_4  g08793(new_n9169, new_n9136, new_n9170);
not_8  g08794(new_n9170, new_n9171);
and_5  g08795(new_n8925, new_n8900, new_n9172);
and_5  g08796(new_n8926, new_n8898, new_n9173);
nor_5  g08797(new_n9173, new_n9172, new_n9174);
xor_4  g08798(new_n9174, new_n9171, new_n9175);
not_8  g08799(new_n9175, new_n9176);
nand_5 g08800(new_n9003, new_n8999, new_n9177);
and_5  g08801(new_n8993, new_n8990, new_n9178);
or_5   g08802(new_n8992, new_n8991, new_n9179);
not_8  g08803(new_n9179, new_n9180);
or_5   g08804(new_n8998, new_n8995, new_n9181);
not_8  g08805(new_n9181, new_n9182);
xor_4  g08806(new_n9182, new_n9180, new_n9183);
or_5   g08807(new_n9183, new_n9178, new_n9184);
or_5   g08808(new_n8982, new_n8981, new_n9185);
not_8  g08809(new_n9185, new_n9186);
nand_5 g08810(n7160, n2802, new_n9187);
not_8  g08811(new_n9187, new_n9188);
xor_4  g08812(new_n9188, new_n9186, new_n9189_1);
nand_5 g08813(n2515, n1512, new_n9190);
not_8  g08814(new_n9190, new_n9191);
nand_5 g08815(n1564, n1199, new_n9192);
nand_5 g08816(n4828, n533, new_n9193);
xor_4  g08817(new_n9193, new_n9192, new_n9194);
xor_4  g08818(new_n9194, new_n9191, new_n9195_1);
xor_4  g08819(new_n9195_1, new_n9189_1, new_n9196);
nor_5  g08820(new_n8984, new_n8980, new_n9197);
and_5  g08821(new_n8989, new_n8985, new_n9198);
or_5   g08822(new_n9198, new_n9197, new_n9199);
not_8  g08823(new_n9199, new_n9200);
nand_5 g08824(n12391, n5069, new_n9201);
not_8  g08825(new_n9201, new_n9202);
nand_5 g08826(n7891, n6806, new_n9203);
nand_5 g08827(n12069, n12044, new_n9204);
xor_4  g08828(new_n9204, new_n9203, new_n9205);
not_8  g08829(new_n9205, new_n9206);
xor_4  g08830(new_n9206, new_n9202, new_n9207);
xor_4  g08831(new_n9207, new_n9200, new_n9208);
xor_4  g08832(new_n9208, new_n9196, new_n9209);
xor_4  g08833(new_n9209, new_n9184, new_n9210);
not_8  g08834(new_n9210, new_n9211);
xor_4  g08835(new_n9211, new_n9177, new_n9212);
not_8  g08836(new_n9212, new_n9213);
nor_5  g08837(new_n9005, new_n8979, new_n9214);
and_5  g08838(new_n9005, new_n8979, new_n9215);
nor_5  g08839(new_n9215, new_n8978, new_n9216);
nor_5  g08840(new_n9216, new_n9214, new_n9217);
xor_4  g08841(new_n9217, new_n9213, new_n9218);
xor_4  g08842(new_n8926, new_n8897, new_n9219);
and_5  g08843(new_n9007, new_n9219, new_n9220);
nor_5  g08844(new_n9048, new_n9008, new_n9221);
nor_5  g08845(new_n9221, new_n9220, new_n9222);
xor_4  g08846(new_n9222, new_n9218, new_n9223);
not_8  g08847(new_n9223, new_n9224);
xor_4  g08848(new_n9224, new_n9176, new_n9225);
xor_4  g08849(new_n9225, new_n9135, new_n9226);
xor_4  g08850(new_n9226, new_n9093, new_n9227);
and_5  g08851(new_n9227, new_n8763, new_n9228);
xor_4  g08852(new_n8723, new_n8721, new_n9229);
xor_4  g08853(new_n8720, new_n8719, new_n9230);
xor_4  g08854(new_n9088, new_n9057, new_n9231);
nor_5  g08855(new_n9231, new_n9230, new_n9232);
xor_4  g08856(new_n8718, new_n8713, new_n9233);
xor_4  g08857(new_n9086, new_n9063, new_n9234);
nor_5  g08858(new_n9234, new_n9233, new_n9235);
not_8  g08859(new_n9233, new_n9236);
xor_4  g08860(new_n9234, new_n9236, new_n9237);
not_8  g08861(new_n9237, new_n9238);
xor_4  g08862(new_n9084, new_n9074, new_n9239);
not_8  g08863(new_n9239, new_n9240);
not_8  g08864(new_n8690, new_n9241_1);
and_5  g08865(new_n9241_1, new_n377, new_n9242);
nor_5  g08866(new_n9242, new_n8714, new_n9243);
or_5   g08867(new_n8688, new_n8687, new_n9244);
and_5  g08868(new_n9242, new_n9244, new_n9245);
or_5   g08869(new_n9245, new_n9243, new_n9246);
not_8  g08870(new_n9246, new_n9247);
nor_5  g08871(new_n9247, new_n9240, new_n9248);
xor_4  g08872(new_n9246, new_n9240, new_n9249);
nand_5 g08873(new_n384, new_n378, new_n9250);
xnor_4 g08874(new_n8716, new_n8715, new_n9251);
and_5  g08875(new_n9251, new_n9250, new_n9252);
xor_4  g08876(new_n9081, new_n9080_1, new_n9253);
xor_4  g08877(new_n9251, new_n9250, new_n9254);
not_8  g08878(new_n9254, new_n9255);
nor_5  g08879(new_n9255, new_n9253, new_n9256);
or_5   g08880(new_n9256, new_n9252, new_n9257);
not_8  g08881(new_n9257, new_n9258);
nor_5  g08882(new_n9258, new_n9249, new_n9259);
or_5   g08883(new_n9259, new_n9248, new_n9260);
and_5  g08884(new_n9260, new_n9238, new_n9261);
or_5   g08885(new_n9261, new_n9235, new_n9262);
not_8  g08886(new_n9230, new_n9263);
xor_4  g08887(new_n9231, new_n9263, new_n9264);
not_8  g08888(new_n9264, new_n9265);
and_5  g08889(new_n9265, new_n9262, new_n9266);
nor_5  g08890(new_n9266, new_n9232, new_n9267);
nor_5  g08891(new_n9267, new_n9229, new_n9268);
xor_4  g08892(new_n9090, new_n9052, new_n9269);
not_8  g08893(new_n9269, new_n9270);
not_8  g08894(new_n9229, new_n9271);
xor_4  g08895(new_n9267, new_n9271, new_n9272);
not_8  g08896(new_n9272, new_n9273);
and_5  g08897(new_n9273, new_n9270, new_n9274);
or_5   g08898(new_n9274, new_n9268, new_n9275);
xor_4  g08899(new_n9227, new_n8762, new_n9276);
not_8  g08900(new_n9276, new_n9277);
and_5  g08901(new_n9277, new_n9275, new_n9278);
nor_5  g08902(new_n9278, new_n9228, new_n9279);
or_5   g08903(new_n9222, new_n9218, new_n9280);
or_5   g08904(new_n9224, new_n9175, new_n9281);
nand_5 g08905(new_n9281, new_n9280, new_n9282);
nor_5  g08906(new_n9225, new_n9135, new_n9283);
and_5  g08907(new_n9226, new_n9093, new_n9284);
nor_5  g08908(new_n9284, new_n9283, new_n9285);
xor_4  g08909(new_n9285, new_n9282, new_n9286);
nor_5  g08910(new_n9129, new_n9094, new_n9287);
and_5  g08911(new_n9134, new_n9130, new_n9288);
nor_5  g08912(new_n9288, new_n9287, new_n9289);
and_5  g08913(new_n9182, new_n9180, new_n9290);
and_5  g08914(new_n9209, new_n9184, new_n9291);
or_5   g08915(new_n9291, new_n9290, new_n9292);
and_5  g08916(new_n9152, new_n9150, new_n9293);
and_5  g08917(new_n9159, new_n9153, new_n9294);
nor_5  g08918(new_n9294, new_n9293, new_n9295);
nor_5  g08919(new_n9193, new_n9192, new_n9296);
and_5  g08920(new_n9193, new_n9192, new_n9297);
nor_5  g08921(new_n9297, new_n9190, new_n9298);
nor_5  g08922(new_n9298, new_n9296, new_n9299);
xor_4  g08923(new_n9299, new_n9295, new_n9300);
and_5  g08924(n8028, n4817, new_n9301);
and_5  g08925(n7523, n7354, new_n9302);
xor_4  g08926(new_n9302, new_n9301, new_n9303);
and_5  g08927(n10848, n9457, new_n9304);
and_5  g08928(n11222, n1906, new_n9305);
xor_4  g08929(new_n9305, new_n9304, new_n9306);
and_5  g08930(n6986, n4928, new_n9307);
and_5  g08931(n4141, n2226, new_n9308);
xor_4  g08932(new_n9308, new_n9307, new_n9309);
xor_4  g08933(new_n9309, new_n9306, new_n9310);
xor_4  g08934(new_n9310, new_n9303, new_n9311);
nor_5  g08935(new_n8747, new_n8746, new_n9312);
and_5  g08936(new_n8747, new_n8746, new_n9313);
nor_5  g08937(new_n9313, new_n8745, new_n9314);
or_5   g08938(new_n9314, new_n9312, new_n9315);
nand_5 g08939(n4516, n2509, new_n9316);
and_5  g08940(n12704, n996, new_n9317);
and_5  g08941(n12720, n3627, new_n9318);
xor_4  g08942(new_n9318, new_n9317, new_n9319);
xor_4  g08943(new_n9319, new_n9316, new_n9320);
xor_4  g08944(new_n9320, new_n9315, new_n9321);
xor_4  g08945(new_n9321, new_n9311, new_n9322);
and_5  g08946(n2515, n533, new_n9323);
nand_5 g08947(n1512, n1199, new_n9324);
and_5  g08948(n12391, n12044, new_n9325);
xor_4  g08949(new_n9325, new_n9324, new_n9326);
xor_4  g08950(new_n9326, new_n9323, new_n9327);
xor_4  g08951(new_n9327, new_n9322, new_n9328);
xor_4  g08952(new_n9328, new_n9300, new_n9329);
or_5   g08953(new_n9147, new_n9139, new_n9330);
not_8  g08954(new_n9160, new_n9331);
nand_5 g08955(new_n9331, new_n9148, new_n9332);
and_5  g08956(new_n9332, new_n9330, new_n9333);
and_5  g08957(new_n9156, new_n9155, new_n9334);
not_8  g08958(new_n9154, new_n9335);
nor_5  g08959(new_n9158, new_n9335, new_n9336);
or_5   g08960(new_n9336, new_n9334, new_n9337);
and_5  g08961(n12069, n5694, new_n9338);
and_5  g08962(n11153, n4903, new_n9339);
xor_4  g08963(new_n9339, new_n9338, new_n9340);
nand_5 g08964(n7294, n5767, new_n9341);
and_5  g08965(n8336, n783, new_n9342);
xor_4  g08966(new_n9342, new_n9341, new_n9343);
xor_4  g08967(new_n9343, new_n9340, new_n9344);
xor_4  g08968(new_n9344, new_n9337, new_n9345);
nand_5 g08969(n4189, n4005, new_n9346);
and_5  g08970(n5814, n5314, new_n9347);
xor_4  g08971(new_n9347, new_n9346, new_n9348);
xor_4  g08972(new_n9348, new_n9345, new_n9349);
xor_4  g08973(new_n9349, new_n9333, new_n9350);
xor_4  g08974(new_n9350, new_n9329, new_n9351);
xor_4  g08975(new_n9351, new_n9292, new_n9352);
xor_4  g08976(new_n9352, new_n9289, new_n9353);
nor_5  g08977(new_n9211, new_n9177, new_n9354);
nor_5  g08978(new_n9217, new_n9213, new_n9355);
nor_5  g08979(new_n9355, new_n9354, new_n9356);
nor_5  g08980(new_n9169, new_n9136, new_n9357);
nor_5  g08981(new_n9174, new_n9171, new_n9358);
nor_5  g08982(new_n9358, new_n9357, new_n9359);
nor_5  g08983(new_n8739, new_n8731, new_n9360);
and_5  g08984(new_n8751, new_n8740, new_n9361);
or_5   g08985(new_n9361, new_n9360, new_n9362);
and_5  g08986(new_n8735, new_n8734, new_n9363);
nor_5  g08987(new_n8737, new_n8733, new_n9364);
nor_5  g08988(new_n9364, new_n9363, new_n9365);
xor_4  g08989(new_n9365, new_n9362, new_n9366);
and_5  g08990(new_n9143, new_n9142, new_n9367);
nor_5  g08991(new_n9145, new_n9141, new_n9368);
or_5   g08992(new_n9368, new_n9367, new_n9369);
and_5  g08993(new_n9204, new_n9203, new_n9370);
nor_5  g08994(new_n9206, new_n9202, new_n9371);
nor_5  g08995(new_n9371, new_n9370, new_n9372);
xor_4  g08996(new_n9372, new_n9369, new_n9373);
xor_4  g08997(new_n9373, new_n9366, new_n9374);
xor_4  g08998(new_n9374, new_n9359, new_n9375);
nor_5  g08999(new_n8759_1, new_n8727, new_n9376);
nor_5  g09000(new_n8761, new_n8726, new_n9377);
or_5   g09001(new_n9377, new_n9376, new_n9378);
and_5  g09002(new_n9207, new_n9200, new_n9379);
not_8  g09003(new_n9196, new_n9380);
and_5  g09004(new_n9208, new_n9380, new_n9381);
nor_5  g09005(new_n9381, new_n9379, new_n9382);
and_5  g09006(n6578, n1564, new_n9383);
xor_4  g09007(new_n9383, new_n9382, new_n9384);
xor_4  g09008(new_n9384, new_n9378, new_n9385);
xor_4  g09009(new_n9385, new_n9375, new_n9386);
nor_5  g09010(new_n9165, new_n9164, new_n9387_1);
nor_5  g09011(new_n9167, new_n9162, new_n9388);
nor_5  g09012(new_n9388, new_n9387_1, new_n9389);
and_5  g09013(new_n9110, new_n9108, new_n9390);
and_5  g09014(new_n9117, new_n9111_1, new_n9391);
nor_5  g09015(new_n9391, new_n9390, new_n9392);
and_5  g09016(new_n9102, new_n9101, new_n9393);
nor_5  g09017(new_n9104, new_n9100, new_n9394);
or_5   g09018(new_n9394, new_n9393, new_n9395);
and_5  g09019(n5319, n1980, new_n9396);
nand_5 g09020(n9920, n2508, new_n9397);
and_5  g09021(n10678, n1209, new_n9398);
xor_4  g09022(new_n9398, new_n9397, new_n9399);
xor_4  g09023(new_n9399, new_n9396, new_n9400_1);
xor_4  g09024(new_n9400_1, new_n9395, new_n9401);
xor_4  g09025(new_n9401, new_n9392, new_n9402);
xor_4  g09026(new_n9402, new_n9389, new_n9403);
nand_5 g09027(new_n9105, new_n9098, new_n9404);
not_8  g09028(new_n9118, new_n9405);
nand_5 g09029(new_n9405, new_n9106, new_n9406);
nand_5 g09030(new_n9406, new_n9404, new_n9407);
and_5  g09031(new_n9114, new_n9113, new_n9408);
not_8  g09032(new_n9112, new_n9409);
nor_5  g09033(new_n9116, new_n9409, new_n9410);
or_5   g09034(new_n9410, new_n9408, new_n9411);
nand_5 g09035(n4828, n2802, new_n9412);
nand_5 g09036(n10928, n8236, new_n9413);
and_5  g09037(n5105, n1094, new_n9414);
xor_4  g09038(new_n9414, new_n9413, new_n9415);
xor_4  g09039(new_n9415, new_n9412, new_n9416);
xor_4  g09040(new_n9416, new_n9411, new_n9417);
xor_4  g09041(new_n9417, new_n9407, new_n9418);
xor_4  g09042(new_n9418, new_n9403, new_n9419);
and_5  g09043(new_n9188, new_n9186, new_n9420);
and_5  g09044(new_n9195_1, new_n9189_1, new_n9421);
or_5   g09045(new_n9421, new_n9420, new_n9422);
nand_5 g09046(n7891, n5069, new_n9423);
and_5  g09047(n6038, n2087, new_n9424);
xor_4  g09048(new_n9424, new_n9423, new_n9425);
xor_4  g09049(new_n9425, new_n9422, new_n9426);
and_5  g09050(n7160, n6806, new_n9427);
and_5  g09051(n6687, n615, new_n9428);
xor_4  g09052(new_n9428, new_n9427, new_n9429);
xor_4  g09053(new_n9429, new_n9426, new_n9430);
xor_4  g09054(new_n9430, new_n9419, new_n9431);
nor_5  g09055(new_n8755, new_n8754, new_n9432);
nor_5  g09056(new_n8757, new_n8752, new_n9433);
nor_5  g09057(new_n9433, new_n9432, new_n9434);
and_5  g09058(new_n9125, new_n9123, new_n9435);
nor_5  g09059(new_n9127, new_n9120, new_n9436);
nor_5  g09060(new_n9436, new_n9435, new_n9437);
nor_5  g09061(new_n8743, new_n8742, new_n9438);
and_5  g09062(new_n8749, new_n8744, new_n9439);
or_5   g09063(new_n9439, new_n9438, new_n9440);
and_5  g09064(n7500, n7320, new_n9441);
nand_5 g09065(n12706, n2564, new_n9442);
and_5  g09066(n6770, n2585, new_n9443);
xor_4  g09067(new_n9443, new_n9442, new_n9444);
xor_4  g09068(new_n9444, new_n9441, new_n9445);
xor_4  g09069(new_n9445, new_n9440, new_n9446);
xor_4  g09070(new_n9446, new_n9437, new_n9447);
xor_4  g09071(new_n9447, new_n9434, new_n9448);
xor_4  g09072(new_n9448, new_n9431, new_n9449);
xor_4  g09073(new_n9449, new_n9386, new_n9450);
xor_4  g09074(new_n9450, new_n9356, new_n9451);
xor_4  g09075(new_n9451, new_n9353, new_n9452);
xor_4  g09076(new_n9452, new_n9286, new_n9453);
xor_4  g09077(new_n9453, new_n9279, n3654);
xor_4  g09078(new_n9273, new_n9269, n3661);
nand_5 g09079(n7456, n5305, new_n9456);
nand_5 g09080(n5964, n3932, new_n9457_1);
nand_5 g09081(n1798, n1097, new_n9458);
nand_5 g09082(n12591, n5305, new_n9459);
nand_5 g09083(new_n9459, new_n9458, new_n9460);
not_8  g09084(new_n9460, new_n9461);
nor_5  g09085(new_n9461, new_n9457_1, new_n9462);
nor_5  g09086(new_n9459, new_n9458, new_n9463);
nor_5  g09087(new_n9463, new_n9462, new_n9464);
xor_4  g09088(new_n9464, new_n9456, new_n9465);
not_8  g09089(new_n9465, new_n9466);
nand_5 g09090(n3932, n1097, new_n9467);
not_8  g09091(new_n9467, new_n9468);
nand_5 g09092(n4312, n1798, new_n9469);
nand_5 g09093(n12591, n5964, new_n9470);
xor_4  g09094(new_n9470, new_n9469, new_n9471);
not_8  g09095(new_n9471, new_n9472);
xor_4  g09096(new_n9472, new_n9468, new_n9473);
xor_4  g09097(new_n9473, new_n9466, new_n9474);
or_5   g09098(new_n6004, new_n6003, new_n9475);
xor_4  g09099(new_n9459, new_n9458, new_n9476);
or_5   g09100(new_n9476, new_n9475, new_n9477);
not_8  g09101(new_n9477, new_n9478);
nand_5 g09102(new_n9478, new_n9474, new_n9479);
not_8  g09103(new_n9479, new_n9480);
nand_5 g09104(n11662, n5305, new_n9481);
not_8  g09105(new_n9481, new_n9482);
nand_5 g09106(n7456, n5964, new_n9483);
nand_5 g09107(n4312, n3932, new_n9484);
not_8  g09108(new_n9484, new_n9485);
nand_5 g09109(n12591, n1097, new_n9486);
nand_5 g09110(n12705, n1798, new_n9487);
xor_4  g09111(new_n9487, new_n9486, new_n9488);
not_8  g09112(new_n9488, new_n9489);
xor_4  g09113(new_n9489, new_n9485, new_n9490);
xor_4  g09114(new_n9490, new_n9483, new_n9491);
and_5  g09115(new_n9470, new_n9469, new_n9492);
nor_5  g09116(new_n9472, new_n9468, new_n9493);
or_5   g09117(new_n9493, new_n9492, new_n9494);
not_8  g09118(new_n9494, new_n9495);
xor_4  g09119(new_n9495, new_n9491, new_n9496);
xor_4  g09120(new_n9496, new_n9482, new_n9497);
not_8  g09121(new_n9497, new_n9498);
nor_5  g09122(new_n9464, new_n9456, new_n9499);
nor_5  g09123(new_n9473, new_n9466, new_n9500);
nor_5  g09124(new_n9500, new_n9499, new_n9501);
xor_4  g09125(new_n9501, new_n9498, new_n9502);
xor_4  g09126(new_n9502, new_n9480, new_n9503);
not_8  g09127(new_n9503, new_n9504);
xor_4  g09128(new_n9478, new_n9474, new_n9505);
not_8  g09129(new_n9505, new_n9506);
nand_5 g09130(n11023, n8759, new_n9507);
not_8  g09131(new_n9507, new_n9508);
and_5  g09132(n8759, n3022, new_n9509);
and_5  g09133(n12299, n6703, new_n9510);
nor_5  g09134(new_n9510, new_n9509, new_n9511);
nand_5 g09135(n12299, n3022, new_n9512);
nor_5  g09136(new_n9512, new_n5996, new_n9513);
nand_5 g09137(n9640, n6776, new_n9514);
not_8  g09138(new_n9514, new_n9515);
nor_5  g09139(new_n9515, new_n9513, new_n9516);
or_5   g09140(new_n9516, new_n9511, new_n9517);
not_8  g09141(new_n9517, new_n9518);
and_5  g09142(new_n9518, new_n9508, new_n9519);
nor_5  g09143(new_n9518, new_n9508, new_n9520);
or_5   g09144(new_n9520, new_n9519, new_n9521);
nand_5 g09145(n12299, n9640, new_n9522);
not_8  g09146(new_n9522, new_n9523);
nand_5 g09147(n6776, n3022, new_n9524);
nand_5 g09148(n7436, n6703, new_n9525);
xor_4  g09149(new_n9525, new_n9524, new_n9526);
xor_4  g09150(new_n9526, new_n9523, new_n9527);
not_8  g09151(new_n9527, new_n9528);
xor_4  g09152(new_n9528, new_n9521, new_n9529);
not_8  g09153(new_n5996, new_n9530);
or_5   g09154(new_n9514, new_n9530, new_n9531);
not_8  g09155(new_n9531, new_n9532);
nor_5  g09156(new_n9513, new_n9511, new_n9533);
or_5   g09157(new_n9533, new_n9532, new_n9534);
not_8  g09158(new_n9534, new_n9535);
nand_5 g09159(new_n9535, new_n9515, new_n9536);
not_8  g09160(new_n9536, new_n9537);
xor_4  g09161(new_n9537, new_n9529, new_n9538);
not_8  g09162(new_n9538, new_n9539);
nand_5 g09163(n11922, n5331, new_n9540);
nand_5 g09164(n2530, n1067, new_n9541);
not_8  g09165(new_n9541, new_n9542);
nand_5 g09166(n8665, n8476, new_n9543);
nand_5 g09167(n12648, n5645, new_n9544);
xor_4  g09168(new_n9544, new_n9543, new_n9545);
xor_4  g09169(new_n9545, new_n9542, new_n9546);
not_8  g09170(new_n9546, new_n9547);
xor_4  g09171(new_n9547, new_n9540, new_n9548);
and_5  g09172(n8665, n5331, new_n9549);
and_5  g09173(n5645, n2530, new_n9550);
or_5   g09174(new_n9550, new_n9549, new_n9551);
not_8  g09175(new_n9551, new_n9552);
nand_5 g09176(n8476, n1067, new_n9553);
not_8  g09177(new_n9553, new_n9554);
nand_5 g09178(n8665, n2530, new_n9555);
nor_5  g09179(new_n9555, new_n5997, new_n9556);
nor_5  g09180(new_n9556, new_n9554, new_n9557);
or_5   g09181(new_n9557, new_n9552, new_n9558);
not_8  g09182(new_n9558, new_n9559);
xor_4  g09183(new_n9559, new_n9548, new_n9560);
nor_5  g09184(new_n6022, new_n6021, new_n9561);
or_5   g09185(new_n9556, new_n9552, new_n9562);
and_5  g09186(new_n9562, new_n9561, new_n9563);
xor_4  g09187(new_n9563, new_n9560, new_n9564);
nand_5 g09188(n7965, n2749, new_n9565);
not_8  g09189(new_n9565, new_n9566);
and_5  g09190(n7965, n3754, new_n9567);
and_5  g09191(n11892, n11876, new_n9568);
nor_5  g09192(new_n9568, new_n9567, new_n9569);
nand_5 g09193(n11892, n3754, new_n9570);
nor_5  g09194(new_n9570, new_n5998, new_n9571_1);
and_5  g09195(n10898, n7388, new_n9572);
nor_5  g09196(new_n9572, new_n9571_1, new_n9573);
or_5   g09197(new_n9573, new_n9569, new_n9574);
not_8  g09198(new_n9574, new_n9575);
and_5  g09199(new_n9575, new_n9566, new_n9576);
nor_5  g09200(new_n9575, new_n9566, new_n9577);
or_5   g09201(new_n9577, new_n9576, new_n9578_1);
nand_5 g09202(n11892, n10898, new_n9579);
nand_5 g09203(n7388, n3754, new_n9580);
nand_5 g09204(n11876, n2393, new_n9581);
xnor_4 g09205(new_n9581, new_n9580, new_n9582);
not_8  g09206(new_n9582, new_n9583_1);
xor_4  g09207(new_n9583_1, new_n9579, new_n9584);
xor_4  g09208(new_n9584, new_n9578_1, new_n9585);
not_8  g09209(new_n9572, new_n9586);
nand_5 g09210(new_n9572, new_n5998, new_n9587);
not_8  g09211(new_n9587, new_n9588);
nor_5  g09212(new_n9571_1, new_n9569, new_n9589);
nor_5  g09213(new_n9589, new_n9588, new_n9590);
not_8  g09214(new_n9590, new_n9591);
or_5   g09215(new_n9591, new_n9586, new_n9592);
xnor_4 g09216(new_n9592, new_n9585, new_n9593);
xor_4  g09217(new_n9593, new_n9564, new_n9594);
not_8  g09218(new_n9594, new_n9595);
or_5   g09219(new_n9587, new_n9569, new_n9596);
and_5  g09220(new_n9596, new_n9591, new_n9597);
nor_5  g09221(new_n6019, new_n6014, new_n9598);
nor_5  g09222(new_n6024, new_n6020, new_n9599);
or_5   g09223(new_n9599, new_n9598, new_n9600);
nor_5  g09224(new_n9600, new_n9597, new_n9601);
not_8  g09225(new_n9600, new_n9602);
xor_4  g09226(new_n9602, new_n9597, new_n9603);
not_8  g09227(new_n5997, new_n9604);
or_5   g09228(new_n9553, new_n9604, new_n9605);
nor_5  g09229(new_n9605, new_n9551, new_n9606);
not_8  g09230(new_n9605, new_n9607);
nor_5  g09231(new_n9607, new_n9562, new_n9608);
or_5   g09232(new_n9608, new_n9606, new_n9609);
nor_5  g09233(new_n9609, new_n9603, new_n9610);
nor_5  g09234(new_n9610, new_n9601, new_n9611);
xor_4  g09235(new_n9611, new_n9595, new_n9612);
not_8  g09236(new_n9612, new_n9613);
xor_4  g09237(new_n9613, new_n9539, new_n9614);
nor_5  g09238(new_n9531, new_n9511, new_n9615);
or_5   g09239(new_n9615, new_n9535, new_n9616);
nor_5  g09240(new_n6012, new_n6009, new_n9617);
and_5  g09241(new_n6025, new_n6013, new_n9618);
or_5   g09242(new_n9618, new_n9617, new_n9619);
not_8  g09243(new_n9619, new_n9620);
and_5  g09244(new_n9620, new_n9616, new_n9621);
xor_4  g09245(new_n9609, new_n9603, new_n9622);
xor_4  g09246(new_n9620, new_n9616, new_n9623);
and_5  g09247(new_n9623, new_n9622, new_n9624);
nor_5  g09248(new_n9624, new_n9621, new_n9625);
xor_4  g09249(new_n9625, new_n9614, new_n9626);
nor_5  g09250(new_n9626, new_n9506, new_n9627);
xor_4  g09251(new_n9626, new_n9506, new_n9628);
not_8  g09252(new_n9628, new_n9629);
not_8  g09253(new_n9622, new_n9630);
xnor_4 g09254(new_n9623, new_n9630, new_n9631);
not_8  g09255(new_n9457_1, new_n9632);
and_5  g09256(new_n9632, new_n5994, new_n9633);
and_5  g09257(new_n9633, new_n9461, new_n9634);
not_8  g09258(new_n9476, new_n9635);
nor_5  g09259(new_n9633, new_n9635, new_n9636);
or_5   g09260(new_n9636, new_n9634, new_n9637_1);
not_8  g09261(new_n9637_1, new_n9638);
and_5  g09262(new_n9638, new_n9631, new_n9639);
nor_5  g09263(new_n6006, new_n6002, new_n9640_1);
nor_5  g09264(new_n6027, new_n6008, new_n9641);
or_5   g09265(new_n9641, new_n9640_1, new_n9642);
xor_4  g09266(new_n9638, new_n9631, new_n9643);
not_8  g09267(new_n9643, new_n9644);
nor_5  g09268(new_n9644, new_n9642, new_n9645);
or_5   g09269(new_n9645, new_n9639, new_n9646);
nor_5  g09270(new_n9646, new_n9629, new_n9647);
nor_5  g09271(new_n9647, new_n9627, new_n9648);
xor_4  g09272(new_n9648, new_n9504, new_n9649);
not_8  g09273(new_n9649, new_n9650);
nand_5 g09274(new_n9537, new_n9529, new_n9651);
nand_5 g09275(n10451, n8759, new_n9652);
not_8  g09276(new_n9652, new_n9653);
nand_5 g09277(n11023, n6776, new_n9654);
not_8  g09278(new_n9654, new_n9655);
and_5  g09279(new_n9525, new_n9524, new_n9656);
nor_5  g09280(new_n9525, new_n9524, new_n9657);
nor_5  g09281(new_n9657, new_n9523, new_n9658);
nor_5  g09282(new_n9658, new_n9656, new_n9659);
not_8  g09283(new_n9659, new_n9660);
xor_4  g09284(new_n9660, new_n9655, new_n9661);
nand_5 g09285(n9640, n7436, new_n9662);
not_8  g09286(new_n9662, new_n9663);
nand_5 g09287(n8276, n6703, new_n9664);
xor_4  g09288(new_n9664, new_n9512, new_n9665);
xor_4  g09289(new_n9665, new_n9663, new_n9666);
not_8  g09290(new_n9666, new_n9667);
xor_4  g09291(new_n9667, new_n9661, new_n9668);
xor_4  g09292(new_n9668, new_n9653, new_n9669);
not_8  g09293(new_n9669, new_n9670);
nor_5  g09294(new_n9528, new_n9521, new_n9671);
nor_5  g09295(new_n9671, new_n9519, new_n9672);
xor_4  g09296(new_n9672, new_n9670, new_n9673);
not_8  g09297(new_n9673, new_n9674);
xor_4  g09298(new_n9674, new_n9651, new_n9675);
not_8  g09299(new_n9675, new_n9676);
not_8  g09300(new_n9592, new_n9677);
nand_5 g09301(new_n9677, new_n9585, new_n9678);
not_8  g09302(new_n9678, new_n9679);
nand_5 g09303(n7965, n159, new_n9680);
not_8  g09304(new_n9680, new_n9681);
nor_5  g09305(new_n9584, new_n9578_1, new_n9682);
nor_5  g09306(new_n9682, new_n9576, new_n9683);
xor_4  g09307(new_n9683, new_n9681, new_n9684);
not_8  g09308(new_n9684, new_n9685);
nand_5 g09309(n7388, n2749, new_n9686);
not_8  g09310(new_n9686, new_n9687);
and_5  g09311(new_n9581, new_n9580, new_n9688);
and_5  g09312(new_n9583_1, new_n9579, new_n9689);
or_5   g09313(new_n9689, new_n9688, new_n9690);
not_8  g09314(new_n9690, new_n9691);
xor_4  g09315(new_n9691, new_n9687, new_n9692);
nand_5 g09316(n11876, n5860, new_n9693);
nand_5 g09317(n10898, n2393, new_n9694);
xor_4  g09318(new_n9694, new_n9693, new_n9695);
not_8  g09319(new_n9695, new_n9696);
xor_4  g09320(new_n9696, new_n9570, new_n9697);
xor_4  g09321(new_n9697, new_n9692, new_n9698);
xor_4  g09322(new_n9698, new_n9685, new_n9699);
xor_4  g09323(new_n9699, new_n9679, new_n9700);
nand_5 g09324(new_n9563, new_n9560, new_n9701);
nand_5 g09325(n5331, n2551, new_n9702);
not_8  g09326(new_n9702, new_n9703);
nand_5 g09327(n11922, n8476, new_n9704);
and_5  g09328(new_n9544, new_n9543, new_n9705);
nor_5  g09329(new_n9544, new_n9543, new_n9706_1);
nor_5  g09330(new_n9706_1, new_n9542, new_n9707);
nor_5  g09331(new_n9707, new_n9705, new_n9708);
not_8  g09332(new_n9708, new_n9709);
xor_4  g09333(new_n9709, new_n9704, new_n9710);
nand_5 g09334(n12648, n1067, new_n9711);
not_8  g09335(new_n9711, new_n9712);
nand_5 g09336(n10545, n5645, new_n9713);
xor_4  g09337(new_n9713, new_n9555, new_n9714);
xor_4  g09338(new_n9714, new_n9712, new_n9715);
xor_4  g09339(new_n9715, new_n9710, new_n9716);
xor_4  g09340(new_n9716, new_n9703, new_n9717);
nor_5  g09341(new_n9547, new_n9540, new_n9718);
and_5  g09342(new_n9559, new_n9548, new_n9719);
or_5   g09343(new_n9719, new_n9718, new_n9720);
xor_4  g09344(new_n9720, new_n9717, new_n9721);
not_8  g09345(new_n9721, new_n9722);
xor_4  g09346(new_n9722, new_n9701, new_n9723);
not_8  g09347(new_n9723, new_n9724);
xor_4  g09348(new_n9724, new_n9700, new_n9725_1);
nor_5  g09349(new_n9593, new_n9564, new_n9726);
nor_5  g09350(new_n9611, new_n9595, new_n9727);
nor_5  g09351(new_n9727, new_n9726, new_n9728);
xor_4  g09352(new_n9728, new_n9725_1, new_n9729);
xor_4  g09353(new_n9729, new_n9676, new_n9730);
not_8  g09354(new_n9730, new_n9731);
nor_5  g09355(new_n9613, new_n9538, new_n9732);
nor_5  g09356(new_n9625, new_n9614, new_n9733);
or_5   g09357(new_n9733, new_n9732, new_n9734);
not_8  g09358(new_n9734, new_n9735);
xnor_4 g09359(new_n9735, new_n9731, new_n9736);
xnor_4 g09360(new_n9736, new_n9650, n3677);
not_8  g09361(new_n8448, new_n9738);
xor_4  g09362(new_n8450, new_n9738, n3849);
xor_4  g09363(new_n5989, new_n5987, n4088);
xor_4  g09364(new_n1136_1, new_n1052, n4155);
xor_4  g09365(new_n2875, new_n2873, n4159);
xor_4  g09366(new_n5977, new_n5823, n4226);
nand_5 g09367(n12591, n4312, new_n9744);
not_8  g09368(new_n9744, new_n9745);
and_5  g09369(new_n9487, new_n9486, new_n9746);
nor_5  g09370(new_n9489, new_n9485, new_n9747);
nor_5  g09371(new_n9747, new_n9746, new_n9748);
xor_4  g09372(new_n9748, new_n9745, new_n9749);
not_8  g09373(new_n9749, new_n9750);
nand_5 g09374(n12705, n3932, new_n9751);
nand_5 g09375(n12025, n1798, new_n9752);
xor_4  g09376(new_n9752, new_n9751, new_n9753);
xor_4  g09377(new_n9753, new_n9750, new_n9754);
nand_5 g09378(n11662, n5964, new_n9755);
nand_5 g09379(n7456, n1097, new_n9756_1);
xor_4  g09380(new_n9756_1, new_n9755, new_n9757);
not_8  g09381(new_n9757, new_n9758);
xor_4  g09382(new_n9758, new_n9754, new_n9759);
nor_5  g09383(new_n9490, new_n9483, new_n9760);
and_5  g09384(new_n9495, new_n9491, new_n9761);
or_5   g09385(new_n9761, new_n9760, new_n9762);
not_8  g09386(new_n9762, new_n9763_1);
xor_4  g09387(new_n9763_1, new_n9759, new_n9764);
and_5  g09388(new_n9496, new_n9482, new_n9765);
nor_5  g09389(new_n9501, new_n9498, new_n9766);
nor_5  g09390(new_n9766, new_n9765, new_n9767_1);
or_5   g09391(new_n9767_1, new_n9764, new_n9768);
not_8  g09392(new_n9768, new_n9769);
nor_5  g09393(new_n9748, new_n9745, new_n9770);
nor_5  g09394(new_n9753, new_n9750, new_n9771);
or_5   g09395(new_n9771, new_n9770, new_n9772);
nand_5 g09396(n10327, n5964, new_n9773);
not_8  g09397(new_n9773, new_n9774);
nand_5 g09398(n11662, n1097, new_n9775);
nand_5 g09399(n9583, n5305, new_n9776);
xor_4  g09400(new_n9776, new_n9775, new_n9777);
not_8  g09401(new_n9777, new_n9778);
xor_4  g09402(new_n9778, new_n9774, new_n9779);
xor_4  g09403(new_n9779, new_n9772, new_n9780);
not_8  g09404(new_n9780, new_n9781);
or_5   g09405(new_n9752, new_n9751, new_n9782);
not_8  g09406(new_n9782, new_n9783);
and_5  g09407(n7456, n4312, new_n9784);
xor_4  g09408(new_n9784, new_n9783, new_n9785);
nand_5 g09409(n12025, n3932, new_n9786);
not_8  g09410(new_n9786, new_n9787);
nand_5 g09411(n12705, n12591, new_n9788);
nand_5 g09412(n11257, n1798, new_n9789);
xor_4  g09413(new_n9789, new_n9788, new_n9790);
not_8  g09414(new_n9790, new_n9791);
xor_4  g09415(new_n9791, new_n9787, new_n9792);
xor_4  g09416(new_n9792, new_n9785, new_n9793);
not_8  g09417(new_n9793, new_n9794);
xor_4  g09418(new_n9794, new_n9781, new_n9795);
nor_5  g09419(new_n9758, new_n9754, new_n9796);
or_5   g09420(new_n9756_1, new_n9755, new_n9797);
not_8  g09421(new_n9797, new_n9798);
nand_5 g09422(new_n9762, new_n9759, new_n9799);
not_8  g09423(new_n9799, new_n9800);
xor_4  g09424(new_n9800, new_n9798, new_n9801);
nor_5  g09425(new_n9801, new_n9796, new_n9802);
xor_4  g09426(new_n9802, new_n9795, new_n9803);
not_8  g09427(new_n9803, new_n9804);
xor_4  g09428(new_n9804, new_n9769, new_n9805);
nand_5 g09429(n10327, n5305, new_n9806);
not_8  g09430(new_n9806, new_n9807);
xor_4  g09431(new_n9767_1, new_n9764, new_n9808);
or_5   g09432(new_n9808, new_n9807, new_n9809);
and_5  g09433(new_n9502, new_n9480, new_n9810);
xor_4  g09434(new_n9808, new_n9807, new_n9811);
not_8  g09435(new_n9811, new_n9812);
or_5   g09436(new_n9812, new_n9810, new_n9813);
nand_5 g09437(new_n9813, new_n9809, new_n9814);
xor_4  g09438(new_n9814, new_n9805, new_n9815);
nor_5  g09439(new_n9660, new_n9654, new_n9816);
nor_5  g09440(new_n9667, new_n9661, new_n9817);
or_5   g09441(new_n9817, new_n9816, new_n9818);
nand_5 g09442(n10451, n6776, new_n9819);
nand_5 g09443(n12299, n11023, new_n9820_1);
xor_4  g09444(new_n9820_1, new_n9819, new_n9821);
xor_4  g09445(new_n9821, new_n9818, new_n9822);
not_8  g09446(new_n9822, new_n9823);
nand_5 g09447(n7436, n3022, new_n9824);
nand_5 g09448(n9640, n8276, new_n9825);
nand_5 g09449(n9241, n6703, new_n9826);
xor_4  g09450(new_n9826, new_n9825, new_n9827);
xor_4  g09451(new_n9827, new_n9824, new_n9828);
and_5  g09452(new_n9664, new_n9512, new_n9829);
nor_5  g09453(new_n9664, new_n9512, new_n9830);
nor_5  g09454(new_n9830, new_n9663, new_n9831);
nor_5  g09455(new_n9831, new_n9829, new_n9832);
xor_4  g09456(new_n9832, new_n9828, new_n9833);
xor_4  g09457(new_n9833, new_n9823, new_n9834);
not_8  g09458(new_n9834, new_n9835);
and_5  g09459(new_n9668, new_n9653, new_n9836);
nor_5  g09460(new_n9672, new_n9670, new_n9837);
nor_5  g09461(new_n9837, new_n9836, new_n9838);
or_5   g09462(new_n9838, new_n9835, new_n9839);
not_8  g09463(new_n9839, new_n9840);
not_8  g09464(new_n9824, new_n9841);
nor_5  g09465(new_n9827, new_n9841, new_n9842);
nor_5  g09466(new_n9832, new_n9828, new_n9843);
or_5   g09467(new_n9843, new_n9842, new_n9844);
not_8  g09468(new_n9844, new_n9845);
nand_5 g09469(n10278, n6776, new_n9846);
not_8  g09470(new_n9846, new_n9847);
nand_5 g09471(n12299, n10451, new_n9848);
nand_5 g09472(n11423, n8759, new_n9849);
xor_4  g09473(new_n9849, new_n9848, new_n9850);
not_8  g09474(new_n9850, new_n9851);
xor_4  g09475(new_n9851, new_n9847, new_n9852);
not_8  g09476(new_n9852, new_n9853);
nor_5  g09477(new_n9853, new_n9845, new_n9854);
and_5  g09478(new_n9853, new_n9845, new_n9855);
or_5   g09479(new_n9855, new_n9854, new_n9856);
or_5   g09480(new_n9826, new_n9825, new_n9857);
nand_5 g09481(n11023, n7436, new_n9858);
not_8  g09482(new_n9858, new_n9859);
xor_4  g09483(new_n9859, new_n9857, new_n9860);
nand_5 g09484(n9640, n9241, new_n9861);
not_8  g09485(new_n9861, new_n9862);
nand_5 g09486(n8276, n3022, new_n9863);
nand_5 g09487(n10510, n6703, new_n9864);
xor_4  g09488(new_n9864, new_n9863, new_n9865);
not_8  g09489(new_n9865, new_n9866);
xor_4  g09490(new_n9866, new_n9862, new_n9867);
xor_4  g09491(new_n9867, new_n9860, new_n9868);
xor_4  g09492(new_n9868, new_n9856, new_n9869);
and_5  g09493(new_n9821, new_n9818, new_n9870);
or_5   g09494(new_n9820_1, new_n9819, new_n9871);
or_5   g09495(new_n9833, new_n9823, new_n9872);
xor_4  g09496(new_n9872, new_n9871, new_n9873);
nor_5  g09497(new_n9873, new_n9870, new_n9874);
xor_4  g09498(new_n9874, new_n9869, new_n9875);
not_8  g09499(new_n9875, new_n9876);
xor_4  g09500(new_n9876, new_n9840, new_n9877);
nand_5 g09501(n10278, n8759, new_n9878);
xor_4  g09502(new_n9838, new_n9835, new_n9879);
not_8  g09503(new_n9879, new_n9880);
nor_5  g09504(new_n9880, new_n9878, new_n9881);
or_5   g09505(new_n9674, new_n9651, new_n9882);
not_8  g09506(new_n9882, new_n9883);
xor_4  g09507(new_n9880, new_n9878, new_n9884);
and_5  g09508(new_n9884, new_n9883, new_n9885);
nor_5  g09509(new_n9885, new_n9881, new_n9886);
xor_4  g09510(new_n9886, new_n9877, new_n9887);
nand_5 g09511(n12648, n8665, new_n9888);
nand_5 g09512(n10545, n1067, new_n9889);
nand_5 g09513(n7690, n5645, new_n9890);
xor_4  g09514(new_n9890, new_n9889, new_n9891);
not_8  g09515(new_n9891, new_n9892);
xor_4  g09516(new_n9892, new_n9888, new_n9893);
and_5  g09517(new_n9713, new_n9555, new_n9894);
nor_5  g09518(new_n9713, new_n9555, new_n9895);
nor_5  g09519(new_n9895, new_n9712, new_n9896);
or_5   g09520(new_n9896, new_n9894, new_n9897);
not_8  g09521(new_n9897, new_n9898);
xor_4  g09522(new_n9898, new_n9893, new_n9899);
nand_5 g09523(n8476, n2551, new_n9900);
nand_5 g09524(n11922, n2530, new_n9901);
xor_4  g09525(new_n9901, new_n9900, new_n9902);
xor_4  g09526(new_n9902, new_n9899, new_n9903);
nor_5  g09527(new_n9709, new_n9704, new_n9904);
and_5  g09528(new_n9715, new_n9710, new_n9905);
or_5   g09529(new_n9905, new_n9904, new_n9906);
xnor_4 g09530(new_n9906, new_n9903, new_n9907);
and_5  g09531(new_n9716, new_n9703, new_n9908);
and_5  g09532(new_n9720, new_n9717, new_n9909);
nor_5  g09533(new_n9909, new_n9908, new_n9910);
or_5   g09534(new_n9910, new_n9907, new_n9911);
not_8  g09535(new_n9911, new_n9912);
or_5   g09536(new_n9890, new_n9889, new_n9913);
not_8  g09537(new_n9913, new_n9914);
nand_5 g09538(n12648, n11922, new_n9915);
not_8  g09539(new_n9915, new_n9916);
xor_4  g09540(new_n9916, new_n9914, new_n9917);
nand_5 g09541(n7690, n1067, new_n9918);
nand_5 g09542(n10545, n8665, new_n9919);
nand_5 g09543(n5645, n3616, new_n9920_1);
xor_4  g09544(new_n9920_1, new_n9919, new_n9921);
not_8  g09545(new_n9921, new_n9922);
xor_4  g09546(new_n9922, new_n9918, new_n9923);
xor_4  g09547(new_n9923, new_n9917, new_n9924);
not_8  g09548(new_n9924, new_n9925);
nor_5  g09549(new_n9892, new_n9888, new_n9926);
and_5  g09550(new_n9898, new_n9893, new_n9927);
or_5   g09551(new_n9927, new_n9926, new_n9928);
nand_5 g09552(n12826, n8476, new_n9929);
not_8  g09553(new_n9929, new_n9930);
nand_5 g09554(n2551, n2530, new_n9931);
nand_5 g09555(n5331, n4094, new_n9932);
xor_4  g09556(new_n9932, new_n9931, new_n9933);
not_8  g09557(new_n9933, new_n9934);
xor_4  g09558(new_n9934, new_n9930, new_n9935);
not_8  g09559(new_n9935, new_n9936);
xor_4  g09560(new_n9936, new_n9928, new_n9937);
xor_4  g09561(new_n9937, new_n9925, new_n9938_1);
and_5  g09562(new_n9902, new_n9899, new_n9939);
or_5   g09563(new_n9901, new_n9900, new_n9940);
not_8  g09564(new_n9940, new_n9941);
nand_5 g09565(new_n9906, new_n9903, new_n9942);
not_8  g09566(new_n9942, new_n9943);
xor_4  g09567(new_n9943, new_n9941, new_n9944);
nor_5  g09568(new_n9944, new_n9939, new_n9945);
xor_4  g09569(new_n9945, new_n9938_1, new_n9946);
not_8  g09570(new_n9946, new_n9947);
xor_4  g09571(new_n9947, new_n9912, new_n9948);
nand_5 g09572(n12826, n5331, new_n9949);
not_8  g09573(new_n9949, new_n9950);
xor_4  g09574(new_n9910, new_n9907, new_n9951);
nor_5  g09575(new_n9951, new_n9950, new_n9952);
or_5   g09576(new_n9722, new_n9701, new_n9953);
not_8  g09577(new_n9953, new_n9954);
xor_4  g09578(new_n9951, new_n9950, new_n9955);
not_8  g09579(new_n9955, new_n9956_1);
nor_5  g09580(new_n9956_1, new_n9954, new_n9957);
or_5   g09581(new_n9957, new_n9952, new_n9958);
xor_4  g09582(new_n9958, new_n9948, new_n9959);
not_8  g09583(new_n9959, new_n9960);
nand_5 g09584(n7965, n1510, new_n9961);
and_5  g09585(new_n9691, new_n9687, new_n9962);
and_5  g09586(new_n9697, new_n9692, new_n9963);
or_5   g09587(new_n9963, new_n9962, new_n9964);
not_8  g09588(new_n9964, new_n9965);
nand_5 g09589(n7388, n159, new_n9966);
nand_5 g09590(n11892, n2749, new_n9967);
xnor_4 g09591(new_n9967, new_n9966, new_n9968);
xor_4  g09592(new_n9968, new_n9965, new_n9969);
nand_5 g09593(n3754, n2393, new_n9970);
nand_5 g09594(n10898, n5860, new_n9971);
nand_5 g09595(n11876, n3986, new_n9972);
xor_4  g09596(new_n9972, new_n9971, new_n9973);
not_8  g09597(new_n9973, new_n9974);
xor_4  g09598(new_n9974, new_n9970, new_n9975);
and_5  g09599(new_n9694, new_n9693, new_n9976);
not_8  g09600(new_n9570, new_n9977);
nor_5  g09601(new_n9696, new_n9977, new_n9978);
or_5   g09602(new_n9978, new_n9976, new_n9979);
not_8  g09603(new_n9979, new_n9980);
xnor_4 g09604(new_n9980, new_n9975, new_n9981);
xor_4  g09605(new_n9981, new_n9969, new_n9982);
nor_5  g09606(new_n9683, new_n9680, new_n9983);
and_5  g09607(new_n9698, new_n9685, new_n9984);
nor_5  g09608(new_n9984, new_n9983, new_n9985);
xor_4  g09609(new_n9985, new_n9982, new_n9986);
not_8  g09610(new_n9986, new_n9987);
nor_5  g09611(new_n9987, new_n9961, new_n9988);
nand_5 g09612(new_n9699, new_n9679, new_n9989);
not_8  g09613(new_n9989, new_n9990);
xor_4  g09614(new_n9987, new_n9961, new_n9991);
and_5  g09615(new_n9991, new_n9990, new_n9992);
or_5   g09616(new_n9992, new_n9988, new_n9993);
not_8  g09617(new_n9993, new_n9994);
or_5   g09618(new_n9985, new_n9982, new_n9995);
not_8  g09619(new_n9995, new_n9996);
or_5   g09620(new_n9967, new_n9966, new_n9997);
not_8  g09621(new_n9997, new_n9998);
and_5  g09622(new_n9968, new_n9965, new_n9999);
and_5  g09623(new_n9981, new_n9969, new_n10000);
or_5   g09624(new_n10000, new_n9999, new_n10001);
not_8  g09625(new_n10001, new_n10002);
xor_4  g09626(new_n10002, new_n9998, new_n10003);
nand_5 g09627(n7388, n1510, new_n10004);
nand_5 g09628(n11892, n159, new_n10005);
and_5  g09629(n12247, n7965, new_n10006);
xor_4  g09630(new_n10006, new_n10005, new_n10007);
not_8  g09631(new_n10007, new_n10008);
xor_4  g09632(new_n10008, new_n10004, new_n10009);
nor_5  g09633(new_n9974, new_n9970, new_n10010);
and_5  g09634(new_n9980, new_n9975, new_n10011);
or_5   g09635(new_n10011, new_n10010, new_n10012);
not_8  g09636(new_n10012, new_n10013);
xor_4  g09637(new_n10013, new_n10009, new_n10014);
or_5   g09638(new_n9972, new_n9971, new_n10015);
nand_5 g09639(n2749, n2393, new_n10016);
not_8  g09640(new_n10016, new_n10017);
xor_4  g09641(new_n10017, new_n10015, new_n10018);
nand_5 g09642(n10898, n3986, new_n10019);
not_8  g09643(new_n10019, new_n10020);
nand_5 g09644(n11876, n5857, new_n10021);
nand_5 g09645(n5860, n3754, new_n10022_1);
xor_4  g09646(new_n10022_1, new_n10021, new_n10023);
not_8  g09647(new_n10023, new_n10024);
xor_4  g09648(new_n10024, new_n10020, new_n10025);
xor_4  g09649(new_n10025, new_n10018, new_n10026);
xor_4  g09650(new_n10026, new_n10014, new_n10027);
xor_4  g09651(new_n10027, new_n10003, new_n10028);
not_8  g09652(new_n10028, new_n10029);
xor_4  g09653(new_n10029, new_n9996, new_n10030);
xnor_4 g09654(new_n10030, new_n9994, new_n10031);
xor_4  g09655(new_n10031, new_n9960, new_n10032);
not_8  g09656(new_n10032, new_n10033);
xor_4  g09657(new_n9991, new_n9990, new_n10034);
and_5  g09658(new_n9956_1, new_n9954, new_n10035);
or_5   g09659(new_n10035, new_n9957, new_n10036);
nor_5  g09660(new_n10036, new_n10034, new_n10037);
nor_5  g09661(new_n9723, new_n9700, new_n10038);
nor_5  g09662(new_n9728, new_n9725_1, new_n10039);
or_5   g09663(new_n10039, new_n10038, new_n10040);
not_8  g09664(new_n10040, new_n10041);
xor_4  g09665(new_n10036, new_n10034, new_n10042);
not_8  g09666(new_n10042, new_n10043);
nor_5  g09667(new_n10043, new_n10041, new_n10044);
nor_5  g09668(new_n10044, new_n10037, new_n10045);
xor_4  g09669(new_n10045, new_n10033, new_n10046);
not_8  g09670(new_n10046, new_n10047);
xor_4  g09671(new_n10047, new_n9887, new_n10048);
xor_4  g09672(new_n9884, new_n9883, new_n10049);
not_8  g09673(new_n10049, new_n10050);
xor_4  g09674(new_n10043, new_n10041, new_n10051);
and_5  g09675(new_n10051, new_n10050, new_n10052);
nor_5  g09676(new_n9729, new_n9676, new_n10053);
nor_5  g09677(new_n9734, new_n9731, new_n10054);
or_5   g09678(new_n10054, new_n10053, new_n10055);
xor_4  g09679(new_n10051, new_n10050, new_n10056);
not_8  g09680(new_n10056, new_n10057);
nor_5  g09681(new_n10057, new_n10055, new_n10058);
or_5   g09682(new_n10058, new_n10052, new_n10059);
xor_4  g09683(new_n10059, new_n10048, new_n10060);
not_8  g09684(new_n10060, new_n10061);
nor_5  g09685(new_n10061, new_n9815, new_n10062);
xor_4  g09686(new_n10061, new_n9815, new_n10063);
nand_5 g09687(new_n9502, new_n9480, new_n10064);
xor_4  g09688(new_n9812, new_n10064, new_n10065);
not_8  g09689(new_n10065, new_n10066);
xor_4  g09690(new_n10057, new_n10055, new_n10067);
and_5  g09691(new_n10067, new_n10066, new_n10068);
xor_4  g09692(new_n10067, new_n10065, new_n10069);
nor_5  g09693(new_n9648, new_n9504, new_n10070);
not_8  g09694(new_n9736, new_n10071);
nor_5  g09695(new_n10071, new_n9650, new_n10072);
or_5   g09696(new_n10072, new_n10070, new_n10073);
nor_5  g09697(new_n10073, new_n10069, new_n10074);
or_5   g09698(new_n10074, new_n10068, new_n10075);
and_5  g09699(new_n10075, new_n10063, new_n10076);
or_5   g09700(new_n10076, new_n10062, new_n10077);
nor_5  g09701(new_n9876, new_n9839, new_n10078);
nor_5  g09702(new_n9886, new_n9877, new_n10079);
nor_5  g09703(new_n10079, new_n10078, new_n10080);
nor_5  g09704(new_n10047, new_n9887, new_n10081);
and_5  g09705(new_n10059, new_n10048, new_n10082);
nor_5  g09706(new_n10082, new_n10081, new_n10083);
nor_5  g09707(new_n9784, new_n9783, new_n10084);
and_5  g09708(new_n9792, new_n9785, new_n10085);
nor_5  g09709(new_n10085, new_n10084, new_n10086);
and_5  g09710(n11662, n4312, new_n10087);
xor_4  g09711(new_n10087, new_n10086, new_n10088);
nor_5  g09712(new_n9858, new_n9857, new_n10089);
nor_5  g09713(new_n9867, new_n9860, new_n10090);
nor_5  g09714(new_n10090, new_n10089, new_n10091);
and_5  g09715(n12299, n10278, new_n10092);
xor_4  g09716(new_n10092, new_n10091, new_n10093);
and_5  g09717(new_n9849, new_n9848, new_n10094);
nor_5  g09718(new_n9851, new_n9847, new_n10095);
nor_5  g09719(new_n10095, new_n10094, new_n10096);
nand_5 g09720(n10451, n7436, new_n10097);
and_5  g09721(n9241, n3022, new_n10098);
xor_4  g09722(new_n10098, new_n10097, new_n10099);
nand_5 g09723(n11257, n3932, new_n10100);
and_5  g09724(n10327, n1097, new_n10101);
xor_4  g09725(new_n10101, new_n10100, new_n10102);
xor_4  g09726(new_n10102, new_n10099, new_n10103);
xor_4  g09727(new_n10103, new_n10096, new_n10104);
and_5  g09728(new_n10022_1, new_n10021, new_n10105);
nor_5  g09729(new_n10024, new_n10020, new_n10106);
nor_5  g09730(new_n10106, new_n10105, new_n10107);
nand_5 g09731(n2393, n159, new_n10108);
and_5  g09732(n5860, n2749, new_n10109);
xor_4  g09733(new_n10109, new_n10108, new_n10110);
xor_4  g09734(new_n10110, new_n10107, new_n10111);
xor_4  g09735(new_n10111, new_n10104, new_n10112);
xor_4  g09736(new_n10112, new_n10093, new_n10113);
xor_4  g09737(new_n10113, new_n10088, new_n10114);
nor_5  g09738(new_n9947, new_n9911, new_n10115);
nor_5  g09739(new_n9958, new_n9948, new_n10116);
nor_5  g09740(new_n10116, new_n10115, new_n10117);
xor_4  g09741(new_n10117, new_n10114, new_n10118);
and_5  g09742(new_n10002, new_n9998, new_n10119);
and_5  g09743(new_n10027, new_n10003, new_n10120);
or_5   g09744(new_n10120, new_n10119, new_n10121);
and_5  g09745(new_n10008, new_n10004, new_n10122);
or_5   g09746(new_n10122, new_n10005, new_n10123);
not_8  g09747(new_n10123, new_n10124);
and_5  g09748(n12247, n7388, new_n10125);
and_5  g09749(new_n10125, new_n10124, new_n10126);
and_5  g09750(new_n10125, new_n9961, new_n10127);
nor_5  g09751(new_n10127, new_n10124, new_n10128);
or_5   g09752(new_n10128, new_n10126, new_n10129);
nand_5 g09753(n10898, n5857, new_n10130);
nand_5 g09754(n12591, n12025, new_n10131);
and_5  g09755(n11876, n45, new_n10132);
xor_4  g09756(new_n10132, new_n10131, new_n10133);
xor_4  g09757(new_n10133, new_n10130, new_n10134);
xor_4  g09758(new_n10134, new_n10129, new_n10135);
xor_4  g09759(new_n10135, new_n10121, new_n10136);
and_5  g09760(new_n9864, new_n9863, new_n10137);
nor_5  g09761(new_n9866, new_n9862, new_n10138);
nor_5  g09762(new_n10138, new_n10137, new_n10139);
nand_5 g09763(n12705, n7456, new_n10140);
and_5  g09764(n11023, n8276, new_n10141);
xor_4  g09765(new_n10141, new_n10140, new_n10142);
xor_4  g09766(new_n10142, new_n10139, new_n10143);
nand_5 g09767(n9583, n5964, new_n10144);
and_5  g09768(n12511, n7965, new_n10145);
xor_4  g09769(new_n10145, new_n10144, new_n10146);
xor_4  g09770(new_n10146, new_n10143, new_n10147);
nor_5  g09771(new_n9872, new_n9871, new_n10148);
nor_5  g09772(new_n9874, new_n9869, new_n10149);
nor_5  g09773(new_n10149, new_n10148, new_n10150);
nor_5  g09774(new_n9868, new_n9856, new_n10151);
nor_5  g09775(new_n10151, new_n9854, new_n10152);
xor_4  g09776(new_n10152, new_n10150, new_n10153);
xor_4  g09777(new_n10153, new_n10147, new_n10154);
xor_4  g09778(new_n10154, new_n10136, new_n10155);
nor_5  g09779(new_n10029, new_n9995, new_n10156);
nor_5  g09780(new_n10030, new_n9994, new_n10157);
nor_5  g09781(new_n10157, new_n10156, new_n10158);
and_5  g09782(new_n9943, new_n9941, new_n10159);
nor_5  g09783(new_n9945, new_n9938_1, new_n10160);
or_5   g09784(new_n10160, new_n10159, new_n10161);
and_5  g09785(new_n9779, new_n9772, new_n10162);
nor_5  g09786(new_n9794, new_n9781, new_n10163);
nor_5  g09787(new_n10163, new_n10162, new_n10164);
xor_4  g09788(new_n10164, new_n10161, new_n10165);
nand_5 g09789(n3986, n3754, new_n10166);
and_5  g09790(n11423, n6776, new_n10167);
xor_4  g09791(new_n10167, new_n10166, new_n10168);
nand_5 g09792(n8759, n2278, new_n10169);
and_5  g09793(n10510, n9640, new_n10170);
xor_4  g09794(new_n10170, new_n10169, new_n10171);
xor_4  g09795(new_n10171, new_n10168, new_n10172);
and_5  g09796(n8476, n4094, new_n10173);
and_5  g09797(n5305, n753, new_n10174_1);
xor_4  g09798(new_n10174_1, new_n10173, new_n10175);
and_5  g09799(n3616, n1067, new_n10176);
and_5  g09800(n10644, n6703, new_n10177);
xor_4  g09801(new_n10177, new_n10176, new_n10178);
xor_4  g09802(new_n10178, new_n10175, new_n10179);
xor_4  g09803(new_n10179, new_n10172, new_n10180);
and_5  g09804(new_n9776, new_n9775, new_n10181);
nor_5  g09805(new_n9778, new_n9774, new_n10182);
or_5   g09806(new_n10182, new_n10181, new_n10183);
and_5  g09807(new_n9789, new_n9788, new_n10184);
nor_5  g09808(new_n9791, new_n9787, new_n10185);
nor_5  g09809(new_n10185, new_n10184, new_n10186);
xor_4  g09810(new_n10186, new_n10183, new_n10187);
xor_4  g09811(new_n10187, new_n10180, new_n10188);
xor_4  g09812(new_n10188, new_n10165, new_n10189);
and_5  g09813(new_n9800, new_n9798, new_n10190);
nor_5  g09814(new_n9802, new_n9795, new_n10191);
nor_5  g09815(new_n10191, new_n10190, new_n10192);
and_5  g09816(new_n10013, new_n10009, new_n10193);
nor_5  g09817(new_n9972, new_n9971, new_n10194);
xor_4  g09818(new_n10017, new_n10194, new_n10195);
xor_4  g09819(new_n10025, new_n10195, new_n10196);
and_5  g09820(new_n10196, new_n10014, new_n10197);
or_5   g09821(new_n10197, new_n10193, new_n10198);
nor_5  g09822(new_n10016, new_n10015, new_n10199);
nor_5  g09823(new_n10025, new_n10018, new_n10200);
or_5   g09824(new_n10200, new_n10199, new_n10201);
and_5  g09825(new_n9920_1, new_n9919, new_n10202);
not_8  g09826(new_n9918, new_n10203);
nor_5  g09827(new_n9922, new_n10203, new_n10204);
or_5   g09828(new_n10204, new_n10202, new_n10205);
and_5  g09829(n10547, n1798, new_n10206);
and_5  g09830(n8665, n7690, new_n10207);
xor_4  g09831(new_n10207, new_n10206, new_n10208);
nand_5 g09832(n12826, n2530, new_n10209);
and_5  g09833(n11892, n1510, new_n10210);
xor_4  g09834(new_n10210, new_n10209, new_n10211);
xor_4  g09835(new_n10211, new_n10208, new_n10212);
xor_4  g09836(new_n10212, new_n10205, new_n10213);
xor_4  g09837(new_n10213, new_n10201, new_n10214);
xor_4  g09838(new_n10214, new_n10198, new_n10215);
nand_5 g09839(n11922, n10545, new_n10216);
nor_5  g09840(new_n9936, new_n9928, new_n10217_1);
and_5  g09841(new_n9937, new_n9925, new_n10218);
nor_5  g09842(new_n10218, new_n10217_1, new_n10219);
xor_4  g09843(new_n10219, new_n10216, new_n10220);
and_5  g09844(new_n9916, new_n9914, new_n10221);
and_5  g09845(new_n9923, new_n9917, new_n10222);
or_5   g09846(new_n10222, new_n10221, new_n10223_1);
and_5  g09847(new_n9932, new_n9931, new_n10224);
nor_5  g09848(new_n9934, new_n9930, new_n10225);
nor_5  g09849(new_n10225, new_n10224, new_n10226);
xor_4  g09850(new_n10226, new_n10223_1, new_n10227);
and_5  g09851(n12648, n2551, new_n10228);
nand_5 g09852(n10685, n5331, new_n10229);
and_5  g09853(n5645, n4499, new_n10230);
xor_4  g09854(new_n10230, new_n10229, new_n10231);
xor_4  g09855(new_n10231, new_n10228, new_n10232);
xor_4  g09856(new_n10232, new_n10227, new_n10233);
xor_4  g09857(new_n10233, new_n10220, new_n10234);
xor_4  g09858(new_n10234, new_n10215, new_n10235);
xor_4  g09859(new_n10235, new_n10192, new_n10236);
xor_4  g09860(new_n10236, new_n10189, new_n10237);
xor_4  g09861(new_n10237, new_n10158, new_n10238);
xor_4  g09862(new_n10238, new_n10155, new_n10239);
xor_4  g09863(new_n10239, new_n10118, new_n10240);
nor_5  g09864(new_n9804, new_n9768, new_n10241);
nor_5  g09865(new_n9814, new_n9805, new_n10242);
nor_5  g09866(new_n10242, new_n10241, new_n10243);
and_5  g09867(new_n10031, new_n9960, new_n10244);
nor_5  g09868(new_n10045, new_n10033, new_n10245);
nor_5  g09869(new_n10245, new_n10244, new_n10246);
xor_4  g09870(new_n10246, new_n10243, new_n10247);
xor_4  g09871(new_n10247, new_n10240, new_n10248);
xor_4  g09872(new_n10248, new_n10083, new_n10249);
xor_4  g09873(new_n10249, new_n10080, new_n10250);
xor_4  g09874(new_n10250, new_n10077, n4230);
nor_5  g09875(new_n5791, new_n5779, new_n10252);
xor_4  g09876(new_n5795, new_n10252, n4300);
xor_4  g09877(new_n3533, new_n3532, n4326);
not_8  g09878(new_n1264, new_n10255);
nand_5 g09879(new_n10255, new_n1257, new_n10256);
not_8  g09880(new_n10256, new_n10257);
nand_5 g09881(n6687, n5320, new_n10258);
nor_5  g09882(new_n1248, new_n1237, new_n10259);
nor_5  g09883(new_n1256, new_n1249, new_n10260);
nor_5  g09884(new_n10260, new_n10259, new_n10261);
xor_4  g09885(new_n10261, new_n10258, new_n10262);
not_8  g09886(new_n10262, new_n10263);
nand_5 g09887(n4370, n2564, new_n10264);
not_8  g09888(new_n10264, new_n10265);
and_5  g09889(new_n1253, new_n1252, new_n10266);
nor_5  g09890(new_n1255, new_n1251, new_n10267);
or_5   g09891(new_n10267, new_n10266, new_n10268);
not_8  g09892(new_n10268, new_n10269);
xor_4  g09893(new_n10269, new_n10265, new_n10270);
nand_5 g09894(n6770, n5212, new_n10271);
nand_5 g09895(n11877, n4189, new_n10272);
nand_5 g09896(n11407, n9920, new_n10273);
xor_4  g09897(new_n10273, new_n10272, new_n10274);
not_8  g09898(new_n10274, new_n10275);
xor_4  g09899(new_n10275, new_n10271, new_n10276);
xor_4  g09900(new_n10276, new_n10270, new_n10277);
not_8  g09901(new_n10277, new_n10278_1);
xor_4  g09902(new_n10278_1, new_n10263, new_n10279);
xor_4  g09903(new_n10279, new_n10257, new_n10280);
not_8  g09904(new_n10280, new_n10281);
or_5   g09905(new_n1376, new_n1375, new_n10282);
not_8  g09906(new_n10282, new_n10283);
nand_5 g09907(n8336, n2433, new_n10284);
not_8  g09908(new_n10284, new_n10285);
nand_5 g09909(n10928, n8819, new_n10286);
not_8  g09910(new_n10286, new_n10287);
and_5  g09911(new_n1367, new_n1366, new_n10288);
nor_5  g09912(new_n1367, new_n1366, new_n10289);
nor_5  g09913(new_n10289, new_n1365, new_n10290);
or_5   g09914(new_n10290, new_n10288, new_n10291);
not_8  g09915(new_n10291, new_n10292);
and_5  g09916(new_n10292, new_n10287, new_n10293);
nor_5  g09917(new_n10292, new_n10287, new_n10294);
or_5   g09918(new_n10294, new_n10293, new_n10295);
nand_5 g09919(n11728, n2226, new_n10296);
not_8  g09920(new_n10296, new_n10297);
nand_5 g09921(n12709, n1094, new_n10298);
xor_4  g09922(new_n10298, new_n1297, new_n10299);
xor_4  g09923(new_n10299, new_n10297, new_n10300);
not_8  g09924(new_n10300, new_n10301);
xor_4  g09925(new_n10301, new_n10295, new_n10302);
xor_4  g09926(new_n10302, new_n10285, new_n10303);
not_8  g09927(new_n10303, new_n10304);
nor_5  g09928(new_n1370, new_n1363, new_n10305);
and_5  g09929(new_n1373, new_n1371, new_n10306);
nor_5  g09930(new_n10306, new_n10305, new_n10307);
xor_4  g09931(new_n10307, new_n10304, new_n10308);
xor_4  g09932(new_n10308, new_n10283, new_n10309);
not_8  g09933(new_n10309, new_n10310);
not_8  g09934(new_n1377, new_n10311);
nor_5  g09935(new_n1418, new_n10311, new_n10312);
nor_5  g09936(new_n1421, new_n1419, new_n10313);
nor_5  g09937(new_n10313, new_n10312, new_n10314);
xor_4  g09938(new_n10314, new_n10310, new_n10315);
not_8  g09939(new_n10315, new_n10316);
nand_5 g09940(new_n1391, new_n1390, new_n10317);
nand_5 g09941(n12069, n11967, new_n10318);
not_8  g09942(new_n10318, new_n10319);
nand_5 g09943(n12391, n6254, new_n10320);
not_8  g09944(new_n10320, new_n10321);
and_5  g09945(new_n1386, new_n1385, new_n10322);
not_8  g09946(new_n1384, new_n10323);
nor_5  g09947(new_n1388, new_n10323, new_n10324);
nor_5  g09948(new_n10324, new_n10322, new_n10325);
xor_4  g09949(new_n10325, new_n10321, new_n10326);
not_8  g09950(new_n10326, new_n10327_1);
nand_5 g09951(n7160, n7159, new_n10328);
not_8  g09952(new_n10328, new_n10329);
nand_5 g09953(n12777, n7891, new_n10330);
nand_5 g09954(n12489, n4828, new_n10331);
xor_4  g09955(new_n10331, new_n10330, new_n10332);
xor_4  g09956(new_n10332, new_n10329, new_n10333);
not_8  g09957(new_n10333, new_n10334);
xor_4  g09958(new_n10334, new_n10327_1, new_n10335);
xor_4  g09959(new_n10335, new_n10319, new_n10336);
or_5   g09960(new_n1382, new_n1378, new_n10337);
not_8  g09961(new_n10337, new_n10338);
and_5  g09962(new_n1389, new_n1383, new_n10339);
or_5   g09963(new_n10339, new_n10338, new_n10340);
xor_4  g09964(new_n10340, new_n10336, new_n10341);
not_8  g09965(new_n10341, new_n10342);
xor_4  g09966(new_n10342, new_n10317, new_n10343);
nand_5 g09967(new_n1410, new_n1408, new_n10344);
nand_5 g09968(n12947, n11222, new_n10345);
not_8  g09969(new_n10345, new_n10346);
nand_5 g09970(n11791, n11153, new_n10347);
not_8  g09971(new_n10347, new_n10348);
and_5  g09972(new_n1404, new_n1403, new_n10349);
nor_5  g09973(new_n1406, new_n1402, new_n10350);
nor_5  g09974(new_n10350, new_n10349, new_n10351);
xor_4  g09975(new_n10351, new_n10348, new_n10352);
not_8  g09976(new_n10352, new_n10353);
nand_5 g09977(n5760, n996, new_n10354);
not_8  g09978(new_n10354, new_n10355);
nand_5 g09979(n5314, n1478, new_n10356);
nand_5 g09980(n10990, n5767, new_n10357);
xor_4  g09981(new_n10357, new_n10356, new_n10358);
xor_4  g09982(new_n10358, new_n10355, new_n10359);
not_8  g09983(new_n10359, new_n10360);
xor_4  g09984(new_n10360, new_n10353, new_n10361);
xor_4  g09985(new_n10361, new_n10346, new_n10362);
nor_5  g09986(new_n1399, new_n1393, new_n10363);
nor_5  g09987(new_n1407, new_n1400, new_n10364);
or_5   g09988(new_n10364, new_n10363, new_n10365);
xor_4  g09989(new_n10365, new_n10362, new_n10366);
not_8  g09990(new_n10366, new_n10367);
xor_4  g09991(new_n10367, new_n10344, new_n10368);
nor_5  g09992(new_n1411, new_n1392, new_n10369);
and_5  g09993(new_n1417, new_n1412, new_n10370);
or_5   g09994(new_n10370, new_n10369, new_n10371);
not_8  g09995(new_n10371, new_n10372);
xor_4  g09996(new_n10372, new_n10368, new_n10373);
xor_4  g09997(new_n10373, new_n10343, new_n10374);
xnor_4 g09998(new_n10374, new_n10316, new_n10375);
xor_4  g09999(new_n10375, new_n10281, new_n10376);
and_5  g10000(new_n1361, new_n1266, new_n10377);
not_8  g10001(new_n1423, new_n10378);
and_5  g10002(new_n10378, new_n1362, new_n10379);
nor_5  g10003(new_n10379, new_n10377, new_n10380);
xor_4  g10004(new_n10380, new_n10376, n4333);
nand_5 g10005(n11877, n11757, new_n10382);
not_8  g10006(new_n10382, new_n10383);
nand_5 g10007(n5240, n5212, new_n10384);
nand_5 g10008(n11821, n11407, new_n10385);
xor_4  g10009(new_n10385, new_n10384, new_n10386);
xor_4  g10010(new_n10386, new_n10383, new_n10387);
not_8  g10011(new_n10387, new_n10388);
nand_5 g10012(n11407, n5240, new_n10389);
nand_5 g10013(n11877, n3172, new_n10390);
and_5  g10014(new_n10390, new_n10389, new_n10391_1);
nand_5 g10015(n11757, n5212, new_n10392);
not_8  g10016(new_n10392, new_n10393);
xor_4  g10017(new_n10390, new_n10389, new_n10394);
not_8  g10018(new_n10394, new_n10395);
nor_5  g10019(new_n10395, new_n10393, new_n10396);
nor_5  g10020(new_n10396, new_n10391_1, new_n10397);
xor_4  g10021(new_n10397, new_n10388, new_n10398);
nand_5 g10022(n5320, n1333, new_n10399);
nand_5 g10023(n4370, n3172, new_n10400);
xor_4  g10024(new_n10400, new_n10399, new_n10401);
xor_4  g10025(new_n10401, new_n10398, new_n10402);
nand_5 g10026(n4370, n1333, new_n10403);
not_8  g10027(new_n10403, new_n10404);
nand_5 g10028(n11877, n1333, new_n10405);
nand_5 g10029(n11757, n11407, new_n10406);
and_5  g10030(new_n10406, new_n10405, new_n10407);
nand_5 g10031(n5212, n3172, new_n10408);
not_8  g10032(new_n10408, new_n10409);
xor_4  g10033(new_n10406, new_n10405, new_n10410);
not_8  g10034(new_n10410, new_n10411);
nor_5  g10035(new_n10411, new_n10409, new_n10412);
or_5   g10036(new_n10412, new_n10407, new_n10413);
not_8  g10037(new_n10413, new_n10414);
and_5  g10038(new_n10414, new_n10404, new_n10415);
xor_4  g10039(new_n10414, new_n10403, new_n10416);
xor_4  g10040(new_n10395, new_n10393, new_n10417);
nor_5  g10041(new_n10417, new_n10416, new_n10418);
nor_5  g10042(new_n10418, new_n10415, new_n10419);
xor_4  g10043(new_n10419, new_n10402, new_n10420);
nand_5 g10044(n7862, n5320, new_n10421);
not_8  g10045(new_n10421, new_n10422);
xor_4  g10046(new_n10417, new_n10416, new_n10423);
nor_5  g10047(new_n10423, new_n10422, new_n10424);
xor_4  g10048(new_n10423, new_n10422, new_n10425);
not_8  g10049(new_n10425, new_n10426);
nand_5 g10050(n7862, n4370, new_n10427);
not_8  g10051(new_n10427, new_n10428);
and_5  g10052(n11407, n3172, new_n10429);
and_5  g10053(n11877, n7862, new_n10430);
or_5   g10054(new_n10430, new_n10429, new_n10431);
not_8  g10055(new_n10431, new_n10432);
nand_5 g10056(n11407, n7862, new_n10433);
nor_5  g10057(new_n10433, new_n10390, new_n10434);
nand_5 g10058(n5212, n1333, new_n10435);
not_8  g10059(new_n10435, new_n10436);
nor_5  g10060(new_n10436, new_n10434, new_n10437);
or_5   g10061(new_n10437, new_n10432, new_n10438);
not_8  g10062(new_n10438, new_n10439_1);
and_5  g10063(new_n10439_1, new_n10428, new_n10440);
xor_4  g10064(new_n10439_1, new_n10428, new_n10441);
xor_4  g10065(new_n10411, new_n10408, new_n10442);
and_5  g10066(new_n10442, new_n10441, new_n10443);
or_5   g10067(new_n10443, new_n10440, new_n10444);
nor_5  g10068(new_n10444, new_n10426, new_n10445);
or_5   g10069(new_n10445, new_n10424, new_n10446);
not_8  g10070(new_n10446, new_n10447);
nand_5 g10071(new_n10447, new_n10420, new_n10448);
not_8  g10072(new_n10401, new_n10449);
or_5   g10073(new_n10449, new_n10398, new_n10450);
or_5   g10074(new_n10400, new_n10399, new_n10451_1);
or_5   g10075(new_n10419, new_n10402, new_n10452);
not_8  g10076(new_n10452, new_n10453);
xor_4  g10077(new_n10453, new_n10451_1, new_n10454);
nand_5 g10078(new_n10454, new_n10450, new_n10455);
or_5   g10079(new_n10385, new_n10384, new_n10456);
not_8  g10080(new_n10456, new_n10457);
and_5  g10081(n11757, n4370, new_n10458);
xor_4  g10082(new_n10458, new_n10457, new_n10459);
nand_5 g10083(n11821, n5212, new_n10460);
not_8  g10084(new_n10460, new_n10461);
nand_5 g10085(n11877, n5240, new_n10462);
nand_5 g10086(n11407, n9080, new_n10463);
xor_4  g10087(new_n10463, new_n10462, new_n10464);
not_8  g10088(new_n10464, new_n10465);
xor_4  g10089(new_n10465, new_n10461, new_n10466);
xor_4  g10090(new_n10466, new_n10459, new_n10467);
not_8  g10091(new_n10467, new_n10468);
nor_5  g10092(new_n10386, new_n10383, new_n10469);
nor_5  g10093(new_n10397, new_n10388, new_n10470);
or_5   g10094(new_n10470, new_n10469, new_n10471);
not_8  g10095(new_n10471, new_n10472);
nand_5 g10096(n12000, n1333, new_n10473);
not_8  g10097(new_n10473, new_n10474);
nand_5 g10098(n5320, n3172, new_n10475);
nand_5 g10099(n9725, n7862, new_n10476_1);
xor_4  g10100(new_n10476_1, new_n10475, new_n10477);
not_8  g10101(new_n10477, new_n10478);
xor_4  g10102(new_n10478, new_n10474, new_n10479);
not_8  g10103(new_n10479, new_n10480);
xor_4  g10104(new_n10480, new_n10472, new_n10481);
xor_4  g10105(new_n10481, new_n10468, new_n10482);
xor_4  g10106(new_n10482, new_n10455, new_n10483);
xnor_4 g10107(new_n10483, new_n10448, new_n10484);
nand_5 g10108(n12000, n7862, new_n10485);
not_8  g10109(new_n10485, new_n10486);
xor_4  g10110(new_n10447, new_n10420, new_n10487);
nor_5  g10111(new_n10487, new_n10486, new_n10488);
xor_4  g10112(new_n10442, new_n10441, new_n10489);
or_5   g10113(new_n10434, new_n10432, new_n10490);
nand_5 g10114(n11407, n1333, new_n10491);
nand_5 g10115(n7862, n5212, new_n10492);
nor_5  g10116(new_n10492, new_n10491, new_n10493);
and_5  g10117(new_n10493, new_n10490, new_n10494);
nand_5 g10118(new_n10494, new_n10489, new_n10495);
not_8  g10119(new_n10444, new_n10496);
xnor_4 g10120(new_n10496, new_n10426, new_n10497);
or_5   g10121(new_n10497, new_n10495, new_n10498);
xor_4  g10122(new_n10487, new_n10486, new_n10499);
and_5  g10123(new_n10499, new_n10498, new_n10500);
or_5   g10124(new_n10500, new_n10488, new_n10501);
not_8  g10125(new_n10501, new_n10502);
and_5  g10126(new_n10502, new_n10484, new_n10503);
nor_5  g10127(new_n10502, new_n10484, new_n10504);
or_5   g10128(new_n10504, new_n10503, new_n10505);
not_8  g10129(new_n10505, new_n10506);
nand_5 g10130(n8819, n6877, new_n10507);
nand_5 g10131(n12709, n2464, new_n10508);
nand_5 g10132(n6877, n6429, new_n10509);
nor_5  g10133(new_n10509, new_n10508, new_n10510_1);
and_5  g10134(new_n10509, new_n10508, new_n10511);
nand_5 g10135(n11728, n9400, new_n10512);
nor_5  g10136(new_n10512, new_n10511, new_n10513);
nor_5  g10137(new_n10513, new_n10510_1, new_n10514);
xor_4  g10138(new_n10514, new_n10507, new_n10515);
not_8  g10139(new_n10515, new_n10516);
nand_5 g10140(n11728, n2464, new_n10517);
not_8  g10141(new_n10517, new_n10518);
nand_5 g10142(n12709, n11311, new_n10519);
nand_5 g10143(n9400, n6429, new_n10520);
xor_4  g10144(new_n10520, new_n10519, new_n10521);
xor_4  g10145(new_n10521, new_n10518, new_n10522);
not_8  g10146(new_n10522, new_n10523);
nor_5  g10147(new_n10523, new_n10516, new_n10524);
and_5  g10148(new_n10523, new_n10516, new_n10525);
or_5   g10149(new_n10525, new_n10524, new_n10526);
xor_4  g10150(new_n10509, new_n10508, new_n10527);
nand_5 g10151(n12709, n9400, new_n10528);
nand_5 g10152(n11728, n6877, new_n10529);
or_5   g10153(new_n10529, new_n10528, new_n10530);
or_5   g10154(new_n10530, new_n10527, new_n10531);
or_5   g10155(new_n10531, new_n10526, new_n10532);
not_8  g10156(new_n10532, new_n10533);
nand_5 g10157(n6877, n2433, new_n10534);
not_8  g10158(new_n10534, new_n10535);
nand_5 g10159(n9400, n8819, new_n10536);
not_8  g10160(new_n10536, new_n10537);
and_5  g10161(new_n10520, new_n10519, new_n10538);
nor_5  g10162(new_n10520, new_n10519, new_n10539);
nor_5  g10163(new_n10539, new_n10518, new_n10540);
or_5   g10164(new_n10540, new_n10538, new_n10541);
not_8  g10165(new_n10541, new_n10542);
and_5  g10166(new_n10542, new_n10537, new_n10543);
nor_5  g10167(new_n10542, new_n10537, new_n10544);
or_5   g10168(new_n10544, new_n10543, new_n10545_1);
nand_5 g10169(n11728, n11311, new_n10546);
not_8  g10170(new_n10546, new_n10547_1);
nand_5 g10171(n6429, n2464, new_n10548);
nand_5 g10172(n12709, n4187, new_n10549);
xor_4  g10173(new_n10549, new_n10548, new_n10550);
not_8  g10174(new_n10550, new_n10551);
xor_4  g10175(new_n10551, new_n10547_1, new_n10552);
xor_4  g10176(new_n10552, new_n10545_1, new_n10553);
xor_4  g10177(new_n10553, new_n10535, new_n10554);
not_8  g10178(new_n10554, new_n10555);
nor_5  g10179(new_n10514, new_n10507, new_n10556);
nor_5  g10180(new_n10524, new_n10556, new_n10557);
xor_4  g10181(new_n10557, new_n10555, new_n10558);
nand_5 g10182(new_n10558, new_n10533, new_n10559);
not_8  g10183(new_n10559, new_n10560);
nand_5 g10184(n8717, n6877, new_n10561);
nand_5 g10185(n11311, n6429, new_n10562);
nand_5 g10186(n12709, n4203, new_n10563);
nand_5 g10187(n11728, n4187, new_n10564);
xor_4  g10188(new_n10564, new_n10563, new_n10565);
not_8  g10189(new_n10565, new_n10566);
xor_4  g10190(new_n10566, new_n10562, new_n10567);
and_5  g10191(new_n10549, new_n10548, new_n10568);
nor_5  g10192(new_n10551, new_n10547_1, new_n10569);
or_5   g10193(new_n10569, new_n10568, new_n10570);
not_8  g10194(new_n10570, new_n10571);
xor_4  g10195(new_n10571, new_n10567, new_n10572);
nand_5 g10196(n9400, n2433, new_n10573);
nand_5 g10197(n8819, n2464, new_n10574);
xor_4  g10198(new_n10574, new_n10573, new_n10575);
xor_4  g10199(new_n10575, new_n10572, new_n10576);
not_8  g10200(new_n10576, new_n10577);
nor_5  g10201(new_n10552, new_n10545_1, new_n10578);
nor_5  g10202(new_n10578, new_n10543, new_n10579);
xor_4  g10203(new_n10579, new_n10577, new_n10580);
not_8  g10204(new_n10580, new_n10581);
and_5  g10205(new_n10553, new_n10535, new_n10582);
nor_5  g10206(new_n10557, new_n10555, new_n10583);
nor_5  g10207(new_n10583, new_n10582, new_n10584);
xor_4  g10208(new_n10584, new_n10581, new_n10585);
not_8  g10209(new_n10585, new_n10586);
xor_4  g10210(new_n10586, new_n10561, new_n10587);
xor_4  g10211(new_n10587, new_n10560, new_n10588);
xor_4  g10212(new_n10558, new_n10533, new_n10589_1);
not_8  g10213(new_n10589_1, new_n10590);
xor_4  g10214(new_n10531, new_n10526, new_n10591);
not_8  g10215(new_n10591, new_n10592);
nand_5 g10216(n12489, n4805, new_n10593);
nand_5 g10217(n10990, n7236, new_n10594);
or_5   g10218(new_n10594, new_n10593, new_n10595);
not_8  g10219(new_n10595, new_n10596);
and_5  g10220(n12489, n11478, new_n10597);
and_5  g10221(n7159, n4805, new_n10598);
xor_4  g10222(new_n10598, new_n10597, new_n10599);
nor_5  g10223(new_n10599, new_n10596, new_n10600);
xor_4  g10224(new_n10599, new_n10595, new_n10601);
not_8  g10225(new_n10601, new_n10602);
nand_5 g10226(n10990, n3992, new_n10603);
and_5  g10227(n7236, n5760, new_n10604);
xor_4  g10228(new_n10604, new_n10603, new_n10605);
and_5  g10229(new_n10605, new_n10602, new_n10606);
or_5   g10230(new_n10606, new_n10600, new_n10607);
not_8  g10231(new_n10607, new_n10608);
nand_5 g10232(n10990, n8384, new_n10609);
nand_5 g10233(n7236, n1478, new_n10610);
nor_5  g10234(new_n10610, new_n10609, new_n10611);
not_8  g10235(new_n10594, new_n10612);
nand_5 g10236(n5760, n3992, new_n10613);
or_5   g10237(new_n10613, new_n10612, new_n10614);
nand_5 g10238(new_n10610, new_n10609, new_n10615);
not_8  g10239(new_n10615, new_n10616);
and_5  g10240(new_n10616, new_n10614, new_n10617);
or_5   g10241(new_n10617, new_n10611, new_n10618);
not_8  g10242(new_n10618, new_n10619);
or_5   g10243(new_n10616, new_n10614, new_n10620);
and_5  g10244(new_n10620, new_n10619, new_n10621);
nor_5  g10245(new_n10621, new_n10608, new_n10622);
xor_4  g10246(new_n10621, new_n10607, new_n10623);
nand_5 g10247(n11478, n7159, new_n10624);
not_8  g10248(new_n10624, new_n10625);
and_5  g10249(new_n10625, new_n10593, new_n10626);
nand_5 g10250(n12489, n5283, new_n10627);
nand_5 g10251(n12777, n4805, new_n10628);
xor_4  g10252(new_n10628, new_n10627, new_n10629);
nor_5  g10253(new_n10629, new_n10626, new_n10630);
nand_5 g10254(new_n10628, new_n10627, new_n10631);
and_5  g10255(new_n10631, new_n10626, new_n10632);
nor_5  g10256(new_n10632, new_n10630, new_n10633);
nor_5  g10257(new_n10633, new_n10623, new_n10634);
or_5   g10258(new_n10634, new_n10622, new_n10635);
not_8  g10259(new_n10635, new_n10636);
nand_5 g10260(n6254, n4805, new_n10637);
nor_5  g10261(new_n10628, new_n10627, new_n10638);
and_5  g10262(new_n10628, new_n10627, new_n10639);
nor_5  g10263(new_n10639, new_n10624, new_n10640);
nor_5  g10264(new_n10640, new_n10638, new_n10641);
xor_4  g10265(new_n10641, new_n10637, new_n10642);
not_8  g10266(new_n10642, new_n10643);
nand_5 g10267(n7159, n5283, new_n10644_1);
nand_5 g10268(n12489, n137, new_n10645);
nand_5 g10269(n12777, n11478, new_n10646);
xnor_4 g10270(new_n10646, new_n10645, new_n10647);
not_8  g10271(new_n10647, new_n10648);
xor_4  g10272(new_n10648, new_n10644_1, new_n10649);
nor_5  g10273(new_n10649, new_n10643, new_n10650);
and_5  g10274(new_n10649, new_n10643, new_n10651);
or_5   g10275(new_n10651, new_n10650, new_n10652);
nand_5 g10276(new_n10598, new_n10597, new_n10653);
or_5   g10277(new_n10629, new_n10653, new_n10654);
xor_4  g10278(new_n10654, new_n10652, new_n10655);
nand_5 g10279(n11791, n7236, new_n10656);
not_8  g10280(new_n10613, new_n10657);
nor_5  g10281(new_n10657, new_n10611, new_n10658);
or_5   g10282(new_n10658, new_n10616, new_n10659);
not_8  g10283(new_n10659, new_n10660);
xor_4  g10284(new_n10660, new_n10656, new_n10661);
nand_5 g10285(n8384, n5760, new_n10662);
nand_5 g10286(n10990, n6358, new_n10663);
nand_5 g10287(n3992, n1478, new_n10664);
xnor_4 g10288(new_n10664, new_n10663, new_n10665);
not_8  g10289(new_n10665, new_n10666);
xor_4  g10290(new_n10666, new_n10662, new_n10667);
xor_4  g10291(new_n10667, new_n10661, new_n10668);
nor_5  g10292(new_n10619, new_n10613, new_n10669);
xor_4  g10293(new_n10669, new_n10668, new_n10670);
xor_4  g10294(new_n10670, new_n10655, new_n10671);
not_8  g10295(new_n10671, new_n10672);
xor_4  g10296(new_n10672, new_n10636, new_n10673);
nor_5  g10297(new_n10673, new_n10592, new_n10674);
xor_4  g10298(new_n10673, new_n10591, new_n10675);
xor_4  g10299(new_n10633, new_n10623, new_n10676);
not_8  g10300(new_n10676, new_n10677);
not_8  g10301(new_n10512, new_n10678_1);
nand_5 g10302(n12709, n6877, new_n10679);
and_5  g10303(new_n10679, new_n10678_1, new_n10680);
nor_5  g10304(new_n10680, new_n10527, new_n10681);
nand_5 g10305(new_n10509, new_n10508, new_n10682);
and_5  g10306(new_n10680, new_n10682, new_n10683);
or_5   g10307(new_n10683, new_n10681, new_n10684);
not_8  g10308(new_n10684, new_n10685_1);
and_5  g10309(new_n10685_1, new_n10677, new_n10686);
xor_4  g10310(new_n10684, new_n10677, new_n10687);
xor_4  g10311(new_n10605, new_n10602, new_n10688);
xor_4  g10312(new_n10529, new_n10528, new_n10689);
not_8  g10313(new_n10689, new_n10690);
nor_5  g10314(new_n10690, new_n10688, new_n10691);
xor_4  g10315(new_n10594, new_n10593, new_n10692);
not_8  g10316(new_n10692, new_n10693);
or_5   g10317(new_n10693, new_n10679, new_n10694);
not_8  g10318(new_n10694, new_n10695_1);
xor_4  g10319(new_n10690, new_n10688, new_n10696);
and_5  g10320(new_n10696, new_n10695_1, new_n10697);
nor_5  g10321(new_n10697, new_n10691, new_n10698);
nor_5  g10322(new_n10698, new_n10687, new_n10699);
nor_5  g10323(new_n10699, new_n10686, new_n10700);
nor_5  g10324(new_n10700, new_n10675, new_n10701);
or_5   g10325(new_n10701, new_n10674, new_n10702);
not_8  g10326(new_n10702, new_n10703);
and_5  g10327(new_n10703, new_n10590, new_n10704);
nor_5  g10328(new_n10703, new_n10590, new_n10705);
or_5   g10329(new_n10705, new_n10704, new_n10706);
or_5   g10330(new_n10654, new_n10652, new_n10707);
nand_5 g10331(n7159, n137, new_n10708);
not_8  g10332(new_n10708, new_n10709);
nand_5 g10333(n12777, n5283, new_n10710);
nand_5 g10334(n12489, n6294, new_n10711);
xor_4  g10335(new_n10711, new_n10710, new_n10712);
not_8  g10336(new_n10712, new_n10713);
xor_4  g10337(new_n10713, new_n10709, new_n10714);
not_8  g10338(new_n10714, new_n10715);
nand_5 g10339(n11478, n6254, new_n10716);
not_8  g10340(new_n10716, new_n10717);
and_5  g10341(new_n10646, new_n10645, new_n10718);
and_5  g10342(new_n10648, new_n10644_1, new_n10719);
or_5   g10343(new_n10719, new_n10718, new_n10720);
not_8  g10344(new_n10720, new_n10721);
xor_4  g10345(new_n10721, new_n10717, new_n10722);
xor_4  g10346(new_n10722, new_n10715, new_n10723);
nand_5 g10347(n11967, n4805, new_n10724);
not_8  g10348(new_n10724, new_n10725);
nor_5  g10349(new_n10641, new_n10637, new_n10726);
or_5   g10350(new_n10650, new_n10726, new_n10727);
xor_4  g10351(new_n10727, new_n10725, new_n10728);
not_8  g10352(new_n10728, new_n10729);
xor_4  g10353(new_n10729, new_n10723, new_n10730);
xor_4  g10354(new_n10730, new_n10707, new_n10731);
nand_5 g10355(new_n10669, new_n10668, new_n10732);
nand_5 g10356(n6358, n5760, new_n10733);
not_8  g10357(new_n10733, new_n10734);
nand_5 g10358(n8384, n1478, new_n10735);
nand_5 g10359(n10990, n5198, new_n10736);
xor_4  g10360(new_n10736, new_n10735, new_n10737);
not_8  g10361(new_n10737, new_n10738);
xor_4  g10362(new_n10738, new_n10734, new_n10739);
not_8  g10363(new_n10739, new_n10740);
nand_5 g10364(n11791, n3992, new_n10741);
not_8  g10365(new_n10741, new_n10742);
and_5  g10366(new_n10664, new_n10663, new_n10743);
and_5  g10367(new_n10666, new_n10662, new_n10744);
or_5   g10368(new_n10744, new_n10743, new_n10745);
not_8  g10369(new_n10745, new_n10746);
xor_4  g10370(new_n10746, new_n10742, new_n10747);
xor_4  g10371(new_n10747, new_n10740, new_n10748);
not_8  g10372(new_n10748, new_n10749);
nand_5 g10373(n12947, n7236, new_n10750);
not_8  g10374(new_n10750, new_n10751);
not_8  g10375(new_n10656, new_n10752);
and_5  g10376(new_n10660, new_n10752, new_n10753);
nor_5  g10377(new_n10667, new_n10661, new_n10754);
nor_5  g10378(new_n10754, new_n10753, new_n10755);
not_8  g10379(new_n10755, new_n10756);
xor_4  g10380(new_n10756, new_n10751, new_n10757);
xor_4  g10381(new_n10757, new_n10749, new_n10758);
xor_4  g10382(new_n10758, new_n10732, new_n10759);
not_8  g10383(new_n10759, new_n10760);
xor_4  g10384(new_n10760, new_n10731, new_n10761);
nor_5  g10385(new_n10670, new_n10655, new_n10762);
nor_5  g10386(new_n10672, new_n10636, new_n10763);
or_5   g10387(new_n10763, new_n10762, new_n10764);
xor_4  g10388(new_n10764, new_n10761, new_n10765);
nor_5  g10389(new_n10765, new_n10706, new_n10766);
nor_5  g10390(new_n10766, new_n10704, new_n10767);
nor_5  g10391(new_n10767, new_n10588, new_n10768);
or_5   g10392(new_n10758, new_n10732, new_n10769);
not_8  g10393(new_n10769, new_n10770);
nand_5 g10394(n7236, n6441, new_n10771);
not_8  g10395(new_n10771, new_n10772);
and_5  g10396(new_n10746, new_n10742, new_n10773);
and_5  g10397(new_n10747, new_n10740, new_n10774);
or_5   g10398(new_n10774, new_n10773, new_n10775);
not_8  g10399(new_n10775, new_n10776);
nand_5 g10400(n12947, n3992, new_n10777);
nand_5 g10401(n11791, n8384, new_n10778);
xor_4  g10402(new_n10778, new_n10777, new_n10779);
not_8  g10403(new_n10779, new_n10780);
xor_4  g10404(new_n10780, new_n10776, new_n10781);
nand_5 g10405(n6358, n1478, new_n10782);
nand_5 g10406(n5760, n5198, new_n10783);
nand_5 g10407(n10990, n1471, new_n10784);
xor_4  g10408(new_n10784, new_n10783, new_n10785);
not_8  g10409(new_n10785, new_n10786);
xor_4  g10410(new_n10786, new_n10782, new_n10787);
and_5  g10411(new_n10736, new_n10735, new_n10788);
nor_5  g10412(new_n10738, new_n10734, new_n10789_1);
or_5   g10413(new_n10789_1, new_n10788, new_n10790);
not_8  g10414(new_n10790, new_n10791);
xor_4  g10415(new_n10791, new_n10787, new_n10792);
xor_4  g10416(new_n10792, new_n10781, new_n10793);
not_8  g10417(new_n10793, new_n10794);
nor_5  g10418(new_n10756, new_n10751, new_n10795);
and_5  g10419(new_n10757, new_n10749, new_n10796);
nor_5  g10420(new_n10796, new_n10795, new_n10797);
not_8  g10421(new_n10797, new_n10798);
xor_4  g10422(new_n10798, new_n10794, new_n10799);
xor_4  g10423(new_n10799, new_n10772, new_n10800);
xor_4  g10424(new_n10800, new_n10770, new_n10801);
or_5   g10425(new_n10730, new_n10707, new_n10802);
not_8  g10426(new_n10802, new_n10803);
nand_5 g10427(n4805, n447, new_n10804);
not_8  g10428(new_n10804, new_n10805);
and_5  g10429(new_n10721, new_n10717, new_n10806);
and_5  g10430(new_n10722, new_n10715, new_n10807);
or_5   g10431(new_n10807, new_n10806, new_n10808);
not_8  g10432(new_n10808, new_n10809);
nand_5 g10433(n11967, n11478, new_n10810);
nand_5 g10434(n6254, n5283, new_n10811);
xor_4  g10435(new_n10811, new_n10810, new_n10812);
not_8  g10436(new_n10812, new_n10813);
xor_4  g10437(new_n10813, new_n10809, new_n10814);
nand_5 g10438(n12777, n137, new_n10815);
nand_5 g10439(n7159, n6294, new_n10816);
nand_5 g10440(n12489, n6797, new_n10817);
xor_4  g10441(new_n10817, new_n10816, new_n10818);
not_8  g10442(new_n10818, new_n10819);
xor_4  g10443(new_n10819, new_n10815, new_n10820);
and_5  g10444(new_n10711, new_n10710, new_n10821);
nor_5  g10445(new_n10713, new_n10709, new_n10822);
or_5   g10446(new_n10822, new_n10821, new_n10823);
not_8  g10447(new_n10823, new_n10824);
xor_4  g10448(new_n10824, new_n10820, new_n10825);
xor_4  g10449(new_n10825, new_n10814, new_n10826);
not_8  g10450(new_n10826, new_n10827);
nor_5  g10451(new_n10727, new_n10725, new_n10828);
nor_5  g10452(new_n10729, new_n10723, new_n10829);
nor_5  g10453(new_n10829, new_n10828, new_n10830);
not_8  g10454(new_n10830, new_n10831);
xor_4  g10455(new_n10831, new_n10827, new_n10832);
xor_4  g10456(new_n10832, new_n10805, new_n10833);
xor_4  g10457(new_n10833, new_n10803, new_n10834);
not_8  g10458(new_n10834, new_n10835);
not_8  g10459(new_n10731, new_n10836);
nor_5  g10460(new_n10760, new_n10836, new_n10837);
nor_5  g10461(new_n10764, new_n10761, new_n10838);
or_5   g10462(new_n10838, new_n10837, new_n10839);
not_8  g10463(new_n10839, new_n10840);
xor_4  g10464(new_n10840, new_n10835, new_n10841);
xor_4  g10465(new_n10841, new_n10801, new_n10842);
xor_4  g10466(new_n10767, new_n10588, new_n10843);
not_8  g10467(new_n10843, new_n10844);
nor_5  g10468(new_n10844, new_n10842, new_n10845);
or_5   g10469(new_n10845, new_n10768, new_n10846);
or_5   g10470(new_n10584, new_n10581, new_n10847);
not_8  g10471(new_n10847, new_n10848_1);
and_5  g10472(new_n10575, new_n10572, new_n10849);
or_5   g10473(new_n10574, new_n10573, new_n10850);
not_8  g10474(new_n10850, new_n10851_1);
or_5   g10475(new_n10579, new_n10577, new_n10852);
not_8  g10476(new_n10852, new_n10853);
xor_4  g10477(new_n10853, new_n10851_1, new_n10854);
or_5   g10478(new_n10854, new_n10849, new_n10855);
nor_5  g10479(new_n10566, new_n10562, new_n10856);
and_5  g10480(new_n10571, new_n10567, new_n10857);
or_5   g10481(new_n10857, new_n10856, new_n10858);
not_8  g10482(new_n10858, new_n10859);
nand_5 g10483(n9400, n8717, new_n10860);
not_8  g10484(new_n10860, new_n10861);
nand_5 g10485(n2464, n2433, new_n10862);
nand_5 g10486(n7730, n6877, new_n10863);
xor_4  g10487(new_n10863, new_n10862, new_n10864);
not_8  g10488(new_n10864, new_n10865);
xor_4  g10489(new_n10865, new_n10861, new_n10866);
xor_4  g10490(new_n10866, new_n10859, new_n10867);
or_5   g10491(new_n10564, new_n10563, new_n10868);
not_8  g10492(new_n10868, new_n10869);
nand_5 g10493(n11311, n8819, new_n10870);
not_8  g10494(new_n10870, new_n10871);
xor_4  g10495(new_n10871, new_n10869, new_n10872);
nand_5 g10496(n11728, n4203, new_n10873);
nand_5 g10497(n6429, n4187, new_n10874);
nand_5 g10498(n12753, n12709, new_n10875);
xor_4  g10499(new_n10875, new_n10874, new_n10876);
not_8  g10500(new_n10876, new_n10877);
xor_4  g10501(new_n10877, new_n10873, new_n10878);
xor_4  g10502(new_n10878, new_n10872, new_n10879);
xor_4  g10503(new_n10879, new_n10867, new_n10880);
xor_4  g10504(new_n10880, new_n10855, new_n10881);
not_8  g10505(new_n10881, new_n10882);
xor_4  g10506(new_n10882, new_n10848_1, new_n10883);
nor_5  g10507(new_n10586, new_n10561, new_n10884);
and_5  g10508(new_n10587, new_n10560, new_n10885);
nor_5  g10509(new_n10885, new_n10884, new_n10886);
xor_4  g10510(new_n10886, new_n10883, new_n10887);
or_5   g10511(new_n10831, new_n10827, new_n10888);
nand_5 g10512(n11478, n447, new_n10889);
nand_5 g10513(n11967, n5283, new_n10890);
and_5  g10514(n4805, n1353, new_n10891);
xor_4  g10515(new_n10891, new_n10890, new_n10892);
not_8  g10516(new_n10892, new_n10893);
xor_4  g10517(new_n10893, new_n10889, new_n10894);
nor_5  g10518(new_n10819, new_n10815, new_n10895);
and_5  g10519(new_n10824, new_n10820, new_n10896);
or_5   g10520(new_n10896, new_n10895, new_n10897);
not_8  g10521(new_n10897, new_n10898_1);
xor_4  g10522(new_n10898_1, new_n10894, new_n10899);
or_5   g10523(new_n10817, new_n10816, new_n10900);
not_8  g10524(new_n10900, new_n10901);
nand_5 g10525(n6254, n137, new_n10902);
not_8  g10526(new_n10902, new_n10903);
xor_4  g10527(new_n10903, new_n10901, new_n10904);
and_5  g10528(n7159, n6797, new_n10905);
nand_5 g10529(n12777, n6294, new_n10906);
nand_5 g10530(n12489, n3146, new_n10907);
xor_4  g10531(new_n10907, new_n10906, new_n10908);
xor_4  g10532(new_n10908, new_n10905, new_n10909);
xor_4  g10533(new_n10909, new_n10904, new_n10910);
xor_4  g10534(new_n10910, new_n10899, new_n10911);
not_8  g10535(new_n10911, new_n10912);
nor_5  g10536(new_n10813, new_n10809, new_n10913_1);
or_5   g10537(new_n10811, new_n10810, new_n10914);
nand_5 g10538(new_n10825, new_n10814, new_n10915);
xor_4  g10539(new_n10915, new_n10914, new_n10916);
nor_5  g10540(new_n10916, new_n10913_1, new_n10917);
xor_4  g10541(new_n10917, new_n10912, new_n10918);
not_8  g10542(new_n10918, new_n10919);
xor_4  g10543(new_n10919, new_n10888, new_n10920);
not_8  g10544(new_n10920, new_n10921);
xor_4  g10545(new_n10831, new_n10826, new_n10922);
or_5   g10546(new_n10922, new_n10804, new_n10923);
not_8  g10547(new_n10923, new_n10924);
and_5  g10548(new_n10833, new_n10803, new_n10925);
nor_5  g10549(new_n10925, new_n10924, new_n10926);
xor_4  g10550(new_n10926, new_n10921, new_n10927);
not_8  g10551(new_n10927, new_n10928_1);
or_5   g10552(new_n10798, new_n10794, new_n10929);
nor_5  g10553(new_n10786, new_n10782, new_n10930);
and_5  g10554(new_n10791, new_n10787, new_n10931);
or_5   g10555(new_n10931, new_n10930, new_n10932);
not_8  g10556(new_n10932, new_n10933);
nand_5 g10557(n6441, n3992, new_n10934);
not_8  g10558(new_n10934, new_n10935);
nand_5 g10559(n12947, n8384, new_n10936);
nand_5 g10560(n11999, n7236, new_n10937);
xor_4  g10561(new_n10937, new_n10936, new_n10938);
not_8  g10562(new_n10938, new_n10939);
xor_4  g10563(new_n10939, new_n10935, new_n10940);
xor_4  g10564(new_n10940, new_n10933, new_n10941);
or_5   g10565(new_n10784, new_n10783, new_n10942);
not_8  g10566(new_n10942, new_n10943);
nand_5 g10567(n11791, n6358, new_n10944);
not_8  g10568(new_n10944, new_n10945);
xor_4  g10569(new_n10945, new_n10943, new_n10946);
nand_5 g10570(n5760, n1471, new_n10947);
nand_5 g10571(n5198, n1478, new_n10948);
nand_5 g10572(n10990, n7646, new_n10949_1);
xor_4  g10573(new_n10949_1, new_n10948, new_n10950);
not_8  g10574(new_n10950, new_n10951);
xor_4  g10575(new_n10951, new_n10947, new_n10952);
xor_4  g10576(new_n10952, new_n10946, new_n10953);
xor_4  g10577(new_n10953, new_n10941, new_n10954);
not_8  g10578(new_n10954, new_n10955);
nor_5  g10579(new_n10780, new_n10776, new_n10956);
or_5   g10580(new_n10778, new_n10777, new_n10957);
nand_5 g10581(new_n10792, new_n10781, new_n10958);
xor_4  g10582(new_n10958, new_n10957, new_n10959);
nor_5  g10583(new_n10959, new_n10956, new_n10960);
xor_4  g10584(new_n10960, new_n10955, new_n10961);
not_8  g10585(new_n10961, new_n10962);
xor_4  g10586(new_n10962, new_n10929, new_n10963);
not_8  g10587(new_n10963, new_n10964);
and_5  g10588(new_n10799, new_n10772, new_n10965_1);
and_5  g10589(new_n10800, new_n10770, new_n10966);
nor_5  g10590(new_n10966, new_n10965_1, new_n10967);
xor_4  g10591(new_n10967, new_n10964, new_n10968);
not_8  g10592(new_n10968, new_n10969);
xor_4  g10593(new_n10969, new_n10928_1, new_n10970);
and_5  g10594(new_n10840, new_n10835, new_n10971);
xor_4  g10595(new_n10800, new_n10769, new_n10972);
and_5  g10596(new_n10841, new_n10972, new_n10973);
or_5   g10597(new_n10973, new_n10971, new_n10974);
not_8  g10598(new_n10974, new_n10975);
xor_4  g10599(new_n10975, new_n10970, new_n10976);
xor_4  g10600(new_n10976, new_n10887, new_n10977);
xor_4  g10601(new_n10977, new_n10846, new_n10978);
not_8  g10602(new_n10978, new_n10979);
nor_5  g10603(new_n10979, new_n10506, new_n10980);
xor_4  g10604(new_n10979, new_n10505, new_n10981);
xor_4  g10605(new_n10499, new_n10498, new_n10982);
not_8  g10606(new_n10982, new_n10983);
xor_4  g10607(new_n10497, new_n10495, new_n10984);
not_8  g10608(new_n10984, new_n10985);
xor_4  g10609(new_n10765, new_n10706, new_n10986);
and_5  g10610(new_n10986, new_n10985, new_n10987);
xor_4  g10611(new_n10986, new_n10984, new_n10988);
not_8  g10612(new_n10988, new_n10989);
xor_4  g10613(new_n10494, new_n10489, new_n10990_1);
xor_4  g10614(new_n10700, new_n10675, new_n10991);
nor_5  g10615(new_n10991, new_n10990_1, new_n10992);
xor_4  g10616(new_n10698, new_n10687, new_n10993);
not_8  g10617(new_n10433, new_n10994);
or_5   g10618(new_n10435, new_n10994, new_n10995);
nor_5  g10619(new_n10995, new_n10431, new_n10996);
not_8  g10620(new_n10995, new_n10997);
nor_5  g10621(new_n10997, new_n10490, new_n10998);
or_5   g10622(new_n10998, new_n10996, new_n10999);
nor_5  g10623(new_n10999, new_n10993, new_n11000);
xor_4  g10624(new_n10999, new_n10993, new_n11001);
not_8  g10625(new_n11001, new_n11002);
xor_4  g10626(new_n10693, new_n10679, new_n11003);
nand_5 g10627(new_n11003, new_n10994, new_n11004);
xnor_4 g10628(new_n10492, new_n10491, new_n11005);
and_5  g10629(new_n11005, new_n11004, new_n11006);
xor_4  g10630(new_n10696, new_n10695_1, new_n11007);
xor_4  g10631(new_n11005, new_n11004, new_n11008);
not_8  g10632(new_n11008, new_n11009);
nor_5  g10633(new_n11009, new_n11007, new_n11010);
or_5   g10634(new_n11010, new_n11006, new_n11011);
not_8  g10635(new_n11011, new_n11012);
nor_5  g10636(new_n11012, new_n11002, new_n11013);
or_5   g10637(new_n11013, new_n11000, new_n11014);
not_8  g10638(new_n10990_1, new_n11015);
xor_4  g10639(new_n10991, new_n11015, new_n11016);
not_8  g10640(new_n11016, new_n11017);
and_5  g10641(new_n11017, new_n11014, new_n11018);
or_5   g10642(new_n11018, new_n10992, new_n11019);
and_5  g10643(new_n11019, new_n10989, new_n11020);
nor_5  g10644(new_n11020, new_n10987, new_n11021);
nor_5  g10645(new_n11021, new_n10983, new_n11022);
xor_4  g10646(new_n10844, new_n10842, new_n11023_1);
xor_4  g10647(new_n11021, new_n10982, new_n11024);
not_8  g10648(new_n11024, new_n11025);
and_5  g10649(new_n11025, new_n11023_1, new_n11026);
or_5   g10650(new_n11026, new_n11022, new_n11027);
not_8  g10651(new_n11027, new_n11028);
nor_5  g10652(new_n11028, new_n10981, new_n11029);
nor_5  g10653(new_n11029, new_n10980, new_n11030);
and_5  g10654(new_n10976, new_n10887, new_n11031);
nor_5  g10655(new_n10976, new_n10887, new_n11032);
nor_5  g10656(new_n11032, new_n10846, new_n11033);
nor_5  g10657(new_n11033, new_n11031, new_n11034);
not_8  g10658(new_n10483, new_n11035);
nor_5  g10659(new_n11035, new_n10448, new_n11036);
nor_5  g10660(new_n10503, new_n11036, new_n11037);
nor_5  g10661(new_n10915, new_n10914, new_n11038);
nor_5  g10662(new_n10917, new_n10912, new_n11039);
or_5   g10663(new_n11039, new_n11038, new_n11040);
and_5  g10664(new_n10937, new_n10936, new_n11041);
nor_5  g10665(new_n10939, new_n10935, new_n11042);
nor_5  g10666(new_n11042, new_n11041, new_n11043);
and_5  g10667(n4805, n4436, new_n11044);
nand_5 g10668(n8384, n6441, new_n11045);
and_5  g10669(n11791, n5198, new_n11046);
xor_4  g10670(new_n11046, new_n11045, new_n11047);
xor_4  g10671(new_n11047, new_n11044, new_n11048);
xor_4  g10672(new_n11048, new_n11043, new_n11049);
nand_5 g10673(n7159, n3146, new_n11050);
and_5  g10674(n11967, n137, new_n11051);
xor_4  g10675(new_n11051, new_n11050, new_n11052);
and_5  g10676(n6294, n6254, new_n11053);
and_5  g10677(n12947, n6358, new_n11054);
xor_4  g10678(new_n11054, new_n11053, new_n11055);
and_5  g10679(n11407, n6826, new_n11056);
and_5  g10680(n7862, n6604, new_n11057);
xor_4  g10681(new_n11057, new_n11056, new_n11058);
xor_4  g10682(new_n11058, new_n11055, new_n11059);
xor_4  g10683(new_n11059, new_n11052, new_n11060);
xor_4  g10684(new_n11060, new_n11049, new_n11061);
and_5  g10685(n6429, n4203, new_n11062);
and_5  g10686(new_n10903, new_n10901, new_n11063);
and_5  g10687(new_n10909, new_n10904, new_n11064);
nor_5  g10688(new_n11064, new_n11063, new_n11065);
xor_4  g10689(new_n11065, new_n11062, new_n11066);
xor_4  g10690(new_n11066, new_n11061, new_n11067);
nand_5 g10691(new_n10898_1, new_n10894, new_n11068);
not_8  g10692(new_n10910, new_n11069);
nand_5 g10693(new_n11069, new_n10899, new_n11070);
nand_5 g10694(new_n11070, new_n11068, new_n11071);
nand_5 g10695(new_n10940, new_n10933, new_n11072);
not_8  g10696(new_n10953, new_n11073);
nand_5 g10697(new_n11073, new_n10941, new_n11074);
nand_5 g10698(new_n11074, new_n11072, new_n11075);
and_5  g10699(n11478, n1353, new_n11076);
and_5  g10700(new_n10893, new_n10889, new_n11077);
or_5   g10701(new_n11077, new_n10890, new_n11078);
not_8  g10702(new_n11078, new_n11079);
and_5  g10703(new_n11079, new_n11076, new_n11080);
and_5  g10704(new_n11076, new_n10804, new_n11081);
nor_5  g10705(new_n11081, new_n11079, new_n11082);
or_5   g10706(new_n11082, new_n11080, new_n11083);
nor_5  g10707(new_n10907, new_n10906, new_n11084);
nand_5 g10708(n7159, n6797, new_n11085);
and_5  g10709(new_n10907, new_n10906, new_n11086);
nor_5  g10710(new_n11086, new_n11085, new_n11087);
nor_5  g10711(new_n11087, new_n11084, new_n11088);
xor_4  g10712(new_n11088, new_n11083, new_n11089);
xor_4  g10713(new_n11089, new_n11075, new_n11090);
xor_4  g10714(new_n11090, new_n11071, new_n11091);
xor_4  g10715(new_n11091, new_n11067, new_n11092);
not_8  g10716(new_n10451_1, new_n11093);
nand_5 g10717(new_n10453, new_n11093, new_n11094);
nand_5 g10718(new_n10482, new_n10455, new_n11095);
and_5  g10719(new_n11095, new_n11094, new_n11096);
and_5  g10720(n12777, n6797, new_n11097);
xor_4  g10721(new_n11097, new_n11096, new_n11098);
xor_4  g10722(new_n11098, new_n11092, new_n11099);
xor_4  g10723(new_n11099, new_n11040, new_n11100);
xor_4  g10724(new_n11100, new_n11037, new_n11101);
xor_4  g10725(new_n11101, new_n11034, new_n11102);
nor_5  g10726(new_n10882, new_n10847, new_n11103);
nor_5  g10727(new_n10886, new_n10883, new_n11104);
or_5   g10728(new_n11104, new_n11103, new_n11105);
nor_5  g10729(new_n10919, new_n10888, new_n11106);
nor_5  g10730(new_n10926, new_n10921, new_n11107);
nor_5  g10731(new_n11107, new_n11106, new_n11108);
xor_4  g10732(new_n11108, new_n11105, new_n11109);
nor_5  g10733(new_n10962, new_n10929, new_n11110);
nor_5  g10734(new_n10967, new_n10964, new_n11111);
or_5   g10735(new_n11111, new_n11110, new_n11112);
nor_5  g10736(new_n10866, new_n10859, new_n11113);
and_5  g10737(new_n10879, new_n10867, new_n11114);
or_5   g10738(new_n11114, new_n11113, new_n11115);
and_5  g10739(new_n10863, new_n10862, new_n11116);
nor_5  g10740(new_n10865, new_n10861, new_n11117);
nor_5  g10741(new_n11117, new_n11116, new_n11118);
nand_5 g10742(n5283, n447, new_n11119);
and_5  g10743(n11999, n3992, new_n11120);
xor_4  g10744(new_n11120, new_n11119, new_n11121);
xor_4  g10745(new_n11121, new_n11118, new_n11122);
xor_4  g10746(new_n11122, new_n11115, new_n11123);
nand_5 g10747(n7646, n5760, new_n11124);
and_5  g10748(n10990, n4722, new_n11125);
xor_4  g10749(new_n11125, new_n11124, new_n11126);
xor_4  g10750(new_n11126, new_n11123, new_n11127);
xor_4  g10751(new_n11127, new_n11112, new_n11128);
xor_4  g10752(new_n11128, new_n11109, new_n11129);
nor_5  g10753(new_n10969, new_n10928_1, new_n11130);
and_5  g10754(new_n10975, new_n10970, new_n11131);
nor_5  g10755(new_n11131, new_n11130, new_n11132);
and_5  g10756(new_n10853, new_n10851_1, new_n11133);
and_5  g10757(new_n10880, new_n10855, new_n11134);
or_5   g10758(new_n11134, new_n11133, new_n11135);
nor_5  g10759(new_n10480, new_n10472, new_n11136);
and_5  g10760(new_n10481, new_n10467, new_n11137);
nor_5  g10761(new_n11137, new_n11136, new_n11138);
and_5  g10762(new_n10875, new_n10874, new_n11139);
not_8  g10763(new_n10873, new_n11140);
nor_5  g10764(new_n10877, new_n11140, new_n11141);
or_5   g10765(new_n11141, new_n11139, new_n11142);
nand_5 g10766(n12000, n3172, new_n11143);
nand_5 g10767(n9725, n1333, new_n11144);
and_5  g10768(n12709, n10174, new_n11145);
xor_4  g10769(new_n11145, new_n11144, new_n11146);
xor_4  g10770(new_n11146, new_n11143, new_n11147);
xor_4  g10771(new_n11147, new_n11142, new_n11148);
and_5  g10772(new_n10871, new_n10869, new_n11149);
and_5  g10773(new_n10878, new_n10872, new_n11150);
or_5   g10774(new_n11150, new_n11149, new_n11151);
and_5  g10775(new_n10949_1, new_n10948, new_n11152);
not_8  g10776(new_n10947, new_n11153_1);
nor_5  g10777(new_n10951, new_n11153_1, new_n11154);
nor_5  g10778(new_n11154, new_n11152, new_n11155);
nand_5 g10779(n6877, n1198, new_n11156);
and_5  g10780(n12753, n11728, new_n11157);
xor_4  g10781(new_n11157, new_n11156, new_n11158);
xor_4  g10782(new_n11158, new_n11155, new_n11159);
xor_4  g10783(new_n11159, new_n11151, new_n11160);
xor_4  g10784(new_n11160, new_n11148, new_n11161);
xor_4  g10785(new_n11161, new_n11138, new_n11162);
nand_5 g10786(n12489, n4938, new_n11163);
and_5  g10787(new_n10476_1, new_n10475, new_n11164);
nor_5  g10788(new_n10478, new_n10474, new_n11165);
nor_5  g10789(new_n11165, new_n11164, new_n11166);
and_5  g10790(n11757, n5320, new_n11167);
and_5  g10791(n9080, n5212, new_n11168);
xor_4  g10792(new_n11168, new_n11167, new_n11169);
nand_5 g10793(n11877, n11821, new_n11170);
and_5  g10794(n5240, n4370, new_n11171);
xor_4  g10795(new_n11171, new_n11170, new_n11172);
xor_4  g10796(new_n11172, new_n11169, new_n11173);
xor_4  g10797(new_n11173, new_n11166, new_n11174);
nand_5 g10798(n9400, n7730, new_n11175);
and_5  g10799(n11311, n2433, new_n11176);
xor_4  g10800(new_n11176, new_n11175, new_n11177);
xor_4  g10801(new_n11177, new_n11174, new_n11178);
and_5  g10802(new_n10463, new_n10462, new_n11179);
nor_5  g10803(new_n10465, new_n10461, new_n11180);
nor_5  g10804(new_n11180, new_n11179, new_n11181);
nor_5  g10805(new_n10458, new_n10457, new_n11182);
and_5  g10806(new_n10466, new_n10459, new_n11183);
nor_5  g10807(new_n11183, new_n11182, new_n11184);
xor_4  g10808(new_n11184, new_n11181, new_n11185);
xor_4  g10809(new_n11185, new_n11178, new_n11186);
xor_4  g10810(new_n11186, new_n11163, new_n11187);
xor_4  g10811(new_n11187, new_n11162, new_n11188);
xor_4  g10812(new_n11188, new_n11135, new_n11189);
nor_5  g10813(new_n10958, new_n10957, new_n11190);
nor_5  g10814(new_n10960, new_n10955, new_n11191);
or_5   g10815(new_n11191, new_n11190, new_n11192);
nand_5 g10816(n8819, n4187, new_n11193);
and_5  g10817(n1478, n1471, new_n11194);
xor_4  g10818(new_n11194, new_n11193, new_n11195);
nand_5 g10819(n8717, n2464, new_n11196);
and_5  g10820(n10022, n7236, new_n11197);
xor_4  g10821(new_n11197, new_n11196, new_n11198);
xor_4  g10822(new_n11198, new_n11195, new_n11199);
and_5  g10823(new_n10945, new_n10943, new_n11200);
and_5  g10824(new_n10952, new_n10946, new_n11201);
nor_5  g10825(new_n11201, new_n11200, new_n11202);
xor_4  g10826(new_n11202, new_n11199, new_n11203);
xor_4  g10827(new_n11203, new_n11192, new_n11204);
xor_4  g10828(new_n11204, new_n11189, new_n11205);
xor_4  g10829(new_n11205, new_n11132, new_n11206);
xor_4  g10830(new_n11206, new_n11129, new_n11207);
xor_4  g10831(new_n11207, new_n11102, new_n11208);
xor_4  g10832(new_n11208, new_n11030, n4378);
xor_4  g10833(new_n3806, new_n3805, n4397);
xor_4  g10834(new_n4095, new_n4086_1, n4553);
xor_4  g10835(new_n857, new_n856, n4686);
not_8  g10836(new_n9260, new_n11213);
xor_4  g10837(new_n11213, new_n9238, n4689);
xor_4  g10838(new_n4856, new_n4854, n4733);
not_8  g10839(new_n2044, new_n11216_1);
xor_4  g10840(new_n11216_1, new_n2036, n4757);
nor_5  g10841(new_n4845, new_n4831, new_n11218);
xor_4  g10842(new_n4849, new_n11218, n4971);
or_5   g10843(new_n6472, new_n6470, new_n11220);
xor_4  g10844(new_n6476, new_n11220, n5030);
xor_4  g10845(new_n2870, new_n2839, n5034);
not_8  g10846(new_n2863, new_n11223);
xor_4  g10847(new_n11223, new_n2853, n5094);
and_5  g10848(new_n10269, new_n10265, new_n11225);
and_5  g10849(new_n10276, new_n10270, new_n11226);
or_5   g10850(new_n11226, new_n11225, new_n11227);
not_8  g10851(new_n11227, new_n11228);
nand_5 g10852(n5320, n2564, new_n11229);
nand_5 g10853(n4370, n4189, new_n11230);
xor_4  g10854(new_n11230, new_n11229, new_n11231);
not_8  g10855(new_n11231, new_n11232);
xor_4  g10856(new_n11232, new_n11228, new_n11233);
nand_5 g10857(n11877, n6770, new_n11234);
not_8  g10858(new_n11234, new_n11235);
and_5  g10859(new_n10273, new_n10272, new_n11236);
not_8  g10860(new_n10271, new_n11237);
nor_5  g10861(new_n10275, new_n11237, new_n11238);
or_5   g10862(new_n11238, new_n11236, new_n11239);
not_8  g10863(new_n11239, new_n11240);
xor_4  g10864(new_n11240, new_n11235, new_n11241);
nand_5 g10865(n9920, n5212, new_n11242);
nand_5 g10866(n11407, n3627, new_n11243);
xor_4  g10867(new_n11243, new_n11242, new_n11244);
xor_4  g10868(new_n11244, new_n11241, new_n11245);
xor_4  g10869(new_n11245, new_n11233, new_n11246);
not_8  g10870(new_n11246, new_n11247);
nor_5  g10871(new_n10261, new_n10258, new_n11248);
nor_5  g10872(new_n10278_1, new_n10263, new_n11249);
nor_5  g10873(new_n11249, new_n11248, new_n11250);
or_5   g10874(new_n11250, new_n11247, new_n11251);
not_8  g10875(new_n11251, new_n11252);
and_5  g10876(new_n11240, new_n11235, new_n11253);
and_5  g10877(new_n11244, new_n11241, new_n11254);
or_5   g10878(new_n11254, new_n11253, new_n11255);
not_8  g10879(new_n11255, new_n11256);
nand_5 g10880(n12000, n2564, new_n11257_1);
nand_5 g10881(n5320, n4189, new_n11258);
nand_5 g10882(n9725, n6687, new_n11259);
xor_4  g10883(new_n11259, new_n11258, new_n11260);
xor_4  g10884(new_n11260, new_n11257_1, new_n11261);
xor_4  g10885(new_n11261, new_n11256, new_n11262);
or_5   g10886(new_n11243, new_n11242, new_n11263);
not_8  g10887(new_n11263, new_n11264);
nand_5 g10888(n6770, n4370, new_n11265);
not_8  g10889(new_n11265, new_n11266);
xor_4  g10890(new_n11266, new_n11264, new_n11267);
and_5  g10891(n5212, n3627, new_n11268);
nand_5 g10892(n11877, n9920, new_n11269);
nand_5 g10893(n11407, n4516, new_n11270);
xor_4  g10894(new_n11270, new_n11269, new_n11271);
xor_4  g10895(new_n11271, new_n11268, new_n11272);
xor_4  g10896(new_n11272, new_n11267, new_n11273);
xor_4  g10897(new_n11273, new_n11262, new_n11274);
not_8  g10898(new_n11274, new_n11275);
nor_5  g10899(new_n11232, new_n11228, new_n11276);
or_5   g10900(new_n11230, new_n11229, new_n11277);
nand_5 g10901(new_n11245, new_n11233, new_n11278);
xor_4  g10902(new_n11278, new_n11277, new_n11279);
nor_5  g10903(new_n11279, new_n11276, new_n11280);
xor_4  g10904(new_n11280, new_n11275, new_n11281);
not_8  g10905(new_n11281, new_n11282);
xor_4  g10906(new_n11282, new_n11252, new_n11283);
nand_5 g10907(n12000, n6687, new_n11284);
xor_4  g10908(new_n11250, new_n11247, new_n11285);
not_8  g10909(new_n11285, new_n11286);
nor_5  g10910(new_n11286, new_n11284, new_n11287);
and_5  g10911(new_n10279, new_n10257, new_n11288);
xor_4  g10912(new_n11286, new_n11284, new_n11289);
and_5  g10913(new_n11289, new_n11288, new_n11290);
nor_5  g10914(new_n11290, new_n11287, new_n11291);
xor_4  g10915(new_n11291, new_n11283, new_n11292);
nand_5 g10916(n8717, n8336, new_n11293);
nand_5 g10917(n6429, n2226, new_n11294);
nand_5 g10918(n11728, n1094, new_n11295);
nand_5 g10919(n12709, n10678, new_n11296_1);
xor_4  g10920(new_n11296_1, new_n11295, new_n11297);
not_8  g10921(new_n11297, new_n11298);
xor_4  g10922(new_n11298, new_n11294, new_n11299);
and_5  g10923(new_n10298, new_n1297, new_n11300);
nor_5  g10924(new_n10298, new_n1297, new_n11301);
nor_5  g10925(new_n11301, new_n10297, new_n11302);
or_5   g10926(new_n11302, new_n11300, new_n11303);
not_8  g10927(new_n11303, new_n11304);
xor_4  g10928(new_n11304, new_n11299, new_n11305);
nand_5 g10929(n10928, n2433, new_n11306);
nand_5 g10930(n8819, n6986, new_n11307);
xor_4  g10931(new_n11307, new_n11306, new_n11308);
xor_4  g10932(new_n11308, new_n11305, new_n11309);
not_8  g10933(new_n11309, new_n11310);
nor_5  g10934(new_n10301, new_n10295, new_n11311_1);
nor_5  g10935(new_n11311_1, new_n10293, new_n11312);
xor_4  g10936(new_n11312, new_n11310, new_n11313);
not_8  g10937(new_n11313, new_n11314);
and_5  g10938(new_n10302, new_n10285, new_n11315);
nor_5  g10939(new_n10307, new_n10304, new_n11316);
nor_5  g10940(new_n11316, new_n11315, new_n11317);
xor_4  g10941(new_n11317, new_n11314, new_n11318);
not_8  g10942(new_n11318, new_n11319);
nor_5  g10943(new_n11319, new_n11293, new_n11320);
nand_5 g10944(new_n10308, new_n10283, new_n11321);
not_8  g10945(new_n11321, new_n11322);
xor_4  g10946(new_n11319, new_n11293, new_n11323);
and_5  g10947(new_n11323, new_n11322, new_n11324);
or_5   g10948(new_n11324, new_n11320, new_n11325);
not_8  g10949(new_n11325, new_n11326_1);
or_5   g10950(new_n11317, new_n11314, new_n11327);
not_8  g10951(new_n11327, new_n11328);
nor_5  g10952(new_n11298, new_n11294, new_n11329);
and_5  g10953(new_n11304, new_n11299, new_n11330);
or_5   g10954(new_n11330, new_n11329, new_n11331);
nand_5 g10955(n10928, n8717, new_n11332);
not_8  g10956(new_n11332, new_n11333);
nand_5 g10957(n6986, n2433, new_n11334);
nand_5 g10958(n8336, n7730, new_n11335);
xor_4  g10959(new_n11335, new_n11334, new_n11336);
not_8  g10960(new_n11336, new_n11337);
xor_4  g10961(new_n11337, new_n11333, new_n11338);
not_8  g10962(new_n11338, new_n11339);
xor_4  g10963(new_n11339, new_n11331, new_n11340);
or_5   g10964(new_n11296_1, new_n11295, new_n11341);
not_8  g10965(new_n11341, new_n11342);
nand_5 g10966(n8819, n2226, new_n11343);
not_8  g10967(new_n11343, new_n11344);
xor_4  g10968(new_n11344, new_n11342, new_n11345);
nand_5 g10969(n11728, n10678, new_n11346);
nand_5 g10970(n6429, n1094, new_n11347);
nand_5 g10971(n12709, n7320, new_n11348);
xor_4  g10972(new_n11348, new_n11347, new_n11349);
not_8  g10973(new_n11349, new_n11350);
xor_4  g10974(new_n11350, new_n11346, new_n11351);
xor_4  g10975(new_n11351, new_n11345, new_n11352);
xor_4  g10976(new_n11352, new_n11340, new_n11353);
not_8  g10977(new_n11353, new_n11354);
nand_5 g10978(new_n11308, new_n11305, new_n11355);
or_5   g10979(new_n11307, new_n11306, new_n11356);
or_5   g10980(new_n11312, new_n11310, new_n11357);
not_8  g10981(new_n11357, new_n11358);
xor_4  g10982(new_n11358, new_n11356, new_n11359);
and_5  g10983(new_n11359, new_n11355, new_n11360);
xor_4  g10984(new_n11360, new_n11354, new_n11361);
xnor_4 g10985(new_n11361, new_n11328, new_n11362);
xor_4  g10986(new_n11362, new_n11326_1, new_n11363);
not_8  g10987(new_n11363, new_n11364);
xor_4  g10988(new_n11323, new_n11322, new_n11365);
not_8  g10989(new_n11365, new_n11366);
nor_5  g10990(new_n10314, new_n10310, new_n11367);
not_8  g10991(new_n10374, new_n11368);
nor_5  g10992(new_n11368, new_n10316, new_n11369);
or_5   g10993(new_n11369, new_n11367, new_n11370);
not_8  g10994(new_n11370, new_n11371);
and_5  g10995(new_n11371, new_n11366, new_n11372);
or_5   g10996(new_n10367, new_n10344, new_n11373);
not_8  g10997(new_n11373, new_n11374);
nand_5 g10998(n11222, n6441, new_n11375);
and_5  g10999(new_n10351, new_n10348, new_n11376);
nor_5  g11000(new_n10360, new_n10353, new_n11377);
or_5   g11001(new_n11377, new_n11376, new_n11378);
nand_5 g11002(n12947, n11153, new_n11379);
nand_5 g11003(n11791, n5314, new_n11380);
xor_4  g11004(new_n11380, new_n11379, new_n11381);
xor_4  g11005(new_n11381, new_n11378, new_n11382);
not_8  g11006(new_n11382, new_n11383);
nand_5 g11007(n1478, n996, new_n11384);
nand_5 g11008(n10990, n5319, new_n11385);
nand_5 g11009(n5767, n5760, new_n11386);
xor_4  g11010(new_n11386, new_n11385, new_n11387);
not_8  g11011(new_n11387, new_n11388);
xor_4  g11012(new_n11388, new_n11384, new_n11389);
and_5  g11013(new_n10357, new_n10356, new_n11390);
nor_5  g11014(new_n10357, new_n10356, new_n11391);
nor_5  g11015(new_n11391, new_n10355, new_n11392);
or_5   g11016(new_n11392, new_n11390, new_n11393);
not_8  g11017(new_n11393, new_n11394);
xor_4  g11018(new_n11394, new_n11389, new_n11395);
not_8  g11019(new_n11395, new_n11396);
xor_4  g11020(new_n11396, new_n11383, new_n11397);
and_5  g11021(new_n10361, new_n10346, new_n11398);
and_5  g11022(new_n10365, new_n10362, new_n11399);
or_5   g11023(new_n11399, new_n11398, new_n11400);
xor_4  g11024(new_n11400, new_n11397, new_n11401);
not_8  g11025(new_n11401, new_n11402);
xor_4  g11026(new_n11402, new_n11375, new_n11403);
xor_4  g11027(new_n11403, new_n11374, new_n11404);
not_8  g11028(new_n11404, new_n11405);
or_5   g11029(new_n10342, new_n10317, new_n11406);
not_8  g11030(new_n11406, new_n11407_1);
nand_5 g11031(n12069, n447, new_n11408);
not_8  g11032(new_n11408, new_n11409);
nand_5 g11033(n12777, n7160, new_n11410);
nand_5 g11034(n7159, n4828, new_n11411);
nand_5 g11035(n12489, n2515, new_n11412);
xor_4  g11036(new_n11412, new_n11411, new_n11413);
not_8  g11037(new_n11413, new_n11414);
xor_4  g11038(new_n11414, new_n11410, new_n11415);
and_5  g11039(new_n10331, new_n10330, new_n11416);
nor_5  g11040(new_n10331, new_n10330, new_n11417);
nor_5  g11041(new_n11417, new_n10329, new_n11418);
or_5   g11042(new_n11418, new_n11416, new_n11419);
not_8  g11043(new_n11419, new_n11420);
xor_4  g11044(new_n11420, new_n11415, new_n11421);
nand_5 g11045(n12391, n11967, new_n11422);
nand_5 g11046(n7891, n6254, new_n11423_1);
xor_4  g11047(new_n11423_1, new_n11422, new_n11424);
xor_4  g11048(new_n11424, new_n11421, new_n11425);
not_8  g11049(new_n11425, new_n11426);
and_5  g11050(new_n10325, new_n10321, new_n11427);
nor_5  g11051(new_n10334, new_n10327_1, new_n11428);
or_5   g11052(new_n11428, new_n11427, new_n11429);
xor_4  g11053(new_n11429, new_n11426, new_n11430);
and_5  g11054(new_n10335, new_n10319, new_n11431);
and_5  g11055(new_n10340, new_n10336, new_n11432);
nor_5  g11056(new_n11432, new_n11431, new_n11433);
xor_4  g11057(new_n11433, new_n11430, new_n11434);
xor_4  g11058(new_n11434, new_n11409, new_n11435);
not_8  g11059(new_n11435, new_n11436);
and_5  g11060(new_n11436, new_n11407_1, new_n11437);
nor_5  g11061(new_n11436, new_n11407_1, new_n11438);
or_5   g11062(new_n11438, new_n11437, new_n11439);
not_8  g11063(new_n11439, new_n11440);
and_5  g11064(new_n10372, new_n10368, new_n11441);
and_5  g11065(new_n10373, new_n10343, new_n11442);
nor_5  g11066(new_n11442, new_n11441, new_n11443);
xor_4  g11067(new_n11443, new_n11440, new_n11444);
not_8  g11068(new_n11444, new_n11445);
xor_4  g11069(new_n11445, new_n11405, new_n11446);
xor_4  g11070(new_n11371, new_n11365, new_n11447);
nor_5  g11071(new_n11447, new_n11446, new_n11448);
nor_5  g11072(new_n11448, new_n11372, new_n11449);
not_8  g11073(new_n11449, new_n11450);
xor_4  g11074(new_n11450, new_n11364, new_n11451);
nand_5 g11075(new_n11400, new_n11397, new_n11452);
nor_5  g11076(new_n11388, new_n11384, new_n11453);
and_5  g11077(new_n11394, new_n11389, new_n11454);
or_5   g11078(new_n11454, new_n11453, new_n11455);
nand_5 g11079(n11153, n6441, new_n11456);
not_8  g11080(new_n11456, new_n11457);
nand_5 g11081(n12947, n5314, new_n11458);
nand_5 g11082(n11999, n11222, new_n11459);
xor_4  g11083(new_n11459, new_n11458, new_n11460);
not_8  g11084(new_n11460, new_n11461);
xor_4  g11085(new_n11461, new_n11457, new_n11462);
not_8  g11086(new_n11462, new_n11463);
xor_4  g11087(new_n11463, new_n11455, new_n11464);
or_5   g11088(new_n11386, new_n11385, new_n11465);
not_8  g11089(new_n11465, new_n11466);
nand_5 g11090(n11791, n996, new_n11467);
not_8  g11091(new_n11467, new_n11468);
xor_4  g11092(new_n11468, new_n11466, new_n11469);
nand_5 g11093(n5760, n5319, new_n11470);
nand_5 g11094(n5767, n1478, new_n11471);
nand_5 g11095(n10990, n9457, new_n11472);
xor_4  g11096(new_n11472, new_n11471, new_n11473);
not_8  g11097(new_n11473, new_n11474);
xor_4  g11098(new_n11474, new_n11470, new_n11475);
xor_4  g11099(new_n11475, new_n11469, new_n11476);
xor_4  g11100(new_n11476, new_n11464, new_n11477);
not_8  g11101(new_n11477, new_n11478_1);
and_5  g11102(new_n11381, new_n11378, new_n11479);
or_5   g11103(new_n11380, new_n11379, new_n11480);
or_5   g11104(new_n11396, new_n11383, new_n11481);
xor_4  g11105(new_n11481, new_n11480, new_n11482);
nor_5  g11106(new_n11482, new_n11479, new_n11483);
xor_4  g11107(new_n11483, new_n11478_1, new_n11484);
not_8  g11108(new_n11484, new_n11485);
xor_4  g11109(new_n11485, new_n11452, new_n11486);
nor_5  g11110(new_n11402, new_n11375, new_n11487);
and_5  g11111(new_n11403, new_n11374, new_n11488);
or_5   g11112(new_n11488, new_n11487, new_n11489);
xor_4  g11113(new_n11489, new_n11486, new_n11490);
not_8  g11114(new_n11490, new_n11491);
or_5   g11115(new_n11433, new_n11430, new_n11492);
not_8  g11116(new_n11492, new_n11493);
nor_5  g11117(new_n11414, new_n11410, new_n11494);
and_5  g11118(new_n11420, new_n11415, new_n11495);
or_5   g11119(new_n11495, new_n11494, new_n11496);
nand_5 g11120(n12391, n447, new_n11497);
nand_5 g11121(n11967, n7891, new_n11498);
nand_5 g11122(n12069, n1353, new_n11499);
xor_4  g11123(new_n11499, new_n11498, new_n11500);
xor_4  g11124(new_n11500, new_n11497, new_n11501);
not_8  g11125(new_n11501, new_n11502);
xor_4  g11126(new_n11502, new_n11496, new_n11503);
or_5   g11127(new_n11412, new_n11411, new_n11504);
not_8  g11128(new_n11504, new_n11505);
nand_5 g11129(n7160, n6254, new_n11506);
not_8  g11130(new_n11506, new_n11507);
xor_4  g11131(new_n11507, new_n11505, new_n11508);
and_5  g11132(n7159, n2515, new_n11509);
nand_5 g11133(n12777, n4828, new_n11510);
nand_5 g11134(n12489, n1199, new_n11511);
xor_4  g11135(new_n11511, new_n11510, new_n11512);
xor_4  g11136(new_n11512, new_n11509, new_n11513);
xor_4  g11137(new_n11513, new_n11508, new_n11514);
xor_4  g11138(new_n11514, new_n11503, new_n11515);
not_8  g11139(new_n11515, new_n11516);
and_5  g11140(new_n11424, new_n11421, new_n11517);
or_5   g11141(new_n11423_1, new_n11422, new_n11518);
not_8  g11142(new_n11518, new_n11519);
nand_5 g11143(new_n11429, new_n11425, new_n11520);
not_8  g11144(new_n11520, new_n11521);
xor_4  g11145(new_n11521, new_n11519, new_n11522);
nor_5  g11146(new_n11522, new_n11517, new_n11523);
xor_4  g11147(new_n11523, new_n11516, new_n11524);
not_8  g11148(new_n11524, new_n11525);
xor_4  g11149(new_n11525, new_n11493, new_n11526);
nor_5  g11150(new_n11434, new_n11409, new_n11527);
or_5   g11151(new_n11438, new_n11527, new_n11528);
xor_4  g11152(new_n11528, new_n11526, new_n11529);
not_8  g11153(new_n11529, new_n11530);
xor_4  g11154(new_n11530, new_n11491, new_n11531);
not_8  g11155(new_n11531, new_n11532);
nor_5  g11156(new_n11443, new_n11440, new_n11533);
nor_5  g11157(new_n11445, new_n11405, new_n11534);
nor_5  g11158(new_n11534, new_n11533, new_n11535);
xor_4  g11159(new_n11535, new_n11532, new_n11536_1);
xor_4  g11160(new_n11536_1, new_n11451, new_n11537);
xor_4  g11161(new_n11537, new_n11292, new_n11538);
xor_4  g11162(new_n11289, new_n11288, new_n11539);
not_8  g11163(new_n11539, new_n11540);
and_5  g11164(new_n10375, new_n10280, new_n11541);
nor_5  g11165(new_n10380, new_n10376, new_n11542);
or_5   g11166(new_n11542, new_n11541, new_n11543);
not_8  g11167(new_n11543, new_n11544);
and_5  g11168(new_n11544, new_n11540, new_n11545);
xor_4  g11169(new_n11544, new_n11540, new_n11546);
xnor_4 g11170(new_n11447, new_n11446, new_n11547);
not_8  g11171(new_n11547, new_n11548);
and_5  g11172(new_n11548, new_n11546, new_n11549);
or_5   g11173(new_n11549, new_n11545, new_n11550);
not_8  g11174(new_n11550, new_n11551);
xor_4  g11175(new_n11551, new_n11538, n5132);
xor_4  g11176(new_n11003, new_n10994, n5191);
nor_5  g11177(new_n3551, new_n3171, new_n11554);
and_5  g11178(new_n3551, new_n3171, new_n11555);
nor_5  g11179(new_n3698, new_n11555, new_n11556);
or_5   g11180(new_n11556, new_n11554, new_n11557);
nor_5  g11181(new_n3689, new_n3596, new_n11558);
or_5   g11182(new_n3696, new_n11558, new_n11559);
nor_5  g11183(new_n3150, new_n3121, new_n11560);
nor_5  g11184(new_n3170, new_n3152, new_n11561);
or_5   g11185(new_n11561, new_n11560, new_n11562);
nor_5  g11186(new_n3146_1, new_n3145, new_n11563);
nor_5  g11187(new_n3148, new_n3143, new_n11564);
or_5   g11188(new_n11564, new_n11563, new_n11565);
and_5  g11189(n11478, n10965, new_n11566);
and_5  g11190(new_n3570, new_n3568, new_n11567);
and_5  g11191(new_n3577, new_n3571, new_n11568);
or_5   g11192(new_n11568, new_n11567, new_n11569);
and_5  g11193(n8433, n4722, new_n11570);
nand_5 g11194(n8065, n2464, new_n11571);
and_5  g11195(n7646, n405, new_n11572);
xor_4  g11196(new_n11572, new_n11571, new_n11573);
xor_4  g11197(new_n11573, new_n11570, new_n11574);
xor_4  g11198(new_n11574, new_n11569, new_n11575);
xor_4  g11199(new_n11575, new_n11566, new_n11576);
xor_4  g11200(new_n11576, new_n11565, new_n11577);
nand_5 g11201(new_n3652, new_n3648, new_n11578);
not_8  g11202(new_n3664, new_n11579);
nand_5 g11203(new_n11579, new_n3653, new_n11580);
nand_5 g11204(new_n11580, new_n11578, new_n11581);
and_5  g11205(new_n3614, new_n3612, new_n11582);
and_5  g11206(new_n3620, new_n3615, new_n11583);
nor_5  g11207(new_n11583, new_n11582, new_n11584);
and_5  g11208(new_n3657, new_n3655, new_n11585);
and_5  g11209(new_n3663, new_n3658, new_n11586);
nor_5  g11210(new_n11586, new_n11585, new_n11587);
xor_4  g11211(new_n11587, new_n11584, new_n11588);
nand_5 g11212(n8384, n6359, new_n11589);
and_5  g11213(n7546, n4805, new_n11590);
xor_4  g11214(new_n11590, new_n11589, new_n11591);
and_5  g11215(n12925, n4938, new_n11592);
and_5  g11216(n11536, n7862, new_n11593);
xor_4  g11217(new_n11593, new_n11592, new_n11594);
nor_5  g11218(new_n3661_1, new_n3660, new_n11595);
nand_5 g11219(n1471, n405, new_n11596);
and_5  g11220(new_n3661_1, new_n3660, new_n11597);
nor_5  g11221(new_n11597, new_n11596, new_n11598);
nor_5  g11222(new_n11598, new_n11595, new_n11599);
xor_4  g11223(new_n11599, new_n11594, new_n11600);
xor_4  g11224(new_n11600, new_n11591, new_n11601);
xor_4  g11225(new_n11601, new_n11588, new_n11602);
xor_4  g11226(new_n11602, new_n11581, new_n11603);
nand_5 g11227(new_n3609, new_n3605, new_n11604);
not_8  g11228(new_n3621, new_n11605);
nand_5 g11229(new_n11605, new_n3610, new_n11606);
nand_5 g11230(new_n11606, new_n11604, new_n11607);
and_5  g11231(new_n3645, new_n3644, new_n11608);
nor_5  g11232(new_n3647, new_n3643, new_n11609);
or_5   g11233(new_n11609, new_n11608, new_n11610);
and_5  g11234(n9956, n6826, new_n11611);
and_5  g11235(n6797, n4826, new_n11612);
xor_4  g11236(new_n11612, new_n11611, new_n11613);
nand_5 g11237(n7610, n6294, new_n11614);
and_5  g11238(n6611, n6358, new_n11615);
xor_4  g11239(new_n11615, new_n11614, new_n11616);
xor_4  g11240(new_n11616, new_n11613, new_n11617);
xor_4  g11241(new_n11617, new_n11610, new_n11618);
nand_5 g11242(n7733, n3146, new_n11619);
and_5  g11243(new_n3602_1, new_n3601, new_n11620);
nor_5  g11244(new_n3604, new_n3600, new_n11621);
nor_5  g11245(new_n11621, new_n11620, new_n11622);
xor_4  g11246(new_n11622, new_n11619, new_n11623);
xor_4  g11247(new_n11623, new_n11618, new_n11624);
nand_5 g11248(n5198, n217, new_n11625);
and_5  g11249(n5283, n503, new_n11626);
xor_4  g11250(new_n11626, new_n11625, new_n11627);
and_5  g11251(n4970, n137, new_n11628);
and_5  g11252(n11296, n3992, new_n11629);
xor_4  g11253(new_n11629, new_n11628, new_n11630);
xor_4  g11254(new_n11630, new_n11627, new_n11631);
nor_5  g11255(new_n3618, new_n3617, new_n11632);
nand_5 g11256(n7733, n6797, new_n11633);
and_5  g11257(new_n3618, new_n3617, new_n11634);
nor_5  g11258(new_n11634, new_n11633, new_n11635);
nor_5  g11259(new_n11635, new_n11632, new_n11636);
nand_5 g11260(n11311, n10439, new_n11637);
and_5  g11261(n6126, n4203, new_n11638);
xor_4  g11262(new_n11638, new_n11637, new_n11639);
xor_4  g11263(new_n11639, new_n11636, new_n11640);
xor_4  g11264(new_n11640, new_n11631, new_n11641);
xor_4  g11265(new_n11641, new_n11624, new_n11642);
xor_4  g11266(new_n11642, new_n11607, new_n11643);
xor_4  g11267(new_n11643, new_n11603, new_n11644);
and_5  g11268(new_n3586, new_n3583, new_n11645);
nor_5  g11269(new_n3588, new_n3580, new_n11646);
nor_5  g11270(new_n11646, new_n11645, new_n11647);
and_5  g11271(new_n3629, new_n3626, new_n11648);
nor_5  g11272(new_n3631, new_n3623, new_n11649);
nor_5  g11273(new_n11649, new_n11648, new_n11650);
xor_4  g11274(new_n11650, new_n11647, new_n11651);
xor_4  g11275(new_n11651, new_n11644, new_n11652);
xor_4  g11276(new_n11652, new_n11577, new_n11653);
xor_4  g11277(new_n11653, new_n11562, new_n11654);
nor_5  g11278(new_n3590, new_n3555, new_n11655);
not_8  g11279(new_n3591, new_n11656);
nor_5  g11280(new_n3594, new_n11656, new_n11657);
nor_5  g11281(new_n11657, new_n11655, new_n11658);
nand_5 g11282(new_n3565, new_n3561, new_n11659);
not_8  g11283(new_n3578, new_n11660);
nand_5 g11284(new_n11660, new_n3566, new_n11661);
and_5  g11285(new_n11661, new_n11659, new_n11662_1);
nand_5 g11286(n4086, n1471, new_n11663);
and_5  g11287(n10391, n9400, new_n11664);
and_5  g11288(new_n3560, new_n3556, new_n11665);
or_5   g11289(new_n11665, new_n3557, new_n11666);
not_8  g11290(new_n11666, new_n11667);
and_5  g11291(new_n11667, new_n11664, new_n11668);
and_5  g11292(new_n11664, new_n3231, new_n11669);
nor_5  g11293(new_n11669, new_n11667, new_n11670);
or_5   g11294(new_n11670, new_n11668, new_n11671);
nand_5 g11295(n11757, n2577, new_n11672);
nand_5 g11296(n9637, n3172, new_n11673);
and_5  g11297(n5240, n3842, new_n11674);
xor_4  g11298(new_n11674, new_n11673, new_n11675);
xor_4  g11299(new_n11675, new_n11672, new_n11676);
nor_5  g11300(new_n3125, new_n3124_1, new_n11677);
and_5  g11301(new_n3125, new_n3124_1, new_n11678);
nor_5  g11302(new_n11678, new_n3123, new_n11679);
nor_5  g11303(new_n11679, new_n11677, new_n11680);
xor_4  g11304(new_n11680, new_n11676, new_n11681);
xor_4  g11305(new_n11681, new_n11671, new_n11682);
xor_4  g11306(new_n11682, new_n11663, new_n11683);
nand_5 g11307(n7236, n1357, new_n11684);
and_5  g11308(new_n3133, new_n3131, new_n11685);
and_5  g11309(new_n3140, new_n3134, new_n11686);
nor_5  g11310(new_n11686, new_n11685, new_n11687);
xor_4  g11311(new_n11687, new_n11684, new_n11688);
xor_4  g11312(new_n11688, new_n11683, new_n11689);
xor_4  g11313(new_n11689, new_n11662_1, new_n11690);
nand_5 g11314(n1835, n1333, new_n11691);
and_5  g11315(n11917, n11821, new_n11692);
xor_4  g11316(new_n11692, new_n11691, new_n11693);
and_5  g11317(n12753, n3602, new_n11694);
and_5  g11318(n8595, n4187, new_n11695);
xor_4  g11319(new_n11695, new_n11694, new_n11696);
and_5  g11320(n6877, n4190, new_n11697);
and_5  g11321(n10174, n3719, new_n11698);
xor_4  g11322(new_n11698, new_n11697, new_n11699);
xor_4  g11323(new_n11699, new_n11696, new_n11700);
xor_4  g11324(new_n11700, new_n11693, new_n11701);
and_5  g11325(new_n3574, new_n3573, new_n11702);
not_8  g11326(new_n3572, new_n11703);
nor_5  g11327(new_n3576, new_n11703, new_n11704);
nor_5  g11328(new_n11704, new_n11702, new_n11705);
and_5  g11329(n9080, n4921, new_n11706);
xor_4  g11330(new_n11706, new_n11705, new_n11707_1);
xor_4  g11331(new_n11707_1, new_n11701, new_n11708);
or_5   g11332(new_n3128, new_n3122, new_n11709);
not_8  g11333(new_n3141, new_n11710);
nand_5 g11334(new_n11710, new_n3129, new_n11711);
and_5  g11335(new_n11711, new_n11709, new_n11712);
xor_4  g11336(new_n11712, new_n11708, new_n11713);
xor_4  g11337(new_n11713, new_n11690, new_n11714);
and_5  g11338(new_n3671, new_n3669, new_n11715);
nor_5  g11339(new_n3673, new_n3666, new_n11716);
nor_5  g11340(new_n11716, new_n11715, new_n11717);
xor_4  g11341(new_n11717, new_n11714, new_n11718);
xor_4  g11342(new_n11718, new_n11658, new_n11719);
nor_5  g11343(new_n3633, new_n3597, new_n11720);
nor_5  g11344(new_n3637, new_n3635, new_n11721);
nor_5  g11345(new_n11721, new_n11720, new_n11722);
xor_4  g11346(new_n11722, new_n11719, new_n11723);
xor_4  g11347(new_n11723, new_n11654, new_n11724);
and_5  g11348(new_n3682, new_n3638, new_n11725);
and_5  g11349(new_n3688, new_n3683, new_n11726);
or_5   g11350(new_n11726, new_n11725, new_n11727);
nor_5  g11351(new_n3675, new_n3640, new_n11728_1);
not_8  g11352(new_n3676, new_n11729);
nor_5  g11353(new_n3680, new_n11729, new_n11730);
or_5   g11354(new_n11730, new_n11728_1, new_n11731);
and_5  g11355(new_n3137, new_n3136, new_n11732);
not_8  g11356(new_n3135, new_n11733);
nor_5  g11357(new_n3139, new_n11733, new_n11734);
nor_5  g11358(new_n11734, new_n11732, new_n11735);
xor_4  g11359(new_n11735, new_n11731, new_n11736);
xor_4  g11360(new_n11736, new_n11727, new_n11737);
xor_4  g11361(new_n11737, new_n11724, new_n11738);
xor_4  g11362(new_n11738, new_n11559, new_n11739);
xor_4  g11363(new_n11739, new_n11557, n5257);
xor_4  g11364(new_n11011, new_n11002, n5411);
xor_4  g11365(new_n3536, new_n3526, n5435);
xor_4  g11366(new_n6001, new_n5995, n5641);
xor_4  g11367(new_n8452, new_n8441, n5670);
nor_5  g11368(new_n4850, new_n4821, new_n11745);
xor_4  g11369(new_n11745, new_n4818, n5693);
not_8  g11370(new_n1358, new_n11747);
xor_4  g11371(new_n11747, new_n1346, n5934);
nor_5  g11372(new_n11013, new_n11000, new_n11749);
xor_4  g11373(new_n11017, new_n11749, n6089);
or_5   g11374(new_n7674, new_n7671, new_n11751);
not_8  g11375(new_n11751, new_n11752);
nor_5  g11376(new_n7657, new_n7653, new_n11753);
and_5  g11377(new_n7662, new_n7658, new_n11754);
or_5   g11378(new_n11754, new_n11753, new_n11755_1);
not_8  g11379(new_n11755_1, new_n11756);
nand_5 g11380(n2564, n2253, new_n11757_1);
nand_5 g11381(n9195, n4189, new_n11758);
nand_5 g11382(n6687, n3865, new_n11759);
xor_4  g11383(new_n11759, new_n11758, new_n11760);
xor_4  g11384(new_n11760, new_n11757_1, new_n11761);
xor_4  g11385(new_n11761, new_n11756, new_n11762);
or_5   g11386(new_n7655, new_n7654, new_n11763);
not_8  g11387(new_n11763, new_n11764);
and_5  g11388(n6770, n4634, new_n11765);
xor_4  g11389(new_n11765, new_n11764, new_n11766);
nand_5 g11390(n3627, n2879, new_n11767);
not_8  g11391(new_n11767, new_n11768);
nand_5 g11392(n10223, n9920, new_n11769);
nand_5 g11393(n7265, n4516, new_n11770);
xor_4  g11394(new_n11770, new_n11769, new_n11771);
not_8  g11395(new_n11771, new_n11772);
xor_4  g11396(new_n11772, new_n11768, new_n11773);
xor_4  g11397(new_n11773, new_n11766, new_n11774);
xor_4  g11398(new_n11774, new_n11762, new_n11775);
and_5  g11399(new_n7666, new_n7663, new_n11776);
or_5   g11400(new_n7665, new_n7664, new_n11777);
not_8  g11401(new_n7667, new_n11778);
or_5   g11402(new_n7670, new_n11778, new_n11779);
xor_4  g11403(new_n11779, new_n11777, new_n11780_1);
nor_5  g11404(new_n11780_1, new_n11776, new_n11781);
xor_4  g11405(new_n11781, new_n11775, new_n11782);
not_8  g11406(new_n11782, new_n11783);
xor_4  g11407(new_n11783, new_n11752, new_n11784);
nor_5  g11408(new_n7675, new_n7652, new_n11785);
or_5   g11409(new_n7679, new_n11785, new_n11786);
xor_4  g11410(new_n11786, new_n11784, new_n11787);
not_8  g11411(new_n7716, new_n11788);
nor_5  g11412(new_n7719, new_n11788, new_n11789);
nor_5  g11413(new_n7799, new_n11789, new_n11790);
nor_5  g11414(new_n7714, new_n7688, new_n11791_1);
and_5  g11415(new_n7715, new_n7687, new_n11792);
or_5   g11416(new_n11792, new_n11791_1, new_n11793);
not_8  g11417(new_n11793, new_n11794);
or_5   g11418(new_n7712, new_n7709, new_n11795);
nor_5  g11419(new_n7693, new_n7689, new_n11796);
and_5  g11420(new_n7698, new_n7694, new_n11797);
or_5   g11421(new_n11797, new_n11796, new_n11798);
not_8  g11422(new_n11798, new_n11799);
nand_5 g11423(n12221, n10928, new_n11800);
nand_5 g11424(n12145, n6986, new_n11801);
nand_5 g11425(n10217, n8336, new_n11802);
xor_4  g11426(new_n11802, new_n11801, new_n11803);
xor_4  g11427(new_n11803, new_n11800, new_n11804);
xor_4  g11428(new_n11804, new_n11799, new_n11805);
or_5   g11429(new_n7691, new_n7690_1, new_n11806);
not_8  g11430(new_n11806, new_n11807);
and_5  g11431(n2522, n2226, new_n11808);
xor_4  g11432(new_n11808, new_n11807, new_n11809);
nand_5 g11433(n10678, n2024, new_n11810);
not_8  g11434(new_n11810, new_n11811);
nand_5 g11435(n9189, n1094, new_n11812);
nand_5 g11436(n7946, n7320, new_n11813);
xor_4  g11437(new_n11813, new_n11812, new_n11814);
not_8  g11438(new_n11814, new_n11815);
xor_4  g11439(new_n11815, new_n11811, new_n11816);
xor_4  g11440(new_n11816, new_n11809, new_n11817);
xor_4  g11441(new_n11817, new_n11805, new_n11818);
and_5  g11442(new_n7702, new_n7699, new_n11819);
or_5   g11443(new_n7701, new_n7700, new_n11820);
or_5   g11444(new_n7707, new_n7704, new_n11821_1);
xor_4  g11445(new_n11821_1, new_n11820, new_n11822);
nor_5  g11446(new_n11822, new_n11819, new_n11823);
xor_4  g11447(new_n11823, new_n11818, new_n11824);
not_8  g11448(new_n11824, new_n11825);
xor_4  g11449(new_n11825, new_n11795, new_n11826);
xor_4  g11450(new_n11826, new_n11794, new_n11827);
nand_5 g11451(new_n7753, new_n7750, new_n11828);
not_8  g11452(new_n11828, new_n11829);
or_5   g11453(new_n7736, new_n7735, new_n11830);
not_8  g11454(new_n11830, new_n11831);
nand_5 g11455(n7160, n521, new_n11832);
not_8  g11456(new_n11832, new_n11833);
xor_4  g11457(new_n11833, new_n11831, new_n11834);
nand_5 g11458(n2515, n2498, new_n11835);
not_8  g11459(new_n11835, new_n11836);
nand_5 g11460(n2558, n1199, new_n11837);
nand_5 g11461(n5579, n4828, new_n11838);
xor_4  g11462(new_n11838, new_n11837, new_n11839);
xor_4  g11463(new_n11839, new_n11836, new_n11840);
xor_4  g11464(new_n11840, new_n11834, new_n11841);
not_8  g11465(new_n11841, new_n11842);
or_5   g11466(new_n7739, new_n7732, new_n11843);
nand_5 g11467(n12391, n5798, new_n11844);
not_8  g11468(new_n11844, new_n11845);
nand_5 g11469(n7891, n6016, new_n11846);
nand_5 g11470(n12069, n2347, new_n11847);
xor_4  g11471(new_n11847, new_n11846, new_n11848);
not_8  g11472(new_n11848, new_n11849);
xor_4  g11473(new_n11849, new_n11845, new_n11850);
xor_4  g11474(new_n11850, new_n11843, new_n11851);
xor_4  g11475(new_n11851, new_n11842, new_n11852);
or_5   g11476(new_n7744, new_n7740, new_n11853);
or_5   g11477(new_n7742, new_n7741, new_n11854);
or_5   g11478(new_n7747, new_n7746, new_n11855);
and_5  g11479(new_n11855, new_n7745, new_n11856);
xor_4  g11480(new_n11856, new_n11854, new_n11857);
and_5  g11481(new_n11857, new_n11853, new_n11858);
xor_4  g11482(new_n11858, new_n11852, new_n11859);
not_8  g11483(new_n11859, new_n11860);
nand_5 g11484(new_n11860, new_n11829, new_n11861);
or_5   g11485(new_n11860, new_n11829, new_n11862);
and_5  g11486(new_n11862, new_n11861, new_n11863);
not_8  g11487(new_n11863, new_n11864);
nor_5  g11488(new_n7755, new_n7724, new_n11865);
and_5  g11489(new_n7756, new_n7723, new_n11866);
nor_5  g11490(new_n11866, new_n11865, new_n11867);
xor_4  g11491(new_n11867, new_n11864, new_n11868);
not_8  g11492(new_n11868, new_n11869);
or_5   g11493(new_n7785, new_n7782, new_n11870);
not_8  g11494(new_n11870, new_n11871);
nor_5  g11495(new_n7767, new_n7763, new_n11872);
and_5  g11496(new_n7773, new_n7768, new_n11873);
or_5   g11497(new_n11873, new_n11872, new_n11874);
nand_5 g11498(n11153, n5153, new_n11875);
not_8  g11499(new_n11875, new_n11876_1);
nand_5 g11500(n7270, n5314, new_n11877_1);
nand_5 g11501(n11222, n2507, new_n11878);
xor_4  g11502(new_n11878, new_n11877_1, new_n11879);
not_8  g11503(new_n11879, new_n11880);
xor_4  g11504(new_n11880, new_n11876_1, new_n11881);
not_8  g11505(new_n11881, new_n11882);
xor_4  g11506(new_n11882, new_n11874, new_n11883);
or_5   g11507(new_n7765, new_n7764, new_n11884);
not_8  g11508(new_n11884, new_n11885);
nand_5 g11509(n996, n806, new_n11886);
not_8  g11510(new_n11886, new_n11887);
xor_4  g11511(new_n11887, new_n11885, new_n11888);
nand_5 g11512(n9111, n5319, new_n11889);
nand_5 g11513(n5767, n3342, new_n11890);
nand_5 g11514(n9763, n9457, new_n11891);
xor_4  g11515(new_n11891, new_n11890, new_n11892_1);
not_8  g11516(new_n11892_1, new_n11893);
xor_4  g11517(new_n11893, new_n11889, new_n11894);
xor_4  g11518(new_n11894, new_n11888, new_n11895);
xor_4  g11519(new_n11895, new_n11883, new_n11896);
not_8  g11520(new_n11896, new_n11897);
and_5  g11521(new_n7777, new_n7774, new_n11898);
or_5   g11522(new_n7776, new_n7775, new_n11899);
not_8  g11523(new_n11899, new_n11900);
nand_5 g11524(new_n7781, new_n7778, new_n11901);
not_8  g11525(new_n11901, new_n11902);
xor_4  g11526(new_n11902, new_n11900, new_n11903);
nor_5  g11527(new_n11903, new_n11898, new_n11904);
xor_4  g11528(new_n11904, new_n11897, new_n11905);
not_8  g11529(new_n11905, new_n11906);
xor_4  g11530(new_n11906, new_n11871, new_n11907);
not_8  g11531(new_n11907, new_n11908);
or_5   g11532(new_n7786, new_n7762, new_n11909);
nand_5 g11533(new_n7790, new_n11909, new_n11910);
xor_4  g11534(new_n11910, new_n11908, new_n11911);
xor_4  g11535(new_n11911, new_n11869, new_n11912);
nor_5  g11536(new_n7791, new_n7758, new_n11913);
and_5  g11537(new_n7797, new_n7792, new_n11914);
or_5   g11538(new_n11914, new_n11913, new_n11915);
not_8  g11539(new_n11915, new_n11916);
xor_4  g11540(new_n11916, new_n11912, new_n11917_1);
xor_4  g11541(new_n11917_1, new_n11827, new_n11918);
xor_4  g11542(new_n11918, new_n11790, new_n11919_1);
not_8  g11543(new_n11919_1, new_n11920);
nor_5  g11544(new_n11920, new_n11787, new_n11921);
and_5  g11545(new_n7683, new_n7680, new_n11922_1);
nor_5  g11546(new_n7801, new_n7684, new_n11923);
or_5   g11547(new_n11923, new_n11922_1, new_n11924);
not_8  g11548(new_n11787, new_n11925);
xor_4  g11549(new_n11920, new_n11925, new_n11926);
nor_5  g11550(new_n11926, new_n11924, new_n11927);
nor_5  g11551(new_n11927, new_n11921, new_n11928);
and_5  g11552(new_n11917_1, new_n11827, new_n11929);
and_5  g11553(new_n11918, new_n11790, new_n11930);
or_5   g11554(new_n11930, new_n11929, new_n11931);
and_5  g11555(new_n11911, new_n11869, new_n11932);
and_5  g11556(new_n11916, new_n11912, new_n11933);
nor_5  g11557(new_n11933, new_n11932, new_n11934);
nor_5  g11558(new_n11821_1, new_n11820, new_n11935);
nor_5  g11559(new_n11823, new_n11818, new_n11936);
or_5   g11560(new_n11936, new_n11935, new_n11937);
and_5  g11561(new_n11761, new_n11756, new_n11938);
and_5  g11562(new_n11774, new_n11762, new_n11939);
or_5   g11563(new_n11939, new_n11938, new_n11940);
nand_5 g11564(n2522, n1094, new_n11941);
and_5  g11565(new_n11878, new_n11877_1, new_n11942);
nor_5  g11566(new_n11880, new_n11876_1, new_n11943);
nor_5  g11567(new_n11943, new_n11942, new_n11944);
xor_4  g11568(new_n11944, new_n11941, new_n11945);
xor_4  g11569(new_n11945, new_n11940, new_n11946);
xor_4  g11570(new_n11946, new_n11937, new_n11947);
and_5  g11571(new_n11804, new_n11799, new_n11948);
and_5  g11572(new_n11817, new_n11805, new_n11949);
or_5   g11573(new_n11949, new_n11948, new_n11950);
and_5  g11574(n10678, n9189, new_n11951);
xor_4  g11575(new_n11951, new_n11950, new_n11952);
and_5  g11576(new_n11813, new_n11812, new_n11953);
nor_5  g11577(new_n11815, new_n11811, new_n11954);
nor_5  g11578(new_n11954, new_n11953, new_n11955);
nand_5 g11579(n7946, n7523, new_n11956);
nand_5 g11580(n10223, n3627, new_n11957);
and_5  g11581(n3865, n2564, new_n11958);
xor_4  g11582(new_n11958, new_n11957, new_n11959);
xor_4  g11583(new_n11959, new_n11956, new_n11960);
xor_4  g11584(new_n11960, new_n11955, new_n11961);
nand_5 g11585(n12221, n6986, new_n11962);
and_5  g11586(n8336, n7823, new_n11963);
xor_4  g11587(new_n11963, new_n11962, new_n11964);
xor_4  g11588(new_n11964, new_n11961, new_n11965);
and_5  g11589(new_n11770, new_n11769, new_n11966);
nor_5  g11590(new_n11772, new_n11768, new_n11967_1);
or_5   g11591(new_n11967_1, new_n11966, new_n11968);
nor_5  g11592(new_n11808, new_n11807, new_n11969);
and_5  g11593(new_n11816, new_n11809, new_n11970);
nor_5  g11594(new_n11970, new_n11969, new_n11971);
xor_4  g11595(new_n11971, new_n11968, new_n11972);
and_5  g11596(new_n11847, new_n11846, new_n11973);
nor_5  g11597(new_n11849, new_n11845, new_n11974);
nor_5  g11598(new_n11974, new_n11973, new_n11975);
nand_5 g11599(n6687, n2512, new_n11976);
nor_5  g11600(new_n11838, new_n11837, new_n11977);
and_5  g11601(new_n11838, new_n11837, new_n11978);
nor_5  g11602(new_n11978, new_n11835, new_n11979);
nor_5  g11603(new_n11979, new_n11977, new_n11980);
xor_4  g11604(new_n11980, new_n11976, new_n11981);
xor_4  g11605(new_n11981, new_n11975, new_n11982);
xor_4  g11606(new_n11982, new_n11972, new_n11983);
xor_4  g11607(new_n11983, new_n11965, new_n11984);
nand_5 g11608(n11153, n2507, new_n11985);
and_5  g11609(n7270, n996, new_n11986);
xor_4  g11610(new_n11986, new_n11985, new_n11987);
nand_5 g11611(n7160, n6016, new_n11988);
and_5  g11612(n5767, n806, new_n11989);
xor_4  g11613(new_n11989, new_n11988, new_n11990);
xor_4  g11614(new_n11990, new_n11987, new_n11991);
nand_5 g11615(n4828, n521, new_n11992);
and_5  g11616(n5579, n2515, new_n11993);
xor_4  g11617(new_n11993, new_n11992, new_n11994);
and_5  g11618(n12069, n1576, new_n11995);
and_5  g11619(n5314, n5153, new_n11996);
xor_4  g11620(new_n11996, new_n11995, new_n11997);
xor_4  g11621(new_n11997, new_n11994, new_n11998);
xor_4  g11622(new_n11998, new_n11991, new_n11999_1);
nor_5  g11623(new_n11759, new_n11758, new_n12000_1);
and_5  g11624(new_n11759, new_n11758, new_n12001);
nor_5  g11625(new_n12001, new_n11757_1, new_n12002);
or_5   g11626(new_n12002, new_n12000_1, new_n12003);
and_5  g11627(n4516, n2879, new_n12004);
nand_5 g11628(n4189, n2253, new_n12005_1);
and_5  g11629(n9920, n4634, new_n12006);
xor_4  g11630(new_n12006, new_n12005_1, new_n12007);
xor_4  g11631(new_n12007, new_n12004, new_n12008);
xor_4  g11632(new_n12008, new_n12003, new_n12009);
xor_4  g11633(new_n12009, new_n11999_1, new_n12010);
nor_5  g11634(new_n11765, new_n11764, new_n12011);
and_5  g11635(new_n11773, new_n11766, new_n12012);
nor_5  g11636(new_n12012, new_n12011, new_n12013);
and_5  g11637(new_n11887, new_n11885, new_n12014_1);
and_5  g11638(new_n11894, new_n11888, new_n12015);
nor_5  g11639(new_n12015, new_n12014_1, new_n12016);
xor_4  g11640(new_n12016, new_n12013, new_n12017);
xor_4  g11641(new_n12017, new_n12010, new_n12018);
xor_4  g11642(new_n12018, new_n11984, new_n12019);
xor_4  g11643(new_n12019, new_n11952, new_n12020_1);
xor_4  g11644(new_n12020_1, new_n11947, new_n12021);
and_5  g11645(new_n11902, new_n11900, new_n12022);
nor_5  g11646(new_n11904, new_n11897, new_n12023);
or_5   g11647(new_n12023, new_n12022, new_n12024);
nand_5 g11648(n12145, n2226, new_n12025_1);
nor_5  g11649(new_n11802, new_n11801, new_n12026);
and_5  g11650(new_n11802, new_n11801, new_n12027);
nor_5  g11651(new_n12027, new_n11800, new_n12028);
or_5   g11652(new_n12028, new_n12026, new_n12029);
and_5  g11653(n9195, n6770, new_n12030);
and_5  g11654(n11222, n6431, new_n12031);
xor_4  g11655(new_n12031, new_n12030, new_n12032);
nand_5 g11656(n10928, n10217, new_n12033);
and_5  g11657(n7320, n2024, new_n12034);
xor_4  g11658(new_n12034, new_n12033, new_n12035);
xor_4  g11659(new_n12035, new_n12032, new_n12036);
and_5  g11660(n5319, n3342, new_n12037);
and_5  g11661(n9457, n9111, new_n12038);
and_5  g11662(n9763, n4817, new_n12039);
xor_4  g11663(new_n12039, new_n12038, new_n12040);
xor_4  g11664(new_n12040, new_n12037, new_n12041);
xor_4  g11665(new_n12041, new_n12036, new_n12042);
xor_4  g11666(new_n12042, new_n12029, new_n12043);
xor_4  g11667(new_n12043, new_n12025_1, new_n12044_1);
xor_4  g11668(new_n12044_1, new_n12024, new_n12045);
xor_4  g11669(new_n12045, new_n12021, new_n12046);
nor_5  g11670(new_n11825, new_n11795, new_n12047);
not_8  g11671(new_n11826, new_n12048);
nor_5  g11672(new_n12048, new_n11794, new_n12049);
nor_5  g11673(new_n12049, new_n12047, new_n12050);
not_8  g11674(new_n11854, new_n12051);
and_5  g11675(new_n11856, new_n12051, new_n12052);
not_8  g11676(new_n11852, new_n12053);
nor_5  g11677(new_n11858, new_n12053, new_n12054);
nor_5  g11678(new_n12054, new_n12052, new_n12055);
nor_5  g11679(new_n11779, new_n11777, new_n12056);
nor_5  g11680(new_n11781, new_n11775, new_n12057);
or_5   g11681(new_n12057, new_n12056, new_n12058);
or_5   g11682(new_n11882, new_n11874, new_n12059);
not_8  g11683(new_n11895, new_n12060);
nand_5 g11684(new_n12060, new_n11883, new_n12061);
nand_5 g11685(new_n12061, new_n12059, new_n12062);
and_5  g11686(new_n11833, new_n11831, new_n12063);
and_5  g11687(new_n11840, new_n11834, new_n12064);
or_5   g11688(new_n12064, new_n12063, new_n12065);
and_5  g11689(n7891, n5798, new_n12066);
xor_4  g11690(new_n12066, new_n12065, new_n12067);
nand_5 g11691(n12391, n2347, new_n12068);
and_5  g11692(n7265, n2087, new_n12069_1);
xor_4  g11693(new_n12069_1, new_n12068, new_n12070);
xor_4  g11694(new_n12070, new_n12067, new_n12071);
xor_4  g11695(new_n12071, new_n12062, new_n12072);
nand_5 g11696(n2498, n1199, new_n12073);
and_5  g11697(n6578, n2558, new_n12074);
xor_4  g11698(new_n12074, new_n12073, new_n12075);
xor_4  g11699(new_n12075, new_n12072, new_n12076_1);
xor_4  g11700(new_n12076_1, new_n12058, new_n12077);
xor_4  g11701(new_n12077, new_n12055, new_n12078);
xor_4  g11702(new_n12078, new_n12050, new_n12079);
xor_4  g11703(new_n12079, new_n12046, new_n12080);
and_5  g11704(new_n11905, new_n11871, new_n12081);
nor_5  g11705(new_n11910, new_n11907, new_n12082);
or_5   g11706(new_n12082, new_n12081, new_n12083);
and_5  g11707(new_n11891, new_n11890, new_n12084);
not_8  g11708(new_n11889, new_n12085);
nor_5  g11709(new_n11893, new_n12085, new_n12086);
or_5   g11710(new_n12086, new_n12084, new_n12087);
not_8  g11711(new_n11850, new_n12088);
nor_5  g11712(new_n12088, new_n11843, new_n12089);
or_5   g11713(new_n11851, new_n11841, new_n12090);
not_8  g11714(new_n12090, new_n12091);
nor_5  g11715(new_n12091, new_n12089, new_n12092);
xor_4  g11716(new_n12092, new_n12087, new_n12093);
xor_4  g11717(new_n12093, new_n12083, new_n12094);
xor_4  g11718(new_n12094, new_n12080, new_n12095);
xor_4  g11719(new_n12095, new_n11934, new_n12096);
nor_5  g11720(new_n11783, new_n11751, new_n12097);
nor_5  g11721(new_n11786, new_n11784, new_n12098);
or_5   g11722(new_n12098, new_n12097, new_n12099);
and_5  g11723(new_n11860, new_n11829, new_n12100);
nor_5  g11724(new_n11867, new_n11864, new_n12101);
nor_5  g11725(new_n12101, new_n12100, new_n12102);
xor_4  g11726(new_n12102, new_n12099, new_n12103);
xor_4  g11727(new_n12103, new_n12096, new_n12104);
xor_4  g11728(new_n12104, new_n11931, new_n12105);
xor_4  g11729(new_n12105, new_n11928, n6192);
xor_4  g11730(new_n872, new_n840, n6273);
not_8  g11731(new_n7457, new_n12108);
xor_4  g11732(new_n7458, new_n12108, n6445);
nor_5  g11733(new_n9261, new_n9235, new_n12110);
xor_4  g11734(new_n9265, new_n12110, n6645);
xor_4  g11735(new_n7836, new_n7835, n6689);
xor_4  g11736(new_n1347, new_n1259, n6742);
xor_4  g11737(new_n2058, new_n2014, n6809);
not_8  g11738(new_n6687_1, new_n12115);
xor_4  g11739(new_n12115, new_n6683, n6822);
xor_4  g11740(new_n11008, new_n11007, n6860);
xor_4  g11741(new_n9257, new_n9249, n7193);
not_8  g11742(new_n7462, new_n12119);
xnor_4 g11743(new_n12119, new_n7461, n7568);
xor_4  g11744(new_n1355, new_n1354, n7676);
not_8  g11745(new_n500, new_n12122);
nor_5  g11746(new_n878, new_n12122, new_n12123);
and_5  g11747(new_n1024, new_n880, new_n12124);
or_5   g11748(new_n12124, new_n12123, new_n12125);
nor_5  g11749(new_n1018, new_n923, new_n12126);
not_8  g11750(new_n1022, new_n12127);
and_5  g11751(new_n12127, new_n1019, new_n12128);
or_5   g11752(new_n12128, new_n12126, new_n12129);
and_5  g11753(new_n1010, new_n968, new_n12130);
and_5  g11754(new_n1017, new_n1011, new_n12131);
nor_5  g11755(new_n12131, new_n12130, new_n12132);
and_5  g11756(n9241, n1209, new_n12133);
not_8  g11757(new_n1002, new_n12134);
nor_5  g11758(new_n12134, new_n969, new_n12135);
and_5  g11759(new_n1009, new_n1003, new_n12136);
nor_5  g11760(new_n12136, new_n12135, new_n12137);
not_8  g11761(new_n997, new_n12138);
nand_5 g11762(new_n999, new_n12138, new_n12139);
not_8  g11763(new_n12139, new_n12140);
nor_5  g11764(new_n1001, new_n995, new_n12141);
or_5   g11765(new_n12141, new_n12140, new_n12142);
nand_5 g11766(new_n458, new_n453, new_n12143);
not_8  g11767(new_n471, new_n12144);
nand_5 g11768(new_n12144, new_n459, new_n12145_1);
and_5  g11769(new_n12145_1, new_n12143, new_n12146);
and_5  g11770(new_n463, new_n461, new_n12147);
and_5  g11771(new_n470, new_n464, new_n12148);
or_5   g11772(new_n12148, new_n12147, new_n12149);
and_5  g11773(n12705, n2508, new_n12150);
nor_5  g11774(new_n456, new_n455, new_n12151);
and_5  g11775(new_n456, new_n455, new_n12152);
nor_5  g11776(new_n12152, new_n454, new_n12153);
nor_5  g11777(new_n12153, new_n12151, new_n12154);
xor_4  g11778(new_n12154, new_n12150, new_n12155);
and_5  g11779(n3986, n1980, new_n12156);
and_5  g11780(n10848, n5857, new_n12157);
xor_4  g11781(new_n12157, new_n12156, new_n12158);
and_5  g11782(n11257, n2509, new_n12159);
and_5  g11783(n4005, n1097, new_n12160);
xor_4  g11784(new_n12160, new_n12159, new_n12161);
xor_4  g11785(new_n12161, new_n12158, new_n12162);
xor_4  g11786(new_n12162, new_n12155, new_n12163);
xor_4  g11787(new_n12163, new_n12149, new_n12164);
nand_5 g11788(n8028, n45, new_n12165);
and_5  g11789(new_n890, new_n889, new_n12166);
nor_5  g11790(new_n892, new_n888, new_n12167);
nor_5  g11791(new_n12167, new_n12166, new_n12168);
xor_4  g11792(new_n12168, new_n12165, new_n12169);
nor_5  g11793(new_n902, new_n901, new_n12170);
nand_5 g11794(n9241, n7500, new_n12171);
and_5  g11795(new_n902, new_n901, new_n12172);
nor_5  g11796(new_n12172, new_n12171, new_n12173);
nor_5  g11797(new_n12173, new_n12170, new_n12174);
xor_4  g11798(new_n12174, new_n12169, new_n12175);
and_5  g11799(n4312, n2585, new_n12176);
and_5  g11800(new_n467, new_n466, new_n12177);
not_8  g11801(new_n465, new_n12178);
nor_5  g11802(new_n469, new_n12178, new_n12179);
or_5   g11803(new_n12179, new_n12177, new_n12180);
and_5  g11804(n10644, n7354, new_n12181);
nand_5 g11805(n12706, n5964, new_n12182);
and_5  g11806(n12720, n12025, new_n12183);
xor_4  g11807(new_n12183, new_n12182, new_n12184);
xor_4  g11808(new_n12184, new_n12181, new_n12185);
xor_4  g11809(new_n12185, new_n12180, new_n12186);
xor_4  g11810(new_n12186, new_n12176, new_n12187);
xor_4  g11811(new_n12187, new_n12175, new_n12188);
xor_4  g11812(new_n12188, new_n12164, new_n12189);
xor_4  g11813(new_n12189, new_n12146, new_n12190);
nand_5 g11814(n7436, n4141, new_n12191);
and_5  g11815(new_n898, new_n896, new_n12192);
and_5  g11816(new_n904, new_n899, new_n12193);
nor_5  g11817(new_n12193, new_n12192, new_n12194);
xor_4  g11818(new_n12194, new_n12191, new_n12195);
xor_4  g11819(new_n12195, new_n12190, new_n12196);
xor_4  g11820(new_n12196, new_n12142, new_n12197);
xor_4  g11821(new_n12197, new_n12137, new_n12198);
xor_4  g11822(new_n12198, new_n12133, new_n12199);
xor_4  g11823(new_n12199, new_n12132, new_n12200);
and_5  g11824(n10547, n6038, new_n12201);
and_5  g11825(new_n933, new_n932, new_n12202);
nor_5  g11826(new_n935, new_n931, new_n12203);
nor_5  g11827(new_n12203, new_n12202, new_n12204);
xor_4  g11828(new_n12204, new_n12201, new_n12205);
and_5  g11829(new_n945, new_n944, new_n12206);
not_8  g11830(new_n943, new_n12207);
nor_5  g11831(new_n947, new_n12207, new_n12208);
nor_5  g11832(new_n12208, new_n12206, new_n12209);
and_5  g11833(n12044, n8476, new_n12210);
nand_5 g11834(n11892, n5814, new_n12211);
and_5  g11835(n3616, n1512, new_n12212);
xor_4  g11836(new_n12212, new_n12211, new_n12213);
xor_4  g11837(new_n12213, new_n12210, new_n12214);
xor_4  g11838(new_n12214, new_n12209, new_n12215);
xor_4  g11839(new_n12215, new_n12205, new_n12216);
nand_5 g11840(n12299, n4928, new_n12217);
and_5  g11841(new_n989, new_n988, new_n12218);
not_8  g11842(new_n987, new_n12219);
nor_5  g11843(new_n991, new_n12219, new_n12220);
nor_5  g11844(new_n12220, new_n12218, new_n12221_1);
xor_4  g11845(new_n12221_1, new_n12217, new_n12222);
nand_5 g11846(n5069, n2530, new_n12223);
and_5  g11847(n10545, n2802, new_n12224);
xor_4  g11848(new_n12224, new_n12223, new_n12225);
xor_4  g11849(new_n12225, new_n12222, new_n12226);
xor_4  g11850(new_n12226, new_n12216, new_n12227);
nand_5 g11851(new_n936, new_n929, new_n12228);
not_8  g11852(new_n949, new_n12229);
nand_5 g11853(new_n12229, new_n937, new_n12230);
nand_5 g11854(new_n12230, new_n12228, new_n12231);
and_5  g11855(new_n985, new_n983, new_n12232);
and_5  g11856(new_n992_1, new_n986, new_n12233);
nor_5  g11857(new_n12233, new_n12232, new_n12234);
and_5  g11858(new_n941, new_n939, new_n12235);
and_5  g11859(new_n948, new_n942, new_n12236);
or_5   g11860(new_n12236, new_n12235, new_n12237);
and_5  g11861(n7690, n533, new_n12238);
xor_4  g11862(new_n12238, new_n12237, new_n12239);
xor_4  g11863(new_n12239, new_n12234, new_n12240);
xor_4  g11864(new_n12240, new_n12231, new_n12241);
xor_4  g11865(new_n12241, new_n12227, new_n12242);
and_5  g11866(n12704, n2393, new_n12243);
and_5  g11867(n7294, n5860, new_n12244);
xor_4  g11868(new_n12244, new_n12243, new_n12245);
nand_5 g11869(n12648, n6806, new_n12246);
and_5  g11870(n4499, n1564, new_n12247_1);
xor_4  g11871(new_n12247_1, new_n12246, new_n12248);
xor_4  g11872(new_n12248, new_n12245, new_n12249);
and_5  g11873(new_n976, new_n975, new_n12250);
nor_5  g11874(new_n978, new_n974, new_n12251);
nor_5  g11875(new_n12251, new_n12250, new_n12252);
and_5  g11876(n5694, n5331, new_n12253);
and_5  g11877(n7388, n4903, new_n12254);
xor_4  g11878(new_n12254, new_n12253, new_n12255);
xor_4  g11879(new_n12255, new_n12252, new_n12256);
xor_4  g11880(new_n12256, new_n12249, new_n12257);
and_5  g11881(n8276, n5105, new_n12258);
and_5  g11882(n5305, n615, new_n12259);
xor_4  g11883(new_n12259, new_n12258, new_n12260);
xor_4  g11884(new_n12260, new_n12257, new_n12261);
xor_4  g11885(new_n12261, new_n12242, new_n12262);
and_5  g11886(new_n912, new_n910, new_n12263);
nor_5  g11887(new_n914, new_n907, new_n12264);
nor_5  g11888(new_n12264, new_n12263, new_n12265);
and_5  g11889(new_n956, new_n954, new_n12266);
nor_5  g11890(new_n958, new_n951, new_n12267);
nor_5  g11891(new_n12267, new_n12266, new_n12268);
xor_4  g11892(new_n12268, new_n12265, new_n12269);
xor_4  g11893(new_n12269, new_n12262, new_n12270);
nand_5 g11894(n8759, n783, new_n12271);
and_5  g11895(n10510, n7500, new_n12272);
xor_4  g11896(new_n12272, new_n12271, new_n12273);
nor_5  g11897(new_n476, new_n475, new_n12274);
nor_5  g11898(new_n478, new_n473, new_n12275);
nor_5  g11899(new_n12275, new_n12274, new_n12276);
or_5   g11900(new_n980, new_n972, new_n12277);
not_8  g11901(new_n993, new_n12278);
nand_5 g11902(new_n12278, new_n981, new_n12279);
and_5  g11903(new_n12279, new_n12277, new_n12280);
xor_4  g11904(new_n12280, new_n12276, new_n12281);
xor_4  g11905(new_n12281, new_n12273, new_n12282);
xor_4  g11906(new_n12282, new_n12270, new_n12283);
nor_5  g11907(new_n960, new_n924, new_n12284);
nor_5  g11908(new_n966, new_n962, new_n12285);
or_5   g11909(new_n12285, new_n12284, new_n12286);
and_5  g11910(n7965, n1906, new_n12287);
xor_4  g11911(new_n12287, new_n12286, new_n12288);
xor_4  g11912(new_n12288, new_n12283, new_n12289);
nor_5  g11913(new_n480, new_n449, new_n12290);
nor_5  g11914(new_n499, new_n482, new_n12291);
or_5   g11915(new_n12291, new_n12290, new_n12292);
nor_5  g11916(new_n916, new_n881, new_n12293);
nor_5  g11917(new_n921, new_n918, new_n12294);
nor_5  g11918(new_n12294, new_n12293, new_n12295);
nand_5 g11919(new_n893, new_n886, new_n12296);
not_8  g11920(new_n905, new_n12297);
nand_5 g11921(new_n12297, new_n894, new_n12298);
nand_5 g11922(new_n12298, new_n12296, new_n12299_1);
and_5  g11923(n8236, n6776, new_n12300);
xor_4  g11924(new_n12300, new_n12299_1, new_n12301);
xor_4  g11925(new_n12301, new_n12295, new_n12302);
xor_4  g11926(new_n12302, new_n12292, new_n12303);
xor_4  g11927(new_n12303, new_n12289, new_n12304);
xor_4  g11928(new_n12304, new_n12200, new_n12305);
xor_4  g11929(new_n12305, new_n12129, new_n12306);
xor_4  g11930(new_n12306, new_n12125, n7966);
not_8  g11931(new_n11924, new_n12308);
xor_4  g11932(new_n11926, new_n12308, n7981);
nor_5  g11933(new_n11537, new_n11292, new_n12310);
and_5  g11934(new_n11550, new_n11538, new_n12311);
or_5   g11935(new_n12311, new_n12310, new_n12312);
nor_5  g11936(new_n11450, new_n11364, new_n12313);
and_5  g11937(new_n11536_1, new_n11451, new_n12314);
or_5   g11938(new_n12314, new_n12313, new_n12315);
nor_5  g11939(new_n11530, new_n11491, new_n12316);
nor_5  g11940(new_n11535, new_n11532, new_n12317);
nor_5  g11941(new_n12317, new_n12316, new_n12318);
and_5  g11942(new_n11524, new_n11493, new_n12319);
nor_5  g11943(new_n11528, new_n11526, new_n12320);
or_5   g11944(new_n12320, new_n12319, new_n12321);
nor_5  g11945(new_n11278, new_n11277, new_n12322);
nor_5  g11946(new_n11280, new_n11275, new_n12323);
nor_5  g11947(new_n12323, new_n12322, new_n12324);
nor_5  g11948(new_n11511, new_n11510, new_n12325);
nand_5 g11949(n7159, n2515, new_n12326);
and_5  g11950(new_n11511, new_n11510, new_n12327);
nor_5  g11951(new_n12327, new_n12326, new_n12328);
or_5   g11952(new_n12328, new_n12325, new_n12329);
and_5  g11953(n8717, n6986, new_n12330);
nand_5 g11954(n11222, n10022, new_n12331);
and_5  g11955(n12391, n1353, new_n12332);
xor_4  g11956(new_n12332, new_n12331, new_n12333);
xor_4  g11957(new_n12333, new_n12330, new_n12334);
xor_4  g11958(new_n12334, new_n12329, new_n12335);
xor_4  g11959(new_n12335, new_n12324, new_n12336);
xor_4  g11960(new_n12336, new_n12321, new_n12337);
xor_4  g11961(new_n12337, new_n12318, new_n12338);
and_5  g11962(new_n11521, new_n11519, new_n12339);
nor_5  g11963(new_n11523, new_n11516, new_n12340);
or_5   g11964(new_n12340, new_n12339, new_n12341);
or_5   g11965(new_n11502, new_n11496, new_n12342);
not_8  g11966(new_n11514, new_n12343);
nand_5 g11967(new_n12343, new_n11503, new_n12344);
nand_5 g11968(new_n12344, new_n12342, new_n12345);
nand_5 g11969(n12069, n4436, new_n12346);
and_5  g11970(n11999, n11153, new_n12347);
xor_4  g11971(new_n12347, new_n12346, new_n12348);
and_5  g11972(n7159, n1199, new_n12349);
and_5  g11973(n11967, n7160, new_n12350);
xor_4  g11974(new_n12350, new_n12349, new_n12351);
xor_4  g11975(new_n12351, new_n12348, new_n12352);
nor_5  g11976(new_n11499, new_n11498, new_n12353);
and_5  g11977(new_n11499, new_n11498, new_n12354);
nor_5  g11978(new_n12354, new_n11497, new_n12355);
nor_5  g11979(new_n12355, new_n12353, new_n12356);
nand_5 g11980(n6254, n4828, new_n12357);
and_5  g11981(n11407, n2087, new_n12358);
xor_4  g11982(new_n12358, new_n12357, new_n12359);
xor_4  g11983(new_n12359, new_n12356, new_n12360);
xor_4  g11984(new_n12360, new_n12352, new_n12361);
xor_4  g11985(new_n12361, new_n12345, new_n12362);
xor_4  g11986(new_n12362, new_n12341, new_n12363);
or_5   g11987(new_n11463, new_n11455, new_n12364);
not_8  g11988(new_n11476, new_n12365);
nand_5 g11989(new_n12365, new_n11464, new_n12366);
nand_5 g11990(new_n12366, new_n12364, new_n12367);
and_5  g11991(n12489, n6578, new_n12368);
nand_5 g11992(n12947, n996, new_n12369);
and_5  g11993(n9457, n5760, new_n12370);
xor_4  g11994(new_n12370, new_n12369, new_n12371);
xor_4  g11995(new_n12371, new_n12368, new_n12372);
xor_4  g11996(new_n12372, new_n12367, new_n12373);
and_5  g11997(new_n11507, new_n11505, new_n12374);
and_5  g11998(new_n11513, new_n11508, new_n12375);
or_5   g11999(new_n12375, new_n12374, new_n12376);
and_5  g12000(n7891, n447, new_n12377);
xor_4  g12001(new_n12377, new_n12376, new_n12378);
nand_5 g12002(n12777, n2515, new_n12379);
and_5  g12003(new_n11472, new_n11471, new_n12380);
not_8  g12004(new_n11470, new_n12381);
nor_5  g12005(new_n11474, new_n12381, new_n12382);
or_5   g12006(new_n12382, new_n12380, new_n12383);
and_5  g12007(new_n11459, new_n11458, new_n12384);
nor_5  g12008(new_n11461, new_n11457, new_n12385);
nor_5  g12009(new_n12385, new_n12384, new_n12386);
xor_4  g12010(new_n12386, new_n12383, new_n12387);
xor_4  g12011(new_n12387, new_n12379, new_n12388);
xor_4  g12012(new_n12388, new_n12378, new_n12389);
and_5  g12013(n6441, n5314, new_n12390);
and_5  g12014(n11791, n5767, new_n12391_1);
xor_4  g12015(new_n12391_1, new_n12390, new_n12392);
and_5  g12016(new_n11468, new_n11466, new_n12393);
and_5  g12017(new_n11475, new_n11469, new_n12394);
nor_5  g12018(new_n12394, new_n12393, new_n12395);
and_5  g12019(n6687, n6604, new_n12396);
xor_4  g12020(new_n12396, new_n12395, new_n12397);
xor_4  g12021(new_n12397, new_n12392, new_n12398);
xor_4  g12022(new_n12398, new_n12389, new_n12399);
xor_4  g12023(new_n12399, new_n12373, new_n12400);
xor_4  g12024(new_n12400, new_n12363, new_n12401);
not_8  g12025(new_n11356, new_n12402);
nand_5 g12026(new_n11358, new_n12402, new_n12403);
not_8  g12027(new_n12403, new_n12404);
nor_5  g12028(new_n11360, new_n11354, new_n12405);
or_5   g12029(new_n12405, new_n12404, new_n12406);
or_5   g12030(new_n11339, new_n11331, new_n12407);
not_8  g12031(new_n11352, new_n12408);
nand_5 g12032(new_n12408, new_n11340, new_n12409);
and_5  g12033(new_n12409, new_n12407, new_n12410);
nand_5 g12034(n10678, n6429, new_n12411);
xor_4  g12035(new_n12411, new_n12410, new_n12412);
and_5  g12036(new_n11344, new_n11342, new_n12413);
and_5  g12037(new_n11351, new_n11345, new_n12414);
nor_5  g12038(new_n12414, new_n12413, new_n12415);
and_5  g12039(n2433, n2226, new_n12416);
nand_5 g12040(n8819, n1094, new_n12417);
and_5  g12041(n10928, n7730, new_n12418);
xor_4  g12042(new_n12418, new_n12417, new_n12419);
xor_4  g12043(new_n12419, new_n12416, new_n12420);
xor_4  g12044(new_n12420, new_n12415, new_n12421);
xor_4  g12045(new_n12421, new_n12412, new_n12422);
xor_4  g12046(new_n12422, new_n12406, new_n12423);
xor_4  g12047(new_n12423, new_n12401, new_n12424);
nor_5  g12048(new_n11481, new_n11480, new_n12425);
nor_5  g12049(new_n11483, new_n11478_1, new_n12426);
nor_5  g12050(new_n12426, new_n12425, new_n12427);
nor_5  g12051(new_n11282, new_n11251, new_n12428);
nor_5  g12052(new_n11291, new_n11283, new_n12429);
nor_5  g12053(new_n12429, new_n12428, new_n12430);
xor_4  g12054(new_n12430, new_n12427, new_n12431);
xor_4  g12055(new_n12431, new_n12424, new_n12432);
nor_5  g12056(new_n11485, new_n11452, new_n12433);
and_5  g12057(new_n11489, new_n11486, new_n12434);
nor_5  g12058(new_n12434, new_n12433, new_n12435);
and_5  g12059(new_n11361, new_n11328, new_n12436);
nor_5  g12060(new_n11362, new_n11326_1, new_n12437);
nor_5  g12061(new_n12437, new_n12436, new_n12438);
nand_5 g12062(new_n11261, new_n11256, new_n12439);
not_8  g12063(new_n11273, new_n12440);
nand_5 g12064(new_n12440, new_n11262, new_n12441);
nand_5 g12065(new_n12441, new_n12439, new_n12442);
nor_5  g12066(new_n11259, new_n11258, new_n12443);
and_5  g12067(new_n11259, new_n11258, new_n12444_1);
nor_5  g12068(new_n12444_1, new_n11257_1, new_n12445);
or_5   g12069(new_n12445, new_n12443, new_n12446);
nand_5 g12070(n12709, n7523, new_n12447);
and_5  g12071(n12000, n4189, new_n12448);
xor_4  g12072(new_n12448, new_n12447, new_n12449);
xor_4  g12073(new_n12449, new_n12446, new_n12450);
nand_5 g12074(n9725, n2564, new_n12451);
and_5  g12075(n9920, n4370, new_n12452);
xor_4  g12076(new_n12452, new_n12451, new_n12453);
and_5  g12077(n5212, n4516, new_n12454);
nand_5 g12078(n6770, n5320, new_n12455);
and_5  g12079(n5319, n1478, new_n12456);
xor_4  g12080(new_n12456, new_n12455, new_n12457);
xor_4  g12081(new_n12457, new_n12454, new_n12458);
xor_4  g12082(new_n12458, new_n12453, new_n12459);
and_5  g12083(n11728, n7320, new_n12460);
and_5  g12084(new_n11348, new_n11347, new_n12461);
not_8  g12085(new_n11346, new_n12462);
nor_5  g12086(new_n11350, new_n12462, new_n12463);
nor_5  g12087(new_n12463, new_n12461, new_n12464);
xor_4  g12088(new_n12464, new_n12460, new_n12465);
xor_4  g12089(new_n12465, new_n12459, new_n12466);
xor_4  g12090(new_n12466, new_n12450, new_n12467);
nor_5  g12091(new_n11270, new_n11269, new_n12468);
nand_5 g12092(n5212, n3627, new_n12469);
and_5  g12093(new_n11270, new_n11269, new_n12470);
nor_5  g12094(new_n12470, new_n12469, new_n12471);
nor_5  g12095(new_n12471, new_n12468, new_n12472);
nand_5 g12096(n10990, n4817, new_n12473);
and_5  g12097(n11877, n3627, new_n12474);
and_5  g12098(n8336, n1198, new_n12475);
xor_4  g12099(new_n12475, new_n12474, new_n12476);
xor_4  g12100(new_n12476, new_n12473, new_n12477);
xor_4  g12101(new_n12477, new_n12472, new_n12478);
and_5  g12102(new_n11266, new_n11264, new_n12479);
and_5  g12103(new_n11272, new_n11267, new_n12480);
or_5   g12104(new_n12480, new_n12479, new_n12481);
and_5  g12105(new_n11335, new_n11334, new_n12482);
nor_5  g12106(new_n11337, new_n11333, new_n12483);
nor_5  g12107(new_n12483, new_n12482, new_n12484);
xor_4  g12108(new_n12484, new_n12481, new_n12485);
xor_4  g12109(new_n12485, new_n12478, new_n12486);
xor_4  g12110(new_n12486, new_n12467, new_n12487);
xor_4  g12111(new_n12487, new_n12442, new_n12488);
xor_4  g12112(new_n12488, new_n12438, new_n12489_1);
xor_4  g12113(new_n12489_1, new_n12435, new_n12490);
xor_4  g12114(new_n12490, new_n12432, new_n12491);
xor_4  g12115(new_n12491, new_n12338, new_n12492);
xor_4  g12116(new_n12492, new_n12315, new_n12493);
xor_4  g12117(new_n12493, new_n12312, n8100);
xor_4  g12118(new_n9254, new_n9253, n8138);
xor_4  g12119(new_n5786, new_n5785, n8202);
xor_4  g12120(new_n3528, new_n3527, n8303);
xor_4  g12121(new_n2860, new_n2859, n8398);
xor_4  g12122(new_n4100, new_n4099, n9137);
xor_4  g12123(new_n6796, new_n6946, new_n12500);
xor_4  g12124(new_n6800, new_n12500, n9387);
xor_4  g12125(new_n10841, new_n10972, new_n12502);
xor_4  g12126(new_n10844, new_n12502, new_n12503);
xor_4  g12127(new_n11025, new_n12503, n9571);
not_8  g12128(new_n874, new_n12505);
xnor_4 g12129(new_n876, new_n12505, n9578);
xor_4  g12130(new_n1150, new_n1147, n9706);
or_5   g12131(new_n4102, new_n4098, new_n12508);
xor_4  g12132(new_n12508, new_n4094_1, n9756);
not_8  g12133(new_n6124, new_n12510);
nor_5  g12134(new_n6461, new_n12510, new_n12511_1);
and_5  g12135(new_n6461, new_n12510, new_n12512);
nor_5  g12136(new_n6481, new_n12512, new_n12513);
or_5   g12137(new_n12513, new_n12511_1, new_n12514);
nand_5 g12138(n12826, n7891, new_n12515);
and_5  g12139(new_n6200, new_n6198, new_n12516);
nor_5  g12140(new_n6202, new_n6195, new_n12517);
nor_5  g12141(new_n12517, new_n12516, new_n12518);
xor_4  g12142(new_n12518, new_n12515, new_n12519);
nor_5  g12143(new_n6437, new_n6221, new_n12520);
and_5  g12144(new_n6459, new_n6438, new_n12521);
or_5   g12145(new_n12521, new_n12520, new_n12522);
and_5  g12146(n8336, n2278, new_n12523);
nor_5  g12147(new_n6110, new_n6079, new_n12524);
nor_5  g12148(new_n6123, new_n6112, new_n12525);
nor_5  g12149(new_n12525, new_n12524, new_n12526);
xor_4  g12150(new_n12526, new_n12523, new_n12527);
nor_5  g12151(new_n6302, new_n6266, new_n12528);
nor_5  g12152(new_n6316, new_n6303, new_n12529);
or_5   g12153(new_n12529, new_n12528, new_n12530);
nor_5  g12154(new_n6093, new_n6092, new_n12531);
nor_5  g12155(new_n6100, new_n6095, new_n12532);
or_5   g12156(new_n12532, new_n12531, new_n12533);
or_5   g12157(new_n6180, new_n6172, new_n12534);
not_8  g12158(new_n6193, new_n12535);
nand_5 g12159(new_n12535, new_n6181, new_n12536);
nand_5 g12160(new_n12536, new_n12534, new_n12537);
and_5  g12161(n11662, n6770, new_n12538);
nand_5 g12162(n10451, n2226, new_n12539);
and_5  g12163(n5319, n3754, new_n12540);
xor_4  g12164(new_n12540, new_n12539, new_n12541);
xor_4  g12165(new_n12541, new_n12538, new_n12542);
and_5  g12166(new_n6189, new_n6188, new_n12543);
not_8  g12167(new_n6187, new_n12544);
nor_5  g12168(new_n6191, new_n12544, new_n12545);
nor_5  g12169(new_n12545, new_n12543, new_n12546);
xor_4  g12170(new_n12546, new_n12542, new_n12547);
nor_5  g12171(new_n6098, new_n6097, new_n12548);
and_5  g12172(new_n6098, new_n6097, new_n12549);
nor_5  g12173(new_n12549, new_n6096, new_n12550);
or_5   g12174(new_n12550, new_n12548, new_n12551);
and_5  g12175(n10278, n6986, new_n12552);
and_5  g12176(n10678, n3022, new_n12553);
xor_4  g12177(new_n12553, new_n12552, new_n12554);
xor_4  g12178(new_n12554, new_n12551, new_n12555);
xor_4  g12179(new_n12555, new_n12547, new_n12556);
and_5  g12180(new_n6185, new_n6183, new_n12557);
and_5  g12181(new_n6192_1, new_n6186, new_n12558);
nor_5  g12182(new_n12558, new_n12557, new_n12559);
and_5  g12183(new_n6176, new_n6175, new_n12560);
nor_5  g12184(new_n6178, new_n6174, new_n12561);
nor_5  g12185(new_n12561, new_n12560, new_n12562);
xor_4  g12186(new_n12562, new_n12559, new_n12563);
xor_4  g12187(new_n12563, new_n12556, new_n12564);
xor_4  g12188(new_n12564, new_n12537, new_n12565);
xor_4  g12189(new_n12565, new_n12533, new_n12566);
and_5  g12190(new_n6086, new_n6085, new_n12567);
nor_5  g12191(new_n6088, new_n6084, new_n12568);
or_5   g12192(new_n12568, new_n12567, new_n12569);
and_5  g12193(n8665, n2515, new_n12570);
nand_5 g12194(n10898, n9457, new_n12571);
and_5  g12195(n12511, n11222, new_n12572);
xor_4  g12196(new_n12572, new_n12571, new_n12573);
xor_4  g12197(new_n12573, new_n12570, new_n12574);
xor_4  g12198(new_n12574, new_n12569, new_n12575);
xor_4  g12199(new_n12575, new_n12566, new_n12576);
and_5  g12200(n12391, n4094, new_n12577);
nor_5  g12201(new_n6090, new_n6082, new_n12578);
nor_5  g12202(new_n6054, new_n6053, new_n12579);
xor_4  g12203(new_n6094, new_n12579, new_n12580);
xor_4  g12204(new_n6100, new_n12580, new_n12581);
and_5  g12205(new_n12581, new_n6091, new_n12582);
or_5   g12206(new_n12582, new_n12578, new_n12583);
nand_5 g12207(n4516, n3932, new_n12584);
and_5  g12208(n7523, n6703, new_n12585);
xor_4  g12209(new_n12585, new_n12584, new_n12586);
nand_5 g12210(n11423, n10928, new_n12587);
and_5  g12211(n12591, n3627, new_n12588);
xor_4  g12212(new_n12588, new_n12587, new_n12589);
xor_4  g12213(new_n12589, new_n12586, new_n12590);
xor_4  g12214(new_n12590, new_n12583, new_n12591_1);
nand_5 g12215(n11876, n4817, new_n12592);
nor_5  g12216(new_n6287, new_n6286, new_n12593);
nand_5 g12217(n2515, n1067, new_n12594);
and_5  g12218(new_n6287, new_n6286, new_n12595);
nor_5  g12219(new_n12595, new_n12594, new_n12596);
or_5   g12220(new_n12596, new_n12593, new_n12597);
nand_5 g12221(n10327, n4189, new_n12598);
and_5  g12222(n9920, n7456, new_n12599);
xor_4  g12223(new_n12599, new_n12598, new_n12600);
xor_4  g12224(new_n12600, new_n12597, new_n12601);
xor_4  g12225(new_n12601, new_n12592, new_n12602);
xor_4  g12226(new_n12602, new_n12591_1, new_n12603);
xor_4  g12227(new_n12603, new_n12577, new_n12604);
xor_4  g12228(new_n12604, new_n12576, new_n12605);
xor_4  g12229(new_n12605, new_n12530, new_n12606);
xor_4  g12230(new_n12606, new_n12527, new_n12607);
nor_5  g12231(new_n6106, new_n6105, new_n12608);
nor_5  g12232(new_n6108, new_n6103, new_n12609);
nor_5  g12233(new_n12609, new_n12608, new_n12610);
and_5  g12234(new_n6298, new_n6295, new_n12611);
nor_5  g12235(new_n6300, new_n6292, new_n12612);
nor_5  g12236(new_n12612, new_n12611, new_n12613);
xor_4  g12237(new_n12613, new_n12610, new_n12614);
and_5  g12238(new_n6371, new_n6368, new_n12615);
and_5  g12239(new_n6398, new_n6373, new_n12616);
or_5   g12240(new_n12616, new_n12615, new_n12617);
and_5  g12241(n11023, n1094, new_n12618);
xor_4  g12242(new_n12618, new_n12617, new_n12619);
nor_5  g12243(new_n6384, new_n6377, new_n12620);
and_5  g12244(new_n6397, new_n6385, new_n12621);
or_5   g12245(new_n12621, new_n12620, new_n12622);
and_5  g12246(new_n6283, new_n6281, new_n12623);
and_5  g12247(new_n6289, new_n6284, new_n12624);
nor_5  g12248(new_n12624, new_n12623, new_n12625);
and_5  g12249(new_n6381, new_n6380, new_n12626);
nor_5  g12250(new_n6383, new_n6379, new_n12627);
or_5   g12251(new_n12627, new_n12626, new_n12628);
and_5  g12252(new_n6393, new_n6392, new_n12629);
not_8  g12253(new_n6391, new_n12630);
nor_5  g12254(new_n6395, new_n12630, new_n12631);
nor_5  g12255(new_n12631, new_n12629, new_n12632);
xor_4  g12256(new_n12632, new_n12628, new_n12633);
nand_5 g12257(n12069, n10685, new_n12634);
and_5  g12258(n6578, n5645, new_n12635);
xor_4  g12259(new_n12635, new_n12634, new_n12636);
nand_5 g12260(n5767, n2749, new_n12637);
and_5  g12261(n996, n159, new_n12638);
and_5  g12262(n5314, n1510, new_n12639);
xor_4  g12263(new_n12639, new_n12638, new_n12640);
xor_4  g12264(new_n12640, new_n12637, new_n12641);
xor_4  g12265(new_n12641, new_n12636, new_n12642);
xor_4  g12266(new_n12642, new_n12633, new_n12643);
and_5  g12267(new_n6389, new_n6387, new_n12644);
and_5  g12268(new_n6396, new_n6390, new_n12645);
nor_5  g12269(new_n12645, new_n12644, new_n12646);
and_5  g12270(n7160, n2551, new_n12647);
nand_5 g12271(n9583, n2564, new_n12648_1);
and_5  g12272(n9640, n7320, new_n12649);
xor_4  g12273(new_n12649, new_n12648_1, new_n12650);
xor_4  g12274(new_n12650, new_n12647, new_n12651);
nand_5 g12275(n1199, n1067, new_n12652);
and_5  g12276(n12247, n11153, new_n12653);
xor_4  g12277(new_n12653, new_n12652, new_n12654);
xor_4  g12278(new_n12654, new_n12651, new_n12655);
xor_4  g12279(new_n12655, new_n12646, new_n12656);
xor_4  g12280(new_n12656, new_n12643, new_n12657);
xor_4  g12281(new_n12657, new_n12625, new_n12658);
nand_5 g12282(new_n6278, new_n6271, new_n12659);
not_8  g12283(new_n6290, new_n12660);
nand_5 g12284(new_n12660, new_n6279, new_n12661);
and_5  g12285(new_n12661, new_n12659, new_n12662);
and_5  g12286(new_n6275, new_n6274, new_n12663);
nor_5  g12287(new_n6277, new_n6273_1, new_n12664);
or_5   g12288(new_n12664, new_n12663, new_n12665);
and_5  g12289(n6687, n753, new_n12666);
and_5  g12290(n2087, n1798, new_n12667);
xor_4  g12291(new_n12667, new_n12666, new_n12668);
xor_4  g12292(new_n12668, new_n12665, new_n12669);
xor_4  g12293(new_n12669, new_n12662, new_n12670);
xor_4  g12294(new_n12670, new_n12658, new_n12671);
xor_4  g12295(new_n12671, new_n12622, new_n12672);
xor_4  g12296(new_n12672, new_n12619, new_n12673);
xor_4  g12297(new_n12673, new_n12614, new_n12674);
nor_5  g12298(new_n6400, new_n6364, new_n12675);
nor_5  g12299(new_n6415, new_n6401, new_n12676);
nor_5  g12300(new_n12676, new_n12675, new_n12677);
nor_5  g12301(new_n6204, new_n6168, new_n12678);
nor_5  g12302(new_n6219, new_n6205, new_n12679);
nor_5  g12303(new_n12679, new_n12678, new_n12680);
xor_4  g12304(new_n12680, new_n12677, new_n12681);
xor_4  g12305(new_n12681, new_n12674, new_n12682);
xor_4  g12306(new_n12682, new_n12607, new_n12683);
nand_5 g12307(n11922, n4828, new_n12684);
nor_5  g12308(new_n6435, new_n6416, new_n12685);
and_5  g12309(new_n6436, new_n6318, new_n12686);
nor_5  g12310(new_n12686, new_n12685, new_n12687);
xor_4  g12311(new_n12687, new_n12684, new_n12688);
xor_4  g12312(new_n12688, new_n12683, new_n12689);
xor_4  g12313(new_n12689, new_n12522, new_n12690);
xor_4  g12314(new_n12690, new_n12519, new_n12691);
xor_4  g12315(new_n12691, new_n12514, n9767);
xor_4  g12316(new_n2041, new_n2040, n9820);
xor_4  g12317(new_n9276, new_n9275, n9938);
not_8  g12318(new_n869, new_n12695);
xnor_4 g12319(new_n870, new_n12695, n10476);
xor_4  g12320(new_n866, new_n855, n10589);
xor_4  g12321(new_n1143, new_n1142, n10695);
xor_4  g12322(new_n3503, new_n3173, new_n12699);
xor_4  g12323(new_n12699, new_n3548, n10789);
xor_4  g12324(new_n2855, new_n2854, n10851);
not_8  g12325(new_n4844, new_n12702);
xor_4  g12326(new_n12702, new_n4834, n10913);
xor_4  g12327(new_n6949, new_n6806_1, n10949);
xor_4  g12328(new_n11027, new_n10981, n11216);
xor_4  g12329(new_n4836, new_n4835, n11326);
nor_5  g12330(new_n5361, new_n5141, new_n12707);
nor_5  g12331(new_n5495, new_n5362, new_n12708);
or_5   g12332(new_n12708, new_n12707, new_n12709_1);
not_8  g12333(new_n5402, new_n12710);
nor_5  g12334(new_n5406, new_n12710, new_n12711);
nor_5  g12335(new_n5494, new_n5407, new_n12712);
or_5   g12336(new_n12712, new_n12711, new_n12713);
nor_5  g12337(new_n5400, new_n5367, new_n12714);
and_5  g12338(new_n5401, new_n5366, new_n12715);
or_5   g12339(new_n12715, new_n12714, new_n12716);
and_5  g12340(new_n5396, new_n5393, new_n12717);
nor_5  g12341(new_n5398, new_n5390, new_n12718);
nor_5  g12342(new_n12718, new_n12717, new_n12719);
nand_5 g12343(n9763, n45, new_n12720_1);
and_5  g12344(n8759, n7823, new_n12721);
xor_4  g12345(new_n12721, new_n12720_1, new_n12722);
xor_4  g12346(new_n12722, new_n12719, new_n12723);
and_5  g12347(new_n5115, new_n5114, new_n12724);
not_8  g12348(new_n5113, new_n12725);
nor_5  g12349(new_n5117, new_n12725, new_n12726);
nor_5  g12350(new_n12726, new_n12724, new_n12727);
and_5  g12351(n9241, n9189, new_n12728);
xor_4  g12352(new_n12728, new_n12727, new_n12729);
and_5  g12353(n12705, n4634, new_n12730);
and_5  g12354(n12145, n7436, new_n12731);
xor_4  g12355(new_n12731, new_n12730, new_n12732);
and_5  g12356(n9195, n4312, new_n12733);
and_5  g12357(n10217, n6776, new_n12734);
xor_4  g12358(new_n12734, new_n12733, new_n12735);
xor_4  g12359(new_n12735, new_n12732, new_n12736);
xor_4  g12360(new_n12736, new_n12729, new_n12737);
and_5  g12361(new_n5381, new_n5379, new_n12738);
and_5  g12362(new_n5387, new_n5382, new_n12739);
nor_5  g12363(new_n12739, new_n12738, new_n12740);
and_5  g12364(new_n5372, new_n5371, new_n12741);
nor_5  g12365(new_n5374, new_n5370, new_n12742);
nor_5  g12366(new_n12742, new_n12741, new_n12743);
xor_4  g12367(new_n12743, new_n12740, new_n12744);
xor_4  g12368(new_n12744, new_n12737, new_n12745);
nor_5  g12369(new_n5385, new_n5384, new_n12746);
nand_5 g12370(n9241, n2024, new_n12747);
and_5  g12371(new_n5385, new_n5384, new_n12748);
nor_5  g12372(new_n12748, new_n12747, new_n12749);
nor_5  g12373(new_n12749, new_n12746, new_n12750);
xor_4  g12374(new_n12750, new_n12745, new_n12751);
nand_5 g12375(n3986, n3342, new_n12752);
nand_5 g12376(n8276, n2522, new_n12753_1);
and_5  g12377(n12299, n12221, new_n12754);
xor_4  g12378(new_n12754, new_n12753_1, new_n12755);
xor_4  g12379(new_n12755, new_n12752, new_n12756);
xor_4  g12380(new_n12756, new_n12751, new_n12757);
or_5   g12381(new_n5376, new_n5368, new_n12758);
not_8  g12382(new_n5388, new_n12759);
nand_5 g12383(new_n12759, new_n5377, new_n12760);
and_5  g12384(new_n12760, new_n12758, new_n12761);
not_8  g12385(new_n5478, new_n12762);
nand_5 g12386(new_n5481, new_n12762, new_n12763);
or_5   g12387(new_n5483, new_n5476, new_n12764);
and_5  g12388(new_n12764, new_n12763, new_n12765);
xor_4  g12389(new_n12765, new_n12761, new_n12766);
xor_4  g12390(new_n12766, new_n12757, new_n12767);
xor_4  g12391(new_n12767, new_n12723, new_n12768);
xor_4  g12392(new_n12768, new_n12716, new_n12769);
and_5  g12393(n12025, n10223, new_n12770);
and_5  g12394(new_n5111, new_n5109, new_n12771);
and_5  g12395(new_n5118, new_n5112, new_n12772);
nor_5  g12396(new_n12772, new_n12771, new_n12773);
xor_4  g12397(new_n12773, new_n12770, new_n12774);
xor_4  g12398(new_n12774, new_n12769, new_n12775);
or_5   g12399(new_n5461, new_n5453, new_n12776);
not_8  g12400(new_n5474, new_n12777_1);
nand_5 g12401(new_n12777_1, new_n5462, new_n12778);
nand_5 g12402(new_n12778, new_n12776, new_n12779);
nand_5 g12403(n7690, n5579, new_n12780);
and_5  g12404(n7388, n2507, new_n12781);
xor_4  g12405(new_n12781, new_n12780, new_n12782);
nand_5 g12406(n7270, n2393, new_n12783);
and_5  g12407(n5331, n1576, new_n12784);
xor_4  g12408(new_n12784, new_n12783, new_n12785);
xor_4  g12409(new_n12785, new_n12782, new_n12786);
nand_5 g12410(n3616, n2498, new_n12787);
and_5  g12411(n12648, n6016, new_n12788);
xor_4  g12412(new_n12788, new_n12787, new_n12789);
xor_4  g12413(new_n12789, new_n12786, new_n12790);
and_5  g12414(n5798, n2530, new_n12791);
and_5  g12415(n10644, n7946, new_n12792);
xor_4  g12416(new_n12792, new_n12791, new_n12793);
and_5  g12417(new_n5457, new_n5456, new_n12794);
nor_5  g12418(new_n5459, new_n5455, new_n12795);
nor_5  g12419(new_n12795, new_n12794, new_n12796);
and_5  g12420(new_n5102, new_n5101, new_n12797);
nor_5  g12421(new_n5104, new_n5100, new_n12798);
nor_5  g12422(new_n12798, new_n12797, new_n12799);
xor_4  g12423(new_n12799, new_n12796, new_n12800);
xor_4  g12424(new_n12800, new_n12793, new_n12801);
xor_4  g12425(new_n12801, new_n12790, new_n12802);
xor_4  g12426(new_n12802, new_n12779, new_n12803);
not_8  g12427(new_n5436, new_n12804);
nand_5 g12428(new_n5438, new_n12804, new_n12805);
or_5   g12429(new_n5440, new_n5434, new_n12806);
nand_5 g12430(new_n12806, new_n12805, new_n12807_1);
and_5  g12431(new_n5470, new_n5469, new_n12808);
not_8  g12432(new_n5468, new_n12809);
nor_5  g12433(new_n5472, new_n12809, new_n12810);
or_5   g12434(new_n12810, new_n12808, new_n12811);
and_5  g12435(new_n5466, new_n5464, new_n12812);
and_5  g12436(new_n5473, new_n5467, new_n12813);
or_5   g12437(new_n12813, new_n12812, new_n12814);
nand_5 g12438(n7965, n6431, new_n12815);
and_5  g12439(n9111, n5857, new_n12816);
xor_4  g12440(new_n12816, new_n12815, new_n12817);
and_5  g12441(n11892, n5153, new_n12818);
and_5  g12442(n5860, n806, new_n12819);
xor_4  g12443(new_n12819, new_n12818, new_n12820);
and_5  g12444(n10545, n521, new_n12821);
and_5  g12445(n10547, n7265, new_n12822);
xor_4  g12446(new_n12822, new_n12821, new_n12823);
xor_4  g12447(new_n12823, new_n12820, new_n12824);
xor_4  g12448(new_n12824, new_n12817, new_n12825);
xor_4  g12449(new_n12825, new_n12814, new_n12826_1);
xor_4  g12450(new_n12826_1, new_n12811, new_n12827);
xor_4  g12451(new_n12827, new_n12807_1, new_n12828);
or_5   g12452(new_n5106, new_n5098, new_n12829);
not_8  g12453(new_n5119, new_n12830);
nand_5 g12454(new_n12830, new_n5107, new_n12831);
and_5  g12455(new_n12831, new_n12829, new_n12832);
and_5  g12456(new_n5424, new_n5422, new_n12833);
and_5  g12457(new_n5431, new_n5425, new_n12834);
nor_5  g12458(new_n12834, new_n12833, new_n12835);
xor_4  g12459(new_n12835, new_n12832, new_n12836);
xor_4  g12460(new_n12836, new_n12828, new_n12837);
xor_4  g12461(new_n12837, new_n12803, new_n12838);
and_5  g12462(new_n5441, new_n5409, new_n12839);
nor_5  g12463(new_n5446, new_n5443, new_n12840);
nor_5  g12464(new_n12840, new_n12839, new_n12841);
nor_5  g12465(new_n5124, new_n5123, new_n12842);
nor_5  g12466(new_n5126, new_n5121, new_n12843);
or_5   g12467(new_n12843, new_n12842, new_n12844);
or_5   g12468(new_n5419, new_n5416, new_n12845);
not_8  g12469(new_n5432, new_n12846);
nand_5 g12470(new_n12846, new_n5420, new_n12847);
nand_5 g12471(new_n12847, new_n12845, new_n12848);
and_5  g12472(new_n5428, new_n5427, new_n12849);
not_8  g12473(new_n5426, new_n12850);
nor_5  g12474(new_n5430, new_n12850, new_n12851);
or_5   g12475(new_n12851, new_n12849, new_n12852);
nand_5 g12476(n4499, n2558, new_n12853);
and_5  g12477(n5305, n2512, new_n12854);
xor_4  g12478(new_n12854, new_n12853, new_n12855);
xor_4  g12479(new_n12855, new_n12852, new_n12856);
and_5  g12480(new_n5414, new_n5410, new_n12857);
or_5   g12481(new_n12857, new_n5411_1, new_n12858);
not_8  g12482(new_n12858, new_n12859);
and_5  g12483(n8476, n2347, new_n12860);
and_5  g12484(new_n12860, new_n12859, new_n12861);
and_5  g12485(new_n12860, new_n5273, new_n12862);
nor_5  g12486(new_n12862, new_n12859, new_n12863);
or_5   g12487(new_n12863, new_n12861, new_n12864);
and_5  g12488(n2253, n1097, new_n12865);
and_5  g12489(n5964, n3865, new_n12866);
xor_4  g12490(new_n12866, new_n12865, new_n12867);
xor_4  g12491(new_n12867, new_n12864, new_n12868);
xor_4  g12492(new_n12868, new_n12856, new_n12869);
xor_4  g12493(new_n12869, new_n12848, new_n12870);
nand_5 g12494(n10510, n2024, new_n12871);
and_5  g12495(n11257, n2879, new_n12872);
xor_4  g12496(new_n12872, new_n12871, new_n12873);
xor_4  g12497(new_n12873, new_n12870, new_n12874);
xor_4  g12498(new_n12874, new_n12844, new_n12875);
xor_4  g12499(new_n12875, new_n12841, new_n12876);
xor_4  g12500(new_n12876, new_n12838, new_n12877);
xor_4  g12501(new_n12877, new_n12775, new_n12878);
xor_4  g12502(new_n5488, new_n5485, new_n12879);
and_5  g12503(new_n12879, new_n5448, new_n12880);
nor_5  g12504(new_n5493, new_n5490, new_n12881);
nor_5  g12505(new_n12881, new_n12880, new_n12882);
nor_5  g12506(new_n5128, new_n5097, new_n12883);
and_5  g12507(new_n5140, new_n5129, new_n12884);
nor_5  g12508(new_n12884, new_n12883, new_n12885);
and_5  g12509(new_n5484, new_n5450, new_n12886);
nor_5  g12510(new_n5488, new_n5486, new_n12887);
nor_5  g12511(new_n12887, new_n12886, new_n12888);
xor_4  g12512(new_n12888, new_n12885, new_n12889);
xor_4  g12513(new_n12889, new_n12882, new_n12890);
xor_4  g12514(new_n12890, new_n12878, new_n12891);
xor_4  g12515(new_n12891, new_n12713, new_n12892);
xor_4  g12516(new_n12892, new_n12709_1, n11707);
xor_4  g12517(new_n5984, new_n5983, n11755);
xor_4  g12518(new_n3540, new_n3539, n11780);
not_8  g12519(new_n9642, new_n12896);
xor_4  g12520(new_n9644, new_n12896, n11919);
xor_4  g12521(new_n9646, new_n9629, n12005);
not_8  g12522(new_n10073, new_n12899);
xor_4  g12523(new_n12899, new_n10069, n12014);
not_8  g12524(new_n8458, new_n12901);
xnor_4 g12525(new_n12901, new_n8430, n12020);
nor_5  g12526(new_n11018, new_n10992, new_n12903);
xor_4  g12527(new_n12903, new_n10989, n12076);
xnor_4 g12528(new_n11548, new_n11546, n12111);
nor_5  g12529(new_n10074, new_n10068, new_n12906);
xor_4  g12530(new_n12906, new_n10063, n12444);
nor_5  g12531(new_n5359, new_n5347, new_n12908);
or_5   g12532(new_n12908, new_n5360, n12807);
endmodule


