// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Thu Jun 27 03:00:32 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1, new_n993,
    new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067_1,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094_1, new_n1095, new_n1096, new_n1097_1,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198_1, new_n1199_1, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209_1, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269_1, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333_1, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355, new_n1356,
    new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471_1, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1781, new_n1782,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1794,
    new_n1795, new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1807, new_n1808, new_n1809, new_n1810, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1816, new_n1817, new_n1818,
    new_n1819, new_n1820, new_n1821, new_n1822, new_n1823, new_n1824,
    new_n1825, new_n1826, new_n1827, new_n1828, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848,
    new_n1849, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1,
    new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389,
    new_n2390, new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1,
    new_n2432, new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2479,
    new_n2480, new_n2481, new_n2482, new_n2483, new_n2484, new_n2485,
    new_n2486, new_n2487, new_n2488, new_n2489, new_n2490, new_n2491,
    new_n2492, new_n2493, new_n2494, new_n2495, new_n2496, new_n2497,
    new_n2498_1, new_n2499, new_n2500, new_n2501, new_n2502, new_n2503,
    new_n2504, new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1,
    new_n2510, new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1,
    new_n2516, new_n2517, new_n2518, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3017, new_n3018, new_n3019, new_n3020, new_n3021,
    new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026, new_n3027,
    new_n3028, new_n3029, new_n3030, new_n3031, new_n3032, new_n3033,
    new_n3034, new_n3035, new_n3036, new_n3037, new_n3038, new_n3039,
    new_n3040, new_n3041, new_n3042, new_n3043, new_n3044, new_n3045,
    new_n3046, new_n3047, new_n3048, new_n3049, new_n3050, new_n3051,
    new_n3052, new_n3053, new_n3054, new_n3055, new_n3056, new_n3057,
    new_n3058, new_n3059, new_n3060, new_n3061, new_n3062, new_n3063,
    new_n3064, new_n3065, new_n3066, new_n3067, new_n3068, new_n3069,
    new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074, new_n3075,
    new_n3076, new_n3077, new_n3078, new_n3079, new_n3080, new_n3081,
    new_n3082, new_n3083, new_n3084, new_n3085, new_n3086, new_n3087,
    new_n3088, new_n3089, new_n3090, new_n3091, new_n3092, new_n3093,
    new_n3094, new_n3095, new_n3096, new_n3097, new_n3098, new_n3099,
    new_n3100, new_n3101, new_n3102, new_n3103, new_n3104, new_n3105,
    new_n3106, new_n3107, new_n3108, new_n3109, new_n3110, new_n3111,
    new_n3112, new_n3113, new_n3114, new_n3115, new_n3116, new_n3117,
    new_n3118, new_n3119, new_n3120, new_n3121, new_n3122, new_n3123,
    new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128, new_n3129,
    new_n3130, new_n3131, new_n3132, new_n3133, new_n3134, new_n3135,
    new_n3136, new_n3137, new_n3138, new_n3139, new_n3140, new_n3141,
    new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1, new_n3147,
    new_n3148, new_n3149, new_n3150, new_n3151, new_n3152, new_n3153,
    new_n3154, new_n3155, new_n3156, new_n3157, new_n3158, new_n3159,
    new_n3160, new_n3161, new_n3162, new_n3163, new_n3165, new_n3166,
    new_n3167, new_n3168, new_n3169, new_n3170, new_n3171, new_n3172_1,
    new_n3173, new_n3174, new_n3175, new_n3176, new_n3177, new_n3178,
    new_n3179, new_n3180, new_n3181, new_n3182, new_n3183, new_n3184,
    new_n3185, new_n3186, new_n3187, new_n3188, new_n3189, new_n3190,
    new_n3191, new_n3192, new_n3193, new_n3194, new_n3195, new_n3196,
    new_n3197, new_n3198, new_n3199, new_n3200, new_n3201, new_n3202,
    new_n3203, new_n3204, new_n3205, new_n3206, new_n3207, new_n3208,
    new_n3209, new_n3210, new_n3211, new_n3212, new_n3213, new_n3214_1,
    new_n3215, new_n3216, new_n3217, new_n3218, new_n3219, new_n3220,
    new_n3221, new_n3222, new_n3223, new_n3224, new_n3225, new_n3226,
    new_n3227, new_n3228, new_n3229, new_n3230_1, new_n3231, new_n3232,
    new_n3233, new_n3234, new_n3235, new_n3236, new_n3237, new_n3238,
    new_n3239, new_n3240, new_n3241, new_n3242, new_n3243, new_n3244,
    new_n3245, new_n3246, new_n3247, new_n3248, new_n3249, new_n3250,
    new_n3251, new_n3252, new_n3253, new_n3254, new_n3255, new_n3256,
    new_n3257, new_n3258, new_n3259, new_n3260, new_n3261, new_n3262,
    new_n3263, new_n3264, new_n3265, new_n3266, new_n3267, new_n3268,
    new_n3269, new_n3270, new_n3271, new_n3272_1, new_n3273, new_n3274,
    new_n3275, new_n3276, new_n3277, new_n3278, new_n3279, new_n3280,
    new_n3281, new_n3282, new_n3283, new_n3284, new_n3285, new_n3286,
    new_n3287_1, new_n3288, new_n3289, new_n3290, new_n3291, new_n3292,
    new_n3293, new_n3294, new_n3295, new_n3296, new_n3297, new_n3298,
    new_n3299, new_n3300, new_n3301, new_n3302, new_n3303, new_n3304,
    new_n3305, new_n3306, new_n3307, new_n3308, new_n3309, new_n3310,
    new_n3311, new_n3312, new_n3313, new_n3314, new_n3315, new_n3316,
    new_n3317, new_n3318, new_n3319, new_n3320, new_n3321, new_n3322,
    new_n3323, new_n3324, new_n3325, new_n3326, new_n3327, new_n3328,
    new_n3329, new_n3330, new_n3331, new_n3332, new_n3333, new_n3334,
    new_n3335, new_n3336, new_n3337, new_n3338, new_n3339_1, new_n3340,
    new_n3341, new_n3342_1, new_n3343, new_n3344, new_n3345, new_n3346,
    new_n3347, new_n3348, new_n3349, new_n3350, new_n3351, new_n3352,
    new_n3353, new_n3354, new_n3355, new_n3356, new_n3357, new_n3358,
    new_n3359, new_n3360, new_n3361, new_n3362, new_n3363, new_n3364,
    new_n3365, new_n3366, new_n3367, new_n3368, new_n3369, new_n3370,
    new_n3371, new_n3372, new_n3373, new_n3374, new_n3375, new_n3376,
    new_n3377, new_n3378, new_n3379, new_n3380, new_n3381, new_n3382,
    new_n3383, new_n3384, new_n3385, new_n3386, new_n3387, new_n3388,
    new_n3389, new_n3390, new_n3391, new_n3392, new_n3393, new_n3394,
    new_n3395, new_n3396, new_n3397, new_n3398, new_n3399, new_n3400,
    new_n3401, new_n3402, new_n3403, new_n3404, new_n3405, new_n3406,
    new_n3407, new_n3408, new_n3410, new_n3411, new_n3412, new_n3413,
    new_n3414, new_n3415, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627_1, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758,
    new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782,
    new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794,
    new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849_1, new_n3850, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866,
    new_n3867, new_n3868, new_n3869, new_n3870, new_n3871, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878,
    new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884,
    new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909, new_n3910, new_n3911, new_n3912, new_n3913, new_n3914,
    new_n3915, new_n3916, new_n3917, new_n3918, new_n3919, new_n3920,
    new_n3921, new_n3922, new_n3923, new_n3924, new_n3925, new_n3926,
    new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1,
    new_n3933, new_n3934, new_n3935, new_n3936, new_n3937, new_n3938,
    new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944,
    new_n3945, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950,
    new_n3951, new_n3952, new_n3953, new_n3954, new_n3955, new_n3956,
    new_n3957, new_n3958, new_n3959, new_n3960, new_n3961, new_n3962,
    new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968,
    new_n3969, new_n3970, new_n3971, new_n3972, new_n3973, new_n3974,
    new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980,
    new_n3981, new_n3982, new_n3983, new_n3984, new_n3985, new_n3986_1,
    new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3992_1,
    new_n3993, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998,
    new_n3999, new_n4000, new_n4001, new_n4002, new_n4003, new_n4004,
    new_n4005_1, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010,
    new_n4011, new_n4012, new_n4013, new_n4014, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034,
    new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040,
    new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046,
    new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052,
    new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058,
    new_n4059, new_n4060, new_n4061, new_n4062, new_n4063, new_n4064,
    new_n4065, new_n4066, new_n4067, new_n4068, new_n4069, new_n4070,
    new_n4071, new_n4072, new_n4073, new_n4074, new_n4075, new_n4076,
    new_n4077, new_n4078, new_n4079, new_n4080, new_n4081, new_n4082,
    new_n4083, new_n4084, new_n4085, new_n4086_1, new_n4087, new_n4088_1,
    new_n4089, new_n4090, new_n4091, new_n4093, new_n4094_1, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101,
    new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4120, new_n4121, new_n4122, new_n4123, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143,
    new_n4144, new_n4145, new_n4146, new_n4147, new_n4148, new_n4149,
    new_n4150, new_n4151, new_n4152, new_n4153, new_n4154, new_n4155_1,
    new_n4156, new_n4157, new_n4158, new_n4159_1, new_n4160, new_n4161,
    new_n4162, new_n4163, new_n4164, new_n4165, new_n4166, new_n4167,
    new_n4168, new_n4169, new_n4170, new_n4171, new_n4172, new_n4173,
    new_n4174, new_n4175, new_n4176, new_n4177, new_n4178, new_n4179,
    new_n4180, new_n4181, new_n4182, new_n4183, new_n4184, new_n4185,
    new_n4186, new_n4187_1, new_n4188, new_n4189_1, new_n4190_1, new_n4191,
    new_n4192, new_n4193, new_n4194, new_n4195, new_n4196, new_n4197,
    new_n4198, new_n4199, new_n4200, new_n4201, new_n4202, new_n4203_1,
    new_n4204, new_n4205, new_n4206, new_n4207, new_n4208, new_n4209,
    new_n4210, new_n4211, new_n4212, new_n4213, new_n4214, new_n4215,
    new_n4216, new_n4217, new_n4218, new_n4219, new_n4220, new_n4221,
    new_n4222, new_n4223, new_n4224, new_n4225, new_n4226_1, new_n4227,
    new_n4228, new_n4229, new_n4230_1, new_n4231, new_n4232, new_n4233,
    new_n4234, new_n4235, new_n4236, new_n4237, new_n4238, new_n4239,
    new_n4240, new_n4241, new_n4242, new_n4243, new_n4244, new_n4245,
    new_n4246, new_n4247, new_n4248, new_n4249, new_n4250, new_n4251,
    new_n4252, new_n4253, new_n4254, new_n4255, new_n4256, new_n4257,
    new_n4258, new_n4259, new_n4260, new_n4261, new_n4262, new_n4263,
    new_n4264, new_n4265, new_n4266, new_n4267, new_n4268, new_n4269,
    new_n4270, new_n4271, new_n4272, new_n4273, new_n4274, new_n4275,
    new_n4276, new_n4277, new_n4278, new_n4279, new_n4280, new_n4281,
    new_n4282, new_n4283, new_n4284, new_n4285, new_n4286, new_n4287,
    new_n4288, new_n4289, new_n4290, new_n4291, new_n4292, new_n4293,
    new_n4294, new_n4295, new_n4296, new_n4297, new_n4298, new_n4299,
    new_n4300_1, new_n4301, new_n4302, new_n4303, new_n4304, new_n4305,
    new_n4306, new_n4307, new_n4308, new_n4309, new_n4310, new_n4311,
    new_n4312_1, new_n4313, new_n4314, new_n4315, new_n4316, new_n4317,
    new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4324, new_n4325, new_n4326_1, new_n4327, new_n4328, new_n4329,
    new_n4330, new_n4331, new_n4332, new_n4333_1, new_n4334, new_n4335,
    new_n4336, new_n4337, new_n4338, new_n4339, new_n4340, new_n4341,
    new_n4342, new_n4343, new_n4344, new_n4345, new_n4346, new_n4347,
    new_n4348, new_n4349, new_n4350, new_n4351, new_n4352, new_n4353,
    new_n4354, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359,
    new_n4360, new_n4361, new_n4362, new_n4363, new_n4364, new_n4365,
    new_n4366, new_n4367, new_n4368, new_n4369, new_n4370_1, new_n4371,
    new_n4372, new_n4373, new_n4374, new_n4375, new_n4376, new_n4377,
    new_n4378_1, new_n4379, new_n4380, new_n4381, new_n4382, new_n4383,
    new_n4384, new_n4385, new_n4386, new_n4387, new_n4388, new_n4389,
    new_n4390, new_n4391, new_n4392, new_n4393, new_n4394, new_n4395,
    new_n4396, new_n4397_1, new_n4398, new_n4399, new_n4400, new_n4401,
    new_n4402, new_n4403, new_n4404, new_n4405, new_n4406, new_n4407,
    new_n4408, new_n4409, new_n4410, new_n4411, new_n4412, new_n4413,
    new_n4414, new_n4415, new_n4416, new_n4417, new_n4418, new_n4419,
    new_n4420, new_n4421, new_n4422, new_n4423, new_n4424, new_n4425,
    new_n4426, new_n4427, new_n4428, new_n4429, new_n4430, new_n4431,
    new_n4432, new_n4433, new_n4434, new_n4435, new_n4436_1, new_n4437,
    new_n4439, new_n4440, new_n4441, new_n4442, new_n4443, new_n4444,
    new_n4445, new_n4446, new_n4447, new_n4448, new_n4449, new_n4450,
    new_n4451, new_n4452, new_n4453, new_n4454, new_n4455, new_n4456,
    new_n4457, new_n4458, new_n4459, new_n4460, new_n4461, new_n4462,
    new_n4463, new_n4464, new_n4465, new_n4466, new_n4467, new_n4468,
    new_n4469, new_n4470, new_n4471, new_n4472, new_n4473, new_n4474,
    new_n4475, new_n4476, new_n4477, new_n4478, new_n4479, new_n4480,
    new_n4481, new_n4482, new_n4483, new_n4484, new_n4485, new_n4486,
    new_n4487, new_n4488, new_n4489, new_n4490, new_n4491, new_n4492,
    new_n4493, new_n4494, new_n4495, new_n4496, new_n4497, new_n4498,
    new_n4499_1, new_n4500, new_n4501, new_n4502, new_n4503, new_n4504,
    new_n4505, new_n4506, new_n4507, new_n4508, new_n4509, new_n4510,
    new_n4511, new_n4512, new_n4513, new_n4514, new_n4515, new_n4516_1,
    new_n4517, new_n4518, new_n4519, new_n4520, new_n4521, new_n4522,
    new_n4523, new_n4524, new_n4525, new_n4526, new_n4527, new_n4528,
    new_n4529, new_n4530, new_n4531, new_n4532, new_n4533, new_n4534,
    new_n4535, new_n4536, new_n4537, new_n4538, new_n4539, new_n4540,
    new_n4541, new_n4542, new_n4543, new_n4544, new_n4545, new_n4546,
    new_n4547, new_n4548, new_n4549, new_n4550, new_n4551, new_n4552,
    new_n4553_1, new_n4554, new_n4555, new_n4556, new_n4557, new_n4558,
    new_n4559, new_n4560, new_n4561, new_n4562, new_n4563, new_n4564,
    new_n4565, new_n4566, new_n4567, new_n4568, new_n4569, new_n4570,
    new_n4571, new_n4572, new_n4573, new_n4574, new_n4575, new_n4576,
    new_n4577, new_n4578, new_n4579, new_n4580, new_n4581, new_n4582,
    new_n4583, new_n4584, new_n4585, new_n4586, new_n4587, new_n4588,
    new_n4589, new_n4590, new_n4591, new_n4592, new_n4593, new_n4594,
    new_n4595, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618,
    new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624,
    new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630,
    new_n4631, new_n4632, new_n4633, new_n4634_1, new_n4635, new_n4636,
    new_n4637, new_n4638, new_n4639, new_n4640, new_n4641, new_n4642,
    new_n4643, new_n4644, new_n4645, new_n4646, new_n4647, new_n4648,
    new_n4649, new_n4650, new_n4651, new_n4652, new_n4653, new_n4654,
    new_n4655, new_n4656, new_n4657, new_n4658, new_n4659, new_n4660,
    new_n4661, new_n4662, new_n4663, new_n4664, new_n4665, new_n4666,
    new_n4667, new_n4668, new_n4669, new_n4670, new_n4671, new_n4672,
    new_n4673, new_n4674, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686_1, new_n4687, new_n4688, new_n4689_1, new_n4690, new_n4691,
    new_n4692, new_n4693, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703,
    new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709,
    new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715,
    new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721,
    new_n4722_1, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727,
    new_n4728, new_n4729, new_n4730, new_n4731, new_n4732, new_n4733_1,
    new_n4734, new_n4735, new_n4736, new_n4737, new_n4738, new_n4739,
    new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745,
    new_n4746, new_n4747, new_n4748, new_n4749, new_n4750, new_n4751,
    new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757_1,
    new_n4758, new_n4759, new_n4760, new_n4761, new_n4762, new_n4763,
    new_n4764, new_n4765, new_n4766, new_n4767, new_n4768, new_n4769,
    new_n4770, new_n4771, new_n4772, new_n4773, new_n4774, new_n4775,
    new_n4776, new_n4777, new_n4778, new_n4779, new_n4780, new_n4781,
    new_n4782, new_n4783, new_n4784, new_n4785, new_n4786, new_n4787,
    new_n4788, new_n4789, new_n4790, new_n4791, new_n4792, new_n4793,
    new_n4794, new_n4795, new_n4796, new_n4797, new_n4798, new_n4799,
    new_n4800, new_n4801, new_n4802, new_n4803, new_n4804, new_n4805_1,
    new_n4806, new_n4807, new_n4808, new_n4809, new_n4810, new_n4811,
    new_n4812, new_n4813, new_n4814, new_n4815, new_n4816, new_n4817_1,
    new_n4818, new_n4819, new_n4820, new_n4821, new_n4822, new_n4823,
    new_n4825, new_n4826_1, new_n4827, new_n4828_1, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1,
    new_n4971_1, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000,
    new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012,
    new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018,
    new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024,
    new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1,
    new_n5031, new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048,
    new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054,
    new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060,
    new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066,
    new_n5067, new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072,
    new_n5073, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078,
    new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084,
    new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090,
    new_n5091, new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114,
    new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120,
    new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126,
    new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1,
    new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144,
    new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150,
    new_n5151, new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156,
    new_n5157, new_n5158, new_n5159, new_n5160, new_n5161, new_n5162,
    new_n5163, new_n5164, new_n5165, new_n5166, new_n5167, new_n5168,
    new_n5169, new_n5170, new_n5171, new_n5172, new_n5173, new_n5174,
    new_n5175, new_n5176, new_n5177, new_n5178, new_n5179, new_n5180,
    new_n5181, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186,
    new_n5187, new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192,
    new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1,
    new_n5199, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212_1,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314_1,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1, new_n5320_1,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643, new_n5644,
    new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5730, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859, new_n5860_1,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934_1, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6005, new_n6006, new_n6007, new_n6008, new_n6009, new_n6010,
    new_n6011, new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1,
    new_n6017, new_n6018, new_n6019, new_n6020, new_n6021, new_n6022,
    new_n6023, new_n6024, new_n6025, new_n6026, new_n6027, new_n6028,
    new_n6029, new_n6030, new_n6031, new_n6032, new_n6033, new_n6034,
    new_n6035, new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040,
    new_n6041, new_n6042, new_n6043, new_n6044, new_n6045, new_n6046,
    new_n6047, new_n6048, new_n6049, new_n6050, new_n6051, new_n6052,
    new_n6053, new_n6054, new_n6055, new_n6056, new_n6057, new_n6058,
    new_n6059, new_n6060, new_n6061, new_n6062, new_n6063, new_n6064,
    new_n6065, new_n6066, new_n6067, new_n6068, new_n6069, new_n6070,
    new_n6071, new_n6072, new_n6073, new_n6074, new_n6075, new_n6076,
    new_n6077, new_n6078, new_n6079, new_n6080, new_n6081, new_n6082,
    new_n6083, new_n6084, new_n6085, new_n6086, new_n6087, new_n6088,
    new_n6089_1, new_n6090, new_n6091, new_n6092, new_n6093, new_n6094,
    new_n6095, new_n6096, new_n6097, new_n6098, new_n6099, new_n6100,
    new_n6101, new_n6102, new_n6103, new_n6104, new_n6105, new_n6106,
    new_n6107, new_n6108, new_n6109, new_n6110, new_n6111, new_n6112,
    new_n6113, new_n6114, new_n6115, new_n6116, new_n6117, new_n6118,
    new_n6119, new_n6120, new_n6121, new_n6122, new_n6123, new_n6124,
    new_n6125, new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130,
    new_n6131, new_n6132, new_n6133, new_n6134, new_n6135, new_n6136,
    new_n6137, new_n6138, new_n6139, new_n6140, new_n6141, new_n6142,
    new_n6143, new_n6144, new_n6145, new_n6146, new_n6147, new_n6148,
    new_n6149, new_n6150, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254_1, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273_1, new_n6274, new_n6278,
    new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6286,
    new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292,
    new_n6293, new_n6294_1, new_n6295, new_n6296, new_n6297, new_n6298,
    new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304,
    new_n6305, new_n6306, new_n6307, new_n6308, new_n6309, new_n6310,
    new_n6311, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316,
    new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322,
    new_n6323, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328,
    new_n6329, new_n6330, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354, new_n6355, new_n6356, new_n6357, new_n6358_1,
    new_n6359_1, new_n6360, new_n6364, new_n6365, new_n6366, new_n6367,
    new_n6368, new_n6369, new_n6370, new_n6371, new_n6372, new_n6373,
    new_n6374, new_n6375, new_n6376, new_n6377, new_n6378, new_n6379,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429_1, new_n6430, new_n6431_1, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441_1, new_n6442, new_n6443, new_n6444, new_n6445_1,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469,
    new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475,
    new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6562, new_n6563, new_n6564, new_n6565,
    new_n6566, new_n6567, new_n6568, new_n6569, new_n6570, new_n6571,
    new_n6572, new_n6573, new_n6574, new_n6575, new_n6576, new_n6577,
    new_n6578_1, new_n6579, new_n6580, new_n6581, new_n6582, new_n6583,
    new_n6584, new_n6585, new_n6586, new_n6587, new_n6588, new_n6589,
    new_n6590, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604_1, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611_1, new_n6612, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625,
    new_n6626, new_n6627, new_n6628, new_n6629, new_n6630, new_n6631,
    new_n6632, new_n6633, new_n6634, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645_1, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6650, new_n6651, new_n6652, new_n6653, new_n6654, new_n6655,
    new_n6656, new_n6657, new_n6658, new_n6659, new_n6660, new_n6661,
    new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667,
    new_n6668, new_n6669, new_n6670, new_n6671, new_n6672, new_n6673,
    new_n6674, new_n6675, new_n6676, new_n6677, new_n6678, new_n6679,
    new_n6680, new_n6681, new_n6682, new_n6683, new_n6684, new_n6685,
    new_n6686, new_n6687_1, new_n6688, new_n6689_1, new_n6690, new_n6691,
    new_n6692, new_n6693, new_n6694, new_n6695, new_n6696, new_n6697,
    new_n6698, new_n6699, new_n6700, new_n6701, new_n6702, new_n6703_1,
    new_n6704, new_n6705, new_n6706, new_n6707, new_n6708, new_n6709,
    new_n6710, new_n6711, new_n6712, new_n6713, new_n6714, new_n6715,
    new_n6716, new_n6717, new_n6718, new_n6719, new_n6720, new_n6721,
    new_n6722, new_n6723, new_n6724, new_n6725, new_n6726, new_n6727,
    new_n6728, new_n6729, new_n6730, new_n6731, new_n6732, new_n6733,
    new_n6734, new_n6735, new_n6736, new_n6737, new_n6738, new_n6739,
    new_n6740, new_n6741, new_n6742_1, new_n6743, new_n6744, new_n6745,
    new_n6746, new_n6747, new_n6748, new_n6749, new_n6750, new_n6751,
    new_n6752, new_n6753, new_n6754, new_n6755, new_n6756, new_n6757,
    new_n6758, new_n6759, new_n6760, new_n6761, new_n6762, new_n6763,
    new_n6764, new_n6765, new_n6766, new_n6767, new_n6768, new_n6769,
    new_n6770_1, new_n6771, new_n6772, new_n6773, new_n6774, new_n6775,
    new_n6776_1, new_n6777, new_n6778, new_n6779, new_n6780, new_n6781,
    new_n6782, new_n6783, new_n6784, new_n6785, new_n6786, new_n6787,
    new_n6788, new_n6789, new_n6790, new_n6791, new_n6792, new_n6793,
    new_n6794, new_n6795, new_n6796, new_n6797_1, new_n6798, new_n6799,
    new_n6800, new_n6801, new_n6802, new_n6803, new_n6804, new_n6805,
    new_n6806_1, new_n6807, new_n6808, new_n6809_1, new_n6810, new_n6811,
    new_n6812, new_n6813, new_n6814, new_n6815, new_n6816, new_n6817,
    new_n6818, new_n6819, new_n6820, new_n6821, new_n6822_1, new_n6823,
    new_n6824, new_n6825, new_n6826_1, new_n6827, new_n6828, new_n6829,
    new_n6830, new_n6831, new_n6832, new_n6833, new_n6834, new_n6835,
    new_n6836, new_n6837, new_n6838, new_n6839, new_n6840, new_n6841,
    new_n6842, new_n6843, new_n6844, new_n6845, new_n6846, new_n6847,
    new_n6848, new_n6849, new_n6850, new_n6851, new_n6852, new_n6853,
    new_n6854, new_n6855, new_n6856, new_n6857, new_n6858, new_n6859,
    new_n6860_1, new_n6861, new_n6862, new_n6863, new_n6864, new_n6865,
    new_n6866, new_n6867, new_n6868, new_n6869, new_n6870, new_n6871,
    new_n6872, new_n6873, new_n6874, new_n6875, new_n6876, new_n6877_1,
    new_n6878, new_n6879, new_n6880, new_n6881, new_n6882, new_n6883,
    new_n6884, new_n6885, new_n6886, new_n6887, new_n6888, new_n6889,
    new_n6890, new_n6891, new_n6892, new_n6893, new_n6894, new_n6895,
    new_n6896, new_n6897, new_n6898, new_n6899, new_n6900, new_n6901,
    new_n6902, new_n6903, new_n6904, new_n6905, new_n6906, new_n6907,
    new_n6908, new_n6909, new_n6910, new_n6911, new_n6912, new_n6913,
    new_n6914, new_n6915, new_n6916, new_n6917, new_n6918, new_n6919,
    new_n6920, new_n6921, new_n6922, new_n6923, new_n6924, new_n6925,
    new_n6926, new_n6927, new_n6928, new_n6929, new_n6930, new_n6931,
    new_n6932, new_n6933, new_n6934, new_n6935, new_n6936, new_n6937,
    new_n6938, new_n6939, new_n6940, new_n6941, new_n6942, new_n6943,
    new_n6944, new_n6945, new_n6946, new_n6947, new_n6948, new_n6949,
    new_n6950, new_n6951, new_n6952, new_n6953, new_n6954, new_n6958,
    new_n6959, new_n6960, new_n6961, new_n6962, new_n6963, new_n6964,
    new_n6965, new_n6966, new_n6967, new_n6968, new_n6969, new_n6970,
    new_n6971, new_n6972, new_n6973, new_n6974, new_n6975, new_n6976,
    new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982,
    new_n6983, new_n6984, new_n6985, new_n6986_1, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072,
    new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078,
    new_n7079, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084,
    new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090,
    new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096,
    new_n7097, new_n7098, new_n7099, new_n7100, new_n7101, new_n7102,
    new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108,
    new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114,
    new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120,
    new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159_1, new_n7160_1, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190, new_n7191, new_n7192,
    new_n7193_1, new_n7194, new_n7195, new_n7196, new_n7197, new_n7198,
    new_n7199, new_n7200, new_n7201, new_n7202, new_n7203, new_n7204,
    new_n7205, new_n7206, new_n7207, new_n7208, new_n7209, new_n7210,
    new_n7211, new_n7212, new_n7213, new_n7214, new_n7215, new_n7216,
    new_n7217, new_n7218, new_n7219, new_n7220, new_n7221, new_n7222,
    new_n7223, new_n7224, new_n7225, new_n7226, new_n7227, new_n7228,
    new_n7229, new_n7230, new_n7231, new_n7232, new_n7233, new_n7234,
    new_n7235, new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240,
    new_n7241, new_n7242, new_n7243, new_n7244, new_n7245, new_n7246,
    new_n7247, new_n7248, new_n7249, new_n7250, new_n7251, new_n7252,
    new_n7253, new_n7254, new_n7255, new_n7256, new_n7257, new_n7258,
    new_n7259, new_n7260, new_n7261, new_n7262, new_n7263, new_n7264,
    new_n7265_1, new_n7266, new_n7267, new_n7268, new_n7269, new_n7270_1,
    new_n7271, new_n7272, new_n7273, new_n7274, new_n7275, new_n7276,
    new_n7277, new_n7278, new_n7279, new_n7280, new_n7281, new_n7282,
    new_n7283, new_n7284, new_n7285, new_n7286, new_n7287, new_n7288,
    new_n7289, new_n7290, new_n7291, new_n7292, new_n7293, new_n7294_1,
    new_n7295, new_n7296, new_n7297, new_n7298, new_n7299, new_n7300,
    new_n7301, new_n7302, new_n7303, new_n7304, new_n7305, new_n7306,
    new_n7307, new_n7308, new_n7309, new_n7310, new_n7311, new_n7312,
    new_n7313, new_n7314, new_n7315, new_n7316, new_n7317, new_n7318,
    new_n7319, new_n7320_1, new_n7321, new_n7322, new_n7323, new_n7324,
    new_n7325, new_n7326, new_n7327, new_n7328, new_n7329, new_n7330,
    new_n7331, new_n7332, new_n7333, new_n7334, new_n7335, new_n7336,
    new_n7337, new_n7338, new_n7339, new_n7340, new_n7341, new_n7342,
    new_n7343, new_n7344, new_n7345, new_n7346, new_n7347, new_n7348,
    new_n7349, new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1,
    new_n7355, new_n7356, new_n7357, new_n7358, new_n7359, new_n7360,
    new_n7361, new_n7362, new_n7363, new_n7364, new_n7365, new_n7366,
    new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372,
    new_n7373, new_n7374, new_n7375, new_n7376, new_n7377, new_n7378,
    new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384,
    new_n7385, new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390,
    new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396,
    new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402,
    new_n7403, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408,
    new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7414,
    new_n7415, new_n7416, new_n7417, new_n7418, new_n7419, new_n7420,
    new_n7421, new_n7422, new_n7423, new_n7424, new_n7425, new_n7426,
    new_n7427, new_n7428, new_n7429, new_n7430, new_n7431, new_n7432,
    new_n7433, new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438,
    new_n7439, new_n7440, new_n7441, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1,
    new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523_1, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570,
    new_n7571, new_n7572, new_n7573, new_n7574, new_n7575, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585, new_n7586, new_n7587, new_n7588,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607, new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616, new_n7617, new_n7618,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028_1,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076,
    new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082,
    new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088,
    new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094,
    new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100_1,
    new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106,
    new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112,
    new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118,
    new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124,
    new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130,
    new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136,
    new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141, new_n8142,
    new_n8143, new_n8144, new_n8145, new_n8146, new_n8147, new_n8148,
    new_n8149, new_n8150, new_n8151, new_n8152, new_n8153, new_n8154,
    new_n8155, new_n8156, new_n8157, new_n8158, new_n8159, new_n8160,
    new_n8161, new_n8162, new_n8163, new_n8164, new_n8165, new_n8166,
    new_n8167, new_n8168, new_n8169, new_n8170, new_n8171, new_n8172,
    new_n8173, new_n8174, new_n8175, new_n8176, new_n8177, new_n8178,
    new_n8179, new_n8180, new_n8181, new_n8182, new_n8183, new_n8184,
    new_n8185, new_n8186, new_n8187, new_n8188, new_n8189, new_n8190,
    new_n8191, new_n8192, new_n8193, new_n8194, new_n8195, new_n8196,
    new_n8197, new_n8198, new_n8199, new_n8200, new_n8201, new_n8202_1,
    new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208,
    new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214,
    new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220,
    new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8272, new_n8273, new_n8274, new_n8275, new_n8276_1, new_n8277,
    new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283,
    new_n8284, new_n8285, new_n8286, new_n8287, new_n8288, new_n8289,
    new_n8290, new_n8291, new_n8292, new_n8293, new_n8294, new_n8295,
    new_n8296, new_n8297, new_n8298, new_n8299, new_n8300, new_n8301,
    new_n8302, new_n8303_1, new_n8304, new_n8305, new_n8306, new_n8307,
    new_n8308, new_n8309, new_n8310, new_n8311, new_n8312, new_n8313,
    new_n8314, new_n8315, new_n8316, new_n8317, new_n8318, new_n8319,
    new_n8320, new_n8321, new_n8322, new_n8323, new_n8324, new_n8325,
    new_n8326, new_n8327, new_n8328, new_n8329, new_n8330, new_n8331,
    new_n8332, new_n8333, new_n8334, new_n8335, new_n8336_1, new_n8337,
    new_n8338, new_n8339, new_n8340, new_n8341, new_n8342, new_n8343,
    new_n8344, new_n8345, new_n8346, new_n8347, new_n8348, new_n8349,
    new_n8350, new_n8351, new_n8352, new_n8353, new_n8354, new_n8355,
    new_n8356, new_n8357, new_n8358, new_n8359, new_n8360, new_n8361,
    new_n8363, new_n8364, new_n8365, new_n8366, new_n8367, new_n8368,
    new_n8369, new_n8370, new_n8371, new_n8372, new_n8373, new_n8374,
    new_n8375, new_n8376, new_n8377, new_n8378, new_n8379, new_n8380,
    new_n8381, new_n8382, new_n8383, new_n8384_1, new_n8385, new_n8386,
    new_n8387, new_n8388, new_n8389, new_n8390, new_n8391, new_n8392,
    new_n8393, new_n8394, new_n8395, new_n8396, new_n8397, new_n8398_1,
    new_n8399, new_n8400, new_n8401, new_n8402, new_n8403, new_n8404,
    new_n8405, new_n8406, new_n8407, new_n8408, new_n8409, new_n8410,
    new_n8411, new_n8412, new_n8413, new_n8414, new_n8415, new_n8416,
    new_n8417, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422,
    new_n8423, new_n8424, new_n8425, new_n8426, new_n8427, new_n8428,
    new_n8429, new_n8430, new_n8431, new_n8432, new_n8433_1, new_n8434,
    new_n8435, new_n8436, new_n8437, new_n8438, new_n8439, new_n8440,
    new_n8441, new_n8442, new_n8443, new_n8444, new_n8445, new_n8446,
    new_n8447, new_n8448, new_n8449, new_n8450, new_n8451, new_n8452,
    new_n8453, new_n8454, new_n8455, new_n8456, new_n8457, new_n8458,
    new_n8459, new_n8460, new_n8461, new_n8462, new_n8463, new_n8464,
    new_n8465, new_n8466, new_n8467, new_n8468, new_n8469, new_n8470,
    new_n8471, new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1,
    new_n8477, new_n8478, new_n8479, new_n8480, new_n8481, new_n8482,
    new_n8483, new_n8484, new_n8485, new_n8486, new_n8487, new_n8488,
    new_n8489, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494,
    new_n8495, new_n8496, new_n8497, new_n8498, new_n8499, new_n8500,
    new_n8501, new_n8502, new_n8503, new_n8504, new_n8505, new_n8506,
    new_n8507, new_n8508, new_n8509, new_n8510, new_n8511, new_n8512,
    new_n8513, new_n8514, new_n8515, new_n8516, new_n8517, new_n8518,
    new_n8519, new_n8520, new_n8521, new_n8522, new_n8523, new_n8524,
    new_n8525, new_n8526, new_n8527, new_n8528, new_n8529, new_n8530,
    new_n8531, new_n8532, new_n8533, new_n8534, new_n8535, new_n8536,
    new_n8537, new_n8538, new_n8539, new_n8540, new_n8541, new_n8542,
    new_n8543, new_n8544, new_n8545, new_n8546, new_n8547, new_n8548,
    new_n8549, new_n8550, new_n8551, new_n8552, new_n8553, new_n8554,
    new_n8555, new_n8556, new_n8557, new_n8558, new_n8559, new_n8560,
    new_n8561, new_n8562, new_n8563, new_n8564, new_n8565, new_n8566,
    new_n8567, new_n8568, new_n8569, new_n8570, new_n8571, new_n8572,
    new_n8573, new_n8574, new_n8575, new_n8576, new_n8577, new_n8578,
    new_n8579, new_n8580, new_n8581, new_n8582, new_n8583, new_n8584,
    new_n8585, new_n8586, new_n8587, new_n8588, new_n8589, new_n8590,
    new_n8591, new_n8592, new_n8593, new_n8594, new_n8595_1, new_n8596,
    new_n8597, new_n8598, new_n8599, new_n8600, new_n8601, new_n8602,
    new_n8603, new_n8604, new_n8605, new_n8606, new_n8607, new_n8608,
    new_n8609, new_n8610, new_n8611, new_n8612, new_n8613, new_n8614,
    new_n8615, new_n8616, new_n8617, new_n8618, new_n8619, new_n8620,
    new_n8621, new_n8622, new_n8623, new_n8624, new_n8625, new_n8626,
    new_n8627, new_n8628, new_n8629, new_n8630, new_n8631, new_n8632,
    new_n8633, new_n8634, new_n8635, new_n8636, new_n8637, new_n8638,
    new_n8639, new_n8640, new_n8641, new_n8642, new_n8643, new_n8644,
    new_n8645, new_n8646, new_n8647, new_n8648, new_n8649, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662,
    new_n8663, new_n8664, new_n8665_1, new_n8666, new_n8667, new_n8668,
    new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674,
    new_n8675, new_n8676, new_n8677, new_n8678, new_n8679, new_n8680,
    new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686,
    new_n8687, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692,
    new_n8693, new_n8694, new_n8695, new_n8696, new_n8697, new_n8698,
    new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704,
    new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710,
    new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716,
    new_n8717_1, new_n8718, new_n8719, new_n8720, new_n8721, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744, new_n8745, new_n8746,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759_1, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803, new_n8804, new_n8805, new_n8806,
    new_n8807, new_n8808, new_n8809, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819_1, new_n8820, new_n8821, new_n8822, new_n8823, new_n8824,
    new_n8825, new_n8826, new_n8827, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861, new_n8862, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884,
    new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890,
    new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896,
    new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902,
    new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908,
    new_n8909, new_n8910, new_n8911, new_n8912, new_n8913, new_n8914,
    new_n8915, new_n8916, new_n8917, new_n8918, new_n8919, new_n8920,
    new_n8921, new_n8922, new_n8923, new_n8924, new_n8925, new_n8926,
    new_n8927, new_n8928, new_n8929, new_n8930, new_n8931, new_n8932,
    new_n8933, new_n8934, new_n8935, new_n8936, new_n8937, new_n8938,
    new_n8939, new_n8940, new_n8941, new_n8942, new_n8943, new_n8944,
    new_n8945, new_n8946, new_n8947, new_n8948, new_n8949, new_n8950,
    new_n8951, new_n8952, new_n8953, new_n8954, new_n8955, new_n8956,
    new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962,
    new_n8963, new_n8964, new_n8965, new_n8966, new_n8967, new_n8968,
    new_n8969, new_n8970, new_n8971, new_n8972, new_n8973, new_n8974,
    new_n8975, new_n8976, new_n8977, new_n8978, new_n8979, new_n8980,
    new_n8981, new_n8982, new_n8983, new_n8984, new_n8985, new_n8986,
    new_n8987, new_n8988, new_n8989, new_n8990, new_n8991, new_n8992,
    new_n8993, new_n8994, new_n8995, new_n8996, new_n8997, new_n8998,
    new_n8999, new_n9000, new_n9001, new_n9002, new_n9003, new_n9004,
    new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010,
    new_n9011, new_n9012, new_n9013, new_n9014, new_n9015, new_n9016,
    new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022,
    new_n9023, new_n9024, new_n9025, new_n9026, new_n9027, new_n9028,
    new_n9029, new_n9030, new_n9042, new_n9043, new_n9044, new_n9045,
    new_n9046, new_n9047, new_n9048, new_n9049, new_n9050, new_n9051,
    new_n9052, new_n9053, new_n9054, new_n9055, new_n9056, new_n9057,
    new_n9058, new_n9059, new_n9060, new_n9061, new_n9062, new_n9063,
    new_n9064, new_n9065, new_n9066, new_n9067, new_n9068, new_n9069,
    new_n9070, new_n9071, new_n9072, new_n9073, new_n9074, new_n9075,
    new_n9076, new_n9077, new_n9078, new_n9079, new_n9080_1, new_n9081,
    new_n9082, new_n9083, new_n9084, new_n9085, new_n9086, new_n9087,
    new_n9088, new_n9089, new_n9090, new_n9091, new_n9092, new_n9093,
    new_n9094, new_n9095, new_n9096, new_n9097, new_n9098, new_n9099,
    new_n9100, new_n9101, new_n9102, new_n9103, new_n9104, new_n9105,
    new_n9106, new_n9107, new_n9108, new_n9109, new_n9110, new_n9111_1,
    new_n9112, new_n9113, new_n9114, new_n9115, new_n9116, new_n9117,
    new_n9118, new_n9119, new_n9120, new_n9121, new_n9122, new_n9123,
    new_n9124, new_n9125, new_n9126, new_n9127, new_n9128, new_n9129,
    new_n9130, new_n9131, new_n9132, new_n9133, new_n9134, new_n9135,
    new_n9136, new_n9137_1, new_n9138, new_n9139, new_n9140, new_n9141,
    new_n9142, new_n9143, new_n9144, new_n9145, new_n9146, new_n9147,
    new_n9148, new_n9149, new_n9150, new_n9151, new_n9152, new_n9153,
    new_n9154, new_n9155, new_n9156, new_n9157, new_n9158, new_n9159,
    new_n9160, new_n9161, new_n9162, new_n9163, new_n9164, new_n9165,
    new_n9166, new_n9167, new_n9168, new_n9169, new_n9170, new_n9171,
    new_n9172, new_n9173, new_n9174, new_n9175, new_n9176, new_n9177,
    new_n9178, new_n9179, new_n9180, new_n9181, new_n9182, new_n9183,
    new_n9184, new_n9185, new_n9186, new_n9187, new_n9188, new_n9189_1,
    new_n9190, new_n9191, new_n9192, new_n9193, new_n9194, new_n9195_1,
    new_n9196, new_n9197, new_n9198, new_n9199, new_n9200, new_n9201,
    new_n9202, new_n9203, new_n9204, new_n9205, new_n9206, new_n9207,
    new_n9208, new_n9209, new_n9210, new_n9211, new_n9212, new_n9213,
    new_n9214, new_n9215, new_n9216, new_n9217, new_n9218, new_n9219,
    new_n9220, new_n9221, new_n9222, new_n9223, new_n9224, new_n9225,
    new_n9226, new_n9227, new_n9228, new_n9229, new_n9230, new_n9231,
    new_n9232, new_n9233, new_n9234, new_n9235, new_n9236, new_n9237,
    new_n9238, new_n9239, new_n9240, new_n9241_1, new_n9242, new_n9243,
    new_n9244, new_n9245, new_n9246, new_n9247, new_n9248, new_n9249,
    new_n9250, new_n9251, new_n9252, new_n9253, new_n9254, new_n9255,
    new_n9256, new_n9257, new_n9258, new_n9259, new_n9260, new_n9261,
    new_n9262, new_n9263, new_n9264, new_n9265, new_n9266, new_n9267,
    new_n9268, new_n9269, new_n9270, new_n9271, new_n9272, new_n9273,
    new_n9274, new_n9275, new_n9276, new_n9277, new_n9278, new_n9279,
    new_n9280, new_n9281, new_n9282, new_n9283, new_n9284, new_n9285,
    new_n9286, new_n9287, new_n9288, new_n9289, new_n9290, new_n9291,
    new_n9292, new_n9293, new_n9294, new_n9295, new_n9296, new_n9297,
    new_n9298, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387_1, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400_1, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457_1, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9485, new_n9486, new_n9487,
    new_n9488, new_n9489, new_n9490, new_n9491, new_n9492, new_n9493,
    new_n9494, new_n9495, new_n9496, new_n9497, new_n9498, new_n9499,
    new_n9500, new_n9501, new_n9502, new_n9503, new_n9504, new_n9505,
    new_n9506, new_n9507, new_n9508, new_n9509, new_n9510, new_n9511,
    new_n9512, new_n9513, new_n9514, new_n9515, new_n9516, new_n9517,
    new_n9518, new_n9519, new_n9520, new_n9521, new_n9522, new_n9523,
    new_n9524, new_n9525, new_n9526, new_n9527, new_n9528, new_n9529,
    new_n9530, new_n9531, new_n9532, new_n9533, new_n9534, new_n9535,
    new_n9536, new_n9537, new_n9538, new_n9539, new_n9540, new_n9541,
    new_n9542, new_n9543, new_n9544, new_n9545, new_n9546, new_n9547,
    new_n9548, new_n9549, new_n9550, new_n9551, new_n9552, new_n9553,
    new_n9554, new_n9555, new_n9556, new_n9557, new_n9558, new_n9559,
    new_n9560, new_n9561, new_n9562, new_n9563, new_n9564, new_n9565,
    new_n9566, new_n9567, new_n9568, new_n9569, new_n9570, new_n9571_1,
    new_n9572, new_n9573, new_n9574, new_n9575, new_n9576, new_n9577,
    new_n9578_1, new_n9579, new_n9580, new_n9581, new_n9582, new_n9583_1,
    new_n9584, new_n9585, new_n9586, new_n9587, new_n9588, new_n9589,
    new_n9590, new_n9591, new_n9592, new_n9593, new_n9594, new_n9595,
    new_n9596, new_n9597, new_n9598, new_n9599, new_n9600, new_n9601,
    new_n9602, new_n9603, new_n9604, new_n9605, new_n9606, new_n9607,
    new_n9608, new_n9609, new_n9610, new_n9611, new_n9612, new_n9613,
    new_n9614, new_n9615, new_n9616, new_n9617, new_n9618, new_n9619,
    new_n9620, new_n9621, new_n9622, new_n9623, new_n9624, new_n9625,
    new_n9626, new_n9627, new_n9628, new_n9629, new_n9630, new_n9631,
    new_n9632, new_n9633, new_n9634, new_n9635, new_n9636, new_n9637_1,
    new_n9638, new_n9639, new_n9640_1, new_n9641, new_n9642, new_n9643,
    new_n9644, new_n9645, new_n9646, new_n9647, new_n9648, new_n9649,
    new_n9650, new_n9651, new_n9652, new_n9653, new_n9654, new_n9655,
    new_n9656, new_n9657, new_n9658, new_n9659, new_n9660, new_n9661,
    new_n9662, new_n9663, new_n9664, new_n9665, new_n9666, new_n9667,
    new_n9668, new_n9669, new_n9670, new_n9671, new_n9672, new_n9673,
    new_n9674, new_n9675, new_n9676, new_n9677, new_n9678, new_n9679,
    new_n9680, new_n9681, new_n9682, new_n9683, new_n9684, new_n9685,
    new_n9686, new_n9687, new_n9688, new_n9689, new_n9690, new_n9691,
    new_n9692, new_n9693, new_n9694, new_n9695, new_n9696, new_n9697,
    new_n9698, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703,
    new_n9704, new_n9705, new_n9706_1, new_n9707, new_n9708, new_n9709,
    new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715,
    new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725_1, new_n9726, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739,
    new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753, new_n9754, new_n9755, new_n9756_1, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763_1,
    new_n9764, new_n9765, new_n9766, new_n9767_1, new_n9768, new_n9769,
    new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9808, new_n9809, new_n9810, new_n9811,
    new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817,
    new_n9818, new_n9819, new_n9820_1, new_n9821, new_n9822, new_n9823,
    new_n9824, new_n9825, new_n9826, new_n9827, new_n9828, new_n9829,
    new_n9830, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835,
    new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841,
    new_n9842, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889,
    new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920_1, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938_1, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956_1, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009, new_n10010, new_n10011,
    new_n10012, new_n10013, new_n10014, new_n10015, new_n10016, new_n10017,
    new_n10018, new_n10019, new_n10020, new_n10021, new_n10022_1,
    new_n10023, new_n10024, new_n10025, new_n10026, new_n10027, new_n10028,
    new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034,
    new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10048, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053, new_n10054, new_n10055, new_n10056, new_n10057, new_n10058,
    new_n10059, new_n10060, new_n10061, new_n10062, new_n10063, new_n10064,
    new_n10065, new_n10066, new_n10067, new_n10068, new_n10069, new_n10070,
    new_n10071, new_n10072, new_n10073, new_n10074, new_n10075, new_n10076,
    new_n10077, new_n10078, new_n10079, new_n10080, new_n10081, new_n10082,
    new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088,
    new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094,
    new_n10095, new_n10096, new_n10097, new_n10098, new_n10099, new_n10100,
    new_n10101, new_n10102, new_n10103, new_n10104, new_n10105, new_n10106,
    new_n10107, new_n10108, new_n10109, new_n10110, new_n10111, new_n10112,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117, new_n10118,
    new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125, new_n10126, new_n10127, new_n10128, new_n10129, new_n10130,
    new_n10131, new_n10132, new_n10133, new_n10134, new_n10135, new_n10136,
    new_n10137, new_n10138, new_n10139, new_n10140, new_n10141, new_n10142,
    new_n10143, new_n10144, new_n10145, new_n10146, new_n10147, new_n10148,
    new_n10149, new_n10150, new_n10151, new_n10152, new_n10153, new_n10154,
    new_n10155, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174_1, new_n10175, new_n10176,
    new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182,
    new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188,
    new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194,
    new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206,
    new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212,
    new_n10213, new_n10214, new_n10215, new_n10216, new_n10217_1,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222,
    new_n10223_1, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251,
    new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275,
    new_n10276, new_n10277, new_n10278_1, new_n10279, new_n10280,
    new_n10281, new_n10282, new_n10283, new_n10284, new_n10285, new_n10286,
    new_n10287, new_n10288, new_n10289, new_n10290, new_n10291, new_n10292,
    new_n10293, new_n10294, new_n10295, new_n10296, new_n10297, new_n10298,
    new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304,
    new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310,
    new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316,
    new_n10317, new_n10318, new_n10319, new_n10320, new_n10321, new_n10322,
    new_n10323, new_n10324, new_n10325, new_n10326, new_n10327_1,
    new_n10328, new_n10329, new_n10330, new_n10331, new_n10332, new_n10333,
    new_n10334, new_n10335, new_n10336, new_n10337, new_n10338, new_n10339,
    new_n10346, new_n10353, new_n10354, new_n10355, new_n10356, new_n10357,
    new_n10358, new_n10359, new_n10360, new_n10361, new_n10362, new_n10363,
    new_n10364, new_n10365, new_n10366, new_n10367, new_n10368, new_n10369,
    new_n10370, new_n10371, new_n10372, new_n10373, new_n10374, new_n10375,
    new_n10376, new_n10377, new_n10378, new_n10379, new_n10380, new_n10381,
    new_n10382, new_n10383, new_n10384, new_n10385, new_n10386, new_n10387,
    new_n10388, new_n10389, new_n10390, new_n10391_1, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439_1,
    new_n10440, new_n10441, new_n10442, new_n10443, new_n10444, new_n10445,
    new_n10446, new_n10447, new_n10448, new_n10449, new_n10450,
    new_n10451_1, new_n10452, new_n10453, new_n10454, new_n10455,
    new_n10456, new_n10457, new_n10458, new_n10459, new_n10460, new_n10461,
    new_n10462, new_n10463, new_n10464, new_n10465, new_n10466, new_n10467,
    new_n10468, new_n10469, new_n10470, new_n10471, new_n10472, new_n10473,
    new_n10474, new_n10475, new_n10476_1, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484,
    new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490,
    new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496,
    new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502,
    new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508,
    new_n10509, new_n10510_1, new_n10511, new_n10512, new_n10513,
    new_n10514, new_n10515, new_n10516, new_n10517, new_n10518, new_n10519,
    new_n10520, new_n10521, new_n10522, new_n10523, new_n10524, new_n10525;
and_5  g00000(n6687, n6038, new_n377);
and_5  g00001(n8336, n7354, new_n378);
and_5  g00002(n11222, n8028, new_n379);
and_5  g00003(n12069, n1564, new_n380);
xnor_4 g00004(new_n380, new_n379, new_n381_1);
xnor_4 g00005(new_n381_1, new_n378, new_n382);
xor_4  g00006(new_n382, new_n377, n112);
nand_5 g00007(n12720, n4312, new_n384);
and_5  g00008(n12025, n6038, new_n385);
and_5  g00009(n12705, n2509, new_n386);
xnor_4 g00010(new_n386, new_n385, new_n387);
xnor_4 g00011(new_n387, new_n384, new_n388);
and_5  g00012(n12705, n6038, new_n389);
and_5  g00013(n12720, n1097, new_n390);
nor_5  g00014(new_n390, new_n389, new_n391);
and_5  g00015(n4312, n2509, new_n392);
xnor_4 g00016(new_n390, new_n389, new_n393);
nor_5  g00017(new_n393, new_n392, new_n394);
or_5   g00018(new_n394, new_n391, new_n395);
xnor_4 g00019(new_n395, new_n388, new_n396);
and_5  g00020(n2508, n1097, new_n397_1);
and_5  g00021(n5964, n2585, new_n398);
xnor_4 g00022(new_n398, new_n397_1, new_n399);
xnor_4 g00023(new_n399, new_n396, new_n400);
and_5  g00024(n5964, n2508, new_n401);
xnor_4 g00025(new_n393, new_n392, new_n402);
nor_5  g00026(new_n402, new_n401, new_n403);
xnor_4 g00027(new_n402, new_n401, new_n404);
and_5  g00028(n6038, n4312, new_n405_1);
and_5  g00029(n12720, n5964, new_n406);
nor_5  g00030(new_n406, new_n405_1, new_n407);
nand_5 g00031(new_n406, new_n405_1, new_n408);
nand_5 g00032(n2509, n1097, new_n409);
and_5  g00033(new_n409, new_n408, new_n410);
nor_5  g00034(new_n410, new_n407, new_n411);
nor_5  g00035(new_n411, new_n404, new_n412);
or_5   g00036(new_n412, new_n403, new_n413);
xnor_4 g00037(new_n413, new_n400, new_n414);
nand_5 g00038(n5305, n2585, new_n415);
xor_4  g00039(new_n411, new_n404, new_n416);
and_5  g00040(new_n416, new_n415, new_n417);
xnor_4 g00041(new_n416, new_n415, new_n418);
nand_5 g00042(n5305, n2508, new_n419);
and_5  g00043(n6038, n1097, new_n420);
and_5  g00044(n12720, n5305, new_n421);
nand_5 g00045(new_n421, new_n420, new_n422);
nor_5  g00046(new_n421, new_n420, new_n423);
nand_5 g00047(n5964, n2509, new_n424);
or_5   g00048(new_n424, new_n423, new_n425);
and_5  g00049(new_n425, new_n422, new_n426);
nor_5  g00050(new_n426, new_n419, new_n427);
xnor_4 g00051(new_n426, new_n419, new_n428);
xnor_4 g00052(new_n406, new_n405_1, new_n429);
xnor_4 g00053(new_n429, new_n409, new_n430);
nor_5  g00054(new_n430, new_n428, new_n431);
or_5   g00055(new_n431, new_n427, new_n432);
nor_5  g00056(new_n432, new_n418, new_n433);
or_5   g00057(new_n433, new_n417, new_n434);
nor_5  g00058(new_n434, new_n414, new_n435);
nor_5  g00059(new_n387, new_n384, new_n436);
nor_5  g00060(new_n395, new_n388, new_n437);
or_5   g00061(new_n437, new_n436, new_n438);
nand_5 g00062(n5964, n4005, new_n439);
and_5  g00063(n2585, n1097, new_n440);
and_5  g00064(n12706, n5305, new_n441);
xnor_4 g00065(new_n441, new_n440, new_n442);
xor_4  g00066(new_n442, new_n439, new_n443);
xnor_4 g00067(new_n443, new_n438, new_n444);
and_5  g00068(new_n386, new_n385, new_n445);
and_5  g00069(n4312, n2508, new_n446);
xnor_4 g00070(new_n446, new_n445, new_n447_1);
and_5  g00071(n12025, n2509, new_n448);
and_5  g00072(n12720, n12705, new_n449);
and_5  g00073(n11257, n6038, new_n450);
xnor_4 g00074(new_n450, new_n449, new_n451);
xor_4  g00075(new_n451, new_n448, new_n452);
xor_4  g00076(new_n452, new_n447_1, new_n453);
xor_4  g00077(new_n453, new_n444, new_n454);
nor_5  g00078(new_n399, new_n396, new_n455);
nand_5 g00079(new_n398, new_n397_1, new_n456);
or_5   g00080(new_n413, new_n400, new_n457);
xor_4  g00081(new_n457, new_n456, new_n458);
nor_5  g00082(new_n458, new_n455, new_n459);
xor_4  g00083(new_n459, new_n454, new_n460);
xnor_4 g00084(new_n460, new_n435, new_n461);
and_5  g00085(n5305, n4005, new_n462);
xor_4  g00086(new_n434, new_n414, new_n463);
and_5  g00087(new_n463, new_n462, new_n464);
nor_5  g00088(new_n463, new_n462, new_n465);
xnor_4 g00089(new_n430, new_n428, new_n466);
xor_4  g00090(new_n421, new_n420, new_n467);
and_5  g00091(n6038, n5964, new_n468);
and_5  g00092(n5305, n2509, new_n469);
nand_5 g00093(new_n469, new_n468, new_n470);
or_5   g00094(new_n470, new_n467, new_n471);
or_5   g00095(new_n471, new_n466, new_n472);
xor_4  g00096(new_n432, new_n418, new_n473);
or_5   g00097(new_n473, new_n472, new_n474);
nor_5  g00098(new_n474, new_n465, new_n475);
nor_5  g00099(new_n475, new_n464, new_n476);
xnor_4 g00100(new_n476, new_n461, new_n477);
nand_5 g00101(n8759, n5105, new_n478);
and_5  g00102(n12299, n7354, new_n479);
and_5  g00103(n8759, n1209, new_n480);
nor_5  g00104(new_n480, new_n479, new_n481);
and_5  g00105(new_n480, new_n479, new_n482);
and_5  g00106(n7500, n6776, new_n483);
nor_5  g00107(new_n483, new_n482, new_n484);
or_5   g00108(new_n484, new_n481, new_n485);
xnor_4 g00109(new_n485, new_n478, new_n486);
and_5  g00110(n12299, n7500, new_n487);
and_5  g00111(n7436, n7354, new_n488);
and_5  g00112(n6776, n1209, new_n489);
xnor_4 g00113(new_n489, new_n488, new_n490);
xor_4  g00114(new_n490, new_n487, new_n491);
xnor_4 g00115(new_n491, new_n486, new_n492);
nand_5 g00116(n7500, n6776, new_n493);
and_5  g00117(n8759, n7354, new_n494);
or_5   g00118(new_n494, new_n493, new_n495);
and_5  g00119(new_n495, new_n481, new_n496);
nor_5  g00120(new_n496, new_n482, new_n497);
or_5   g00121(new_n497, new_n493, new_n498);
or_5   g00122(new_n498, new_n492, new_n499);
nand_5 g00123(n8759, n4141, new_n500);
and_5  g00124(n6776, n5105, new_n501);
nor_5  g00125(new_n489, new_n488, new_n502);
nor_5  g00126(new_n490, new_n487, new_n503_1);
nor_5  g00127(new_n503_1, new_n502, new_n504);
xnor_4 g00128(new_n504, new_n501, new_n505);
and_5  g00129(n7500, n7436, new_n506);
and_5  g00130(n12299, n1209, new_n507);
and_5  g00131(n8276, n7354, new_n508);
xnor_4 g00132(new_n508, new_n507, new_n509);
xor_4  g00133(new_n509, new_n506, new_n510);
xnor_4 g00134(new_n510, new_n505, new_n511);
xnor_4 g00135(new_n511, new_n500, new_n512);
nor_5  g00136(new_n485, new_n478, new_n513);
nor_5  g00137(new_n491, new_n486, new_n514);
nor_5  g00138(new_n514, new_n513, new_n515);
xnor_4 g00139(new_n515, new_n512, new_n516);
or_5   g00140(new_n516, new_n499, new_n517);
nand_5 g00141(n8759, n4928, new_n518);
nand_5 g00142(n7436, n1209, new_n519);
and_5  g00143(n8276, n7500, new_n520);
and_5  g00144(n9241, n7354, new_n521_1);
xnor_4 g00145(new_n521_1, new_n520, new_n522);
xnor_4 g00146(new_n522, new_n519, new_n523);
nor_5  g00147(new_n508, new_n507, new_n524);
nor_5  g00148(new_n509, new_n506, new_n525);
or_5   g00149(new_n525, new_n524, new_n526);
xnor_4 g00150(new_n526, new_n523, new_n527);
and_5  g00151(n6776, n4141, new_n528);
and_5  g00152(n12299, n5105, new_n529);
xnor_4 g00153(new_n529, new_n528, new_n530);
xnor_4 g00154(new_n530, new_n527, new_n531);
and_5  g00155(new_n504, new_n501, new_n532);
nor_5  g00156(new_n510, new_n505, new_n533_1);
nor_5  g00157(new_n533_1, new_n532, new_n534);
xnor_4 g00158(new_n534, new_n531, new_n535);
nor_5  g00159(new_n511, new_n500, new_n536);
nor_5  g00160(new_n515, new_n512, new_n537);
nor_5  g00161(new_n537, new_n536, new_n538);
xnor_4 g00162(new_n538, new_n535, new_n539);
xnor_4 g00163(new_n539, new_n518, new_n540);
xor_4  g00164(new_n540, new_n517, new_n541);
xor_4  g00165(new_n516, new_n499, new_n542);
xor_4  g00166(new_n498, new_n492, new_n543);
nand_5 g00167(n8759, n7354, new_n544);
and_5  g00168(n5331, n1564, new_n545);
and_5  g00169(n8028, n7965, new_n546);
xnor_4 g00170(new_n546, new_n545, new_n547);
nor_5  g00171(new_n547, new_n544, new_n548);
and_5  g00172(n7354, n6776, new_n549);
and_5  g00173(n8759, n7500, new_n550);
xor_4  g00174(new_n550, new_n549, new_n551);
nor_5  g00175(new_n551, new_n548, new_n552);
and_5  g00176(new_n546, new_n545, new_n553);
and_5  g00177(n5331, n1512, new_n554);
and_5  g00178(n8476, n1564, new_n555);
xor_4  g00179(new_n555, new_n554, new_n556);
xnor_4 g00180(new_n556, new_n553, new_n557);
and_5  g00181(n8028, n7388, new_n558);
and_5  g00182(n10848, n7965, new_n559);
xnor_4 g00183(new_n559, new_n558, new_n560);
xor_4  g00184(new_n560, new_n557, new_n561);
xnor_4 g00185(new_n551, new_n548, new_n562);
nor_5  g00186(new_n562, new_n561, new_n563);
nor_5  g00187(new_n563, new_n552, new_n564);
or_5   g00188(new_n495, new_n481, new_n565);
and_5  g00189(new_n565, new_n497, new_n566);
nor_5  g00190(new_n566, new_n564, new_n567);
nand_5 g00191(n10848, n7388, new_n568);
nor_5  g00192(new_n568, new_n546, new_n569);
and_5  g00193(n11892, n8028, new_n570);
and_5  g00194(n7965, n1980, new_n571);
nor_5  g00195(new_n571, new_n570, new_n572);
and_5  g00196(n11892, n1980, new_n573);
and_5  g00197(new_n573, new_n546, new_n574);
nor_5  g00198(new_n574, new_n572, new_n575);
or_5   g00199(new_n575, new_n569, new_n576);
or_5   g00200(new_n568, new_n546, new_n577);
or_5   g00201(new_n572, new_n577, new_n578);
nand_5 g00202(new_n578, new_n576, new_n579);
nand_5 g00203(n8476, n1512, new_n580);
or_5   g00204(new_n580, new_n545, new_n581);
and_5  g00205(n2530, n1564, new_n582);
and_5  g00206(n5331, n533, new_n583);
nor_5  g00207(new_n583, new_n582, new_n584);
and_5  g00208(new_n584, new_n581, new_n585);
and_5  g00209(new_n583, new_n582, new_n586);
nor_5  g00210(new_n586, new_n585, new_n587);
or_5   g00211(new_n584, new_n581, new_n588);
nand_5 g00212(new_n588, new_n587, new_n589);
xnor_4 g00213(new_n589, new_n579, new_n590);
and_5  g00214(new_n556, new_n553, new_n591);
nor_5  g00215(new_n560, new_n557, new_n592);
nor_5  g00216(new_n592, new_n591, new_n593);
xnor_4 g00217(new_n593, new_n590, new_n594);
xor_4  g00218(new_n566, new_n564, new_n595);
and_5  g00219(new_n595, new_n594, new_n596);
nor_5  g00220(new_n596, new_n567, new_n597);
nor_5  g00221(new_n597, new_n543, new_n598);
nand_5 g00222(n5331, n2802, new_n599);
and_5  g00223(n8476, n1512, new_n600);
nor_5  g00224(new_n586, new_n600, new_n601);
or_5   g00225(new_n601, new_n584, new_n602);
xnor_4 g00226(new_n602, new_n599, new_n603);
and_5  g00227(n2530, n1512, new_n604);
and_5  g00228(n12648, n1564, new_n605);
and_5  g00229(n8476, n533, new_n606);
xnor_4 g00230(new_n606, new_n605, new_n607);
xor_4  g00231(new_n607, new_n604, new_n608);
xnor_4 g00232(new_n608, new_n603, new_n609);
or_5   g00233(new_n587, new_n580, new_n610);
xor_4  g00234(new_n610, new_n609, new_n611);
nand_5 g00235(n7965, n7294, new_n612);
and_5  g00236(n10848, n7388, new_n613);
nor_5  g00237(new_n574, new_n613, new_n614);
or_5   g00238(new_n614, new_n572, new_n615_1);
xor_4  g00239(new_n615_1, new_n612, new_n616);
and_5  g00240(n11892, n10848, new_n617);
and_5  g00241(n7388, n1980, new_n618);
and_5  g00242(n8028, n2393, new_n619);
xnor_4 g00243(new_n619, new_n618, new_n620);
xnor_4 g00244(new_n620, new_n617, new_n621);
xnor_4 g00245(new_n621, new_n616, new_n622);
or_5   g00246(new_n576, new_n568, new_n623);
xor_4  g00247(new_n623, new_n622, new_n624);
xor_4  g00248(new_n624, new_n611, new_n625);
nor_5  g00249(new_n589, new_n579, new_n626);
nor_5  g00250(new_n593, new_n590, new_n627);
nor_5  g00251(new_n627, new_n626, new_n628);
xnor_4 g00252(new_n628, new_n625, new_n629);
xnor_4 g00253(new_n597, new_n543, new_n630);
nor_5  g00254(new_n630, new_n629, new_n631);
nor_5  g00255(new_n631, new_n598, new_n632);
nor_5  g00256(new_n632, new_n542, new_n633);
nor_5  g00257(new_n623, new_n622, new_n634);
nor_5  g00258(new_n615_1, new_n612, new_n635);
and_5  g00259(new_n621, new_n616, new_n636);
nor_5  g00260(new_n636, new_n635, new_n637);
and_5  g00261(n12704, n7965, new_n638);
nand_5 g00262(n7388, n7294, new_n639);
nor_5  g00263(new_n619, new_n618, new_n640);
and_5  g00264(new_n619, new_n618, new_n641);
nor_5  g00265(new_n641, new_n617, new_n642);
or_5   g00266(new_n642, new_n640, new_n643);
xnor_4 g00267(new_n643, new_n639, new_n644);
and_5  g00268(n10848, n2393, new_n645);
and_5  g00269(n8028, n5860, new_n646);
xnor_4 g00270(new_n646, new_n573, new_n647);
xor_4  g00271(new_n647, new_n645, new_n648);
xor_4  g00272(new_n648, new_n644, new_n649);
xor_4  g00273(new_n649, new_n638, new_n650);
xnor_4 g00274(new_n650, new_n637, new_n651);
xnor_4 g00275(new_n651, new_n634, new_n652);
or_5   g00276(new_n610, new_n609, new_n653);
nand_5 g00277(n6806, n5331, new_n654);
and_5  g00278(n8476, n2802, new_n655);
nor_5  g00279(new_n606, new_n605, new_n656);
nor_5  g00280(new_n607, new_n604, new_n657);
nor_5  g00281(new_n657, new_n656, new_n658_1);
xnor_4 g00282(new_n658_1, new_n655, new_n659);
and_5  g00283(n12648, n1512, new_n660);
and_5  g00284(n2530, n533, new_n661);
and_5  g00285(n10545, n1564, new_n662);
xnor_4 g00286(new_n662, new_n661, new_n663);
xor_4  g00287(new_n663, new_n660, new_n664);
xnor_4 g00288(new_n664, new_n659, new_n665);
xnor_4 g00289(new_n665, new_n654, new_n666);
nor_5  g00290(new_n602, new_n599, new_n667);
nor_5  g00291(new_n608, new_n603, new_n668);
nor_5  g00292(new_n668, new_n667, new_n669);
xnor_4 g00293(new_n669, new_n666, new_n670);
xor_4  g00294(new_n670, new_n653, new_n671_1);
nor_5  g00295(new_n624, new_n611, new_n672);
and_5  g00296(new_n628, new_n625, new_n673);
nor_5  g00297(new_n673, new_n672, new_n674);
xor_4  g00298(new_n674, new_n671_1, new_n675);
xnor_4 g00299(new_n675, new_n652, new_n676);
xnor_4 g00300(new_n632, new_n542, new_n677);
nor_5  g00301(new_n677, new_n676, new_n678);
nor_5  g00302(new_n678, new_n633, new_n679);
xnor_4 g00303(new_n679, new_n541, new_n680);
nor_5  g00304(new_n674, new_n671_1, new_n681);
and_5  g00305(new_n675, new_n652, new_n682);
nor_5  g00306(new_n682, new_n681, new_n683);
or_5   g00307(new_n670, new_n653, new_n684);
and_5  g00308(n5331, n5069, new_n685);
nand_5 g00309(n12648, n533, new_n686);
and_5  g00310(n10545, n1512, new_n687);
and_5  g00311(n7690, n1564, new_n688);
xnor_4 g00312(new_n688, new_n687, new_n689);
xnor_4 g00313(new_n689, new_n686, new_n690);
nor_5  g00314(new_n662, new_n661, new_n691);
nor_5  g00315(new_n663, new_n660, new_n692);
or_5   g00316(new_n692, new_n691, new_n693);
xnor_4 g00317(new_n693, new_n690, new_n694);
and_5  g00318(n8476, n6806, new_n695);
and_5  g00319(n2802, n2530, new_n696);
xnor_4 g00320(new_n696, new_n695, new_n697);
xnor_4 g00321(new_n697, new_n694, new_n698);
and_5  g00322(new_n658_1, new_n655, new_n699);
nor_5  g00323(new_n664, new_n659, new_n700);
nor_5  g00324(new_n700, new_n699, new_n701);
xnor_4 g00325(new_n701, new_n698, new_n702);
nor_5  g00326(new_n665, new_n654, new_n703);
nor_5  g00327(new_n669, new_n666, new_n704);
nor_5  g00328(new_n704, new_n703, new_n705);
xor_4  g00329(new_n705, new_n702, new_n706);
xor_4  g00330(new_n706, new_n685, new_n707);
xnor_4 g00331(new_n707, new_n684, new_n708);
xnor_4 g00332(new_n708, new_n683, new_n709);
and_5  g00333(new_n651, new_n634, new_n710);
and_5  g00334(n7965, n5814, new_n711);
nand_5 g00335(n2393, n1980, new_n712);
and_5  g00336(n8028, n3986, new_n713);
and_5  g00337(n10848, n5860, new_n714);
xnor_4 g00338(new_n714, new_n713, new_n715);
xnor_4 g00339(new_n715, new_n712, new_n716);
nor_5  g00340(new_n646, new_n573, new_n717);
and_5  g00341(new_n646, new_n573, new_n718);
nor_5  g00342(new_n718, new_n645, new_n719);
or_5   g00343(new_n719, new_n717, new_n720);
xnor_4 g00344(new_n720, new_n716, new_n721);
and_5  g00345(n12704, n7388, new_n722);
and_5  g00346(n11892, n7294, new_n723);
xnor_4 g00347(new_n723, new_n722, new_n724);
xnor_4 g00348(new_n724, new_n721, new_n725);
nor_5  g00349(new_n643, new_n639, new_n726);
nor_5  g00350(new_n648, new_n644, new_n727);
nor_5  g00351(new_n727, new_n726, new_n728);
xnor_4 g00352(new_n728, new_n725, new_n729);
nor_5  g00353(new_n649, new_n638, new_n730);
nand_5 g00354(new_n649, new_n638, new_n731);
and_5  g00355(new_n731, new_n637, new_n732);
or_5   g00356(new_n732, new_n730, new_n733);
xor_4  g00357(new_n733, new_n729, new_n734);
xor_4  g00358(new_n734, new_n711, new_n735);
xnor_4 g00359(new_n735, new_n710, new_n736);
xor_4  g00360(new_n736, new_n709, new_n737);
xor_4  g00361(new_n737, new_n680, new_n738);
xnor_4 g00362(new_n463, new_n462, new_n739);
xnor_4 g00363(new_n739, new_n474, new_n740);
nor_5  g00364(new_n740, new_n738, new_n741);
xnor_4 g00365(new_n473, new_n472, new_n742);
xor_4  g00366(new_n677, new_n676, new_n743);
nor_5  g00367(new_n743, new_n742, new_n744);
xnor_4 g00368(new_n743, new_n742, new_n745);
xnor_4 g00369(new_n471, new_n466, new_n746);
xor_4  g00370(new_n630, new_n629, new_n747);
nor_5  g00371(new_n747, new_n746, new_n748);
xnor_4 g00372(new_n595, new_n594, new_n749);
and_5  g00373(n6038, n5305, new_n750);
nor_5  g00374(new_n750, new_n424, new_n751);
nor_5  g00375(new_n751, new_n467, new_n752);
nor_5  g00376(new_n750, new_n425, new_n753_1);
nor_5  g00377(new_n753_1, new_n752, new_n754);
nor_5  g00378(new_n754, new_n749, new_n755);
xnor_4 g00379(new_n754, new_n749, new_n756);
xnor_4 g00380(new_n547, new_n494, new_n757);
and_5  g00381(new_n757, new_n750, new_n758);
xor_4  g00382(new_n469, new_n468, new_n759);
nor_5  g00383(new_n759, new_n758, new_n760);
xor_4  g00384(new_n562, new_n561, new_n761);
xor_4  g00385(new_n759, new_n758, new_n762);
and_5  g00386(new_n762, new_n761, new_n763);
nor_5  g00387(new_n763, new_n760, new_n764);
nor_5  g00388(new_n764, new_n756, new_n765);
or_5   g00389(new_n765, new_n755, new_n766);
xnor_4 g00390(new_n747, new_n746, new_n767);
nor_5  g00391(new_n767, new_n766, new_n768);
nor_5  g00392(new_n768, new_n748, new_n769);
nor_5  g00393(new_n769, new_n745, new_n770);
nor_5  g00394(new_n770, new_n744, new_n771);
xnor_4 g00395(new_n740, new_n738, new_n772);
nor_5  g00396(new_n772, new_n771, new_n773);
nor_5  g00397(new_n773, new_n741, new_n774);
xnor_4 g00398(new_n774, new_n477, new_n775);
or_5   g00399(new_n538, new_n535, new_n776);
nor_5  g00400(new_n522, new_n519, new_n777);
nor_5  g00401(new_n526, new_n523, new_n778);
or_5   g00402(new_n778, new_n777, new_n779);
and_5  g00403(n6776, n4928, new_n780);
and_5  g00404(n12299, n4141, new_n781);
and_5  g00405(n8759, n8236, new_n782);
xnor_4 g00406(new_n782, new_n781, new_n783_1);
xnor_4 g00407(new_n783_1, new_n780, new_n784);
xnor_4 g00408(new_n784, new_n779, new_n785);
and_5  g00409(new_n521_1, new_n520, new_n786);
and_5  g00410(n7436, n5105, new_n787);
xnor_4 g00411(new_n787, new_n786, new_n788);
nand_5 g00412(n9241, n7500, new_n789);
and_5  g00413(n8276, n1209, new_n790);
and_5  g00414(n10510, n7354, new_n791);
xnor_4 g00415(new_n791, new_n790, new_n792);
xnor_4 g00416(new_n792, new_n789, new_n793);
xor_4  g00417(new_n793, new_n788, new_n794);
xor_4  g00418(new_n794, new_n785, new_n795);
nor_5  g00419(new_n530, new_n527, new_n796);
nand_5 g00420(new_n529, new_n528, new_n797);
or_5   g00421(new_n534, new_n531, new_n798);
xor_4  g00422(new_n798, new_n797, new_n799);
nor_5  g00423(new_n799, new_n796, new_n800);
xnor_4 g00424(new_n800, new_n795, new_n801);
xnor_4 g00425(new_n801, new_n776, new_n802);
nor_5  g00426(new_n539, new_n518, new_n803);
nor_5  g00427(new_n540, new_n517, new_n804);
nor_5  g00428(new_n804, new_n803, new_n805);
xnor_4 g00429(new_n805, new_n802, new_n806_1);
or_5   g00430(new_n705, new_n702, new_n807);
nor_5  g00431(new_n689, new_n686, new_n808);
nor_5  g00432(new_n693, new_n690, new_n809);
or_5   g00433(new_n809, new_n808, new_n810);
and_5  g00434(n8476, n5069, new_n811);
and_5  g00435(n6806, n2530, new_n812);
and_5  g00436(n12044, n5331, new_n813);
xnor_4 g00437(new_n813, new_n812, new_n814);
xnor_4 g00438(new_n814, new_n811, new_n815);
xnor_4 g00439(new_n815, new_n810, new_n816);
and_5  g00440(new_n688, new_n687, new_n817);
and_5  g00441(n12648, n2802, new_n818);
xnor_4 g00442(new_n818, new_n817, new_n819);
and_5  g00443(n7690, n1512, new_n820);
and_5  g00444(n10545, n533, new_n821);
and_5  g00445(n3616, n1564, new_n822);
xnor_4 g00446(new_n822, new_n821, new_n823);
xor_4  g00447(new_n823, new_n820, new_n824);
xor_4  g00448(new_n824, new_n819, new_n825);
xor_4  g00449(new_n825, new_n816, new_n826);
nor_5  g00450(new_n697, new_n694, new_n827);
nand_5 g00451(new_n696, new_n695, new_n828);
or_5   g00452(new_n701, new_n698, new_n829);
xor_4  g00453(new_n829, new_n828, new_n830);
nor_5  g00454(new_n830, new_n827, new_n831);
xnor_4 g00455(new_n831, new_n826, new_n832);
xnor_4 g00456(new_n832, new_n807, new_n833);
and_5  g00457(new_n706, new_n685, new_n834);
nor_5  g00458(new_n706, new_n685, new_n835);
nor_5  g00459(new_n835, new_n684, new_n836);
nor_5  g00460(new_n836, new_n834, new_n837_1);
xor_4  g00461(new_n837_1, new_n833, new_n838);
nor_5  g00462(new_n733, new_n729, new_n839);
nor_5  g00463(new_n715, new_n712, new_n840);
nor_5  g00464(new_n720, new_n716, new_n841);
or_5   g00465(new_n841, new_n840, new_n842);
and_5  g00466(n7388, n5814, new_n843);
and_5  g00467(n12704, n11892, new_n844_1);
and_5  g00468(n7965, n4903, new_n845);
xnor_4 g00469(new_n845, new_n844_1, new_n846);
xnor_4 g00470(new_n846, new_n843, new_n847);
xnor_4 g00471(new_n847, new_n842, new_n848);
and_5  g00472(new_n714, new_n713, new_n849);
and_5  g00473(n7294, n2393, new_n850);
xnor_4 g00474(new_n850, new_n849, new_n851);
and_5  g00475(n10848, n3986, new_n852);
and_5  g00476(n5860, n1980, new_n853);
and_5  g00477(n8028, n5857, new_n854);
xnor_4 g00478(new_n854, new_n853, new_n855);
xor_4  g00479(new_n855, new_n852, new_n856);
xor_4  g00480(new_n856, new_n851, new_n857);
xor_4  g00481(new_n857, new_n848, new_n858);
nor_5  g00482(new_n724, new_n721, new_n859);
nand_5 g00483(new_n723, new_n722, new_n860);
or_5   g00484(new_n728, new_n725, new_n861);
xor_4  g00485(new_n861, new_n860, new_n862);
nor_5  g00486(new_n862, new_n859, new_n863);
xor_4  g00487(new_n863, new_n858, new_n864);
xnor_4 g00488(new_n864, new_n839, new_n865);
nor_5  g00489(new_n734, new_n711, new_n866);
and_5  g00490(new_n734, new_n711, new_n867);
nor_5  g00491(new_n867, new_n710, new_n868);
or_5   g00492(new_n868, new_n866, new_n869);
xor_4  g00493(new_n869, new_n865, new_n870);
xnor_4 g00494(new_n870, new_n838, new_n871);
and_5  g00495(new_n708, new_n683, new_n872);
nor_5  g00496(new_n708, new_n683, new_n873);
nor_5  g00497(new_n736, new_n873, new_n874);
or_5   g00498(new_n874, new_n872, new_n875);
xor_4  g00499(new_n875, new_n871, new_n876);
xnor_4 g00500(new_n876, new_n806_1, new_n877);
nor_5  g00501(new_n679, new_n541, new_n878);
nor_5  g00502(new_n737, new_n680, new_n879);
or_5   g00503(new_n879, new_n878, new_n880);
xnor_4 g00504(new_n880, new_n877, new_n881);
xor_4  g00505(new_n881, new_n775, n226);
nand_5 g00506(n5305, n4634, new_n883);
and_5  g00507(n10223, n5305, new_n884);
and_5  g00508(n7265, n1097, new_n885);
nor_5  g00509(new_n885, new_n884, new_n886);
and_5  g00510(n7265, n5305, new_n887);
and_5  g00511(n10223, n1097, new_n888);
and_5  g00512(new_n888, new_n887, new_n889);
and_5  g00513(n5964, n2879, new_n890);
nor_5  g00514(new_n890, new_n889, new_n891);
or_5   g00515(new_n891, new_n886, new_n892);
xnor_4 g00516(new_n892, new_n883, new_n893);
and_5  g00517(n2879, n1097, new_n894);
and_5  g00518(n10223, n5964, new_n895);
and_5  g00519(n7265, n4312, new_n896);
xnor_4 g00520(new_n896, new_n895, new_n897);
xor_4  g00521(new_n897, new_n894, new_n898);
xnor_4 g00522(new_n898, new_n893, new_n899);
nand_5 g00523(n5964, n2879, new_n900);
or_5   g00524(new_n900, new_n887, new_n901);
or_5   g00525(new_n889, new_n886, new_n902);
and_5  g00526(new_n902, new_n901, new_n903);
nand_5 g00527(new_n903, new_n890, new_n904);
xnor_4 g00528(new_n904, new_n899, new_n905);
nor_5  g00529(new_n901, new_n886, new_n906);
or_5   g00530(new_n906, new_n903, new_n907);
nand_5 g00531(n8759, n7946, new_n908);
and_5  g00532(n5331, n2558, new_n909);
and_5  g00533(n9763, n7965, new_n910);
xnor_4 g00534(new_n910, new_n909, new_n911_1);
nor_5  g00535(new_n911_1, new_n908, new_n912);
and_5  g00536(n7946, n6776, new_n913);
and_5  g00537(n8759, n2024, new_n914);
xor_4  g00538(new_n914, new_n913, new_n915);
and_5  g00539(new_n915, new_n912, new_n916);
and_5  g00540(new_n910, new_n909, new_n917);
and_5  g00541(n9111, n7965, new_n918);
and_5  g00542(n9763, n7388, new_n919);
xor_4  g00543(new_n919, new_n918, new_n920);
xnor_4 g00544(new_n920, new_n917, new_n921);
and_5  g00545(n5331, n2498, new_n922);
and_5  g00546(n8476, n2558, new_n923);
xor_4  g00547(new_n923, new_n922, new_n924);
xor_4  g00548(new_n924, new_n921, new_n925);
xnor_4 g00549(new_n915, new_n912, new_n926);
nor_5  g00550(new_n926, new_n925, new_n927);
nor_5  g00551(new_n927, new_n916, new_n928);
and_5  g00552(n8759, n7946, new_n929);
nand_5 g00553(n6776, n2024, new_n930);
nor_5  g00554(new_n930, new_n929, new_n931);
and_5  g00555(n12299, n7946, new_n932);
and_5  g00556(n9189, n8759, new_n933);
xor_4  g00557(new_n933, new_n932, new_n934);
or_5   g00558(new_n934, new_n931, new_n935);
or_5   g00559(new_n930, new_n929, new_n936);
nor_5  g00560(new_n933, new_n932, new_n937);
or_5   g00561(new_n937, new_n936, new_n938);
nand_5 g00562(new_n938, new_n935, new_n939);
xnor_4 g00563(new_n939, new_n928, new_n940);
nor_5  g00564(new_n920, new_n917, new_n941);
nor_5  g00565(new_n924, new_n921, new_n942);
nor_5  g00566(new_n942, new_n941, new_n943);
nand_5 g00567(n9111, n7388, new_n944);
or_5   g00568(new_n944, new_n910, new_n945);
and_5  g00569(n11892, n3342, new_n946);
and_5  g00570(new_n946, new_n910, new_n947);
and_5  g00571(n11892, n9763, new_n948);
and_5  g00572(n7965, n3342, new_n949);
nor_5  g00573(new_n949, new_n948, new_n950);
or_5   g00574(new_n950, new_n947, new_n951);
nand_5 g00575(new_n951, new_n945, new_n952);
or_5   g00576(new_n950, new_n945, new_n953);
and_5  g00577(new_n953, new_n952, new_n954);
xnor_4 g00578(new_n954, new_n943, new_n955);
nand_5 g00579(n8476, n2498, new_n956);
or_5   g00580(new_n956, new_n909, new_n957);
and_5  g00581(n2558, n2530, new_n958);
and_5  g00582(n5579, n5331, new_n959);
or_5   g00583(new_n959, new_n958, new_n960);
nor_5  g00584(new_n960, new_n957, new_n961);
nor_5  g00585(new_n959, new_n958, new_n962);
and_5  g00586(n5579, n2530, new_n963);
and_5  g00587(new_n963, new_n909, new_n964);
nor_5  g00588(new_n964, new_n962, new_n965);
and_5  g00589(new_n965, new_n957, new_n966);
or_5   g00590(new_n966, new_n961, new_n967);
xnor_4 g00591(new_n967, new_n955, new_n968);
xor_4  g00592(new_n968, new_n940, new_n969);
nor_5  g00593(new_n969, new_n907, new_n970);
xnor_4 g00594(new_n911_1, new_n929, new_n971);
and_5  g00595(new_n971, new_n887, new_n972);
and_5  g00596(n7265, n5964, new_n973);
and_5  g00597(n5305, n2879, new_n974);
xor_4  g00598(new_n974, new_n973, new_n975);
nor_5  g00599(new_n975, new_n972, new_n976);
xnor_4 g00600(new_n926, new_n925, new_n977);
xor_4  g00601(new_n975, new_n972, new_n978);
and_5  g00602(new_n978, new_n977, new_n979);
or_5   g00603(new_n979, new_n976, new_n980);
xnor_4 g00604(new_n969, new_n907, new_n981);
nor_5  g00605(new_n981, new_n980, new_n982);
nor_5  g00606(new_n982, new_n970, new_n983);
xnor_4 g00607(new_n983, new_n905, new_n984);
nand_5 g00608(n8759, n2522, new_n985);
nand_5 g00609(new_n933, new_n932, new_n986);
and_5  g00610(new_n986, new_n930, new_n987);
or_5   g00611(new_n987, new_n937, new_n988);
xnor_4 g00612(new_n988, new_n985, new_n989);
and_5  g00613(n12299, n2024, new_n990);
and_5  g00614(n7946, n7436, new_n991);
and_5  g00615(n9189, n6776, new_n992_1);
xnor_4 g00616(new_n992_1, new_n991, new_n993);
xor_4  g00617(new_n993, new_n990, new_n994);
xnor_4 g00618(new_n994, new_n989, new_n995);
or_5   g00619(new_n935, new_n930, new_n996_1);
xnor_4 g00620(new_n996_1, new_n995, new_n997);
and_5  g00621(new_n939, new_n928, new_n998);
nor_5  g00622(new_n968, new_n940, new_n999);
or_5   g00623(new_n999, new_n998, new_n1000);
xnor_4 g00624(new_n1000, new_n997, new_n1001);
nand_5 g00625(n5331, n521, new_n1002);
and_5  g00626(n8476, n2498, new_n1003);
nor_5  g00627(new_n964, new_n1003, new_n1004);
or_5   g00628(new_n1004, new_n962, new_n1005);
xnor_4 g00629(new_n1005, new_n1002, new_n1006);
and_5  g00630(n2530, n2498, new_n1007);
and_5  g00631(n12648, n2558, new_n1008);
and_5  g00632(n8476, n5579, new_n1009);
xnor_4 g00633(new_n1009, new_n1008, new_n1010);
xor_4  g00634(new_n1010, new_n1007, new_n1011);
xnor_4 g00635(new_n1011, new_n1006, new_n1012);
nand_5 g00636(new_n923, new_n922, new_n1013);
or_5   g00637(new_n965, new_n1013, new_n1014);
xor_4  g00638(new_n1014, new_n1012, new_n1015);
nand_5 g00639(n7965, n806, new_n1016);
nor_5  g00640(new_n950, new_n944, new_n1017);
nor_5  g00641(new_n1017, new_n947, new_n1018);
xnor_4 g00642(new_n1018, new_n1016, new_n1019);
and_5  g00643(n11892, n9111, new_n1020_1);
and_5  g00644(n9763, n2393, new_n1021);
and_5  g00645(n7388, n3342, new_n1022);
xnor_4 g00646(new_n1022, new_n1021, new_n1023);
xor_4  g00647(new_n1023, new_n1020_1, new_n1024);
xnor_4 g00648(new_n1024, new_n1019, new_n1025);
or_5   g00649(new_n952, new_n944, new_n1026);
xor_4  g00650(new_n1026, new_n1025, new_n1027);
xnor_4 g00651(new_n1027, new_n1015, new_n1028);
nor_5  g00652(new_n954, new_n943, new_n1029);
nor_5  g00653(new_n967, new_n955, new_n1030);
nor_5  g00654(new_n1030, new_n1029, new_n1031);
xor_4  g00655(new_n1031, new_n1028, new_n1032);
xnor_4 g00656(new_n1032, new_n1001, new_n1033);
xor_4  g00657(new_n1033, new_n984, n381);
and_5  g00658(n7862, n6038, new_n1035);
and_5  g00659(n7354, n6877, new_n1036);
and_5  g00660(n4805, n1564, new_n1037);
and_5  g00661(n8028, n7236, new_n1038);
xnor_4 g00662(new_n1038, new_n1037, new_n1039);
xnor_4 g00663(new_n1039, new_n1036, new_n1040);
xor_4  g00664(new_n1040, new_n1035, n397);
nand_5 g00665(n6687, n4370, new_n1042);
and_5  g00666(n11407, n4189, new_n1043);
and_5  g00667(n11877, n6687, new_n1044);
nor_5  g00668(new_n1044, new_n1043, new_n1045);
and_5  g00669(new_n1044, new_n1043, new_n1046);
and_5  g00670(n5212, n2564, new_n1047);
nor_5  g00671(new_n1047, new_n1046, new_n1048);
or_5   g00672(new_n1048, new_n1045, new_n1049);
xnor_4 g00673(new_n1049, new_n1042, new_n1050);
and_5  g00674(n5212, n4189, new_n1051);
and_5  g00675(n11407, n6770, new_n1052);
and_5  g00676(n11877, n2564, new_n1053);
xnor_4 g00677(new_n1053, new_n1052, new_n1054);
xor_4  g00678(new_n1054, new_n1051, new_n1055);
xnor_4 g00679(new_n1055, new_n1050, new_n1056);
nand_5 g00680(n5212, n2564, new_n1057);
and_5  g00681(n11407, n6687, new_n1058);
or_5   g00682(new_n1058, new_n1057, new_n1059);
and_5  g00683(new_n1059, new_n1045, new_n1060);
nor_5  g00684(new_n1060, new_n1046, new_n1061);
or_5   g00685(new_n1061, new_n1057, new_n1062);
xor_4  g00686(new_n1062, new_n1056, new_n1063);
nand_5 g00687(n12709, n8336, new_n1064);
and_5  g00688(n11222, n10990, new_n1065);
and_5  g00689(n12489, n12069, new_n1066);
xnor_4 g00690(new_n1066, new_n1065, new_n1067_1);
nor_5  g00691(new_n1067_1, new_n1064, new_n1068);
and_5  g00692(n11728, n8336, new_n1069);
and_5  g00693(n12709, n10928, new_n1070);
xor_4  g00694(new_n1070, new_n1069, new_n1071);
nor_5  g00695(new_n1071, new_n1068, new_n1072);
and_5  g00696(new_n1066, new_n1065, new_n1073);
and_5  g00697(n11222, n5760, new_n1074);
and_5  g00698(n11153, n10990, new_n1075);
xor_4  g00699(new_n1075, new_n1074, new_n1076);
xnor_4 g00700(new_n1076, new_n1073, new_n1077);
and_5  g00701(n12069, n7159, new_n1078);
and_5  g00702(n12489, n12391, new_n1079);
xnor_4 g00703(new_n1079, new_n1078, new_n1080);
xor_4  g00704(new_n1080, new_n1077, new_n1081);
xnor_4 g00705(new_n1071, new_n1068, new_n1082);
nor_5  g00706(new_n1082, new_n1081, new_n1083);
nor_5  g00707(new_n1083, new_n1072, new_n1084);
and_5  g00708(n12709, n8336, new_n1085);
nand_5 g00709(n11728, n10928, new_n1086);
or_5   g00710(new_n1086, new_n1085, new_n1087);
and_5  g00711(n6986, n6429, new_n1088);
and_5  g00712(new_n1088, new_n1085, new_n1089);
and_5  g00713(n12709, n6986, new_n1090);
and_5  g00714(n8336, n6429, new_n1091);
nor_5  g00715(new_n1091, new_n1090, new_n1092);
or_5   g00716(new_n1092, new_n1089, new_n1093);
nand_5 g00717(new_n1093, new_n1087, new_n1094_1);
or_5   g00718(new_n1092, new_n1087, new_n1095);
and_5  g00719(new_n1095, new_n1094_1, new_n1096);
xnor_4 g00720(new_n1096, new_n1084, new_n1097_1);
nand_5 g00721(n12391, n7159, new_n1098);
or_5   g00722(new_n1098, new_n1066, new_n1099);
and_5  g00723(n12489, n7891, new_n1100);
and_5  g00724(n12777, n12069, new_n1101);
nor_5  g00725(new_n1101, new_n1100, new_n1102);
and_5  g00726(new_n1102, new_n1099, new_n1103);
and_5  g00727(new_n1101, new_n1100, new_n1104);
nor_5  g00728(new_n1104, new_n1103, new_n1105);
or_5   g00729(new_n1102, new_n1099, new_n1106);
and_5  g00730(new_n1106, new_n1105, new_n1107);
nand_5 g00731(n11153, n5760, new_n1108);
nor_5  g00732(new_n1108, new_n1065, new_n1109);
and_5  g00733(n10990, n5314, new_n1110);
and_5  g00734(n11222, n1478, new_n1111);
xor_4  g00735(new_n1111, new_n1110, new_n1112);
or_5   g00736(new_n1112, new_n1109, new_n1113);
or_5   g00737(new_n1108, new_n1065, new_n1114);
nor_5  g00738(new_n1111, new_n1110, new_n1115);
or_5   g00739(new_n1115, new_n1114, new_n1116);
and_5  g00740(new_n1116, new_n1113, new_n1117);
xnor_4 g00741(new_n1117, new_n1107, new_n1118);
and_5  g00742(new_n1076, new_n1073, new_n1119);
nor_5  g00743(new_n1080, new_n1077, new_n1120);
nor_5  g00744(new_n1120, new_n1119, new_n1121);
xor_4  g00745(new_n1121, new_n1118, new_n1122);
xnor_4 g00746(new_n1122, new_n1097_1, new_n1123);
or_5   g00747(new_n1059, new_n1045, new_n1124);
and_5  g00748(new_n1124, new_n1061, new_n1125);
nor_5  g00749(new_n1125, new_n1123, new_n1126);
xnor_4 g00750(new_n1125, new_n1123, new_n1127);
xnor_4 g00751(new_n1067_1, new_n1085, new_n1128);
and_5  g00752(new_n1128, new_n1058, new_n1129);
and_5  g00753(n11407, n2564, new_n1130);
and_5  g00754(n6687, n5212, new_n1131);
xor_4  g00755(new_n1131, new_n1130, new_n1132);
nor_5  g00756(new_n1132, new_n1129, new_n1133);
xor_4  g00757(new_n1082, new_n1081, new_n1134);
xor_4  g00758(new_n1132, new_n1129, new_n1135);
and_5  g00759(new_n1135, new_n1134, new_n1136_1);
nor_5  g00760(new_n1136_1, new_n1133, new_n1137);
nor_5  g00761(new_n1137, new_n1127, new_n1138_1);
nor_5  g00762(new_n1138_1, new_n1126, new_n1139);
xnor_4 g00763(new_n1139, new_n1063, new_n1140);
nand_5 g00764(n8819, n8336, new_n1141);
and_5  g00765(n11728, n6986, new_n1142);
and_5  g00766(n10928, n6429, new_n1143);
and_5  g00767(n12709, n2226, new_n1144);
xnor_4 g00768(new_n1144, new_n1143, new_n1145);
xor_4  g00769(new_n1145, new_n1142, new_n1146);
xnor_4 g00770(new_n1146, new_n1141, new_n1147);
nor_5  g00771(new_n1092, new_n1086, new_n1148);
nor_5  g00772(new_n1148, new_n1089, new_n1149);
xnor_4 g00773(new_n1149, new_n1147, new_n1150);
or_5   g00774(new_n1094_1, new_n1086, new_n1151);
xnor_4 g00775(new_n1151, new_n1150, new_n1152);
and_5  g00776(n12069, n6254, new_n1153);
and_5  g00777(n12391, n7159, new_n1154);
nor_5  g00778(new_n1104, new_n1154, new_n1155);
nor_5  g00779(new_n1155, new_n1102, new_n1156);
xnor_4 g00780(new_n1156, new_n1153, new_n1157);
and_5  g00781(n12489, n7160, new_n1158);
and_5  g00782(n12777, n12391, new_n1159);
and_5  g00783(n7891, n7159, new_n1160);
xnor_4 g00784(new_n1160, new_n1159, new_n1161);
xor_4  g00785(new_n1161, new_n1158, new_n1162);
xnor_4 g00786(new_n1162, new_n1157, new_n1163);
or_5   g00787(new_n1105, new_n1098, new_n1164);
xor_4  g00788(new_n1164, new_n1163, new_n1165);
and_5  g00789(n11791, n11222, new_n1166);
nand_5 g00790(new_n1111, new_n1110, new_n1167);
and_5  g00791(new_n1167, new_n1108, new_n1168);
nor_5  g00792(new_n1168, new_n1115, new_n1169);
xnor_4 g00793(new_n1169, new_n1166, new_n1170);
and_5  g00794(n5760, n5314, new_n1171);
and_5  g00795(n10990, n996, new_n1172);
and_5  g00796(n11153, n1478, new_n1173);
xnor_4 g00797(new_n1173, new_n1172, new_n1174);
xor_4  g00798(new_n1174, new_n1171, new_n1175);
xnor_4 g00799(new_n1175, new_n1170, new_n1176);
or_5   g00800(new_n1113, new_n1108, new_n1177);
xor_4  g00801(new_n1177, new_n1176, new_n1178);
xnor_4 g00802(new_n1178, new_n1165, new_n1179);
and_5  g00803(new_n1117, new_n1107, new_n1180);
nor_5  g00804(new_n1121, new_n1118, new_n1181);
or_5   g00805(new_n1181, new_n1180, new_n1182);
xor_4  g00806(new_n1182, new_n1179, new_n1183);
xnor_4 g00807(new_n1183, new_n1152, new_n1184);
nor_5  g00808(new_n1096, new_n1084, new_n1185);
nor_5  g00809(new_n1122, new_n1097_1, new_n1186);
or_5   g00810(new_n1186, new_n1185, new_n1187);
xnor_4 g00811(new_n1187, new_n1184, new_n1188);
xor_4  g00812(new_n1188, new_n1140, n658);
and_5  g00813(n7862, n2585, new_n1190);
nand_5 g00814(n2508, n1333, new_n1191);
and_5  g00815(n11757, n6038, new_n1192);
and_5  g00816(n12720, n1333, new_n1193);
nor_5  g00817(new_n1193, new_n1192, new_n1194);
nand_5 g00818(new_n1193, new_n1192, new_n1195);
nand_5 g00819(n3172, n2509, new_n1196);
and_5  g00820(new_n1196, new_n1195, new_n1197);
or_5   g00821(new_n1197, new_n1194, new_n1198_1);
xnor_4 g00822(new_n1198_1, new_n1191, new_n1199_1);
and_5  g00823(n11757, n2509, new_n1200);
and_5  g00824(n6038, n5240, new_n1201);
and_5  g00825(n12720, n3172, new_n1202);
xnor_4 g00826(new_n1202, new_n1201, new_n1203);
xor_4  g00827(new_n1203, new_n1200, new_n1204);
xor_4  g00828(new_n1204, new_n1199_1, new_n1205);
nor_5  g00829(new_n1205, new_n1190, new_n1206);
xnor_4 g00830(new_n1205, new_n1190, new_n1207);
nand_5 g00831(n7862, n2508, new_n1208);
nand_5 g00832(n2509, n1333, new_n1209_1);
and_5  g00833(n6038, n3172, new_n1210);
and_5  g00834(n12720, n7862, new_n1211);
nor_5  g00835(new_n1211, new_n1210, new_n1212);
or_5   g00836(new_n1212, new_n1209_1, new_n1213);
nand_5 g00837(new_n1211, new_n1210, new_n1214);
and_5  g00838(new_n1214, new_n1213, new_n1215);
nor_5  g00839(new_n1215, new_n1208, new_n1216);
xnor_4 g00840(new_n1215, new_n1208, new_n1217);
xnor_4 g00841(new_n1193, new_n1192, new_n1218);
xnor_4 g00842(new_n1218, new_n1196, new_n1219);
nor_5  g00843(new_n1219, new_n1217, new_n1220);
or_5   g00844(new_n1220, new_n1216, new_n1221);
nor_5  g00845(new_n1221, new_n1207, new_n1222);
or_5   g00846(new_n1222, new_n1206, new_n1223);
nand_5 g00847(n12720, n11757, new_n1224);
and_5  g00848(n5240, n2509, new_n1225);
and_5  g00849(n11821, n6038, new_n1226);
xnor_4 g00850(new_n1226, new_n1225, new_n1227);
xnor_4 g00851(new_n1227, new_n1224, new_n1228);
nor_5  g00852(new_n1202, new_n1201, new_n1229);
nor_5  g00853(new_n1203, new_n1200, new_n1230);
or_5   g00854(new_n1230, new_n1229, new_n1231);
xnor_4 g00855(new_n1231, new_n1228, new_n1232);
nor_5  g00856(new_n1198_1, new_n1191, new_n1233);
nor_5  g00857(new_n1204, new_n1199_1, new_n1234);
nor_5  g00858(new_n1234, new_n1233, new_n1235);
and_5  g00859(n2585, n1333, new_n1236);
and_5  g00860(n3172, n2508, new_n1237);
xnor_4 g00861(new_n1237, new_n1236, new_n1238);
xnor_4 g00862(new_n1238, new_n1235, new_n1239);
xnor_4 g00863(new_n1239, new_n1232, new_n1240);
or_5   g00864(new_n1240, new_n1223, new_n1241);
nor_5  g00865(new_n1238, new_n1235, new_n1242);
nand_5 g00866(new_n1237, new_n1236, new_n1243);
and_5  g00867(new_n1238, new_n1235, new_n1244);
or_5   g00868(new_n1244, new_n1232, new_n1245);
xor_4  g00869(new_n1245, new_n1243, new_n1246);
nor_5  g00870(new_n1246, new_n1242, new_n1247);
and_5  g00871(new_n1226, new_n1225, new_n1248);
and_5  g00872(n11757, n2508, new_n1249);
xnor_4 g00873(new_n1249, new_n1248, new_n1250);
and_5  g00874(n11821, n2509, new_n1251);
and_5  g00875(n12720, n5240, new_n1252);
and_5  g00876(n9080, n6038, new_n1253);
xnor_4 g00877(new_n1253, new_n1252, new_n1254);
xor_4  g00878(new_n1254, new_n1251, new_n1255);
xor_4  g00879(new_n1255, new_n1250, new_n1256);
nor_5  g00880(new_n1227, new_n1224, new_n1257);
nor_5  g00881(new_n1231, new_n1228, new_n1258);
or_5   g00882(new_n1258, new_n1257, new_n1259);
nand_5 g00883(n4005, n1333, new_n1260);
and_5  g00884(n3172, n2585, new_n1261);
and_5  g00885(n12706, n7862, new_n1262);
xnor_4 g00886(new_n1262, new_n1261, new_n1263);
xor_4  g00887(new_n1263, new_n1260, new_n1264);
xnor_4 g00888(new_n1264, new_n1259, new_n1265);
xor_4  g00889(new_n1265, new_n1256, new_n1266);
xnor_4 g00890(new_n1266, new_n1247, new_n1267);
xnor_4 g00891(new_n1267, new_n1241, new_n1268);
and_5  g00892(n7862, n4005, new_n1269_1);
xor_4  g00893(new_n1240, new_n1223, new_n1270);
and_5  g00894(new_n1270, new_n1269_1, new_n1271);
xnor_4 g00895(new_n1219, new_n1217, new_n1272);
xor_4  g00896(new_n1211, new_n1210, new_n1273);
and_5  g00897(n6038, n1333, new_n1274);
and_5  g00898(n7862, n2509, new_n1275);
nand_5 g00899(new_n1275, new_n1274, new_n1276);
or_5   g00900(new_n1276, new_n1273, new_n1277);
or_5   g00901(new_n1277, new_n1272, new_n1278);
xor_4  g00902(new_n1221, new_n1207, new_n1279);
nor_5  g00903(new_n1279, new_n1278, new_n1280);
xor_4  g00904(new_n1270, new_n1269_1, new_n1281);
and_5  g00905(new_n1281, new_n1280, new_n1282);
nor_5  g00906(new_n1282, new_n1271, new_n1283);
xnor_4 g00907(new_n1283, new_n1268, new_n1284);
nand_5 g00908(n6877, n5105, new_n1285);
and_5  g00909(n6877, n1209, new_n1286);
and_5  g00910(n7354, n2464, new_n1287);
and_5  g00911(new_n1287, new_n1286, new_n1288);
nor_5  g00912(new_n1287, new_n1286, new_n1289);
nand_5 g00913(n9400, n7500, new_n1290);
nor_5  g00914(new_n1290, new_n1289, new_n1291);
nor_5  g00915(new_n1291, new_n1288, new_n1292);
xnor_4 g00916(new_n1292, new_n1285, new_n1293);
and_5  g00917(n7500, n2464, new_n1294);
and_5  g00918(n9400, n1209, new_n1295);
and_5  g00919(n11311, n7354, new_n1296);
xnor_4 g00920(new_n1296, new_n1295, new_n1297);
xor_4  g00921(new_n1297, new_n1294, new_n1298);
xnor_4 g00922(new_n1298, new_n1293, new_n1299);
xnor_4 g00923(new_n1287, new_n1286, new_n1300);
and_5  g00924(n9400, n7354, new_n1301);
and_5  g00925(n7500, n6877, new_n1302);
and_5  g00926(new_n1302, new_n1301, new_n1303);
nand_5 g00927(new_n1303, new_n1300, new_n1304);
or_5   g00928(new_n1304, new_n1299, new_n1305);
and_5  g00929(n11311, n7500, new_n1306);
and_5  g00930(n2464, n1209, new_n1307);
and_5  g00931(n7354, n4187, new_n1308);
xnor_4 g00932(new_n1308, new_n1307, new_n1309);
xor_4  g00933(new_n1309, new_n1306, new_n1310);
nand_5 g00934(n9400, n5105, new_n1311);
nor_5  g00935(new_n1296, new_n1295, new_n1312);
and_5  g00936(new_n1296, new_n1295, new_n1313);
nor_5  g00937(new_n1313, new_n1294, new_n1314);
or_5   g00938(new_n1314, new_n1312, new_n1315);
xnor_4 g00939(new_n1315, new_n1311, new_n1316);
xor_4  g00940(new_n1316, new_n1310, new_n1317);
and_5  g00941(n6877, n4141, new_n1318);
nor_5  g00942(new_n1292, new_n1285, new_n1319);
nor_5  g00943(new_n1298, new_n1293, new_n1320);
or_5   g00944(new_n1320, new_n1319, new_n1321);
xnor_4 g00945(new_n1321, new_n1318, new_n1322);
xor_4  g00946(new_n1322, new_n1317, new_n1323);
or_5   g00947(new_n1323, new_n1305, new_n1324);
and_5  g00948(n6877, n4928, new_n1325);
nor_5  g00949(new_n1321, new_n1318, new_n1326);
nor_5  g00950(new_n1322, new_n1317, new_n1327);
or_5   g00951(new_n1327, new_n1326, new_n1328);
nand_5 g00952(n11311, n1209, new_n1329);
and_5  g00953(n7500, n4187, new_n1330);
and_5  g00954(n7354, n4203, new_n1331);
xnor_4 g00955(new_n1331, new_n1330, new_n1332);
xnor_4 g00956(new_n1332, new_n1329, new_n1333_1);
nor_5  g00957(new_n1308, new_n1307, new_n1334);
nor_5  g00958(new_n1309, new_n1306, new_n1335);
or_5   g00959(new_n1335, new_n1334, new_n1336);
xnor_4 g00960(new_n1336, new_n1333_1, new_n1337);
nor_5  g00961(new_n1315, new_n1311, new_n1338);
nor_5  g00962(new_n1316, new_n1310, new_n1339);
nor_5  g00963(new_n1339, new_n1338, new_n1340);
and_5  g00964(n9400, n4141, new_n1341);
and_5  g00965(n5105, n2464, new_n1342);
xnor_4 g00966(new_n1342, new_n1341, new_n1343);
xnor_4 g00967(new_n1343, new_n1340, new_n1344);
xnor_4 g00968(new_n1344, new_n1337, new_n1345);
xor_4  g00969(new_n1345, new_n1328, new_n1346);
xnor_4 g00970(new_n1346, new_n1325, new_n1347);
xnor_4 g00971(new_n1347, new_n1324, new_n1348);
nand_5 g00972(n7294, n7236, new_n1349);
nand_5 g00973(n10848, n3992, new_n1350);
and_5  g00974(n8384, n8028, new_n1351);
and_5  g00975(n7236, n1980, new_n1352);
nor_5  g00976(new_n1352, new_n1351, new_n1353_1);
or_5   g00977(new_n1353_1, new_n1350, new_n1354);
nand_5 g00978(new_n1352, new_n1351, new_n1355);
and_5  g00979(new_n1355, new_n1354, new_n1356);
xnor_4 g00980(new_n1356, new_n1349, new_n1357_1);
and_5  g00981(n8028, n6358, new_n1358);
and_5  g00982(n10848, n8384, new_n1359);
and_5  g00983(n3992, n1980, new_n1360);
xnor_4 g00984(new_n1360, new_n1359, new_n1361);
xor_4  g00985(new_n1361, new_n1358, new_n1362);
xnor_4 g00986(new_n1362, new_n1357_1, new_n1363);
xor_4  g00987(new_n1352, new_n1351, new_n1364);
and_5  g00988(n10848, n7236, new_n1365);
and_5  g00989(n8028, n3992, new_n1366);
nand_5 g00990(new_n1366, new_n1365, new_n1367);
or_5   g00991(new_n1367, new_n1364, new_n1368);
or_5   g00992(new_n1368, new_n1363, new_n1369);
and_5  g00993(n10848, n6358, new_n1370);
and_5  g00994(n8384, n1980, new_n1371);
and_5  g00995(n8028, n5198, new_n1372);
xnor_4 g00996(new_n1372, new_n1371, new_n1373);
xor_4  g00997(new_n1373, new_n1370, new_n1374);
and_5  g00998(n7294, n3992, new_n1375);
nor_5  g00999(new_n1360, new_n1359, new_n1376);
nor_5  g01000(new_n1361, new_n1358, new_n1377);
nor_5  g01001(new_n1377, new_n1376, new_n1378);
xnor_4 g01002(new_n1378, new_n1375, new_n1379);
xor_4  g01003(new_n1379, new_n1374, new_n1380);
nand_5 g01004(n12704, n7236, new_n1381);
nor_5  g01005(new_n1356, new_n1349, new_n1382);
nor_5  g01006(new_n1362, new_n1357_1, new_n1383);
nor_5  g01007(new_n1383, new_n1382, new_n1384);
xnor_4 g01008(new_n1384, new_n1381, new_n1385);
xor_4  g01009(new_n1385, new_n1380, new_n1386);
or_5   g01010(new_n1386, new_n1369, new_n1387);
and_5  g01011(n7236, n5814, new_n1388);
and_5  g01012(new_n1378, new_n1375, new_n1389);
nor_5  g01013(new_n1379, new_n1374, new_n1390);
nor_5  g01014(new_n1390, new_n1389, new_n1391);
and_5  g01015(n8384, n7294, new_n1392);
and_5  g01016(n12704, n3992, new_n1393);
xnor_4 g01017(new_n1393, new_n1392, new_n1394);
xnor_4 g01018(new_n1394, new_n1391, new_n1395);
and_5  g01019(n6358, n1980, new_n1396);
nor_5  g01020(new_n1372, new_n1371, new_n1397);
nor_5  g01021(new_n1373, new_n1370, new_n1398);
nor_5  g01022(new_n1398, new_n1397, new_n1399);
xnor_4 g01023(new_n1399, new_n1396, new_n1400);
and_5  g01024(n10848, n5198, new_n1401);
and_5  g01025(n8028, n1471, new_n1402);
xor_4  g01026(new_n1402, new_n1401, new_n1403);
xor_4  g01027(new_n1403, new_n1400, new_n1404);
xnor_4 g01028(new_n1404, new_n1395, new_n1405);
and_5  g01029(new_n1384, new_n1381, new_n1406);
nor_5  g01030(new_n1385, new_n1380, new_n1407);
or_5   g01031(new_n1407, new_n1406, new_n1408);
xor_4  g01032(new_n1408, new_n1405, new_n1409);
xnor_4 g01033(new_n1409, new_n1388, new_n1410);
xor_4  g01034(new_n1410, new_n1387, new_n1411);
nand_5 g01035(n4805, n2802, new_n1412);
and_5  g01036(n5283, n1564, new_n1413);
and_5  g01037(n4805, n533, new_n1414);
nand_5 g01038(new_n1414, new_n1413, new_n1415);
nor_5  g01039(new_n1414, new_n1413, new_n1416);
nand_5 g01040(n11478, n1512, new_n1417);
or_5   g01041(new_n1417, new_n1416, new_n1418);
and_5  g01042(new_n1418, new_n1415, new_n1419);
xnor_4 g01043(new_n1419, new_n1412, new_n1420);
and_5  g01044(n1564, n137, new_n1421);
and_5  g01045(n5283, n1512, new_n1422);
and_5  g01046(n11478, n533, new_n1423);
xnor_4 g01047(new_n1423, new_n1422, new_n1424);
xor_4  g01048(new_n1424, new_n1421, new_n1425);
xnor_4 g01049(new_n1425, new_n1420, new_n1426);
xor_4  g01050(new_n1414, new_n1413, new_n1427);
and_5  g01051(n4805, n1512, new_n1428);
and_5  g01052(n11478, n1564, new_n1429);
nand_5 g01053(new_n1429, new_n1428, new_n1430);
or_5   g01054(new_n1430, new_n1427, new_n1431);
or_5   g01055(new_n1431, new_n1426, new_n1432);
and_5  g01056(n6806, n4805, new_n1433);
and_5  g01057(n11478, n2802, new_n1434);
nor_5  g01058(new_n1423, new_n1422, new_n1435);
nor_5  g01059(new_n1424, new_n1421, new_n1436);
nor_5  g01060(new_n1436, new_n1435, new_n1437);
xnor_4 g01061(new_n1437, new_n1434, new_n1438);
and_5  g01062(n1512, n137, new_n1439);
and_5  g01063(n5283, n533, new_n1440);
and_5  g01064(n6294, n1564, new_n1441);
xnor_4 g01065(new_n1441, new_n1440, new_n1442);
xor_4  g01066(new_n1442, new_n1439, new_n1443);
xor_4  g01067(new_n1443, new_n1438, new_n1444);
xnor_4 g01068(new_n1444, new_n1433, new_n1445);
nor_5  g01069(new_n1419, new_n1412, new_n1446);
nor_5  g01070(new_n1425, new_n1420, new_n1447);
or_5   g01071(new_n1447, new_n1446, new_n1448);
xor_4  g01072(new_n1448, new_n1445, new_n1449);
or_5   g01073(new_n1449, new_n1432, new_n1450);
and_5  g01074(n5069, n4805, new_n1451);
nand_5 g01075(n533, n137, new_n1452);
and_5  g01076(n6294, n1512, new_n1453);
and_5  g01077(n6797, n1564, new_n1454);
xnor_4 g01078(new_n1454, new_n1453, new_n1455);
xnor_4 g01079(new_n1455, new_n1452, new_n1456);
nor_5  g01080(new_n1441, new_n1440, new_n1457);
nor_5  g01081(new_n1442, new_n1439, new_n1458);
or_5   g01082(new_n1458, new_n1457, new_n1459);
xnor_4 g01083(new_n1459, new_n1456, new_n1460);
and_5  g01084(n11478, n6806, new_n1461);
and_5  g01085(n5283, n2802, new_n1462);
xnor_4 g01086(new_n1462, new_n1461, new_n1463);
xnor_4 g01087(new_n1463, new_n1460, new_n1464);
and_5  g01088(new_n1437, new_n1434, new_n1465);
nor_5  g01089(new_n1443, new_n1438, new_n1466);
nor_5  g01090(new_n1466, new_n1465, new_n1467);
xnor_4 g01091(new_n1467, new_n1464, new_n1468);
nor_5  g01092(new_n1444, new_n1433, new_n1469);
nor_5  g01093(new_n1448, new_n1445, new_n1470);
or_5   g01094(new_n1470, new_n1469, new_n1471_1);
xor_4  g01095(new_n1471_1, new_n1468, new_n1472);
xnor_4 g01096(new_n1472, new_n1451, new_n1473);
xor_4  g01097(new_n1473, new_n1450, new_n1474);
xnor_4 g01098(new_n1474, new_n1411, new_n1475);
xor_4  g01099(new_n1386, new_n1369, new_n1476);
xor_4  g01100(new_n1431, new_n1426, new_n1477);
xor_4  g01101(new_n1368, new_n1363, new_n1478_1);
nor_5  g01102(new_n1478_1, new_n1477, new_n1479);
and_5  g01103(new_n1038, new_n1037, new_n1480);
xor_4  g01104(new_n1429, new_n1428, new_n1481);
nor_5  g01105(new_n1481, new_n1480, new_n1482);
xnor_4 g01106(new_n1481, new_n1480, new_n1483);
xor_4  g01107(new_n1366, new_n1365, new_n1484);
nor_5  g01108(new_n1484, new_n1483, new_n1485);
nor_5  g01109(new_n1485, new_n1482, new_n1486);
nor_5  g01110(new_n1417, new_n1037, new_n1487);
nor_5  g01111(new_n1487, new_n1427, new_n1488);
nor_5  g01112(new_n1418, new_n1037, new_n1489);
nor_5  g01113(new_n1489, new_n1488, new_n1490);
nor_5  g01114(new_n1490, new_n1486, new_n1491);
xnor_4 g01115(new_n1490, new_n1486, new_n1492);
nor_5  g01116(new_n1350, new_n1038, new_n1493);
nor_5  g01117(new_n1493, new_n1364, new_n1494);
nor_5  g01118(new_n1354, new_n1038, new_n1495);
nor_5  g01119(new_n1495, new_n1494, new_n1496);
nor_5  g01120(new_n1496, new_n1492, new_n1497);
nor_5  g01121(new_n1497, new_n1491, new_n1498);
xnor_4 g01122(new_n1478_1, new_n1477, new_n1499);
nor_5  g01123(new_n1499, new_n1498, new_n1500);
nor_5  g01124(new_n1500, new_n1479, new_n1501);
nor_5  g01125(new_n1501, new_n1476, new_n1502);
xor_4  g01126(new_n1449, new_n1432, new_n1503);
xnor_4 g01127(new_n1501, new_n1476, new_n1504);
nor_5  g01128(new_n1504, new_n1503, new_n1505);
nor_5  g01129(new_n1505, new_n1502, new_n1506);
xor_4  g01130(new_n1506, new_n1475, new_n1507);
and_5  g01131(new_n1507, new_n1348, new_n1508);
xnor_4 g01132(new_n1507, new_n1348, new_n1509);
xnor_4 g01133(new_n1323, new_n1305, new_n1510_1);
xor_4  g01134(new_n1504, new_n1503, new_n1511);
nor_5  g01135(new_n1511, new_n1510_1, new_n1512_1);
xnor_4 g01136(new_n1511, new_n1510_1, new_n1513);
xnor_4 g01137(new_n1304, new_n1299, new_n1514);
xor_4  g01138(new_n1499, new_n1498, new_n1515);
nor_5  g01139(new_n1515, new_n1514, new_n1516);
xnor_4 g01140(new_n1515, new_n1514, new_n1517);
xor_4  g01141(new_n1496, new_n1492, new_n1518);
nor_5  g01142(new_n1290, new_n1036, new_n1519);
and_5  g01143(new_n1519, new_n1289, new_n1520);
nor_5  g01144(new_n1519, new_n1300, new_n1521);
nor_5  g01145(new_n1521, new_n1520, new_n1522);
nor_5  g01146(new_n1522, new_n1518, new_n1523_1);
xnor_4 g01147(new_n1522, new_n1518, new_n1524);
xor_4  g01148(new_n1484, new_n1483, new_n1525);
xnor_4 g01149(new_n1302, new_n1301, new_n1526);
nor_5  g01150(new_n1526, new_n1525, new_n1527);
nand_5 g01151(n7354, n6877, new_n1528);
or_5   g01152(new_n1039, new_n1528, new_n1529);
xnor_4 g01153(new_n1526, new_n1525, new_n1530);
nor_5  g01154(new_n1530, new_n1529, new_n1531);
nor_5  g01155(new_n1531, new_n1527, new_n1532);
nor_5  g01156(new_n1532, new_n1524, new_n1533);
nor_5  g01157(new_n1533, new_n1523_1, new_n1534);
nor_5  g01158(new_n1534, new_n1517, new_n1535);
nor_5  g01159(new_n1535, new_n1516, new_n1536);
nor_5  g01160(new_n1536, new_n1513, new_n1537);
or_5   g01161(new_n1537, new_n1512_1, new_n1538);
nor_5  g01162(new_n1538, new_n1509, new_n1539);
nor_5  g01163(new_n1539, new_n1508, new_n1540);
or_5   g01164(new_n1345, new_n1328, new_n1541);
nor_5  g01165(new_n1332, new_n1329, new_n1542);
nor_5  g01166(new_n1336, new_n1333_1, new_n1543);
or_5   g01167(new_n1543, new_n1542, new_n1544);
nand_5 g01168(n9400, n4928, new_n1545);
and_5  g01169(n4141, n2464, new_n1546);
and_5  g01170(n8236, n6877, new_n1547);
xnor_4 g01171(new_n1547, new_n1546, new_n1548);
xor_4  g01172(new_n1548, new_n1545, new_n1549);
xnor_4 g01173(new_n1549, new_n1544, new_n1550);
and_5  g01174(new_n1331, new_n1330, new_n1551);
and_5  g01175(n11311, n5105, new_n1552);
xnor_4 g01176(new_n1552, new_n1551, new_n1553);
and_5  g01177(n7500, n4203, new_n1554);
and_5  g01178(n4187, n1209, new_n1555);
and_5  g01179(n12753, n7354, new_n1556);
xnor_4 g01180(new_n1556, new_n1555, new_n1557);
xor_4  g01181(new_n1557, new_n1554, new_n1558);
xor_4  g01182(new_n1558, new_n1553, new_n1559);
xor_4  g01183(new_n1559, new_n1550, new_n1560);
nor_5  g01184(new_n1343, new_n1340, new_n1561);
nand_5 g01185(new_n1342, new_n1341, new_n1562);
and_5  g01186(new_n1343, new_n1340, new_n1563);
or_5   g01187(new_n1563, new_n1337, new_n1564_1);
xor_4  g01188(new_n1564_1, new_n1562, new_n1565);
nor_5  g01189(new_n1565, new_n1561, new_n1566);
xnor_4 g01190(new_n1566, new_n1560, new_n1567);
xnor_4 g01191(new_n1567, new_n1541, new_n1568);
and_5  g01192(new_n1346, new_n1325, new_n1569);
nor_5  g01193(new_n1347, new_n1324, new_n1570);
nor_5  g01194(new_n1570, new_n1569, new_n1571);
xor_4  g01195(new_n1571, new_n1568, new_n1572);
or_5   g01196(new_n1408, new_n1405, new_n1573);
nor_5  g01197(new_n1399, new_n1396, new_n1574);
nor_5  g01198(new_n1403, new_n1400, new_n1575);
nor_5  g01199(new_n1575, new_n1574, new_n1576_1);
and_5  g01200(n5814, n3992, new_n1577);
and_5  g01201(n12704, n8384, new_n1578);
and_5  g01202(n7236, n4903, new_n1579);
xnor_4 g01203(new_n1579, new_n1578, new_n1580);
xnor_4 g01204(new_n1580, new_n1577, new_n1581);
xnor_4 g01205(new_n1581, new_n1576_1, new_n1582);
and_5  g01206(new_n1402, new_n1401, new_n1583);
and_5  g01207(n7294, n6358, new_n1584);
xnor_4 g01208(new_n1584, new_n1583, new_n1585);
and_5  g01209(n10848, n1471, new_n1586);
and_5  g01210(n5198, n1980, new_n1587);
and_5  g01211(n8028, n7646, new_n1588);
xnor_4 g01212(new_n1588, new_n1587, new_n1589);
xor_4  g01213(new_n1589, new_n1586, new_n1590);
xor_4  g01214(new_n1590, new_n1585, new_n1591);
xor_4  g01215(new_n1591, new_n1582, new_n1592);
nor_5  g01216(new_n1394, new_n1391, new_n1593);
nand_5 g01217(new_n1393, new_n1392, new_n1594);
or_5   g01218(new_n1404, new_n1395, new_n1595);
xor_4  g01219(new_n1595, new_n1594, new_n1596);
nor_5  g01220(new_n1596, new_n1593, new_n1597);
xnor_4 g01221(new_n1597, new_n1592, new_n1598);
xnor_4 g01222(new_n1598, new_n1573, new_n1599);
and_5  g01223(new_n1409, new_n1388, new_n1600);
nor_5  g01224(new_n1410, new_n1387, new_n1601);
nor_5  g01225(new_n1601, new_n1600, new_n1602);
xor_4  g01226(new_n1602, new_n1599, new_n1603);
and_5  g01227(new_n1472, new_n1451, new_n1604);
nor_5  g01228(new_n1473, new_n1450, new_n1605);
nor_5  g01229(new_n1605, new_n1604, new_n1606);
or_5   g01230(new_n1471_1, new_n1468, new_n1607);
nor_5  g01231(new_n1455, new_n1452, new_n1608);
nor_5  g01232(new_n1459, new_n1456, new_n1609);
or_5   g01233(new_n1609, new_n1608, new_n1610);
nand_5 g01234(n11478, n5069, new_n1611);
and_5  g01235(n6806, n5283, new_n1612);
and_5  g01236(n12044, n4805, new_n1613);
xnor_4 g01237(new_n1613, new_n1612, new_n1614);
xor_4  g01238(new_n1614, new_n1611, new_n1615);
xnor_4 g01239(new_n1615, new_n1610, new_n1616);
and_5  g01240(new_n1454, new_n1453, new_n1617);
and_5  g01241(n2802, n137, new_n1618);
xnor_4 g01242(new_n1618, new_n1617, new_n1619);
and_5  g01243(n6797, n1512, new_n1620);
and_5  g01244(n6294, n533, new_n1621);
and_5  g01245(n3146, n1564, new_n1622);
xnor_4 g01246(new_n1622, new_n1621, new_n1623);
xor_4  g01247(new_n1623, new_n1620, new_n1624);
xor_4  g01248(new_n1624, new_n1619, new_n1625);
xor_4  g01249(new_n1625, new_n1616, new_n1626);
nor_5  g01250(new_n1463, new_n1460, new_n1627);
nand_5 g01251(new_n1462, new_n1461, new_n1628);
or_5   g01252(new_n1467, new_n1464, new_n1629);
xor_4  g01253(new_n1629, new_n1628, new_n1630);
nor_5  g01254(new_n1630, new_n1627, new_n1631);
xnor_4 g01255(new_n1631, new_n1626, new_n1632);
xnor_4 g01256(new_n1632, new_n1607, new_n1633);
xor_4  g01257(new_n1633, new_n1606, new_n1634);
xnor_4 g01258(new_n1634, new_n1603, new_n1635);
nor_5  g01259(new_n1474, new_n1411, new_n1636);
nor_5  g01260(new_n1506, new_n1475, new_n1637);
nor_5  g01261(new_n1637, new_n1636, new_n1638);
xnor_4 g01262(new_n1638, new_n1635, new_n1639);
xnor_4 g01263(new_n1639, new_n1572, new_n1640);
xor_4  g01264(new_n1640, new_n1540, new_n1641);
nor_5  g01265(new_n1641, new_n1284, new_n1642);
xnor_4 g01266(new_n1641, new_n1284, new_n1643);
xnor_4 g01267(new_n1281, new_n1280, new_n1644);
xor_4  g01268(new_n1538, new_n1509, new_n1645);
nor_5  g01269(new_n1645, new_n1644, new_n1646);
xor_4  g01270(new_n1279, new_n1278, new_n1647);
xor_4  g01271(new_n1536, new_n1513, new_n1648);
nor_5  g01272(new_n1648, new_n1647, new_n1649);
xnor_4 g01273(new_n1648, new_n1647, new_n1650);
xor_4  g01274(new_n1277, new_n1272, new_n1651);
xor_4  g01275(new_n1534, new_n1517, new_n1652);
nor_5  g01276(new_n1652, new_n1651, new_n1653);
xor_4  g01277(new_n1532, new_n1524, new_n1654);
nor_5  g01278(new_n1209_1, new_n1035, new_n1655);
nor_5  g01279(new_n1655, new_n1273, new_n1656);
nor_5  g01280(new_n1213, new_n1035, new_n1657);
nor_5  g01281(new_n1657, new_n1656, new_n1658_1);
nor_5  g01282(new_n1658_1, new_n1654, new_n1659);
xnor_4 g01283(new_n1658_1, new_n1654, new_n1660);
and_5  g01284(new_n1040, new_n1035, new_n1661);
xor_4  g01285(new_n1275, new_n1274, new_n1662);
nor_5  g01286(new_n1662, new_n1661, new_n1663);
xnor_4 g01287(new_n1530, new_n1529, new_n1664);
xor_4  g01288(new_n1662, new_n1661, new_n1665);
and_5  g01289(new_n1665, new_n1664, new_n1666);
nor_5  g01290(new_n1666, new_n1663, new_n1667);
nor_5  g01291(new_n1667, new_n1660, new_n1668);
nor_5  g01292(new_n1668, new_n1659, new_n1669);
xnor_4 g01293(new_n1652, new_n1651, new_n1670);
nor_5  g01294(new_n1670, new_n1669, new_n1671);
nor_5  g01295(new_n1671, new_n1653, new_n1672);
nor_5  g01296(new_n1672, new_n1650, new_n1673);
or_5   g01297(new_n1673, new_n1649, new_n1674);
xnor_4 g01298(new_n1645, new_n1644, new_n1675);
nor_5  g01299(new_n1675, new_n1674, new_n1676);
nor_5  g01300(new_n1676, new_n1646, new_n1677);
nor_5  g01301(new_n1677, new_n1643, new_n1678);
nor_5  g01302(new_n1678, new_n1642, new_n1679);
nor_5  g01303(new_n1639, new_n1572, new_n1680);
nor_5  g01304(new_n1640, new_n1540, new_n1681);
nor_5  g01305(new_n1681, new_n1680, new_n1682);
nor_5  g01306(new_n1634, new_n1603, new_n1683);
nor_5  g01307(new_n1638, new_n1635, new_n1684);
nor_5  g01308(new_n1684, new_n1683, new_n1685);
nor_5  g01309(new_n1267, new_n1241, new_n1686);
nor_5  g01310(new_n1283, new_n1268, new_n1687);
nor_5  g01311(new_n1687, new_n1686, new_n1688);
nor_5  g01312(new_n1598, new_n1573, new_n1689);
nor_5  g01313(new_n1602, new_n1599, new_n1690);
or_5   g01314(new_n1690, new_n1689, new_n1691);
xnor_4 g01315(new_n1691, new_n1688, new_n1692);
nor_5  g01316(new_n1595, new_n1594, new_n1693);
nor_5  g01317(new_n1597, new_n1592, new_n1694);
nor_5  g01318(new_n1694, new_n1693, new_n1695);
and_5  g01319(new_n1618, new_n1617, new_n1696);
nor_5  g01320(new_n1624, new_n1619, new_n1697);
nor_5  g01321(new_n1697, new_n1696, new_n1698);
and_5  g01322(n7862, n615, new_n1699);
and_5  g01323(n4903, n3992, new_n1700);
and_5  g01324(n6806, n137, new_n1701);
xnor_4 g01325(new_n1701, new_n1700, new_n1702);
xnor_4 g01326(new_n1702, new_n1699, new_n1703);
xnor_4 g01327(new_n1703, new_n1698, new_n1704);
and_5  g01328(n6797, n533, new_n1705);
and_5  g01329(n8384, n5814, new_n1706);
xnor_4 g01330(new_n1706, new_n1705, new_n1707);
and_5  g01331(n12044, n11478, new_n1708);
and_5  g01332(n7294, n5198, new_n1709);
xnor_4 g01333(new_n1709, new_n1708, new_n1710);
xor_4  g01334(new_n1710, new_n1707, new_n1711);
and_5  g01335(new_n1613, new_n1612, new_n1712);
nor_5  g01336(new_n1613, new_n1612, new_n1713);
nor_5  g01337(new_n1713, new_n1611, new_n1714);
nor_5  g01338(new_n1714, new_n1712, new_n1715);
xnor_4 g01339(new_n1715, new_n1711, new_n1716);
and_5  g01340(n10174, n7354, new_n1717);
and_5  g01341(n4928, n2464, new_n1718);
and_5  g01342(n11311, n4141, new_n1719);
xnor_4 g01343(new_n1719, new_n1718, new_n1720);
and_5  g01344(n4005, n3172, new_n1721);
and_5  g01345(n7236, n1906, new_n1722);
xnor_4 g01346(new_n1722, new_n1721, new_n1723);
xnor_4 g01347(new_n1723, new_n1720, new_n1724);
xnor_4 g01348(new_n1724, new_n1717, new_n1725);
xnor_4 g01349(new_n1725, new_n1716, new_n1726);
xnor_4 g01350(new_n1726, new_n1704, new_n1727);
xnor_4 g01351(new_n1727, new_n1695, new_n1728);
nor_5  g01352(new_n1581, new_n1576_1, new_n1729);
nor_5  g01353(new_n1591, new_n1582, new_n1730);
nor_5  g01354(new_n1730, new_n1729, new_n1731);
nand_5 g01355(n9080, n2509, new_n1732);
nor_5  g01356(new_n1253, new_n1252, new_n1733);
nor_5  g01357(new_n1254, new_n1251, new_n1734);
nor_5  g01358(new_n1734, new_n1733, new_n1735);
nand_5 g01359(n5240, n2508, new_n1736);
and_5  g01360(n11757, n2585, new_n1737);
and_5  g01361(n12706, n1333, new_n1738);
xnor_4 g01362(new_n1738, new_n1737, new_n1739);
xnor_4 g01363(new_n1739, new_n1736, new_n1740);
xnor_4 g01364(new_n1740, new_n1735, new_n1741);
xnor_4 g01365(new_n1741, new_n1732, new_n1742);
xnor_4 g01366(new_n1742, new_n1731, new_n1743);
xnor_4 g01367(new_n1743, new_n1728, new_n1744);
nor_5  g01368(new_n1564_1, new_n1562, new_n1745);
nor_5  g01369(new_n1566, new_n1560, new_n1746);
nor_5  g01370(new_n1746, new_n1745, new_n1747);
nor_5  g01371(new_n1245, new_n1243, new_n1748);
nor_5  g01372(new_n1266, new_n1247, new_n1749);
nor_5  g01373(new_n1749, new_n1748, new_n1750);
xnor_4 g01374(new_n1750, new_n1747, new_n1751);
nor_5  g01375(new_n1549, new_n1544, new_n1752);
nor_5  g01376(new_n1559, new_n1550, new_n1753);
nor_5  g01377(new_n1753, new_n1752, new_n1754);
and_5  g01378(n12704, n6358, new_n1755);
and_5  g01379(n3146, n1512, new_n1756);
xor_4  g01380(new_n1756, new_n1755, new_n1757);
and_5  g01381(n5105, n4187, new_n1758);
and_5  g01382(n6294, n2802, new_n1759);
xnor_4 g01383(new_n1759, new_n1758, new_n1760);
and_5  g01384(n9400, n8236, new_n1761);
and_5  g01385(n1980, n1471, new_n1762);
xnor_4 g01386(new_n1762, new_n1761, new_n1763);
xnor_4 g01387(new_n1763, new_n1760, new_n1764);
xnor_4 g01388(new_n1764, new_n1757, new_n1765);
nand_5 g01389(n12720, n11821, new_n1766);
and_5  g01390(n4938, n1564, new_n1767);
and_5  g01391(n5694, n4805, new_n1768);
xnor_4 g01392(new_n1768, new_n1767, new_n1769);
xnor_4 g01393(new_n1769, new_n1766, new_n1770);
xnor_4 g01394(new_n1770, new_n1765, new_n1771);
nor_5  g01395(new_n1579, new_n1578, new_n1772);
nor_5  g01396(new_n1580, new_n1577, new_n1773);
or_5   g01397(new_n1773, new_n1772, new_n1774);
and_5  g01398(new_n1249, new_n1248, new_n1775);
nor_5  g01399(new_n1255, new_n1250, new_n1776);
nor_5  g01400(new_n1776, new_n1775, new_n1777);
xnor_4 g01401(new_n1777, new_n1774, new_n1778);
xnor_4 g01402(new_n1778, new_n1771, new_n1779);
xnor_4 g01403(new_n1779, new_n1754, new_n1780);
nor_5  g01404(new_n1629, new_n1628, new_n1781);
nor_5  g01405(new_n1631, new_n1626, new_n1782);
nor_5  g01406(new_n1782, new_n1781, new_n1783);
nor_5  g01407(new_n1615, new_n1610, new_n1784);
nor_5  g01408(new_n1625, new_n1616, new_n1785);
nor_5  g01409(new_n1785, new_n1784, new_n1786);
and_5  g01410(new_n1584, new_n1583, new_n1787);
nor_5  g01411(new_n1590, new_n1585, new_n1788);
nor_5  g01412(new_n1788, new_n1787, new_n1789);
nand_5 g01413(n4203, n1209, new_n1790);
and_5  g01414(n6826, n6038, new_n1791);
and_5  g01415(n5283, n5069, new_n1792);
xnor_4 g01416(new_n1792, new_n1791, new_n1793);
xnor_4 g01417(new_n1793, new_n1790, new_n1794);
xnor_4 g01418(new_n1794, new_n1789, new_n1795);
nor_5  g01419(new_n1622, new_n1621, new_n1796);
nor_5  g01420(new_n1623, new_n1620, new_n1797);
nor_5  g01421(new_n1797, new_n1796, new_n1798_1);
nor_5  g01422(new_n1588, new_n1587, new_n1799);
nor_5  g01423(new_n1589, new_n1586, new_n1800);
nor_5  g01424(new_n1800, new_n1799, new_n1801);
and_5  g01425(new_n1547, new_n1546, new_n1802);
nor_5  g01426(new_n1547, new_n1546, new_n1803);
nor_5  g01427(new_n1803, new_n1545, new_n1804);
nor_5  g01428(new_n1804, new_n1802, new_n1805);
xnor_4 g01429(new_n1805, new_n1801, new_n1806);
xnor_4 g01430(new_n1806, new_n1798_1, new_n1807);
xnor_4 g01431(new_n1807, new_n1795, new_n1808);
xnor_4 g01432(new_n1808, new_n1786, new_n1809);
xnor_4 g01433(new_n1809, new_n1783, new_n1810);
xnor_4 g01434(new_n1810, new_n1780, new_n1811);
xnor_4 g01435(new_n1811, new_n1751, new_n1812);
xnor_4 g01436(new_n1812, new_n1744, new_n1813);
xnor_4 g01437(new_n1813, new_n1692, new_n1814);
xnor_4 g01438(new_n1814, new_n1685, new_n1815);
and_5  g01439(new_n1552, new_n1551, new_n1816);
nor_5  g01440(new_n1558, new_n1553, new_n1817);
nor_5  g01441(new_n1817, new_n1816, new_n1818);
and_5  g01442(n6877, n783, new_n1819);
and_5  g01443(n8028, n4722, new_n1820);
xor_4  g01444(new_n1820, new_n1819, new_n1821);
xnor_4 g01445(new_n1821, new_n1818, new_n1822);
nor_5  g01446(new_n1567, new_n1541, new_n1823);
nor_5  g01447(new_n1571, new_n1568, new_n1824);
nor_5  g01448(new_n1824, new_n1823, new_n1825);
and_5  g01449(n10848, n7646, new_n1826);
xnor_4 g01450(new_n1826, new_n1825, new_n1827);
xnor_4 g01451(new_n1827, new_n1822, new_n1828);
nor_5  g01452(new_n1632, new_n1607, new_n1829);
nor_5  g01453(new_n1633, new_n1606, new_n1830);
nor_5  g01454(new_n1830, new_n1829, new_n1831);
nor_5  g01455(new_n1264, new_n1259, new_n1832);
nor_5  g01456(new_n1265, new_n1256, new_n1833);
nor_5  g01457(new_n1833, new_n1832, new_n1834);
nor_5  g01458(new_n1556, new_n1555, new_n1835_1);
nor_5  g01459(new_n1557, new_n1554, new_n1836);
or_5   g01460(new_n1836, new_n1835_1, new_n1837);
and_5  g01461(n12753, n7500, new_n1838);
and_5  g01462(new_n1262, new_n1261, new_n1839);
nor_5  g01463(new_n1262, new_n1261, new_n1840);
nor_5  g01464(new_n1840, new_n1260, new_n1841);
nor_5  g01465(new_n1841, new_n1839, new_n1842);
xnor_4 g01466(new_n1842, new_n1838, new_n1843);
xnor_4 g01467(new_n1843, new_n1837, new_n1844);
xnor_4 g01468(new_n1844, new_n1834, new_n1845);
xnor_4 g01469(new_n1845, new_n1831, new_n1846);
xnor_4 g01470(new_n1846, new_n1828, new_n1847_1);
xnor_4 g01471(new_n1847_1, new_n1815, new_n1848);
xnor_4 g01472(new_n1848, new_n1682, new_n1849);
xnor_4 g01473(new_n1849, new_n1679, n671);
and_5  g01474(n11917, n4312, new_n1851);
and_5  g01475(n12705, n4921, new_n1852);
and_5  g01476(n12025, n9956, new_n1853);
xor_4  g01477(new_n1853, new_n1852, new_n1854);
xnor_4 g01478(new_n1854, new_n1851, new_n1855);
and_5  g01479(n12705, n9956, new_n1856);
and_5  g01480(n11917, n1097, new_n1857);
nor_5  g01481(new_n1857, new_n1856, new_n1858);
nand_5 g01482(new_n1857, new_n1856, new_n1859);
nand_5 g01483(n4921, n4312, new_n1860);
and_5  g01484(new_n1860, new_n1859, new_n1861);
nor_5  g01485(new_n1861, new_n1858, new_n1862);
xor_4  g01486(new_n1862, new_n1855, new_n1863);
and_5  g01487(n5964, n2577, new_n1864);
and_5  g01488(n3842, n1097, new_n1865);
xnor_4 g01489(new_n1865, new_n1864, new_n1866);
xnor_4 g01490(new_n1866, new_n1863, new_n1867);
nand_5 g01491(n5964, n3842, new_n1868);
and_5  g01492(n9956, n4312, new_n1869);
and_5  g01493(n11917, n5964, new_n1870);
nor_5  g01494(new_n1870, new_n1869, new_n1871);
nand_5 g01495(new_n1870, new_n1869, new_n1872);
nand_5 g01496(n4921, n1097, new_n1873);
and_5  g01497(new_n1873, new_n1872, new_n1874);
or_5   g01498(new_n1874, new_n1871, new_n1875);
nor_5  g01499(new_n1875, new_n1868, new_n1876);
xnor_4 g01500(new_n1875, new_n1868, new_n1877);
xnor_4 g01501(new_n1857, new_n1856, new_n1878);
xnor_4 g01502(new_n1878, new_n1860, new_n1879);
nor_5  g01503(new_n1879, new_n1877, new_n1880);
nor_5  g01504(new_n1880, new_n1876, new_n1881);
xnor_4 g01505(new_n1881, new_n1867, new_n1882);
and_5  g01506(n5305, n2577, new_n1883);
xor_4  g01507(new_n1879, new_n1877, new_n1884);
nor_5  g01508(new_n1884, new_n1883, new_n1885);
xnor_4 g01509(new_n1884, new_n1883, new_n1886);
nand_5 g01510(n5305, n3842, new_n1887);
and_5  g01511(n9956, n1097, new_n1888);
and_5  g01512(n11917, n5305, new_n1889);
and_5  g01513(new_n1889, new_n1888, new_n1890);
nor_5  g01514(new_n1889, new_n1888, new_n1891);
nand_5 g01515(n5964, n4921, new_n1892);
nor_5  g01516(new_n1892, new_n1891, new_n1893);
nor_5  g01517(new_n1893, new_n1890, new_n1894);
nor_5  g01518(new_n1894, new_n1887, new_n1895);
xnor_4 g01519(new_n1894, new_n1887, new_n1896);
xnor_4 g01520(new_n1870, new_n1869, new_n1897);
xnor_4 g01521(new_n1897, new_n1873, new_n1898);
nor_5  g01522(new_n1898, new_n1896, new_n1899);
or_5   g01523(new_n1899, new_n1895, new_n1900);
nor_5  g01524(new_n1900, new_n1886, new_n1901);
or_5   g01525(new_n1901, new_n1885, new_n1902);
or_5   g01526(new_n1902, new_n1882, new_n1903);
nor_5  g01527(new_n1854, new_n1851, new_n1904);
nor_5  g01528(new_n1862, new_n1855, new_n1905);
nor_5  g01529(new_n1905, new_n1904, new_n1906_1);
and_5  g01530(n9637, n5964, new_n1907);
and_5  g01531(n2577, n1097, new_n1908);
and_5  g01532(n5305, n1835, new_n1909);
xnor_4 g01533(new_n1909, new_n1908, new_n1910);
xnor_4 g01534(new_n1910, new_n1907, new_n1911);
xnor_4 g01535(new_n1911, new_n1906_1, new_n1912);
and_5  g01536(new_n1853, new_n1852, new_n1913);
and_5  g01537(n4312, n3842, new_n1914);
xnor_4 g01538(new_n1914, new_n1913, new_n1915);
and_5  g01539(n12025, n4921, new_n1916);
and_5  g01540(n12705, n11917, new_n1917);
and_5  g01541(n11257, n9956, new_n1918);
xnor_4 g01542(new_n1918, new_n1917, new_n1919);
xnor_4 g01543(new_n1919, new_n1916, new_n1920);
xnor_4 g01544(new_n1920, new_n1915, new_n1921);
xor_4  g01545(new_n1921, new_n1912, new_n1922);
nor_5  g01546(new_n1866, new_n1863, new_n1923);
nand_5 g01547(new_n1865, new_n1864, new_n1924);
or_5   g01548(new_n1881, new_n1867, new_n1925);
xor_4  g01549(new_n1925, new_n1924, new_n1926);
nor_5  g01550(new_n1926, new_n1923, new_n1927);
xnor_4 g01551(new_n1927, new_n1922, new_n1928);
xnor_4 g01552(new_n1928, new_n1903, new_n1929);
and_5  g01553(n9637, n5305, new_n1930);
xor_4  g01554(new_n1902, new_n1882, new_n1931);
and_5  g01555(new_n1931, new_n1930, new_n1932);
xnor_4 g01556(new_n1898, new_n1896, new_n1933);
xor_4  g01557(new_n1889, new_n1888, new_n1934);
and_5  g01558(n9956, n5964, new_n1935);
and_5  g01559(n5305, n4921, new_n1936);
nand_5 g01560(new_n1936, new_n1935, new_n1937);
or_5   g01561(new_n1937, new_n1934, new_n1938);
or_5   g01562(new_n1938, new_n1933, new_n1939);
xor_4  g01563(new_n1900, new_n1886, new_n1940);
nor_5  g01564(new_n1940, new_n1939, new_n1941);
xor_4  g01565(new_n1931, new_n1930, new_n1942);
and_5  g01566(new_n1942, new_n1941, new_n1943);
nor_5  g01567(new_n1943, new_n1932, new_n1944);
xnor_4 g01568(new_n1944, new_n1929, new_n1945);
and_5  g01569(n8759, n8065, new_n1946);
nand_5 g01570(n7436, n6126, new_n1947);
and_5  g01571(n9241, n3719, new_n1948);
and_5  g01572(n8276, n3602, new_n1949);
xnor_4 g01573(new_n1949, new_n1948, new_n1950);
xnor_4 g01574(new_n1950, new_n1947, new_n1951);
and_5  g01575(n8276, n3719, new_n1952);
and_5  g01576(n12299, n6126, new_n1953);
nor_5  g01577(new_n1953, new_n1952, new_n1954);
nand_5 g01578(new_n1953, new_n1952, new_n1955);
nand_5 g01579(n7436, n3602, new_n1956);
and_5  g01580(new_n1956, new_n1955, new_n1957);
or_5   g01581(new_n1957, new_n1954, new_n1958);
xnor_4 g01582(new_n1958, new_n1951, new_n1959);
and_5  g01583(n10439, n6776, new_n1960);
and_5  g01584(n12299, n8595, new_n1961);
xnor_4 g01585(new_n1961, new_n1960, new_n1962);
xnor_4 g01586(new_n1962, new_n1959, new_n1963);
nand_5 g01587(n8595, n6776, new_n1964);
and_5  g01588(n7436, n3719, new_n1965);
and_5  g01589(n6776, n6126, new_n1966);
nor_5  g01590(new_n1966, new_n1965, new_n1967);
nand_5 g01591(new_n1966, new_n1965, new_n1968);
nand_5 g01592(n12299, n3602, new_n1969);
and_5  g01593(new_n1969, new_n1968, new_n1970);
or_5   g01594(new_n1970, new_n1967, new_n1971);
nor_5  g01595(new_n1971, new_n1964, new_n1972);
xnor_4 g01596(new_n1971, new_n1964, new_n1973);
xnor_4 g01597(new_n1953, new_n1952, new_n1974);
xnor_4 g01598(new_n1974, new_n1956, new_n1975);
nor_5  g01599(new_n1975, new_n1973, new_n1976);
nor_5  g01600(new_n1976, new_n1972, new_n1977);
xnor_4 g01601(new_n1977, new_n1963, new_n1978);
and_5  g01602(n10439, n8759, new_n1979);
xor_4  g01603(new_n1975, new_n1973, new_n1980_1);
nor_5  g01604(new_n1980_1, new_n1979, new_n1981);
xnor_4 g01605(new_n1980_1, new_n1979, new_n1982);
nand_5 g01606(n8759, n8595, new_n1983);
and_5  g01607(n12299, n3719, new_n1984);
and_5  g01608(n8759, n6126, new_n1985);
and_5  g01609(new_n1985, new_n1984, new_n1986);
nor_5  g01610(new_n1985, new_n1984, new_n1987);
nand_5 g01611(n6776, n3602, new_n1988);
nor_5  g01612(new_n1988, new_n1987, new_n1989);
nor_5  g01613(new_n1989, new_n1986, new_n1990);
nor_5  g01614(new_n1990, new_n1983, new_n1991);
xnor_4 g01615(new_n1990, new_n1983, new_n1992);
xnor_4 g01616(new_n1966, new_n1965, new_n1993);
xnor_4 g01617(new_n1993, new_n1969, new_n1994);
nor_5  g01618(new_n1994, new_n1992, new_n1995);
or_5   g01619(new_n1995, new_n1991, new_n1996);
nor_5  g01620(new_n1996, new_n1982, new_n1997);
or_5   g01621(new_n1997, new_n1981, new_n1998);
xor_4  g01622(new_n1998, new_n1978, new_n1999);
and_5  g01623(new_n1999, new_n1946, new_n2000);
xnor_4 g01624(new_n1994, new_n1992, new_n2001);
xor_4  g01625(new_n1985, new_n1984, new_n2002);
and_5  g01626(n6776, n3719, new_n2003);
and_5  g01627(n8759, n3602, new_n2004);
nand_5 g01628(new_n2004, new_n2003, new_n2005);
or_5   g01629(new_n2005, new_n2002, new_n2006);
or_5   g01630(new_n2006, new_n2001, new_n2007);
xor_4  g01631(new_n1996, new_n1982, new_n2008);
or_5   g01632(new_n2008, new_n2007, new_n2009);
xnor_4 g01633(new_n1999, new_n1946, new_n2010);
nor_5  g01634(new_n2010, new_n2009, new_n2011);
nor_5  g01635(new_n2011, new_n2000, new_n2012);
or_5   g01636(new_n1998, new_n1978, new_n2013);
nor_5  g01637(new_n1950, new_n1947, new_n2014);
nor_5  g01638(new_n1958, new_n1951, new_n2015);
or_5   g01639(new_n2015, new_n2014, new_n2016);
and_5  g01640(n8065, n6776, new_n2017);
and_5  g01641(n12299, n10439, new_n2018);
and_5  g01642(n10391, n8759, new_n2019);
xnor_4 g01643(new_n2019, new_n2018, new_n2020);
xnor_4 g01644(new_n2020, new_n2017, new_n2021);
xnor_4 g01645(new_n2021, new_n2016, new_n2022);
and_5  g01646(new_n1949, new_n1948, new_n2023);
and_5  g01647(n8595, n7436, new_n2024_1);
xnor_4 g01648(new_n2024_1, new_n2023, new_n2025);
nand_5 g01649(n9241, n3602, new_n2026);
and_5  g01650(n8276, n6126, new_n2027);
and_5  g01651(n10510, n3719, new_n2028);
xnor_4 g01652(new_n2028, new_n2027, new_n2029);
xnor_4 g01653(new_n2029, new_n2026, new_n2030);
xor_4  g01654(new_n2030, new_n2025, new_n2031);
xor_4  g01655(new_n2031, new_n2022, new_n2032);
nor_5  g01656(new_n1962, new_n1959, new_n2033);
nand_5 g01657(new_n1961, new_n1960, new_n2034);
or_5   g01658(new_n1977, new_n1963, new_n2035);
xor_4  g01659(new_n2035, new_n2034, new_n2036);
nor_5  g01660(new_n2036, new_n2033, new_n2037);
xnor_4 g01661(new_n2037, new_n2032, new_n2038);
xnor_4 g01662(new_n2038, new_n2013, new_n2039);
xnor_4 g01663(new_n2039, new_n2012, new_n2040);
nand_5 g01664(n12648, n4826, new_n2041);
and_5  g01665(n10545, n7733, new_n2042);
and_5  g01666(n12925, n7690, new_n2043);
xnor_4 g01667(new_n2043, new_n2042, new_n2044);
xnor_4 g01668(new_n2044, new_n2041, new_n2045);
and_5  g01669(n12925, n10545, new_n2046);
and_5  g01670(n4826, n2530, new_n2047);
nor_5  g01671(new_n2047, new_n2046, new_n2048);
and_5  g01672(n12648, n7733, new_n2049);
xnor_4 g01673(new_n2047, new_n2046, new_n2050);
nor_5  g01674(new_n2050, new_n2049, new_n2051);
or_5   g01675(new_n2051, new_n2048, new_n2052);
xnor_4 g01676(new_n2052, new_n2045, new_n2053);
and_5  g01677(n8476, n4970, new_n2054);
and_5  g01678(n7610, n2530, new_n2055);
xnor_4 g01679(new_n2055, new_n2054, new_n2056);
xnor_4 g01680(new_n2056, new_n2053, new_n2057);
and_5  g01681(n8476, n7610, new_n2058);
and_5  g01682(n12925, n12648, new_n2059);
and_5  g01683(n8476, n4826, new_n2060);
nor_5  g01684(new_n2060, new_n2059, new_n2061);
and_5  g01685(n7733, n2530, new_n2062);
xnor_4 g01686(new_n2060, new_n2059, new_n2063);
nor_5  g01687(new_n2063, new_n2062, new_n2064);
nor_5  g01688(new_n2064, new_n2061, new_n2065);
and_5  g01689(new_n2065, new_n2058, new_n2066);
xnor_4 g01690(new_n2065, new_n2058, new_n2067);
xor_4  g01691(new_n2050, new_n2049, new_n2068);
nor_5  g01692(new_n2068, new_n2067, new_n2069);
nor_5  g01693(new_n2069, new_n2066, new_n2070);
xnor_4 g01694(new_n2070, new_n2057, new_n2071);
and_5  g01695(n5331, n4970, new_n2072);
nand_5 g01696(n7610, n5331, new_n2073);
and_5  g01697(n12925, n2530, new_n2074);
and_5  g01698(n5331, n4826, new_n2075);
nor_5  g01699(new_n2075, new_n2074, new_n2076);
and_5  g01700(new_n2075, new_n2074, new_n2077);
and_5  g01701(n8476, n7733, new_n2078);
nor_5  g01702(new_n2078, new_n2077, new_n2079);
or_5   g01703(new_n2079, new_n2076, new_n2080);
nor_5  g01704(new_n2080, new_n2073, new_n2081);
xnor_4 g01705(new_n2080, new_n2073, new_n2082);
xor_4  g01706(new_n2063, new_n2062, new_n2083);
nor_5  g01707(new_n2083, new_n2082, new_n2084);
or_5   g01708(new_n2084, new_n2081, new_n2085);
nor_5  g01709(new_n2085, new_n2072, new_n2086);
xor_4  g01710(new_n2068, new_n2067, new_n2087_1);
xnor_4 g01711(new_n2085, new_n2072, new_n2088);
nor_5  g01712(new_n2088, new_n2087_1, new_n2089);
or_5   g01713(new_n2089, new_n2086, new_n2090);
or_5   g01714(new_n2090, new_n2071, new_n2091);
nor_5  g01715(new_n2056, new_n2053, new_n2092);
nand_5 g01716(new_n2055, new_n2054, new_n2093);
or_5   g01717(new_n2070, new_n2057, new_n2094);
xor_4  g01718(new_n2094, new_n2093, new_n2095);
nor_5  g01719(new_n2095, new_n2092, new_n2096_1);
and_5  g01720(new_n2043, new_n2042, new_n2097);
and_5  g01721(n12648, n7610, new_n2098);
xnor_4 g01722(new_n2098, new_n2097, new_n2099);
and_5  g01723(n7733, n7690, new_n2100);
and_5  g01724(n10545, n4826, new_n2101);
and_5  g01725(n12925, n3616, new_n2102);
xnor_4 g01726(new_n2102, new_n2101, new_n2103);
xor_4  g01727(new_n2103, new_n2100, new_n2104);
xnor_4 g01728(new_n2104, new_n2099, new_n2105);
nor_5  g01729(new_n2044, new_n2041, new_n2106);
nor_5  g01730(new_n2052, new_n2045, new_n2107);
nor_5  g01731(new_n2107, new_n2106, new_n2108);
and_5  g01732(n8476, n503, new_n2109);
and_5  g01733(n4970, n2530, new_n2110);
and_5  g01734(n10965, n5331, new_n2111);
xnor_4 g01735(new_n2111, new_n2110, new_n2112);
xor_4  g01736(new_n2112, new_n2109, new_n2113);
xnor_4 g01737(new_n2113, new_n2108, new_n2114);
xnor_4 g01738(new_n2114, new_n2105, new_n2115);
xnor_4 g01739(new_n2115, new_n2096_1, new_n2116);
xnor_4 g01740(new_n2116, new_n2091, new_n2117);
and_5  g01741(n5331, n503, new_n2118);
xor_4  g01742(new_n2090, new_n2071, new_n2119);
and_5  g01743(new_n2119, new_n2118, new_n2120);
xnor_4 g01744(new_n2083, new_n2082, new_n2121);
nand_5 g01745(n8476, n7733, new_n2122);
and_5  g01746(n12925, n5331, new_n2123);
or_5   g01747(new_n2123, new_n2122, new_n2124);
and_5  g01748(new_n2124, new_n2076, new_n2125);
nor_5  g01749(new_n2125, new_n2077, new_n2126);
or_5   g01750(new_n2126, new_n2122, new_n2127);
or_5   g01751(new_n2127, new_n2121, new_n2128);
xor_4  g01752(new_n2088, new_n2087_1, new_n2129);
or_5   g01753(new_n2129, new_n2128, new_n2130);
xnor_4 g01754(new_n2119, new_n2118, new_n2131_1);
nor_5  g01755(new_n2131_1, new_n2130, new_n2132);
nor_5  g01756(new_n2132, new_n2120, new_n2133);
xor_4  g01757(new_n2133, new_n2117, new_n2134);
nand_5 g01758(n4086, n2393, new_n2135);
and_5  g01759(n5860, n405, new_n2136);
and_5  g01760(n8433, n3986, new_n2137);
xnor_4 g01761(new_n2137, new_n2136, new_n2138);
xnor_4 g01762(new_n2138, new_n2135, new_n2139);
and_5  g01763(n8433, n5860, new_n2140);
and_5  g01764(n11892, n4086, new_n2141);
nor_5  g01765(new_n2141, new_n2140, new_n2142);
and_5  g01766(n2393, n405, new_n2143);
xnor_4 g01767(new_n2141, new_n2140, new_n2144);
nor_5  g01768(new_n2144, new_n2143, new_n2145);
or_5   g01769(new_n2145, new_n2142, new_n2146);
xnor_4 g01770(new_n2146, new_n2139, new_n2147);
and_5  g01771(n7388, n6611, new_n2148);
and_5  g01772(n11892, n217, new_n2149);
xnor_4 g01773(new_n2149, new_n2148, new_n2150);
xnor_4 g01774(new_n2150, new_n2147, new_n2151);
and_5  g01775(n7388, n217, new_n2152);
and_5  g01776(n8433, n2393, new_n2153);
and_5  g01777(n7388, n4086, new_n2154);
nor_5  g01778(new_n2154, new_n2153, new_n2155);
and_5  g01779(n11892, n405, new_n2156);
xnor_4 g01780(new_n2154, new_n2153, new_n2157);
nor_5  g01781(new_n2157, new_n2156, new_n2158);
nor_5  g01782(new_n2158, new_n2155, new_n2159);
and_5  g01783(new_n2159, new_n2152, new_n2160);
xnor_4 g01784(new_n2159, new_n2152, new_n2161);
xor_4  g01785(new_n2144, new_n2143, new_n2162);
nor_5  g01786(new_n2162, new_n2161, new_n2163);
nor_5  g01787(new_n2163, new_n2160, new_n2164);
xnor_4 g01788(new_n2164, new_n2151, new_n2165);
nand_5 g01789(n7965, n6611, new_n2166);
xnor_4 g01790(new_n2162, new_n2161, new_n2167);
nor_5  g01791(new_n2167, new_n2166, new_n2168);
xnor_4 g01792(new_n2167, new_n2166, new_n2169);
nand_5 g01793(n7965, n217, new_n2170);
and_5  g01794(n11892, n8433, new_n2171);
and_5  g01795(n7965, n4086, new_n2172);
and_5  g01796(new_n2172, new_n2171, new_n2173);
nor_5  g01797(new_n2172, new_n2171, new_n2174);
nand_5 g01798(n7388, n405, new_n2175);
nor_5  g01799(new_n2175, new_n2174, new_n2176);
nor_5  g01800(new_n2176, new_n2173, new_n2177);
nor_5  g01801(new_n2177, new_n2170, new_n2178);
xnor_4 g01802(new_n2177, new_n2170, new_n2179);
xor_4  g01803(new_n2157, new_n2156, new_n2180);
nor_5  g01804(new_n2180, new_n2179, new_n2181);
nor_5  g01805(new_n2181, new_n2178, new_n2182);
nor_5  g01806(new_n2182, new_n2169, new_n2183);
nor_5  g01807(new_n2183, new_n2168, new_n2184);
or_5   g01808(new_n2184, new_n2165, new_n2185);
nor_5  g01809(new_n2150, new_n2147, new_n2186);
nand_5 g01810(new_n2149, new_n2148, new_n2187);
or_5   g01811(new_n2164, new_n2151, new_n2188);
xor_4  g01812(new_n2188, new_n2187, new_n2189);
nor_5  g01813(new_n2189, new_n2186, new_n2190);
and_5  g01814(new_n2137, new_n2136, new_n2191);
and_5  g01815(n2393, n217, new_n2192);
xnor_4 g01816(new_n2192, new_n2191, new_n2193);
and_5  g01817(n3986, n405, new_n2194);
and_5  g01818(n5860, n4086, new_n2195);
and_5  g01819(n8433, n5857, new_n2196);
xnor_4 g01820(new_n2196, new_n2195, new_n2197);
xor_4  g01821(new_n2197, new_n2194, new_n2198);
xor_4  g01822(new_n2198, new_n2193, new_n2199);
nor_5  g01823(new_n2138, new_n2135, new_n2200);
nor_5  g01824(new_n2146, new_n2139, new_n2201);
or_5   g01825(new_n2201, new_n2200, new_n2202);
and_5  g01826(n11296, n7965, new_n2203);
and_5  g01827(n11892, n6611, new_n2204);
and_5  g01828(n7388, n6359, new_n2205);
xnor_4 g01829(new_n2205, new_n2204, new_n2206);
xnor_4 g01830(new_n2206, new_n2203, new_n2207);
xnor_4 g01831(new_n2207, new_n2202, new_n2208);
xor_4  g01832(new_n2208, new_n2199, new_n2209);
xnor_4 g01833(new_n2209, new_n2190, new_n2210);
xnor_4 g01834(new_n2210, new_n2185, new_n2211);
nand_5 g01835(n7965, n6359, new_n2212);
xnor_4 g01836(new_n2184, new_n2165, new_n2213);
nor_5  g01837(new_n2213, new_n2212, new_n2214);
xnor_4 g01838(new_n2180, new_n2179, new_n2215);
xor_4  g01839(new_n2172, new_n2171, new_n2216);
and_5  g01840(n8433, n7388, new_n2217);
and_5  g01841(n7965, n405, new_n2218);
nand_5 g01842(new_n2218, new_n2217, new_n2219);
or_5   g01843(new_n2219, new_n2216, new_n2220);
or_5   g01844(new_n2220, new_n2215, new_n2221);
xnor_4 g01845(new_n2182, new_n2169, new_n2222);
or_5   g01846(new_n2222, new_n2221, new_n2223);
xnor_4 g01847(new_n2213, new_n2212, new_n2224);
nor_5  g01848(new_n2224, new_n2223, new_n2225);
nor_5  g01849(new_n2225, new_n2214, new_n2226_1);
xor_4  g01850(new_n2226_1, new_n2211, new_n2227);
xnor_4 g01851(new_n2227, new_n2134, new_n2228);
xor_4  g01852(new_n2131_1, new_n2130, new_n2229);
xor_4  g01853(new_n2224, new_n2223, new_n2230);
nor_5  g01854(new_n2230, new_n2229, new_n2231);
xor_4  g01855(new_n2222, new_n2221, new_n2232);
xor_4  g01856(new_n2127, new_n2121, new_n2233);
xor_4  g01857(new_n2220, new_n2215, new_n2234);
nor_5  g01858(new_n2234, new_n2233, new_n2235);
and_5  g01859(n8433, n7965, new_n2236);
and_5  g01860(new_n2236, new_n2123, new_n2237);
xor_4  g01861(new_n2218, new_n2217, new_n2238);
nor_5  g01862(new_n2238, new_n2237, new_n2239);
xnor_4 g01863(new_n2238, new_n2237, new_n2240);
and_5  g01864(n12925, n8476, new_n2241);
and_5  g01865(n7733, n5331, new_n2242);
xor_4  g01866(new_n2242, new_n2241, new_n2243);
nor_5  g01867(new_n2243, new_n2240, new_n2244);
nor_5  g01868(new_n2244, new_n2239, new_n2245);
or_5   g01869(new_n2124, new_n2076, new_n2246);
and_5  g01870(new_n2246, new_n2126, new_n2247);
nor_5  g01871(new_n2247, new_n2245, new_n2248);
xnor_4 g01872(new_n2247, new_n2245, new_n2249);
nor_5  g01873(new_n2236, new_n2175, new_n2250);
nor_5  g01874(new_n2250, new_n2216, new_n2251);
or_5   g01875(new_n2236, new_n2175, new_n2252);
nor_5  g01876(new_n2252, new_n2174, new_n2253_1);
nor_5  g01877(new_n2253_1, new_n2251, new_n2254);
nor_5  g01878(new_n2254, new_n2249, new_n2255);
nor_5  g01879(new_n2255, new_n2248, new_n2256);
xnor_4 g01880(new_n2234, new_n2233, new_n2257);
nor_5  g01881(new_n2257, new_n2256, new_n2258);
nor_5  g01882(new_n2258, new_n2235, new_n2259);
nor_5  g01883(new_n2259, new_n2232, new_n2260);
xor_4  g01884(new_n2129, new_n2128, new_n2261);
xnor_4 g01885(new_n2259, new_n2232, new_n2262);
nor_5  g01886(new_n2262, new_n2261, new_n2263);
nor_5  g01887(new_n2263, new_n2260, new_n2264);
xnor_4 g01888(new_n2230, new_n2229, new_n2265);
nor_5  g01889(new_n2265, new_n2264, new_n2266);
nor_5  g01890(new_n2266, new_n2231, new_n2267);
xor_4  g01891(new_n2267, new_n2228, new_n2268);
xnor_4 g01892(new_n2268, new_n2040, new_n2269);
xnor_4 g01893(new_n2010, new_n2009, new_n2270);
xor_4  g01894(new_n2265, new_n2264, new_n2271);
and_5  g01895(new_n2271, new_n2270, new_n2272);
xnor_4 g01896(new_n2271, new_n2270, new_n2273);
xnor_4 g01897(new_n2008, new_n2007, new_n2274);
xor_4  g01898(new_n2262, new_n2261, new_n2275);
nor_5  g01899(new_n2275, new_n2274, new_n2276);
xnor_4 g01900(new_n2275, new_n2274, new_n2277);
xnor_4 g01901(new_n2006, new_n2001, new_n2278_1);
xor_4  g01902(new_n2257, new_n2256, new_n2279);
nor_5  g01903(new_n2279, new_n2278_1, new_n2280);
xnor_4 g01904(new_n2279, new_n2278_1, new_n2281);
xor_4  g01905(new_n2254, new_n2249, new_n2282);
and_5  g01906(n8759, n3719, new_n2283);
nor_5  g01907(new_n2283, new_n1988, new_n2284);
nor_5  g01908(new_n2284, new_n2002, new_n2285);
or_5   g01909(new_n2283, new_n1988, new_n2286);
nor_5  g01910(new_n2286, new_n1987, new_n2287);
or_5   g01911(new_n2287, new_n2285, new_n2288);
nor_5  g01912(new_n2288, new_n2282, new_n2289);
xnor_4 g01913(new_n2288, new_n2282, new_n2290);
xor_4  g01914(new_n2243, new_n2240, new_n2291);
xnor_4 g01915(new_n2004, new_n2003, new_n2292);
nor_5  g01916(new_n2292, new_n2291, new_n2293);
nand_5 g01917(n8759, n3719, new_n2294);
xnor_4 g01918(new_n2236, new_n2123, new_n2295);
or_5   g01919(new_n2295, new_n2294, new_n2296);
xnor_4 g01920(new_n2292, new_n2291, new_n2297);
nor_5  g01921(new_n2297, new_n2296, new_n2298);
nor_5  g01922(new_n2298, new_n2293, new_n2299);
nor_5  g01923(new_n2299, new_n2290, new_n2300);
nor_5  g01924(new_n2300, new_n2289, new_n2301_1);
nor_5  g01925(new_n2301_1, new_n2281, new_n2302);
nor_5  g01926(new_n2302, new_n2280, new_n2303);
nor_5  g01927(new_n2303, new_n2277, new_n2304);
or_5   g01928(new_n2304, new_n2276, new_n2305);
nor_5  g01929(new_n2305, new_n2273, new_n2306);
nor_5  g01930(new_n2306, new_n2272, new_n2307);
xor_4  g01931(new_n2307, new_n2269, new_n2308);
nor_5  g01932(new_n2308, new_n1945, new_n2309);
xnor_4 g01933(new_n2308, new_n1945, new_n2310);
xnor_4 g01934(new_n1942, new_n1941, new_n2311);
xor_4  g01935(new_n2305, new_n2273, new_n2312);
nor_5  g01936(new_n2312, new_n2311, new_n2313);
xor_4  g01937(new_n1940, new_n1939, new_n2314);
xor_4  g01938(new_n2303, new_n2277, new_n2315);
nor_5  g01939(new_n2315, new_n2314, new_n2316_1);
xnor_4 g01940(new_n2315, new_n2314, new_n2317);
xor_4  g01941(new_n1938, new_n1933, new_n2318);
xor_4  g01942(new_n2301_1, new_n2281, new_n2319);
nor_5  g01943(new_n2319, new_n2318, new_n2320);
xor_4  g01944(new_n2299, new_n2290, new_n2321);
and_5  g01945(n9956, n5305, new_n2322);
nor_5  g01946(new_n2322, new_n1892, new_n2323);
nor_5  g01947(new_n2323, new_n1934, new_n2324);
or_5   g01948(new_n2322, new_n1892, new_n2325);
nor_5  g01949(new_n2325, new_n1891, new_n2326);
nor_5  g01950(new_n2326, new_n2324, new_n2327);
nor_5  g01951(new_n2327, new_n2321, new_n2328);
xnor_4 g01952(new_n2327, new_n2321, new_n2329);
xnor_4 g01953(new_n2295, new_n2283, new_n2330);
and_5  g01954(new_n2330, new_n2322, new_n2331);
xor_4  g01955(new_n1936, new_n1935, new_n2332);
nor_5  g01956(new_n2332, new_n2331, new_n2333);
xnor_4 g01957(new_n2297, new_n2296, new_n2334);
xor_4  g01958(new_n2332, new_n2331, new_n2335);
and_5  g01959(new_n2335, new_n2334, new_n2336);
nor_5  g01960(new_n2336, new_n2333, new_n2337);
nor_5  g01961(new_n2337, new_n2329, new_n2338);
nor_5  g01962(new_n2338, new_n2328, new_n2339);
xnor_4 g01963(new_n2319, new_n2318, new_n2340);
nor_5  g01964(new_n2340, new_n2339, new_n2341);
nor_5  g01965(new_n2341, new_n2320, new_n2342);
nor_5  g01966(new_n2342, new_n2317, new_n2343);
or_5   g01967(new_n2343, new_n2316_1, new_n2344);
xnor_4 g01968(new_n2312, new_n2311, new_n2345);
nor_5  g01969(new_n2345, new_n2344, new_n2346);
nor_5  g01970(new_n2346, new_n2313, new_n2347_1);
nor_5  g01971(new_n2347_1, new_n2310, new_n2348);
nor_5  g01972(new_n2348, new_n2309, new_n2349);
nor_5  g01973(new_n2268, new_n2040, new_n2350);
or_5   g01974(new_n2306, new_n2272, new_n2351);
nor_5  g01975(new_n2351, new_n2269, new_n2352);
nor_5  g01976(new_n2352, new_n2350, new_n2353);
and_5  g01977(new_n2098, new_n2097, new_n2354);
nor_5  g01978(new_n2104, new_n2099, new_n2355);
nor_5  g01979(new_n2355, new_n2354, new_n2356);
nor_5  g01980(new_n2102, new_n2101, new_n2357);
nor_5  g01981(new_n2103, new_n2100, new_n2358);
nor_5  g01982(new_n2358, new_n2357, new_n2359);
and_5  g01983(n12648, n4970, new_n2360);
and_5  g01984(n11296, n7388, new_n2361);
and_5  g01985(n9241, n6126, new_n2362);
xnor_4 g01986(new_n2362, new_n2361, new_n2363);
xnor_4 g01987(new_n2363, new_n2360, new_n2364);
xnor_4 g01988(new_n2364, new_n2359, new_n2365);
xnor_4 g01989(new_n2365, new_n2356, new_n2366);
nor_5  g01990(new_n2196, new_n2195, new_n2367);
nor_5  g01991(new_n2197, new_n2194, new_n2368);
nor_5  g01992(new_n2368, new_n2367, new_n2369);
nor_5  g01993(new_n2205, new_n2204, new_n2370);
nor_5  g01994(new_n2206, new_n2203, new_n2371);
nor_5  g01995(new_n2371, new_n2370, new_n2372);
xnor_4 g01996(new_n2372, new_n2369, new_n2373);
and_5  g01997(n11892, n6359, new_n2374);
and_5  g01998(n7546, n5331, new_n2375);
xor_4  g01999(new_n2375, new_n2374, new_n2376);
xnor_4 g02000(new_n2376, new_n2373, new_n2377);
and_5  g02001(new_n2024_1, new_n2023, new_n2378);
nor_5  g02002(new_n2030, new_n2025, new_n2379);
nor_5  g02003(new_n2379, new_n2378, new_n2380);
and_5  g02004(n8595, n8276, new_n2381);
and_5  g02005(n6611, n2393, new_n2382);
xnor_4 g02006(new_n2382, new_n2381, new_n2383_1);
and_5  g02007(n12925, n4499, new_n2384);
and_5  g02008(n11536, n5305, new_n2385);
xnor_4 g02009(new_n2385, new_n2384, new_n2386);
xor_4  g02010(new_n2386, new_n2383_1, new_n2387);
xnor_4 g02011(new_n2387, new_n2380, new_n2388);
xnor_4 g02012(new_n2388, new_n2377, new_n2389);
and_5  g02013(new_n2192, new_n2191, new_n2390);
nor_5  g02014(new_n2198, new_n2193, new_n2391);
nor_5  g02015(new_n2391, new_n2390, new_n2392);
nor_5  g02016(new_n2111, new_n2110, new_n2393_1);
nor_5  g02017(new_n2112, new_n2109, new_n2394);
nor_5  g02018(new_n2394, new_n2393_1, new_n2395);
and_5  g02019(n4086, n3986, new_n2396);
and_5  g02020(n7733, n3616, new_n2397);
xor_4  g02021(new_n2397, new_n2396, new_n2398);
xnor_4 g02022(new_n2398, new_n2395, new_n2399);
xnor_4 g02023(new_n2399, new_n2392, new_n2400);
xnor_4 g02024(new_n2400, new_n2389, new_n2401);
xnor_4 g02025(new_n2401, new_n2366, new_n2402);
nor_5  g02026(new_n2210, new_n2185, new_n2403);
nor_5  g02027(new_n2226_1, new_n2211, new_n2404);
nor_5  g02028(new_n2404, new_n2403, new_n2405);
nand_5 g02029(n5860, n217, new_n2406);
xnor_4 g02030(new_n2406, new_n2405, new_n2407);
nor_5  g02031(new_n2038, new_n2013, new_n2408);
nor_5  g02032(new_n2039, new_n2012, new_n2409);
nor_5  g02033(new_n2409, new_n2408, new_n2410);
nor_5  g02034(new_n2113, new_n2108, new_n2411);
nor_5  g02035(new_n2114, new_n2105, new_n2412);
nor_5  g02036(new_n2412, new_n2411, new_n2413);
and_5  g02037(n12299, n8065, new_n2414);
and_5  g02038(n10510, n3602, new_n2415);
xor_4  g02039(new_n2415, new_n2414, new_n2416);
and_5  g02040(n10644, n3719, new_n2417);
and_5  g02041(n7965, n1357, new_n2418);
xnor_4 g02042(new_n2418, new_n2417, new_n2419);
and_5  g02043(n10439, n7436, new_n2420);
and_5  g02044(n8759, n4190, new_n2421);
xnor_4 g02045(new_n2421, new_n2420, new_n2422);
xnor_4 g02046(new_n2422, new_n2419, new_n2423);
xnor_4 g02047(new_n2423, new_n2416, new_n2424);
nor_5  g02048(new_n1909, new_n1908, new_n2425_1);
nor_5  g02049(new_n1910, new_n1907, new_n2426);
nor_5  g02050(new_n2426, new_n2425_1, new_n2427);
nand_5 g02051(n9637, n1097, new_n2428);
xnor_4 g02052(new_n2428, new_n2427, new_n2429);
xnor_4 g02053(new_n2429, new_n2424, new_n2430);
xnor_4 g02054(new_n2430, new_n2413, new_n2431_1);
nor_5  g02055(new_n2021, new_n2016, new_n2432);
nor_5  g02056(new_n2031, new_n2022, new_n2433_1);
nor_5  g02057(new_n2433_1, new_n2432, new_n2434_1);
nor_5  g02058(new_n1911, new_n1906_1, new_n2435);
nor_5  g02059(new_n1921, new_n1912, new_n2436);
nor_5  g02060(new_n2436, new_n2435, new_n2437);
xnor_4 g02061(new_n2437, new_n2434_1, new_n2438);
xnor_4 g02062(new_n2438, new_n2431_1, new_n2439);
nor_5  g02063(new_n2035, new_n2034, new_n2440);
nor_5  g02064(new_n2037, new_n2032, new_n2441);
nor_5  g02065(new_n2441, new_n2440, new_n2442);
nor_5  g02066(new_n2019, new_n2018, new_n2443);
nor_5  g02067(new_n2020, new_n2017, new_n2444);
nor_5  g02068(new_n2444, new_n2443, new_n2445);
and_5  g02069(n4312, n2577, new_n2446);
xnor_4 g02070(new_n2446, new_n2445, new_n2447);
and_5  g02071(new_n2028, new_n2027, new_n2448);
nor_5  g02072(new_n2028, new_n2027, new_n2449);
nor_5  g02073(new_n2449, new_n2026, new_n2450);
nor_5  g02074(new_n2450, new_n2448, new_n2451);
and_5  g02075(n11257, n4921, new_n2452);
and_5  g02076(n12705, n3842, new_n2453);
xor_4  g02077(new_n2453, new_n2452, new_n2454);
xnor_4 g02078(new_n2454, new_n2451, new_n2455);
xnor_4 g02079(new_n2455, new_n2447, new_n2456);
and_5  g02080(n8433, n45, new_n2457);
and_5  g02081(n12025, n11917, new_n2458);
xor_4  g02082(new_n2458, new_n2457, new_n2459);
nor_5  g02083(new_n1918, new_n1917, new_n2460);
nor_5  g02084(new_n1919, new_n1916, new_n2461);
nor_5  g02085(new_n2461, new_n2460, new_n2462);
and_5  g02086(n5964, n1835, new_n2463);
and_5  g02087(n5857, n405, new_n2464_1);
xor_4  g02088(new_n2464_1, new_n2463, new_n2465);
xnor_4 g02089(new_n2465, new_n2462, new_n2466);
xnor_4 g02090(new_n2466, new_n2459, new_n2467);
nor_5  g02091(new_n1914, new_n1913, new_n2468);
nor_5  g02092(new_n1920, new_n1915, new_n2469);
nor_5  g02093(new_n2469, new_n2468, new_n2470);
nand_5 g02094(n10391, n6776, new_n2471);
xnor_4 g02095(new_n2471, new_n2470, new_n2472);
xnor_4 g02096(new_n2472, new_n2467, new_n2473);
xnor_4 g02097(new_n2473, new_n2456, new_n2474);
xnor_4 g02098(new_n2474, new_n2442, new_n2475);
xnor_4 g02099(new_n2475, new_n2439, new_n2476);
xnor_4 g02100(new_n2476, new_n2410, new_n2477);
xnor_4 g02101(new_n2477, new_n2407, new_n2478);
xnor_4 g02102(new_n2478, new_n2402, new_n2479);
nor_5  g02103(new_n2227, new_n2134, new_n2480);
nor_5  g02104(new_n2267, new_n2228, new_n2481);
nor_5  g02105(new_n2481, new_n2480, new_n2482);
nor_5  g02106(new_n2188, new_n2187, new_n2483);
nor_5  g02107(new_n2209, new_n2190, new_n2484);
or_5   g02108(new_n2484, new_n2483, new_n2485);
nor_5  g02109(new_n1925, new_n1924, new_n2486);
nor_5  g02110(new_n1927, new_n1922, new_n2487);
nor_5  g02111(new_n2487, new_n2486, new_n2488);
xnor_4 g02112(new_n2488, new_n2485, new_n2489);
xnor_4 g02113(new_n2489, new_n2482, new_n2490);
xnor_4 g02114(new_n2490, new_n2479, new_n2491);
xnor_4 g02115(new_n2491, new_n2353, new_n2492);
nor_5  g02116(new_n2116, new_n2091, new_n2493);
nor_5  g02117(new_n2133, new_n2117, new_n2494);
nor_5  g02118(new_n2494, new_n2493, new_n2495);
nor_5  g02119(new_n1928, new_n1903, new_n2496);
nor_5  g02120(new_n1944, new_n1929, new_n2497);
nor_5  g02121(new_n2497, new_n2496, new_n2498_1);
xnor_4 g02122(new_n2498_1, new_n2495, new_n2499);
nor_5  g02123(new_n2094, new_n2093, new_n2500);
nor_5  g02124(new_n2115, new_n2096_1, new_n2501);
nor_5  g02125(new_n2501, new_n2500, new_n2502);
nor_5  g02126(new_n2207, new_n2202, new_n2503);
nor_5  g02127(new_n2208, new_n2199, new_n2504);
nor_5  g02128(new_n2504, new_n2503, new_n2505);
nand_5 g02129(n10547, n9956, new_n2506);
and_5  g02130(n10965, n8476, new_n2507_1);
and_5  g02131(n7690, n4826, new_n2508_1);
xnor_4 g02132(new_n2508_1, new_n2507_1, new_n2509_1);
and_5  g02133(n10545, n7610, new_n2510);
and_5  g02134(n2530, n503, new_n2511);
xnor_4 g02135(new_n2511, new_n2510, new_n2512_1);
xnor_4 g02136(new_n2512_1, new_n2509_1, new_n2513);
xnor_4 g02137(new_n2513, new_n2506, new_n2514);
xnor_4 g02138(new_n2514, new_n2505, new_n2515_1);
xor_4  g02139(new_n2515_1, new_n2502, new_n2516);
xnor_4 g02140(new_n2516, new_n2499, new_n2517);
xnor_4 g02141(new_n2517, new_n2492, new_n2518);
xnor_4 g02142(new_n2518, new_n2349, n837);
and_5  g02143(n11917, n11757, new_n2520);
nand_5 g02144(n9956, n5240, new_n2521);
and_5  g02145(n11757, n4921, new_n2522_1);
nand_5 g02146(n11917, n3172, new_n2523);
xnor_4 g02147(new_n2523, new_n2521, new_n2524);
nor_5  g02148(new_n2524, new_n2522_1, new_n2525);
nor_5  g02149(new_n2525, new_n2521, new_n2526);
nor_5  g02150(new_n2526, new_n2520, new_n2527);
and_5  g02151(n4921, n3172, new_n2528);
or_5   g02152(new_n2528, new_n2526, new_n2529);
and_5  g02153(new_n2529, new_n2520, new_n2530_1);
or_5   g02154(new_n2530_1, new_n2527, new_n2531);
and_5  g02155(n5240, n4921, new_n2532);
and_5  g02156(n11821, n9956, new_n2533);
xnor_4 g02157(new_n2533, new_n2532, new_n2534);
xnor_4 g02158(new_n2534, new_n2531, new_n2535);
and_5  g02159(n2577, n1333, new_n2536);
and_5  g02160(n3842, n3172, new_n2537);
xnor_4 g02161(new_n2537, new_n2536, new_n2538);
xnor_4 g02162(new_n2538, new_n2535, new_n2539);
nand_5 g02163(n3842, n1333, new_n2540);
and_5  g02164(n11757, n9956, new_n2541);
and_5  g02165(n11917, n1333, new_n2542);
nor_5  g02166(new_n2542, new_n2541, new_n2543);
and_5  g02167(new_n2542, new_n2541, new_n2544);
nor_5  g02168(new_n2544, new_n2528, new_n2545);
or_5   g02169(new_n2545, new_n2543, new_n2546);
nor_5  g02170(new_n2546, new_n2540, new_n2547);
xnor_4 g02171(new_n2524, new_n2522_1, new_n2548);
xor_4  g02172(new_n2546, new_n2540, new_n2549);
and_5  g02173(new_n2549, new_n2548, new_n2550);
nor_5  g02174(new_n2550, new_n2547, new_n2551_1);
xnor_4 g02175(new_n2551_1, new_n2539, new_n2552);
nand_5 g02176(n7862, n2577, new_n2553);
xnor_4 g02177(new_n2549, new_n2548, new_n2554);
nor_5  g02178(new_n2554, new_n2553, new_n2555);
nand_5 g02179(n7862, n3842, new_n2556);
and_5  g02180(n9956, n3172, new_n2557);
and_5  g02181(n11917, n7862, new_n2558_1);
and_5  g02182(new_n2558_1, new_n2557, new_n2559);
nor_5  g02183(new_n2558_1, new_n2557, new_n2560);
nand_5 g02184(n4921, n1333, new_n2561);
nor_5  g02185(new_n2561, new_n2560, new_n2562);
nor_5  g02186(new_n2562, new_n2559, new_n2563);
nor_5  g02187(new_n2563, new_n2556, new_n2564_1);
xnor_4 g02188(new_n2563, new_n2556, new_n2565);
xnor_4 g02189(new_n2542, new_n2541, new_n2566);
xor_4  g02190(new_n2566, new_n2528, new_n2567);
nor_5  g02191(new_n2567, new_n2565, new_n2568);
nor_5  g02192(new_n2568, new_n2564_1, new_n2569);
xnor_4 g02193(new_n2554, new_n2553, new_n2570);
nor_5  g02194(new_n2570, new_n2569, new_n2571);
nor_5  g02195(new_n2571, new_n2555, new_n2572);
or_5   g02196(new_n2572, new_n2552, new_n2573);
nor_5  g02197(new_n2534, new_n2531, new_n2574);
or_5   g02198(new_n2574, new_n2530_1, new_n2575);
nand_5 g02199(n9637, n1333, new_n2576);
and_5  g02200(n3172, n2577, new_n2577_1);
and_5  g02201(n7862, n1835, new_n2578);
xnor_4 g02202(new_n2578, new_n2577_1, new_n2579);
xor_4  g02203(new_n2579, new_n2576, new_n2580);
xnor_4 g02204(new_n2580, new_n2575, new_n2581_1);
and_5  g02205(new_n2533, new_n2532, new_n2582);
and_5  g02206(n11757, n3842, new_n2583);
xnor_4 g02207(new_n2583, new_n2582, new_n2584);
and_5  g02208(n11821, n4921, new_n2585_1);
and_5  g02209(n9956, n9080, new_n2586);
and_5  g02210(n11917, n5240, new_n2587);
xnor_4 g02211(new_n2587, new_n2586, new_n2588);
xor_4  g02212(new_n2588, new_n2585_1, new_n2589);
xor_4  g02213(new_n2589, new_n2584, new_n2590);
xor_4  g02214(new_n2590, new_n2581_1, new_n2591);
nor_5  g02215(new_n2538, new_n2535, new_n2592);
nand_5 g02216(new_n2537, new_n2536, new_n2593);
or_5   g02217(new_n2551_1, new_n2539, new_n2594);
xor_4  g02218(new_n2594, new_n2593, new_n2595);
nor_5  g02219(new_n2595, new_n2592, new_n2596);
xnor_4 g02220(new_n2596, new_n2591, new_n2597);
xnor_4 g02221(new_n2597, new_n2573, new_n2598);
nand_5 g02222(n9637, n7862, new_n2599);
xnor_4 g02223(new_n2572, new_n2552, new_n2600);
nor_5  g02224(new_n2600, new_n2599, new_n2601);
xnor_4 g02225(new_n2567, new_n2565, new_n2602);
xor_4  g02226(new_n2558_1, new_n2557, new_n2603);
and_5  g02227(n9956, n1333, new_n2604);
and_5  g02228(n7862, n4921, new_n2605);
nand_5 g02229(new_n2605, new_n2604, new_n2606);
or_5   g02230(new_n2606, new_n2603, new_n2607);
or_5   g02231(new_n2607, new_n2602, new_n2608);
xnor_4 g02232(new_n2570, new_n2569, new_n2609);
or_5   g02233(new_n2609, new_n2608, new_n2610);
xnor_4 g02234(new_n2600, new_n2599, new_n2611);
nor_5  g02235(new_n2611, new_n2610, new_n2612);
nor_5  g02236(new_n2612, new_n2601, new_n2613);
xnor_4 g02237(new_n2613, new_n2598, new_n2614);
xnor_4 g02238(new_n2611, new_n2610, new_n2615);
nand_5 g02239(n8595, n6877, new_n2616);
and_5  g02240(n6877, n6126, new_n2617);
and_5  g02241(n3719, n2464, new_n2618);
nor_5  g02242(new_n2618, new_n2617, new_n2619);
and_5  g02243(n6877, n3719, new_n2620);
and_5  g02244(n6126, n2464, new_n2621);
and_5  g02245(new_n2621, new_n2620, new_n2622);
and_5  g02246(n9400, n3602, new_n2623);
nor_5  g02247(new_n2623, new_n2622, new_n2624_1);
or_5   g02248(new_n2624_1, new_n2619, new_n2625);
xnor_4 g02249(new_n2625, new_n2616, new_n2626);
and_5  g02250(n3602, n2464, new_n2627);
and_5  g02251(n9400, n6126, new_n2628);
and_5  g02252(n11311, n3719, new_n2629);
xnor_4 g02253(new_n2629, new_n2628, new_n2630);
xor_4  g02254(new_n2630, new_n2627, new_n2631);
xnor_4 g02255(new_n2631, new_n2626, new_n2632);
nand_5 g02256(n9400, n3602, new_n2633);
nor_5  g02257(new_n2633, new_n2620, new_n2634);
nor_5  g02258(new_n2622, new_n2619, new_n2635);
or_5   g02259(new_n2635, new_n2634, new_n2636);
or_5   g02260(new_n2636, new_n2633, new_n2637);
or_5   g02261(new_n2637, new_n2632, new_n2638);
nand_5 g02262(n10439, n6877, new_n2639);
nand_5 g02263(n9400, n8595, new_n2640);
nor_5  g02264(new_n2629, new_n2628, new_n2641);
and_5  g02265(new_n2629, new_n2628, new_n2642);
nor_5  g02266(new_n2642, new_n2627, new_n2643);
or_5   g02267(new_n2643, new_n2641, new_n2644);
xnor_4 g02268(new_n2644, new_n2640, new_n2645);
and_5  g02269(n11311, n3602, new_n2646);
and_5  g02270(n4187, n3719, new_n2647);
xnor_4 g02271(new_n2647, new_n2621, new_n2648);
xor_4  g02272(new_n2648, new_n2646, new_n2649);
xnor_4 g02273(new_n2649, new_n2645, new_n2650);
xnor_4 g02274(new_n2650, new_n2639, new_n2651);
nor_5  g02275(new_n2625, new_n2616, new_n2652);
nor_5  g02276(new_n2631, new_n2626, new_n2653);
nor_5  g02277(new_n2653, new_n2652, new_n2654);
xnor_4 g02278(new_n2654, new_n2651, new_n2655);
nor_5  g02279(new_n2655, new_n2638, new_n2656);
and_5  g02280(n8065, n6877, new_n2657);
nand_5 g02281(n11311, n6126, new_n2658);
and_5  g02282(n4203, n3719, new_n2659);
and_5  g02283(n4187, n3602, new_n2660);
xnor_4 g02284(new_n2660, new_n2659, new_n2661);
xnor_4 g02285(new_n2661, new_n2658, new_n2662);
nor_5  g02286(new_n2647, new_n2621, new_n2663);
nor_5  g02287(new_n2648, new_n2646, new_n2664);
or_5   g02288(new_n2664, new_n2663, new_n2665);
xnor_4 g02289(new_n2665, new_n2662, new_n2666);
and_5  g02290(n10439, n9400, new_n2667);
and_5  g02291(n8595, n2464, new_n2668);
xnor_4 g02292(new_n2668, new_n2667, new_n2669);
xnor_4 g02293(new_n2669, new_n2666, new_n2670);
nor_5  g02294(new_n2644, new_n2640, new_n2671);
nor_5  g02295(new_n2649, new_n2645, new_n2672);
nor_5  g02296(new_n2672, new_n2671, new_n2673);
xnor_4 g02297(new_n2673, new_n2670, new_n2674);
nor_5  g02298(new_n2650, new_n2639, new_n2675);
nor_5  g02299(new_n2654, new_n2651, new_n2676);
nor_5  g02300(new_n2676, new_n2675, new_n2677);
xor_4  g02301(new_n2677, new_n2674, new_n2678);
xnor_4 g02302(new_n2678, new_n2657, new_n2679_1);
xnor_4 g02303(new_n2679_1, new_n2656, new_n2680);
xnor_4 g02304(new_n2655, new_n2638, new_n2681);
xnor_4 g02305(new_n2637, new_n2632, new_n2682);
or_5   g02306(new_n2633, new_n2620, new_n2683);
or_5   g02307(new_n2683, new_n2619, new_n2684);
nand_5 g02308(new_n2684, new_n2636, new_n2685);
and_5  g02309(n8433, n7236, new_n2686);
and_5  g02310(n12925, n4805, new_n2687);
and_5  g02311(new_n2687, new_n2686, new_n2688);
and_5  g02312(n7733, n4805, new_n2689);
and_5  g02313(n12925, n11478, new_n2690);
xor_4  g02314(new_n2690, new_n2689, new_n2691);
nor_5  g02315(new_n2691, new_n2688, new_n2692);
xnor_4 g02316(new_n2691, new_n2688, new_n2693);
and_5  g02317(n7236, n405, new_n2694);
and_5  g02318(n8433, n3992, new_n2695);
xor_4  g02319(new_n2695, new_n2694, new_n2696);
nor_5  g02320(new_n2696, new_n2693, new_n2697);
nor_5  g02321(new_n2697, new_n2692, new_n2698);
nand_5 g02322(n3992, n405, new_n2699);
nor_5  g02323(new_n2699, new_n2686, new_n2700);
and_5  g02324(n8433, n8384, new_n2701);
and_5  g02325(n7236, n4086, new_n2702);
or_5   g02326(new_n2702, new_n2701, new_n2703);
nor_5  g02327(new_n2703, new_n2700, new_n2704);
and_5  g02328(new_n2702, new_n2701, new_n2705);
or_5   g02329(new_n2705, new_n2704, new_n2706);
and_5  g02330(new_n2703, new_n2700, new_n2707);
nor_5  g02331(new_n2707, new_n2706, new_n2708_1);
xnor_4 g02332(new_n2708_1, new_n2698, new_n2709);
nand_5 g02333(n11478, n7733, new_n2710);
nor_5  g02334(new_n2710, new_n2687, new_n2711);
and_5  g02335(n12925, n5283, new_n2712);
and_5  g02336(n4826, n4805, new_n2713);
nor_5  g02337(new_n2713, new_n2712, new_n2714);
and_5  g02338(new_n2714, new_n2711, new_n2715);
xnor_4 g02339(new_n2713, new_n2712, new_n2716);
nor_5  g02340(new_n2716, new_n2711, new_n2717);
nor_5  g02341(new_n2717, new_n2715, new_n2718);
xnor_4 g02342(new_n2718, new_n2709, new_n2719);
nor_5  g02343(new_n2719, new_n2685, new_n2720);
xnor_4 g02344(new_n2719, new_n2685, new_n2721);
xor_4  g02345(new_n2696, new_n2693, new_n2722);
and_5  g02346(n9400, n3719, new_n2723);
and_5  g02347(n6877, n3602, new_n2724);
xnor_4 g02348(new_n2724, new_n2723, new_n2725);
nor_5  g02349(new_n2725, new_n2722, new_n2726);
nand_5 g02350(n6877, n3719, new_n2727);
xnor_4 g02351(new_n2687, new_n2686, new_n2728);
or_5   g02352(new_n2728, new_n2727, new_n2729);
xnor_4 g02353(new_n2725, new_n2722, new_n2730);
nor_5  g02354(new_n2730, new_n2729, new_n2731);
nor_5  g02355(new_n2731, new_n2726, new_n2732);
nor_5  g02356(new_n2732, new_n2721, new_n2733);
nor_5  g02357(new_n2733, new_n2720, new_n2734);
and_5  g02358(new_n2734, new_n2682, new_n2735);
nand_5 g02359(n7610, n4805, new_n2736);
and_5  g02360(new_n2713, new_n2712, new_n2737);
nor_5  g02361(new_n2714, new_n2710, new_n2738);
nor_5  g02362(new_n2738, new_n2737, new_n2739);
xnor_4 g02363(new_n2739, new_n2736, new_n2740);
and_5  g02364(n7733, n5283, new_n2741);
and_5  g02365(n12925, n137, new_n2742);
and_5  g02366(n11478, n4826, new_n2743);
xnor_4 g02367(new_n2743, new_n2742, new_n2744);
xor_4  g02368(new_n2744, new_n2741, new_n2745);
xnor_4 g02369(new_n2745, new_n2740, new_n2746);
and_5  g02370(new_n2690, new_n2689, new_n2747);
nand_5 g02371(new_n2716, new_n2747, new_n2748);
xor_4  g02372(new_n2748, new_n2746, new_n2749_1);
and_5  g02373(n7236, n217, new_n2750);
and_5  g02374(n3992, n405, new_n2751);
or_5   g02375(new_n2705, new_n2751, new_n2752);
and_5  g02376(new_n2752, new_n2703, new_n2753);
xnor_4 g02377(new_n2753, new_n2750, new_n2754);
and_5  g02378(n8384, n405, new_n2755);
and_5  g02379(n8433, n6358, new_n2756);
and_5  g02380(n4086, n3992, new_n2757);
xnor_4 g02381(new_n2757, new_n2756, new_n2758);
xor_4  g02382(new_n2758, new_n2755, new_n2759);
xnor_4 g02383(new_n2759, new_n2754, new_n2760);
nand_5 g02384(new_n2706, new_n2751, new_n2761);
xor_4  g02385(new_n2761, new_n2760, new_n2762);
xnor_4 g02386(new_n2762, new_n2749_1, new_n2763);
nor_5  g02387(new_n2708_1, new_n2698, new_n2764);
or_5   g02388(new_n2717, new_n2715, new_n2765);
nor_5  g02389(new_n2765, new_n2709, new_n2766);
nor_5  g02390(new_n2766, new_n2764, new_n2767);
xnor_4 g02391(new_n2767, new_n2763, new_n2768);
xnor_4 g02392(new_n2734, new_n2682, new_n2769);
nor_5  g02393(new_n2769, new_n2768, new_n2770);
or_5   g02394(new_n2770, new_n2735, new_n2771);
and_5  g02395(new_n2771, new_n2681, new_n2772);
nor_5  g02396(new_n2771, new_n2681, new_n2773);
or_5   g02397(new_n2761, new_n2760, new_n2774);
nand_5 g02398(n7236, n6611, new_n2775);
and_5  g02399(n3992, n217, new_n2776);
nor_5  g02400(new_n2757, new_n2756, new_n2777);
nor_5  g02401(new_n2758, new_n2755, new_n2778);
nor_5  g02402(new_n2778, new_n2777, new_n2779);
xnor_4 g02403(new_n2779, new_n2776, new_n2780);
and_5  g02404(n6358, n405, new_n2781);
and_5  g02405(n8384, n4086, new_n2782);
and_5  g02406(n8433, n5198, new_n2783);
xnor_4 g02407(new_n2783, new_n2782, new_n2784);
xor_4  g02408(new_n2784, new_n2781, new_n2785);
xnor_4 g02409(new_n2785, new_n2780, new_n2786);
xnor_4 g02410(new_n2786, new_n2775, new_n2787);
and_5  g02411(new_n2753, new_n2750, new_n2788);
nor_5  g02412(new_n2759, new_n2754, new_n2789);
nor_5  g02413(new_n2789, new_n2788, new_n2790);
xnor_4 g02414(new_n2790, new_n2787, new_n2791);
xnor_4 g02415(new_n2791, new_n2774, new_n2792);
or_5   g02416(new_n2748, new_n2746, new_n2793);
nand_5 g02417(n4970, n4805, new_n2794);
and_5  g02418(n11478, n7610, new_n2795);
nor_5  g02419(new_n2743, new_n2742, new_n2796);
nor_5  g02420(new_n2744, new_n2741, new_n2797);
nor_5  g02421(new_n2797, new_n2796, new_n2798);
xnor_4 g02422(new_n2798, new_n2795, new_n2799);
and_5  g02423(n7733, n137, new_n2800);
and_5  g02424(n5283, n4826, new_n2801);
and_5  g02425(n12925, n6294, new_n2802_1);
xnor_4 g02426(new_n2802_1, new_n2801, new_n2803);
xor_4  g02427(new_n2803, new_n2800, new_n2804);
xnor_4 g02428(new_n2804, new_n2799, new_n2805);
xnor_4 g02429(new_n2805, new_n2794, new_n2806);
nor_5  g02430(new_n2739, new_n2736, new_n2807);
nor_5  g02431(new_n2745, new_n2740, new_n2808);
nor_5  g02432(new_n2808, new_n2807, new_n2809);
xnor_4 g02433(new_n2809, new_n2806, new_n2810);
xor_4  g02434(new_n2810, new_n2793, new_n2811);
nor_5  g02435(new_n2762, new_n2749_1, new_n2812);
nor_5  g02436(new_n2767, new_n2763, new_n2813);
nor_5  g02437(new_n2813, new_n2812, new_n2814);
xor_4  g02438(new_n2814, new_n2811, new_n2815);
xnor_4 g02439(new_n2815, new_n2792, new_n2816);
nor_5  g02440(new_n2816, new_n2773, new_n2817);
nor_5  g02441(new_n2817, new_n2772, new_n2818_1);
xnor_4 g02442(new_n2818_1, new_n2680, new_n2819);
nor_5  g02443(new_n2791, new_n2774, new_n2820);
and_5  g02444(n7236, n6359, new_n2821);
and_5  g02445(n6358, n4086, new_n2822);
nor_5  g02446(new_n2783, new_n2782, new_n2823);
nor_5  g02447(new_n2784, new_n2781, new_n2824);
nor_5  g02448(new_n2824, new_n2823, new_n2825);
xnor_4 g02449(new_n2825, new_n2822, new_n2826);
and_5  g02450(n5198, n405, new_n2827);
and_5  g02451(n8433, n1471, new_n2828);
xnor_4 g02452(new_n2828, new_n2827, new_n2829);
xnor_4 g02453(new_n2829, new_n2826, new_n2830);
and_5  g02454(n8384, n217, new_n2831);
and_5  g02455(n6611, n3992, new_n2832);
xnor_4 g02456(new_n2832, new_n2831, new_n2833);
xnor_4 g02457(new_n2833, new_n2830, new_n2834);
and_5  g02458(new_n2779, new_n2776, new_n2835);
nor_5  g02459(new_n2785, new_n2780, new_n2836);
nor_5  g02460(new_n2836, new_n2835, new_n2837);
xnor_4 g02461(new_n2837, new_n2834, new_n2838);
nor_5  g02462(new_n2786, new_n2775, new_n2839);
nor_5  g02463(new_n2790, new_n2787, new_n2840);
nor_5  g02464(new_n2840, new_n2839, new_n2841);
xor_4  g02465(new_n2841, new_n2838, new_n2842);
xnor_4 g02466(new_n2842, new_n2821, new_n2843);
xnor_4 g02467(new_n2843, new_n2820, new_n2844);
nor_5  g02468(new_n2810, new_n2793, new_n2845);
and_5  g02469(n4805, n503, new_n2846);
nand_5 g02470(n4826, n137, new_n2847);
and_5  g02471(n7733, n6294, new_n2848);
and_5  g02472(n12925, n6797, new_n2849);
xnor_4 g02473(new_n2849, new_n2848, new_n2850);
xnor_4 g02474(new_n2850, new_n2847, new_n2851);
nor_5  g02475(new_n2802_1, new_n2801, new_n2852);
nor_5  g02476(new_n2803, new_n2800, new_n2853);
or_5   g02477(new_n2853, new_n2852, new_n2854);
xnor_4 g02478(new_n2854, new_n2851, new_n2855);
and_5  g02479(n11478, n4970, new_n2856);
and_5  g02480(n7610, n5283, new_n2857);
xnor_4 g02481(new_n2857, new_n2856, new_n2858);
xnor_4 g02482(new_n2858, new_n2855, new_n2859);
and_5  g02483(new_n2798, new_n2795, new_n2860);
nor_5  g02484(new_n2804, new_n2799, new_n2861);
nor_5  g02485(new_n2861, new_n2860, new_n2862);
xnor_4 g02486(new_n2862, new_n2859, new_n2863);
nor_5  g02487(new_n2805, new_n2794, new_n2864);
nor_5  g02488(new_n2809, new_n2806, new_n2865);
nor_5  g02489(new_n2865, new_n2864, new_n2866);
xor_4  g02490(new_n2866, new_n2863, new_n2867);
xnor_4 g02491(new_n2867, new_n2846, new_n2868);
xnor_4 g02492(new_n2868, new_n2845, new_n2869);
xnor_4 g02493(new_n2869, new_n2844, new_n2870);
nor_5  g02494(new_n2814, new_n2811, new_n2871);
and_5  g02495(new_n2815, new_n2792, new_n2872);
nor_5  g02496(new_n2872, new_n2871, new_n2873);
xor_4  g02497(new_n2873, new_n2870, new_n2874);
xnor_4 g02498(new_n2874, new_n2819, new_n2875);
and_5  g02499(new_n2875, new_n2615, new_n2876);
nor_5  g02500(new_n2875, new_n2615, new_n2877);
xnor_4 g02501(new_n2609, new_n2608, new_n2878);
xor_4  g02502(new_n2771, new_n2681, new_n2879_1);
xnor_4 g02503(new_n2879_1, new_n2816, new_n2880);
nor_5  g02504(new_n2880, new_n2878, new_n2881);
xnor_4 g02505(new_n2607, new_n2602, new_n2882);
xor_4  g02506(new_n2769, new_n2768, new_n2883);
nor_5  g02507(new_n2883, new_n2882, new_n2884);
xor_4  g02508(new_n2732, new_n2721, new_n2885);
and_5  g02509(n9956, n7862, new_n2886);
nor_5  g02510(new_n2886, new_n2561, new_n2887);
nor_5  g02511(new_n2887, new_n2603, new_n2888);
or_5   g02512(new_n2886, new_n2561, new_n2889);
nor_5  g02513(new_n2889, new_n2560, new_n2890);
nor_5  g02514(new_n2890, new_n2888, new_n2891);
nor_5  g02515(new_n2891, new_n2885, new_n2892);
xnor_4 g02516(new_n2891, new_n2885, new_n2893);
xnor_4 g02517(new_n2728, new_n2620, new_n2894);
and_5  g02518(new_n2894, new_n2886, new_n2895);
xor_4  g02519(new_n2605, new_n2604, new_n2896);
nor_5  g02520(new_n2896, new_n2895, new_n2897);
xnor_4 g02521(new_n2730, new_n2729, new_n2898);
xor_4  g02522(new_n2896, new_n2895, new_n2899);
and_5  g02523(new_n2899, new_n2898, new_n2900);
nor_5  g02524(new_n2900, new_n2897, new_n2901);
nor_5  g02525(new_n2901, new_n2893, new_n2902_1);
or_5   g02526(new_n2902_1, new_n2892, new_n2903);
xnor_4 g02527(new_n2883, new_n2882, new_n2904);
nor_5  g02528(new_n2904, new_n2903, new_n2905);
nor_5  g02529(new_n2905, new_n2884, new_n2906);
xnor_4 g02530(new_n2880, new_n2878, new_n2907);
nor_5  g02531(new_n2907, new_n2906, new_n2908);
or_5   g02532(new_n2908, new_n2881, new_n2909);
nor_5  g02533(new_n2909, new_n2877, new_n2910);
or_5   g02534(new_n2910, new_n2876, new_n2911);
xnor_4 g02535(new_n2911, new_n2614, new_n2912);
or_5   g02536(new_n2677, new_n2674, new_n2913);
and_5  g02537(n9400, n8065, new_n2914);
nand_5 g02538(n10439, n2464, new_n2915);
nand_5 g02539(n10391, n6877, new_n2916);
xnor_4 g02540(new_n2916, new_n2915, new_n2917);
xnor_4 g02541(new_n2917, new_n2914, new_n2918);
nor_5  g02542(new_n2661, new_n2658, new_n2919);
nor_5  g02543(new_n2665, new_n2662, new_n2920);
or_5   g02544(new_n2920, new_n2919, new_n2921);
xnor_4 g02545(new_n2921, new_n2918, new_n2922);
and_5  g02546(new_n2660, new_n2659, new_n2923);
and_5  g02547(n11311, n8595, new_n2924);
xnor_4 g02548(new_n2924, new_n2923, new_n2925);
and_5  g02549(n4203, n3602, new_n2926);
and_5  g02550(n6126, n4187, new_n2927);
and_5  g02551(n12753, n3719, new_n2928);
xnor_4 g02552(new_n2928, new_n2927, new_n2929);
xor_4  g02553(new_n2929, new_n2926, new_n2930);
xor_4  g02554(new_n2930, new_n2925, new_n2931);
xor_4  g02555(new_n2931, new_n2922, new_n2932);
nor_5  g02556(new_n2669, new_n2666, new_n2933);
nand_5 g02557(new_n2668, new_n2667, new_n2934);
or_5   g02558(new_n2673, new_n2670, new_n2935);
xor_4  g02559(new_n2935, new_n2934, new_n2936);
nor_5  g02560(new_n2936, new_n2933, new_n2937);
xnor_4 g02561(new_n2937, new_n2932, new_n2938);
xnor_4 g02562(new_n2938, new_n2913, new_n2939);
nor_5  g02563(new_n2678, new_n2657, new_n2940);
nor_5  g02564(new_n2679_1, new_n2656, new_n2941);
or_5   g02565(new_n2941, new_n2940, new_n2942);
xor_4  g02566(new_n2942, new_n2939, new_n2943);
or_5   g02567(new_n2866, new_n2863, new_n2944);
and_5  g02568(n10965, n4805, new_n2945);
and_5  g02569(n5283, n4970, new_n2946);
and_5  g02570(n11478, n503, new_n2947);
xnor_4 g02571(new_n2947, new_n2946, new_n2948);
xnor_4 g02572(new_n2948, new_n2945, new_n2949);
nor_5  g02573(new_n2850, new_n2847, new_n2950);
nor_5  g02574(new_n2854, new_n2851, new_n2951);
or_5   g02575(new_n2951, new_n2950, new_n2952);
xnor_4 g02576(new_n2952, new_n2949, new_n2953);
and_5  g02577(new_n2849, new_n2848, new_n2954);
and_5  g02578(n7610, n137, new_n2955);
xnor_4 g02579(new_n2955, new_n2954, new_n2956);
nand_5 g02580(n7733, n6797, new_n2957);
and_5  g02581(n6294, n4826, new_n2958);
and_5  g02582(n12925, n3146, new_n2959);
xnor_4 g02583(new_n2959, new_n2958, new_n2960);
xnor_4 g02584(new_n2960, new_n2957, new_n2961);
xor_4  g02585(new_n2961, new_n2956, new_n2962);
xor_4  g02586(new_n2962, new_n2953, new_n2963);
nor_5  g02587(new_n2858, new_n2855, new_n2964);
nand_5 g02588(new_n2857, new_n2856, new_n2965);
or_5   g02589(new_n2862, new_n2859, new_n2966);
xor_4  g02590(new_n2966, new_n2965, new_n2967);
nor_5  g02591(new_n2967, new_n2964, new_n2968);
xnor_4 g02592(new_n2968, new_n2963, new_n2969);
xnor_4 g02593(new_n2969, new_n2944, new_n2970);
nor_5  g02594(new_n2867, new_n2846, new_n2971);
nor_5  g02595(new_n2868, new_n2845, new_n2972);
or_5   g02596(new_n2972, new_n2971, new_n2973);
xor_4  g02597(new_n2973, new_n2970, new_n2974);
or_5   g02598(new_n2841, new_n2838, new_n2975);
and_5  g02599(n11296, n7236, new_n2976);
and_5  g02600(n8384, n6611, new_n2977);
and_5  g02601(n6359, n3992, new_n2978);
xnor_4 g02602(new_n2978, new_n2977, new_n2979);
xnor_4 g02603(new_n2979, new_n2976, new_n2980);
and_5  g02604(new_n2825, new_n2822, new_n2981);
nor_5  g02605(new_n2829, new_n2826, new_n2982);
or_5   g02606(new_n2982, new_n2981, new_n2983);
xnor_4 g02607(new_n2983, new_n2980, new_n2984);
and_5  g02608(new_n2828, new_n2827, new_n2985);
and_5  g02609(n6358, n217, new_n2986);
xnor_4 g02610(new_n2986, new_n2985, new_n2987);
nand_5 g02611(n1471, n405, new_n2988);
and_5  g02612(n5198, n4086, new_n2989);
and_5  g02613(n8433, n7646, new_n2990);
xnor_4 g02614(new_n2990, new_n2989, new_n2991);
xnor_4 g02615(new_n2991, new_n2988, new_n2992);
xor_4  g02616(new_n2992, new_n2987, new_n2993);
xor_4  g02617(new_n2993, new_n2984, new_n2994);
nor_5  g02618(new_n2833, new_n2830, new_n2995);
nand_5 g02619(new_n2832, new_n2831, new_n2996);
or_5   g02620(new_n2837, new_n2834, new_n2997);
xor_4  g02621(new_n2997, new_n2996, new_n2998);
nor_5  g02622(new_n2998, new_n2995, new_n2999);
xnor_4 g02623(new_n2999, new_n2994, new_n3000);
xnor_4 g02624(new_n3000, new_n2975, new_n3001);
nor_5  g02625(new_n2842, new_n2821, new_n3002);
nor_5  g02626(new_n2843, new_n2820, new_n3003);
or_5   g02627(new_n3003, new_n3002, new_n3004);
xor_4  g02628(new_n3004, new_n3001, new_n3005);
xnor_4 g02629(new_n3005, new_n2974, new_n3006);
nor_5  g02630(new_n2869, new_n2844, new_n3007);
nor_5  g02631(new_n2873, new_n2870, new_n3008);
or_5   g02632(new_n3008, new_n3007, new_n3009);
xor_4  g02633(new_n3009, new_n3006, new_n3010);
xnor_4 g02634(new_n3010, new_n2943, new_n3011);
and_5  g02635(new_n2818_1, new_n2680, new_n3012);
nor_5  g02636(new_n2874, new_n2819, new_n3013);
or_5   g02637(new_n3013, new_n3012, new_n3014);
xnor_4 g02638(new_n3014, new_n3011, new_n3015);
xnor_4 g02639(new_n3015, new_n2912, n844);
nand_5 g02640(n7456, n6687, new_n3017);
and_5  g02641(n12591, n6687, new_n3018);
and_5  g02642(n4189, n1798, new_n3019);
nor_5  g02643(new_n3019, new_n3018, new_n3020);
and_5  g02644(n6687, n1798, new_n3021);
and_5  g02645(n12591, n4189, new_n3022_1);
and_5  g02646(new_n3022_1, new_n3021, new_n3023);
and_5  g02647(n3932, n2564, new_n3024);
nor_5  g02648(new_n3024, new_n3023, new_n3025);
or_5   g02649(new_n3025, new_n3020, new_n3026);
xnor_4 g02650(new_n3026, new_n3017, new_n3027);
and_5  g02651(n4189, n3932, new_n3028);
and_5  g02652(n12591, n2564, new_n3029);
and_5  g02653(n6770, n1798, new_n3030);
xnor_4 g02654(new_n3030, new_n3029, new_n3031);
xor_4  g02655(new_n3031, new_n3028, new_n3032);
xnor_4 g02656(new_n3032, new_n3027, new_n3033);
nand_5 g02657(n3932, n2564, new_n3034);
or_5   g02658(new_n3034, new_n3021, new_n3035);
or_5   g02659(new_n3023, new_n3020, new_n3036);
and_5  g02660(new_n3036, new_n3035, new_n3037);
nand_5 g02661(new_n3037, new_n3024, new_n3038);
xnor_4 g02662(new_n3038, new_n3033, new_n3039);
nor_5  g02663(new_n3035, new_n3020, new_n3040);
or_5   g02664(new_n3040, new_n3037, new_n3041);
nand_5 g02665(n8336, n6703, new_n3042);
and_5  g02666(n11876, n11222, new_n3043);
and_5  g02667(n12069, n5645, new_n3044);
xnor_4 g02668(new_n3044, new_n3043, new_n3045);
nor_5  g02669(new_n3045, new_n3042, new_n3046);
and_5  g02670(n9640, n8336, new_n3047);
and_5  g02671(n10928, n6703, new_n3048);
xor_4  g02672(new_n3048, new_n3047, new_n3049);
and_5  g02673(new_n3049, new_n3046, new_n3050);
and_5  g02674(new_n3044, new_n3043, new_n3051);
and_5  g02675(n12391, n5645, new_n3052);
and_5  g02676(n12069, n1067, new_n3053);
xor_4  g02677(new_n3053, new_n3052, new_n3054);
xnor_4 g02678(new_n3054, new_n3051, new_n3055);
and_5  g02679(n11222, n10898, new_n3056);
and_5  g02680(n11876, n11153, new_n3057);
xor_4  g02681(new_n3057, new_n3056, new_n3058);
xor_4  g02682(new_n3058, new_n3055, new_n3059);
xnor_4 g02683(new_n3049, new_n3046, new_n3060);
nor_5  g02684(new_n3060, new_n3059, new_n3061);
nor_5  g02685(new_n3061, new_n3050, new_n3062);
and_5  g02686(n8336, n6703, new_n3063);
nand_5 g02687(n10928, n9640, new_n3064);
or_5   g02688(new_n3064, new_n3063, new_n3065);
and_5  g02689(n6986, n6703, new_n3066);
and_5  g02690(n8336, n3022, new_n3067);
nor_5  g02691(new_n3067, new_n3066, new_n3068);
and_5  g02692(n6986, n3022, new_n3069);
and_5  g02693(new_n3069, new_n3063, new_n3070);
or_5   g02694(new_n3070, new_n3068, new_n3071_1);
and_5  g02695(new_n3071_1, new_n3065, new_n3072);
nor_5  g02696(new_n3068, new_n3065, new_n3073);
or_5   g02697(new_n3073, new_n3072, new_n3074);
xnor_4 g02698(new_n3074, new_n3062, new_n3075);
nand_5 g02699(new_n3053, new_n3052, new_n3076);
and_5  g02700(n12069, n8665, new_n3077);
and_5  g02701(n12391, n1067, new_n3078);
and_5  g02702(n7891, n5645, new_n3079);
xnor_4 g02703(new_n3079, new_n3078, new_n3080);
xor_4  g02704(new_n3080, new_n3077, new_n3081);
xor_4  g02705(new_n3081, new_n3076, new_n3082);
nor_5  g02706(new_n3054, new_n3051, new_n3083);
nor_5  g02707(new_n3058, new_n3055, new_n3084);
nor_5  g02708(new_n3084, new_n3083, new_n3085);
nand_5 g02709(n11153, n10898, new_n3086);
or_5   g02710(new_n3086, new_n3043, new_n3087);
and_5  g02711(n11876, n5314, new_n3088);
and_5  g02712(n11222, n3754, new_n3089);
nor_5  g02713(new_n3089, new_n3088, new_n3090);
and_5  g02714(new_n3090, new_n3087, new_n3091);
and_5  g02715(n5314, n3754, new_n3092);
and_5  g02716(new_n3092, new_n3043, new_n3093);
nor_5  g02717(new_n3093, new_n3091, new_n3094);
or_5   g02718(new_n3090, new_n3087, new_n3095);
and_5  g02719(new_n3095, new_n3094, new_n3096);
xnor_4 g02720(new_n3096, new_n3085, new_n3097);
xnor_4 g02721(new_n3097, new_n3082, new_n3098);
xor_4  g02722(new_n3098, new_n3075, new_n3099);
nor_5  g02723(new_n3099, new_n3041, new_n3100);
xnor_4 g02724(new_n3045, new_n3063, new_n3101);
and_5  g02725(new_n3101, new_n3021, new_n3102);
and_5  g02726(n2564, n1798, new_n3103);
and_5  g02727(n6687, n3932, new_n3104);
xor_4  g02728(new_n3104, new_n3103, new_n3105);
nor_5  g02729(new_n3105, new_n3102, new_n3106);
xnor_4 g02730(new_n3060, new_n3059, new_n3107);
xor_4  g02731(new_n3105, new_n3102, new_n3108);
and_5  g02732(new_n3108, new_n3107, new_n3109);
or_5   g02733(new_n3109, new_n3106, new_n3110);
xnor_4 g02734(new_n3099, new_n3041, new_n3111);
nor_5  g02735(new_n3111, new_n3110, new_n3112);
nor_5  g02736(new_n3112, new_n3100, new_n3113);
xnor_4 g02737(new_n3113, new_n3039, new_n3114);
or_5   g02738(new_n3081, new_n3076, new_n3115);
nand_5 g02739(n12069, n11922, new_n3116);
nor_5  g02740(new_n3079, new_n3078, new_n3117);
nor_5  g02741(new_n3080, new_n3077, new_n3118);
or_5   g02742(new_n3118, new_n3117, new_n3119);
xnor_4 g02743(new_n3119, new_n3116, new_n3120);
and_5  g02744(n7160, n5645, new_n3121);
and_5  g02745(n7891, n1067, new_n3122);
and_5  g02746(n12391, n8665, new_n3123);
xnor_4 g02747(new_n3123, new_n3122, new_n3124_1);
xor_4  g02748(new_n3124_1, new_n3121, new_n3125);
xnor_4 g02749(new_n3125, new_n3120, new_n3126);
xor_4  g02750(new_n3126, new_n3115, new_n3127);
and_5  g02751(n11222, n2749, new_n3128);
and_5  g02752(n11153, n10898, new_n3129);
nor_5  g02753(new_n3093, new_n3129, new_n3130);
nor_5  g02754(new_n3130, new_n3090, new_n3131);
xnor_4 g02755(new_n3131, new_n3128, new_n3132);
and_5  g02756(n10898, n5314, new_n3133);
and_5  g02757(n11153, n3754, new_n3134);
and_5  g02758(n11876, n996, new_n3135);
xnor_4 g02759(new_n3135, new_n3134, new_n3136);
xor_4  g02760(new_n3136, new_n3133, new_n3137);
xnor_4 g02761(new_n3137, new_n3132, new_n3138);
or_5   g02762(new_n3094, new_n3086, new_n3139);
xor_4  g02763(new_n3139, new_n3138, new_n3140);
xnor_4 g02764(new_n3140, new_n3127, new_n3141);
nor_5  g02765(new_n3096, new_n3085, new_n3142);
nor_5  g02766(new_n3097, new_n3082, new_n3143);
nor_5  g02767(new_n3143, new_n3142, new_n3144);
xor_4  g02768(new_n3144, new_n3141, new_n3145);
nand_5 g02769(n11023, n8336, new_n3146_1);
and_5  g02770(n10928, n9640, new_n3147);
nor_5  g02771(new_n3070, new_n3147, new_n3148);
or_5   g02772(new_n3148, new_n3068, new_n3149);
xnor_4 g02773(new_n3149, new_n3146_1, new_n3150);
and_5  g02774(n9640, n6986, new_n3151);
and_5  g02775(n10928, n3022, new_n3152);
and_5  g02776(n6703, n2226, new_n3153);
xnor_4 g02777(new_n3153, new_n3152, new_n3154);
xor_4  g02778(new_n3154, new_n3151, new_n3155);
xnor_4 g02779(new_n3155, new_n3150, new_n3156);
nand_5 g02780(new_n3072, new_n3147, new_n3157);
xnor_4 g02781(new_n3157, new_n3156, new_n3158);
and_5  g02782(new_n3074, new_n3062, new_n3159);
nor_5  g02783(new_n3098, new_n3075, new_n3160);
nor_5  g02784(new_n3160, new_n3159, new_n3161);
xor_4  g02785(new_n3161, new_n3158, new_n3162);
xnor_4 g02786(new_n3162, new_n3145, new_n3163);
xor_4  g02787(new_n3163, new_n3114, n911);
nand_5 g02788(n6687, n3842, new_n3165);
and_5  g02789(n11917, n6687, new_n3166);
and_5  g02790(n9956, n4189, new_n3167);
nor_5  g02791(new_n3167, new_n3166, new_n3168);
and_5  g02792(n9956, n6687, new_n3169);
and_5  g02793(n11917, n4189, new_n3170);
and_5  g02794(new_n3170, new_n3169, new_n3171);
and_5  g02795(n4921, n2564, new_n3172_1);
nor_5  g02796(new_n3172_1, new_n3171, new_n3173);
or_5   g02797(new_n3173, new_n3168, new_n3174);
xor_4  g02798(new_n3174, new_n3165, new_n3175);
and_5  g02799(n4921, n4189, new_n3176);
and_5  g02800(n11917, n2564, new_n3177);
and_5  g02801(n9956, n6770, new_n3178);
xnor_4 g02802(new_n3178, new_n3177, new_n3179);
xnor_4 g02803(new_n3179, new_n3176, new_n3180);
xnor_4 g02804(new_n3180, new_n3175, new_n3181);
nor_5  g02805(new_n3171, new_n3168, new_n3182);
and_5  g02806(n9956, n2564, new_n3183);
and_5  g02807(n6687, n4921, new_n3184);
nand_5 g02808(new_n3184, new_n3183, new_n3185);
or_5   g02809(new_n3185, new_n3182, new_n3186);
or_5   g02810(new_n3186, new_n3181, new_n3187);
nand_5 g02811(n6687, n2577, new_n3188);
nor_5  g02812(new_n3174, new_n3165, new_n3189);
and_5  g02813(new_n3180, new_n3175, new_n3190);
nor_5  g02814(new_n3190, new_n3189, new_n3191);
xnor_4 g02815(new_n3191, new_n3188, new_n3192);
nand_5 g02816(n3842, n2564, new_n3193);
nor_5  g02817(new_n3178, new_n3177, new_n3194);
and_5  g02818(new_n3178, new_n3177, new_n3195);
nor_5  g02819(new_n3195, new_n3176, new_n3196);
or_5   g02820(new_n3196, new_n3194, new_n3197);
xnor_4 g02821(new_n3197, new_n3193, new_n3198);
and_5  g02822(n6770, n4921, new_n3199);
and_5  g02823(n9956, n9920, new_n3200);
xnor_4 g02824(new_n3200, new_n3170, new_n3201);
xor_4  g02825(new_n3201, new_n3199, new_n3202);
xnor_4 g02826(new_n3202, new_n3198, new_n3203);
xnor_4 g02827(new_n3203, new_n3192, new_n3204);
xor_4  g02828(new_n3204, new_n3187, new_n3205);
xor_4  g02829(new_n3186, new_n3181, new_n3206);
nand_5 g02830(n8595, n8336, new_n3207);
and_5  g02831(n8336, n6126, new_n3208);
and_5  g02832(n6986, n3719, new_n3209);
nor_5  g02833(new_n3209, new_n3208, new_n3210);
and_5  g02834(n8336, n3719, new_n3211);
and_5  g02835(n6986, n6126, new_n3212);
and_5  g02836(new_n3212, new_n3211, new_n3213);
and_5  g02837(n10928, n3602, new_n3214_1);
nor_5  g02838(new_n3214_1, new_n3213, new_n3215);
or_5   g02839(new_n3215, new_n3210, new_n3216);
xnor_4 g02840(new_n3216, new_n3207, new_n3217);
and_5  g02841(n6986, n3602, new_n3218);
and_5  g02842(n10928, n6126, new_n3219);
and_5  g02843(n3719, n2226, new_n3220);
xnor_4 g02844(new_n3220, new_n3219, new_n3221);
xor_4  g02845(new_n3221, new_n3218, new_n3222);
xnor_4 g02846(new_n3222, new_n3217, new_n3223);
nand_5 g02847(n10928, n3602, new_n3224);
or_5   g02848(new_n3224, new_n3211, new_n3225);
or_5   g02849(new_n3213, new_n3210, new_n3226);
and_5  g02850(new_n3226, new_n3225, new_n3227);
nand_5 g02851(new_n3227, new_n3214_1, new_n3228);
xnor_4 g02852(new_n3228, new_n3223, new_n3229);
nand_5 g02853(n12069, n7610, new_n3230_1);
and_5  g02854(n12069, n4826, new_n3231);
and_5  g02855(n12925, n7891, new_n3232);
nor_5  g02856(new_n3232, new_n3231, new_n3233);
and_5  g02857(n12925, n12069, new_n3234);
and_5  g02858(n7891, n4826, new_n3235);
and_5  g02859(new_n3235, new_n3234, new_n3236);
and_5  g02860(n12391, n7733, new_n3237);
nor_5  g02861(new_n3237, new_n3236, new_n3238);
or_5   g02862(new_n3238, new_n3233, new_n3239);
xnor_4 g02863(new_n3239, new_n3230_1, new_n3240);
and_5  g02864(n7891, n7733, new_n3241);
and_5  g02865(n12925, n7160, new_n3242);
and_5  g02866(n12391, n4826, new_n3243);
xnor_4 g02867(new_n3243, new_n3242, new_n3244);
xor_4  g02868(new_n3244, new_n3241, new_n3245);
xnor_4 g02869(new_n3245, new_n3240, new_n3246);
nor_5  g02870(new_n3236, new_n3233, new_n3247);
and_5  g02871(n12925, n12391, new_n3248);
and_5  g02872(n12069, n7733, new_n3249);
nand_5 g02873(new_n3249, new_n3248, new_n3250);
or_5   g02874(new_n3250, new_n3247, new_n3251);
xor_4  g02875(new_n3251, new_n3246, new_n3252);
nand_5 g02876(n11222, n217, new_n3253);
and_5  g02877(n8433, n5314, new_n3254);
and_5  g02878(n11222, n4086, new_n3255);
nor_5  g02879(new_n3255, new_n3254, new_n3256);
and_5  g02880(new_n3255, new_n3254, new_n3257);
and_5  g02881(n11153, n405, new_n3258);
nor_5  g02882(new_n3258, new_n3257, new_n3259);
or_5   g02883(new_n3259, new_n3256, new_n3260);
xor_4  g02884(new_n3260, new_n3253, new_n3261);
and_5  g02885(n5314, n405, new_n3262);
and_5  g02886(n8433, n996, new_n3263);
and_5  g02887(n11153, n4086, new_n3264);
xnor_4 g02888(new_n3264, new_n3263, new_n3265);
xnor_4 g02889(new_n3265, new_n3262, new_n3266);
xnor_4 g02890(new_n3266, new_n3261, new_n3267);
nand_5 g02891(n11153, n405, new_n3268);
and_5  g02892(n11222, n8433, new_n3269);
or_5   g02893(new_n3269, new_n3268, new_n3270);
and_5  g02894(new_n3270, new_n3256, new_n3271);
nor_5  g02895(new_n3271, new_n3257, new_n3272_1);
or_5   g02896(new_n3272_1, new_n3268, new_n3273);
xor_4  g02897(new_n3273, new_n3267, new_n3274);
xnor_4 g02898(new_n3274, new_n3252, new_n3275);
and_5  g02899(new_n3269, new_n3234, new_n3276);
and_5  g02900(n11153, n8433, new_n3277);
and_5  g02901(n11222, n405, new_n3278);
xor_4  g02902(new_n3278, new_n3277, new_n3279);
nor_5  g02903(new_n3279, new_n3276, new_n3280);
xnor_4 g02904(new_n3279, new_n3276, new_n3281);
xor_4  g02905(new_n3249, new_n3248, new_n3282);
nor_5  g02906(new_n3282, new_n3281, new_n3283);
nor_5  g02907(new_n3283, new_n3280, new_n3284);
or_5   g02908(new_n3270, new_n3256, new_n3285);
and_5  g02909(new_n3285, new_n3272_1, new_n3286);
nor_5  g02910(new_n3286, new_n3284, new_n3287_1);
xnor_4 g02911(new_n3286, new_n3284, new_n3288);
nand_5 g02912(n12391, n7733, new_n3289);
nor_5  g02913(new_n3289, new_n3234, new_n3290);
nor_5  g02914(new_n3290, new_n3247, new_n3291);
or_5   g02915(new_n3289, new_n3234, new_n3292);
nor_5  g02916(new_n3292, new_n3233, new_n3293);
nor_5  g02917(new_n3293, new_n3291, new_n3294);
nor_5  g02918(new_n3294, new_n3288, new_n3295);
nor_5  g02919(new_n3295, new_n3287_1, new_n3296);
xor_4  g02920(new_n3296, new_n3275, new_n3297);
xnor_4 g02921(new_n3297, new_n3229, new_n3298);
nor_5  g02922(new_n3225, new_n3210, new_n3299);
or_5   g02923(new_n3299, new_n3227, new_n3300);
xor_4  g02924(new_n3294, new_n3288, new_n3301);
nor_5  g02925(new_n3301, new_n3300, new_n3302);
xnor_4 g02926(new_n3301, new_n3300, new_n3303);
xor_4  g02927(new_n3282, new_n3281, new_n3304);
and_5  g02928(n10928, n3719, new_n3305);
and_5  g02929(n8336, n3602, new_n3306);
xnor_4 g02930(new_n3306, new_n3305, new_n3307);
nor_5  g02931(new_n3307, new_n3304, new_n3308);
nand_5 g02932(n8336, n3719, new_n3309);
xnor_4 g02933(new_n3269, new_n3234, new_n3310);
or_5   g02934(new_n3310, new_n3309, new_n3311);
xnor_4 g02935(new_n3307, new_n3304, new_n3312);
nor_5  g02936(new_n3312, new_n3311, new_n3313);
nor_5  g02937(new_n3313, new_n3308, new_n3314);
nor_5  g02938(new_n3314, new_n3303, new_n3315);
nor_5  g02939(new_n3315, new_n3302, new_n3316);
xor_4  g02940(new_n3316, new_n3298, new_n3317);
nor_5  g02941(new_n3317, new_n3206, new_n3318);
xor_4  g02942(new_n3314, new_n3303, new_n3319);
nand_5 g02943(n4921, n2564, new_n3320);
nor_5  g02944(new_n3320, new_n3169, new_n3321);
nor_5  g02945(new_n3321, new_n3182, new_n3322);
or_5   g02946(new_n3320, new_n3169, new_n3323);
nor_5  g02947(new_n3323, new_n3168, new_n3324);
nor_5  g02948(new_n3324, new_n3322, new_n3325);
nor_5  g02949(new_n3325, new_n3319, new_n3326);
xnor_4 g02950(new_n3325, new_n3319, new_n3327);
xnor_4 g02951(new_n3310, new_n3211, new_n3328);
and_5  g02952(new_n3328, new_n3169, new_n3329);
xor_4  g02953(new_n3184, new_n3183, new_n3330);
nor_5  g02954(new_n3330, new_n3329, new_n3331);
xnor_4 g02955(new_n3312, new_n3311, new_n3332);
xor_4  g02956(new_n3330, new_n3329, new_n3333);
and_5  g02957(new_n3333, new_n3332, new_n3334);
nor_5  g02958(new_n3334, new_n3331, new_n3335);
nor_5  g02959(new_n3335, new_n3327, new_n3336);
nor_5  g02960(new_n3336, new_n3326, new_n3337);
xnor_4 g02961(new_n3317, new_n3206, new_n3338);
nor_5  g02962(new_n3338, new_n3337, new_n3339_1);
nor_5  g02963(new_n3339_1, new_n3318, new_n3340);
xnor_4 g02964(new_n3340, new_n3205, new_n3341);
or_5   g02965(new_n3228, new_n3223, new_n3342_1);
nand_5 g02966(n10439, n8336, new_n3343);
nor_5  g02967(new_n3216, new_n3207, new_n3344);
nor_5  g02968(new_n3222, new_n3217, new_n3345);
nor_5  g02969(new_n3345, new_n3344, new_n3346);
xnor_4 g02970(new_n3346, new_n3343, new_n3347);
nand_5 g02971(n10928, n8595, new_n3348);
nor_5  g02972(new_n3220, new_n3219, new_n3349);
and_5  g02973(new_n3220, new_n3219, new_n3350);
nor_5  g02974(new_n3350, new_n3218, new_n3351);
or_5   g02975(new_n3351, new_n3349, new_n3352);
xnor_4 g02976(new_n3352, new_n3348, new_n3353);
and_5  g02977(n3602, n2226, new_n3354);
and_5  g02978(n3719, n1094, new_n3355);
xnor_4 g02979(new_n3355, new_n3212, new_n3356);
xor_4  g02980(new_n3356, new_n3354, new_n3357);
xnor_4 g02981(new_n3357, new_n3353, new_n3358);
xnor_4 g02982(new_n3358, new_n3347, new_n3359);
xnor_4 g02983(new_n3359, new_n3342_1, new_n3360);
or_5   g02984(new_n3273, new_n3267, new_n3361);
and_5  g02985(n11222, n6611, new_n3362);
nand_5 g02986(n11153, n217, new_n3363);
and_5  g02987(n996, n405, new_n3364);
and_5  g02988(n5314, n4086, new_n3365);
and_5  g02989(n8433, n5767, new_n3366);
xnor_4 g02990(new_n3366, new_n3365, new_n3367);
xor_4  g02991(new_n3367, new_n3364, new_n3368);
xnor_4 g02992(new_n3368, new_n3363, new_n3369);
nor_5  g02993(new_n3264, new_n3263, new_n3370);
and_5  g02994(new_n3264, new_n3263, new_n3371);
nor_5  g02995(new_n3371, new_n3262, new_n3372);
or_5   g02996(new_n3372, new_n3370, new_n3373);
xor_4  g02997(new_n3373, new_n3369, new_n3374);
xnor_4 g02998(new_n3374, new_n3362, new_n3375);
nor_5  g02999(new_n3260, new_n3253, new_n3376);
and_5  g03000(new_n3266, new_n3261, new_n3377);
nor_5  g03001(new_n3377, new_n3376, new_n3378);
xnor_4 g03002(new_n3378, new_n3375, new_n3379);
xor_4  g03003(new_n3379, new_n3361, new_n3380);
or_5   g03004(new_n3251, new_n3246, new_n3381);
nand_5 g03005(n12069, n4970, new_n3382);
and_5  g03006(n12391, n7610, new_n3383);
nor_5  g03007(new_n3243, new_n3242, new_n3384);
nor_5  g03008(new_n3244, new_n3241, new_n3385);
nor_5  g03009(new_n3385, new_n3384, new_n3386);
xnor_4 g03010(new_n3386, new_n3383, new_n3387);
and_5  g03011(n7733, n7160, new_n3388);
and_5  g03012(n12925, n4828, new_n3389);
xnor_4 g03013(new_n3389, new_n3235, new_n3390);
xor_4  g03014(new_n3390, new_n3388, new_n3391);
xnor_4 g03015(new_n3391, new_n3387, new_n3392);
xnor_4 g03016(new_n3392, new_n3382, new_n3393);
nor_5  g03017(new_n3239, new_n3230_1, new_n3394);
nor_5  g03018(new_n3245, new_n3240, new_n3395);
nor_5  g03019(new_n3395, new_n3394, new_n3396);
xnor_4 g03020(new_n3396, new_n3393, new_n3397);
xor_4  g03021(new_n3397, new_n3381, new_n3398);
nor_5  g03022(new_n3274, new_n3252, new_n3399);
nor_5  g03023(new_n3296, new_n3275, new_n3400);
nor_5  g03024(new_n3400, new_n3399, new_n3401);
xnor_4 g03025(new_n3401, new_n3398, new_n3402);
xor_4  g03026(new_n3402, new_n3380, new_n3403);
xnor_4 g03027(new_n3403, new_n3360, new_n3404);
nor_5  g03028(new_n3297, new_n3229, new_n3405);
nor_5  g03029(new_n3316, new_n3298, new_n3406);
nor_5  g03030(new_n3406, new_n3405, new_n3407);
xnor_4 g03031(new_n3407, new_n3404, new_n3408);
xor_4  g03032(new_n3408, new_n3341, n992);
and_5  g03033(n7265, n6687, new_n3410);
and_5  g03034(n8336, n7946, new_n3411);
and_5  g03035(n11222, n9763, new_n3412);
and_5  g03036(n12069, n2558, new_n3413);
xnor_4 g03037(new_n3413, new_n3412, new_n3414);
xnor_4 g03038(new_n3414, new_n3411, new_n3415);
xor_4  g03039(new_n3415, new_n3410, n1020);
xor_4  g03040(new_n1675, new_n1674, n1136);
xnor_4 g03041(new_n3338, new_n3337, n1138);
nand_5 g03042(n12591, n11757, new_n3419);
and_5  g03043(n5240, n3932, new_n3420);
and_5  g03044(n11821, n1798, new_n3421);
xnor_4 g03045(new_n3421, new_n3420, new_n3422);
xnor_4 g03046(new_n3422, new_n3419, new_n3423);
and_5  g03047(n5240, n1798, new_n3424);
and_5  g03048(n12591, n3172, new_n3425);
nor_5  g03049(new_n3425, new_n3424, new_n3426);
nand_5 g03050(new_n3425, new_n3424, new_n3427);
nand_5 g03051(n11757, n3932, new_n3428);
and_5  g03052(new_n3428, new_n3427, new_n3429);
or_5   g03053(new_n3429, new_n3426, new_n3430);
xnor_4 g03054(new_n3430, new_n3423, new_n3431);
nand_5 g03055(n7456, n1333, new_n3432);
and_5  g03056(n11757, n1798, new_n3433);
and_5  g03057(n12591, n1333, new_n3434);
nor_5  g03058(new_n3434, new_n3433, new_n3435);
nand_5 g03059(new_n3434, new_n3433, new_n3436);
nand_5 g03060(n3932, n3172, new_n3437);
and_5  g03061(new_n3437, new_n3436, new_n3438);
or_5   g03062(new_n3438, new_n3435, new_n3439);
nor_5  g03063(new_n3439, new_n3432, new_n3440);
xnor_4 g03064(new_n3439, new_n3432, new_n3441);
xnor_4 g03065(new_n3425, new_n3424, new_n3442);
xnor_4 g03066(new_n3442, new_n3428, new_n3443);
nor_5  g03067(new_n3443, new_n3441, new_n3444);
nor_5  g03068(new_n3444, new_n3440, new_n3445);
and_5  g03069(n11662, n1333, new_n3446);
and_5  g03070(n7456, n3172, new_n3447);
xnor_4 g03071(new_n3447, new_n3446, new_n3448);
xnor_4 g03072(new_n3448, new_n3445, new_n3449);
xnor_4 g03073(new_n3449, new_n3431, new_n3450);
and_5  g03074(n11662, n7862, new_n3451);
xor_4  g03075(new_n3443, new_n3441, new_n3452);
nor_5  g03076(new_n3452, new_n3451, new_n3453);
xnor_4 g03077(new_n3452, new_n3451, new_n3454);
nand_5 g03078(n7862, n7456, new_n3455);
and_5  g03079(n3172, n1798, new_n3456_1);
and_5  g03080(n12591, n7862, new_n3457);
and_5  g03081(new_n3457, new_n3456_1, new_n3458);
nor_5  g03082(new_n3457, new_n3456_1, new_n3459);
nand_5 g03083(n3932, n1333, new_n3460);
nor_5  g03084(new_n3460, new_n3459, new_n3461);
nor_5  g03085(new_n3461, new_n3458, new_n3462);
nor_5  g03086(new_n3462, new_n3455, new_n3463);
xnor_4 g03087(new_n3462, new_n3455, new_n3464);
xnor_4 g03088(new_n3434, new_n3433, new_n3465);
xnor_4 g03089(new_n3465, new_n3437, new_n3466);
nor_5  g03090(new_n3466, new_n3464, new_n3467);
or_5   g03091(new_n3467, new_n3463, new_n3468);
nor_5  g03092(new_n3468, new_n3454, new_n3469);
or_5   g03093(new_n3469, new_n3453, new_n3470);
or_5   g03094(new_n3470, new_n3450, new_n3471);
nor_5  g03095(new_n3422, new_n3419, new_n3472);
nor_5  g03096(new_n3430, new_n3423, new_n3473);
or_5   g03097(new_n3473, new_n3472, new_n3474);
and_5  g03098(n10327, n1333, new_n3475);
and_5  g03099(n11662, n3172, new_n3476);
and_5  g03100(n9583, n7862, new_n3477);
xnor_4 g03101(new_n3477, new_n3476, new_n3478);
xnor_4 g03102(new_n3478, new_n3475, new_n3479);
xnor_4 g03103(new_n3479, new_n3474, new_n3480);
and_5  g03104(new_n3421, new_n3420, new_n3481);
and_5  g03105(n11757, n7456, new_n3482);
xnor_4 g03106(new_n3482, new_n3481, new_n3483);
nand_5 g03107(n11821, n3932, new_n3484);
and_5  g03108(n12591, n5240, new_n3485);
and_5  g03109(n9080, n1798, new_n3486);
xnor_4 g03110(new_n3486, new_n3485, new_n3487);
xnor_4 g03111(new_n3487, new_n3484, new_n3488);
xor_4  g03112(new_n3488, new_n3483, new_n3489);
xor_4  g03113(new_n3489, new_n3480, new_n3490);
nor_5  g03114(new_n3448, new_n3445, new_n3491);
nand_5 g03115(new_n3447, new_n3446, new_n3492);
or_5   g03116(new_n3449, new_n3431, new_n3493);
xor_4  g03117(new_n3493, new_n3492, new_n3494);
nor_5  g03118(new_n3494, new_n3491, new_n3495);
xnor_4 g03119(new_n3495, new_n3490, new_n3496);
xnor_4 g03120(new_n3496, new_n3471, new_n3497);
and_5  g03121(n10327, n7862, new_n3498);
xor_4  g03122(new_n3470, new_n3450, new_n3499);
and_5  g03123(new_n3499, new_n3498, new_n3500);
xnor_4 g03124(new_n3466, new_n3464, new_n3501);
xor_4  g03125(new_n3457, new_n3456_1, new_n3502);
and_5  g03126(n1798, n1333, new_n3503);
and_5  g03127(n7862, n3932, new_n3504);
nand_5 g03128(new_n3504, new_n3503, new_n3505);
or_5   g03129(new_n3505, new_n3502, new_n3506);
or_5   g03130(new_n3506, new_n3501, new_n3507);
xor_4  g03131(new_n3468, new_n3454, new_n3508);
or_5   g03132(new_n3508, new_n3507, new_n3509);
xnor_4 g03133(new_n3499, new_n3498, new_n3510);
nor_5  g03134(new_n3510, new_n3509, new_n3511);
nor_5  g03135(new_n3511, new_n3500, new_n3512);
xnor_4 g03136(new_n3512, new_n3497, new_n3513);
nand_5 g03137(n11311, n3022, new_n3514);
and_5  g03138(n9640, n4187, new_n3515);
and_5  g03139(n6703, n4203, new_n3516);
xnor_4 g03140(new_n3516, new_n3515, new_n3517);
xnor_4 g03141(new_n3517, new_n3514, new_n3518);
and_5  g03142(n6703, n4187, new_n3519);
and_5  g03143(n3022, n2464, new_n3520);
nor_5  g03144(new_n3520, new_n3519, new_n3521);
nand_5 g03145(new_n3520, new_n3519, new_n3522);
nand_5 g03146(n11311, n9640, new_n3523);
and_5  g03147(new_n3523, new_n3522, new_n3524);
or_5   g03148(new_n3524, new_n3521, new_n3525);
xnor_4 g03149(new_n3525, new_n3518, new_n3526);
and_5  g03150(n10451, n9400, new_n3527);
and_5  g03151(n11023, n2464, new_n3528);
xnor_4 g03152(new_n3528, new_n3527, new_n3529);
xnor_4 g03153(new_n3529, new_n3526, new_n3530);
nand_5 g03154(n11023, n9400, new_n3531);
and_5  g03155(n11311, n6703, new_n3532);
and_5  g03156(n9400, n3022, new_n3533);
nor_5  g03157(new_n3533, new_n3532, new_n3534);
nand_5 g03158(new_n3533, new_n3532, new_n3535);
nand_5 g03159(n9640, n2464, new_n3536);
and_5  g03160(new_n3536, new_n3535, new_n3537);
or_5   g03161(new_n3537, new_n3534, new_n3538);
nor_5  g03162(new_n3538, new_n3531, new_n3539);
xnor_4 g03163(new_n3538, new_n3531, new_n3540);
xnor_4 g03164(new_n3520, new_n3519, new_n3541);
xnor_4 g03165(new_n3541, new_n3523, new_n3542);
nor_5  g03166(new_n3542, new_n3540, new_n3543);
nor_5  g03167(new_n3543, new_n3539, new_n3544);
xnor_4 g03168(new_n3544, new_n3530, new_n3545);
nand_5 g03169(n10451, n6877, new_n3546);
xnor_4 g03170(new_n3542, new_n3540, new_n3547);
nor_5  g03171(new_n3547, new_n3546, new_n3548);
nand_5 g03172(n11023, n6877, new_n3549);
and_5  g03173(n6703, n2464, new_n3550);
and_5  g03174(n6877, n3022, new_n3551);
nor_5  g03175(new_n3551, new_n3550, new_n3552);
nand_5 g03176(new_n3551, new_n3550, new_n3553);
nand_5 g03177(n9640, n9400, new_n3554);
and_5  g03178(new_n3554, new_n3553, new_n3555);
or_5   g03179(new_n3555, new_n3552, new_n3556);
nor_5  g03180(new_n3556, new_n3549, new_n3557);
xnor_4 g03181(new_n3556, new_n3549, new_n3558);
xnor_4 g03182(new_n3533, new_n3532, new_n3559);
xnor_4 g03183(new_n3559, new_n3536, new_n3560);
nor_5  g03184(new_n3560, new_n3558, new_n3561);
nor_5  g03185(new_n3561, new_n3557, new_n3562);
xnor_4 g03186(new_n3547, new_n3546, new_n3563);
nor_5  g03187(new_n3563, new_n3562, new_n3564);
nor_5  g03188(new_n3564, new_n3548, new_n3565);
or_5   g03189(new_n3565, new_n3545, new_n3566);
nor_5  g03190(new_n3517, new_n3514, new_n3567);
nor_5  g03191(new_n3525, new_n3518, new_n3568);
or_5   g03192(new_n3568, new_n3567, new_n3569);
nand_5 g03193(n10278, n9400, new_n3570);
and_5  g03194(n10451, n2464, new_n3571);
and_5  g03195(n11423, n6877, new_n3572);
xnor_4 g03196(new_n3572, new_n3571, new_n3573);
xor_4  g03197(new_n3573, new_n3570, new_n3574);
xnor_4 g03198(new_n3574, new_n3569, new_n3575);
and_5  g03199(new_n3516, new_n3515, new_n3576);
and_5  g03200(n11311, n11023, new_n3577);
xnor_4 g03201(new_n3577, new_n3576, new_n3578);
nand_5 g03202(n9640, n4203, new_n3579);
and_5  g03203(n4187, n3022, new_n3580);
and_5  g03204(n12753, n6703, new_n3581);
xnor_4 g03205(new_n3581, new_n3580, new_n3582);
xnor_4 g03206(new_n3582, new_n3579, new_n3583);
xor_4  g03207(new_n3583, new_n3578, new_n3584);
xor_4  g03208(new_n3584, new_n3575, new_n3585);
nor_5  g03209(new_n3529, new_n3526, new_n3586);
nand_5 g03210(new_n3528, new_n3527, new_n3587);
or_5   g03211(new_n3544, new_n3530, new_n3588);
xor_4  g03212(new_n3588, new_n3587, new_n3589);
nor_5  g03213(new_n3589, new_n3586, new_n3590);
xnor_4 g03214(new_n3590, new_n3585, new_n3591);
xnor_4 g03215(new_n3591, new_n3566, new_n3592);
nand_5 g03216(n10278, n6877, new_n3593);
xnor_4 g03217(new_n3565, new_n3545, new_n3594);
nor_5  g03218(new_n3594, new_n3593, new_n3595);
xnor_4 g03219(new_n3560, new_n3558, new_n3596);
and_5  g03220(n6877, n6703, new_n3597);
nor_5  g03221(new_n3597, new_n3554, new_n3598);
xor_4  g03222(new_n3551, new_n3550, new_n3599);
or_5   g03223(new_n3599, new_n3598, new_n3600);
or_5   g03224(new_n3600, new_n3554, new_n3601);
or_5   g03225(new_n3601, new_n3596, new_n3602_1);
xnor_4 g03226(new_n3563, new_n3562, new_n3603);
or_5   g03227(new_n3603, new_n3602_1, new_n3604);
xnor_4 g03228(new_n3594, new_n3593, new_n3605);
nor_5  g03229(new_n3605, new_n3604, new_n3606);
nor_5  g03230(new_n3606, new_n3595, new_n3607);
xor_4  g03231(new_n3607, new_n3592, new_n3608);
and_5  g03232(n12826, n4805, new_n3609);
nand_5 g03233(n8665, n137, new_n3610);
and_5  g03234(n6294, n1067, new_n3611);
and_5  g03235(n6797, n5645, new_n3612);
xnor_4 g03236(new_n3612, new_n3611, new_n3613);
xnor_4 g03237(new_n3613, new_n3610, new_n3614);
and_5  g03238(n6294, n5645, new_n3615);
and_5  g03239(n8665, n5283, new_n3616_1);
nor_5  g03240(new_n3616_1, new_n3615, new_n3617);
and_5  g03241(n1067, n137, new_n3618);
xnor_4 g03242(new_n3616_1, new_n3615, new_n3619);
nor_5  g03243(new_n3619, new_n3618, new_n3620);
or_5   g03244(new_n3620, new_n3617, new_n3621);
xnor_4 g03245(new_n3621, new_n3614, new_n3622);
and_5  g03246(n11922, n11478, new_n3623);
and_5  g03247(n5283, n1067, new_n3624);
and_5  g03248(n11478, n8665, new_n3625);
nor_5  g03249(new_n3625, new_n3624, new_n3626);
and_5  g03250(n5645, n137, new_n3627_1);
xnor_4 g03251(new_n3625, new_n3624, new_n3628);
nor_5  g03252(new_n3628, new_n3627_1, new_n3629);
nor_5  g03253(new_n3629, new_n3626, new_n3630);
and_5  g03254(new_n3630, new_n3623, new_n3631);
xor_4  g03255(new_n3619, new_n3618, new_n3632);
xnor_4 g03256(new_n3630, new_n3623, new_n3633);
nor_5  g03257(new_n3633, new_n3632, new_n3634);
nor_5  g03258(new_n3634, new_n3631, new_n3635);
and_5  g03259(n11478, n2551, new_n3636);
and_5  g03260(n11922, n5283, new_n3637);
xnor_4 g03261(new_n3637, new_n3636, new_n3638);
xnor_4 g03262(new_n3638, new_n3635, new_n3639);
xnor_4 g03263(new_n3639, new_n3622, new_n3640);
and_5  g03264(n4805, n2551, new_n3641);
nand_5 g03265(n11922, n4805, new_n3642);
and_5  g03266(n5645, n5283, new_n3643);
and_5  g03267(n8665, n4805, new_n3644);
and_5  g03268(new_n3644, new_n3643, new_n3645);
nor_5  g03269(new_n3644, new_n3643, new_n3646);
nand_5 g03270(n11478, n1067, new_n3647);
nor_5  g03271(new_n3647, new_n3646, new_n3648);
nor_5  g03272(new_n3648, new_n3645, new_n3649);
nor_5  g03273(new_n3649, new_n3642, new_n3650);
xnor_4 g03274(new_n3649, new_n3642, new_n3651);
xor_4  g03275(new_n3628, new_n3627_1, new_n3652);
nor_5  g03276(new_n3652, new_n3651, new_n3653);
or_5   g03277(new_n3653, new_n3650, new_n3654_1);
nor_5  g03278(new_n3654_1, new_n3641, new_n3655);
xor_4  g03279(new_n3633, new_n3632, new_n3656);
xnor_4 g03280(new_n3654_1, new_n3641, new_n3657);
nor_5  g03281(new_n3657, new_n3656, new_n3658);
or_5   g03282(new_n3658, new_n3655, new_n3659);
xor_4  g03283(new_n3659, new_n3640, new_n3660);
and_5  g03284(new_n3660, new_n3609, new_n3661_1);
xnor_4 g03285(new_n3652, new_n3651, new_n3662);
xnor_4 g03286(new_n3644, new_n3643, new_n3663);
and_5  g03287(n4805, n1067, new_n3664);
and_5  g03288(n11478, n5645, new_n3665);
and_5  g03289(new_n3665, new_n3664, new_n3666);
nand_5 g03290(new_n3666, new_n3663, new_n3667);
or_5   g03291(new_n3667, new_n3662, new_n3668);
xor_4  g03292(new_n3657, new_n3656, new_n3669);
or_5   g03293(new_n3669, new_n3668, new_n3670);
xnor_4 g03294(new_n3660, new_n3609, new_n3671);
nor_5  g03295(new_n3671, new_n3670, new_n3672);
nor_5  g03296(new_n3672, new_n3661_1, new_n3673);
or_5   g03297(new_n3659, new_n3640, new_n3674);
and_5  g03298(n12826, n11478, new_n3675);
nand_5 g03299(n5283, n2551, new_n3676);
nand_5 g03300(n4805, n4094, new_n3677_1);
xnor_4 g03301(new_n3677_1, new_n3676, new_n3678);
xnor_4 g03302(new_n3678, new_n3675, new_n3679);
nor_5  g03303(new_n3613, new_n3610, new_n3680);
nor_5  g03304(new_n3621, new_n3614, new_n3681);
or_5   g03305(new_n3681, new_n3680, new_n3682);
xnor_4 g03306(new_n3682, new_n3679, new_n3683);
and_5  g03307(new_n3612, new_n3611, new_n3684);
and_5  g03308(n11922, n137, new_n3685);
xnor_4 g03309(new_n3685, new_n3684, new_n3686);
and_5  g03310(n6797, n1067, new_n3687);
and_5  g03311(n8665, n6294, new_n3688);
and_5  g03312(n5645, n3146, new_n3689);
xnor_4 g03313(new_n3689, new_n3688, new_n3690);
xor_4  g03314(new_n3690, new_n3687, new_n3691);
xor_4  g03315(new_n3691, new_n3686, new_n3692);
xor_4  g03316(new_n3692, new_n3683, new_n3693);
nor_5  g03317(new_n3638, new_n3635, new_n3694);
nand_5 g03318(new_n3637, new_n3636, new_n3695);
or_5   g03319(new_n3639, new_n3622, new_n3696);
xor_4  g03320(new_n3696, new_n3695, new_n3697);
nor_5  g03321(new_n3697, new_n3694, new_n3698);
xnor_4 g03322(new_n3698, new_n3693, new_n3699);
xnor_4 g03323(new_n3699, new_n3674, new_n3700);
xor_4  g03324(new_n3700, new_n3673, new_n3701);
and_5  g03325(n3992, n2749, new_n3702);
and_5  g03326(n11876, n6358, new_n3703);
and_5  g03327(n3992, n3754, new_n3704);
nor_5  g03328(new_n3704, new_n3703, new_n3705);
and_5  g03329(n10898, n8384, new_n3706);
xnor_4 g03330(new_n3704, new_n3703, new_n3707);
nor_5  g03331(new_n3707, new_n3706, new_n3708);
nor_5  g03332(new_n3708, new_n3705, new_n3709);
and_5  g03333(new_n3709, new_n3702, new_n3710);
xnor_4 g03334(new_n3709, new_n3702, new_n3711);
and_5  g03335(n10898, n6358, new_n3712);
and_5  g03336(n11876, n5198, new_n3713);
and_5  g03337(n8384, n3754, new_n3714);
xnor_4 g03338(new_n3714, new_n3713, new_n3715);
xor_4  g03339(new_n3715, new_n3712, new_n3716);
nor_5  g03340(new_n3716, new_n3711, new_n3717);
nor_5  g03341(new_n3717, new_n3710, new_n3718);
and_5  g03342(n8384, n2749, new_n3719_1);
and_5  g03343(n3992, n159, new_n3720);
xnor_4 g03344(new_n3720, new_n3719_1, new_n3721);
xnor_4 g03345(new_n3721, new_n3718, new_n3722);
and_5  g03346(n6358, n3754, new_n3723);
and_5  g03347(n10898, n5198, new_n3724);
and_5  g03348(n11876, n1471, new_n3725);
xor_4  g03349(new_n3725, new_n3724, new_n3726);
xnor_4 g03350(new_n3726, new_n3723, new_n3727);
nor_5  g03351(new_n3714, new_n3713, new_n3728);
nor_5  g03352(new_n3715, new_n3712, new_n3729);
nor_5  g03353(new_n3729, new_n3728, new_n3730);
xor_4  g03354(new_n3730, new_n3727, new_n3731);
xnor_4 g03355(new_n3731, new_n3722, new_n3732);
nand_5 g03356(n7236, n159, new_n3733);
and_5  g03357(n7236, n2749, new_n3734);
and_5  g03358(n11876, n8384, new_n3735);
and_5  g03359(n7236, n3754, new_n3736);
nor_5  g03360(new_n3736, new_n3735, new_n3737);
and_5  g03361(n11876, n7236, new_n3738);
and_5  g03362(new_n3738, new_n3714, new_n3739);
and_5  g03363(n10898, n3992, new_n3740);
nor_5  g03364(new_n3740, new_n3739, new_n3741);
nor_5  g03365(new_n3741, new_n3737, new_n3742);
and_5  g03366(new_n3742, new_n3734, new_n3743);
xnor_4 g03367(new_n3742, new_n3734, new_n3744);
xor_4  g03368(new_n3707, new_n3706, new_n3745);
nor_5  g03369(new_n3745, new_n3744, new_n3746);
nor_5  g03370(new_n3746, new_n3743, new_n3747);
and_5  g03371(new_n3747, new_n3733, new_n3748);
xor_4  g03372(new_n3716, new_n3711, new_n3749);
xnor_4 g03373(new_n3747, new_n3733, new_n3750);
nor_5  g03374(new_n3750, new_n3749, new_n3751);
or_5   g03375(new_n3751, new_n3748, new_n3752);
or_5   g03376(new_n3752, new_n3732, new_n3753);
and_5  g03377(new_n3725, new_n3724, new_n3754_1);
and_5  g03378(n6358, n2749, new_n3755);
xnor_4 g03379(new_n3755, new_n3754_1, new_n3756);
and_5  g03380(n10898, n1471, new_n3757);
and_5  g03381(n5198, n3754, new_n3758);
and_5  g03382(n11876, n7646, new_n3759);
xnor_4 g03383(new_n3759, new_n3758, new_n3760);
xor_4  g03384(new_n3760, new_n3757, new_n3761);
xor_4  g03385(new_n3761, new_n3756, new_n3762);
nor_5  g03386(new_n3726, new_n3723, new_n3763);
nor_5  g03387(new_n3730, new_n3727, new_n3764);
nor_5  g03388(new_n3764, new_n3763, new_n3765);
and_5  g03389(n3992, n1510, new_n3766);
and_5  g03390(n8384, n159, new_n3767);
and_5  g03391(n12247, n7236, new_n3768);
xnor_4 g03392(new_n3768, new_n3767, new_n3769);
xnor_4 g03393(new_n3769, new_n3766, new_n3770);
xnor_4 g03394(new_n3770, new_n3765, new_n3771);
xor_4  g03395(new_n3771, new_n3762, new_n3772);
nor_5  g03396(new_n3721, new_n3718, new_n3773);
nand_5 g03397(new_n3720, new_n3719_1, new_n3774);
or_5   g03398(new_n3731, new_n3722, new_n3775);
xor_4  g03399(new_n3775, new_n3774, new_n3776);
nor_5  g03400(new_n3776, new_n3773, new_n3777);
xnor_4 g03401(new_n3777, new_n3772, new_n3778);
xnor_4 g03402(new_n3778, new_n3753, new_n3779);
and_5  g03403(n7236, n1510, new_n3780);
xor_4  g03404(new_n3752, new_n3732, new_n3781);
and_5  g03405(new_n3781, new_n3780, new_n3782);
xnor_4 g03406(new_n3745, new_n3744, new_n3783);
nor_5  g03407(new_n3739, new_n3737, new_n3784);
and_5  g03408(n11876, n3992, new_n3785);
and_5  g03409(n10898, n7236, new_n3786);
nand_5 g03410(new_n3786, new_n3785, new_n3787);
or_5   g03411(new_n3787, new_n3784, new_n3788);
or_5   g03412(new_n3788, new_n3783, new_n3789);
xor_4  g03413(new_n3750, new_n3749, new_n3790);
or_5   g03414(new_n3790, new_n3789, new_n3791);
xnor_4 g03415(new_n3781, new_n3780, new_n3792);
nor_5  g03416(new_n3792, new_n3791, new_n3793);
nor_5  g03417(new_n3793, new_n3782, new_n3794);
xor_4  g03418(new_n3794, new_n3779, new_n3795);
xnor_4 g03419(new_n3795, new_n3701, new_n3796);
xor_4  g03420(new_n3671, new_n3670, new_n3797);
xor_4  g03421(new_n3792, new_n3791, new_n3798);
nor_5  g03422(new_n3798, new_n3797, new_n3799);
xnor_4 g03423(new_n3798, new_n3797, new_n3800);
xor_4  g03424(new_n3790, new_n3789, new_n3801);
xor_4  g03425(new_n3667, new_n3662, new_n3802);
xor_4  g03426(new_n3788, new_n3783, new_n3803);
nor_5  g03427(new_n3803, new_n3802, new_n3804);
xnor_4 g03428(new_n3786, new_n3785, new_n3805);
xnor_4 g03429(new_n3665, new_n3664, new_n3806);
and_5  g03430(new_n3806, new_n3805, new_n3807);
and_5  g03431(n5645, n4805, new_n3808);
and_5  g03432(new_n3808, new_n3738, new_n3809);
xnor_4 g03433(new_n3806, new_n3805, new_n3810);
nor_5  g03434(new_n3810, new_n3809, new_n3811);
nor_5  g03435(new_n3811, new_n3807, new_n3812);
nor_5  g03436(new_n3808, new_n3647, new_n3813);
and_5  g03437(new_n3813, new_n3646, new_n3814);
nor_5  g03438(new_n3813, new_n3663, new_n3815);
or_5   g03439(new_n3815, new_n3814, new_n3816);
nor_5  g03440(new_n3816, new_n3812, new_n3817);
xnor_4 g03441(new_n3816, new_n3812, new_n3818);
nand_5 g03442(n10898, n3992, new_n3819);
nor_5  g03443(new_n3819, new_n3738, new_n3820);
nor_5  g03444(new_n3820, new_n3784, new_n3821);
or_5   g03445(new_n3819, new_n3738, new_n3822);
nor_5  g03446(new_n3822, new_n3737, new_n3823);
nor_5  g03447(new_n3823, new_n3821, new_n3824);
nor_5  g03448(new_n3824, new_n3818, new_n3825);
nor_5  g03449(new_n3825, new_n3817, new_n3826);
xnor_4 g03450(new_n3803, new_n3802, new_n3827);
nor_5  g03451(new_n3827, new_n3826, new_n3828);
nor_5  g03452(new_n3828, new_n3804, new_n3829);
nor_5  g03453(new_n3829, new_n3801, new_n3830);
xor_4  g03454(new_n3669, new_n3668, new_n3831);
xnor_4 g03455(new_n3829, new_n3801, new_n3832);
nor_5  g03456(new_n3832, new_n3831, new_n3833);
nor_5  g03457(new_n3833, new_n3830, new_n3834);
nor_5  g03458(new_n3834, new_n3800, new_n3835);
nor_5  g03459(new_n3835, new_n3799, new_n3836);
xnor_4 g03460(new_n3836, new_n3796, new_n3837);
xnor_4 g03461(new_n3837, new_n3608, new_n3838);
xor_4  g03462(new_n3605, new_n3604, new_n3839);
xnor_4 g03463(new_n3834, new_n3800, new_n3840);
nor_5  g03464(new_n3840, new_n3839, new_n3841);
xor_4  g03465(new_n3603, new_n3602_1, new_n3842_1);
xnor_4 g03466(new_n3601, new_n3596, new_n3843);
xor_4  g03467(new_n3827, new_n3826, new_n3844);
nor_5  g03468(new_n3844, new_n3843, new_n3845);
xnor_4 g03469(new_n3844, new_n3843, new_n3846);
xor_4  g03470(new_n3824, new_n3818, new_n3847);
or_5   g03471(new_n3597, new_n3554, new_n3848);
or_5   g03472(new_n3848, new_n3552, new_n3849_1);
nand_5 g03473(new_n3849_1, new_n3600, new_n3850);
nor_5  g03474(new_n3850, new_n3847, new_n3851);
xnor_4 g03475(new_n3850, new_n3847, new_n3852);
xor_4  g03476(new_n3810, new_n3809, new_n3853);
and_5  g03477(n9400, n6703, new_n3854);
and_5  g03478(n9640, n6877, new_n3855);
xnor_4 g03479(new_n3855, new_n3854, new_n3856);
nor_5  g03480(new_n3856, new_n3853, new_n3857);
nand_5 g03481(n6877, n6703, new_n3858);
xnor_4 g03482(new_n3808, new_n3738, new_n3859);
or_5   g03483(new_n3859, new_n3858, new_n3860);
xnor_4 g03484(new_n3810, new_n3809, new_n3861);
xor_4  g03485(new_n3856, new_n3861, new_n3862);
nor_5  g03486(new_n3862, new_n3860, new_n3863);
nor_5  g03487(new_n3863, new_n3857, new_n3864);
nor_5  g03488(new_n3864, new_n3852, new_n3865_1);
nor_5  g03489(new_n3865_1, new_n3851, new_n3866);
nor_5  g03490(new_n3866, new_n3846, new_n3867);
or_5   g03491(new_n3867, new_n3845, new_n3868);
nor_5  g03492(new_n3868, new_n3842_1, new_n3869);
xnor_4 g03493(new_n3832, new_n3831, new_n3870);
nor_5  g03494(new_n3867, new_n3845, new_n3871);
xor_4  g03495(new_n3871, new_n3842_1, new_n3872);
nor_5  g03496(new_n3872, new_n3870, new_n3873);
nor_5  g03497(new_n3873, new_n3869, new_n3874);
xnor_4 g03498(new_n3840, new_n3839, new_n3875);
nor_5  g03499(new_n3875, new_n3874, new_n3876);
nor_5  g03500(new_n3876, new_n3841, new_n3877);
xor_4  g03501(new_n3877, new_n3838, new_n3878);
nor_5  g03502(new_n3878, new_n3513, new_n3879);
xnor_4 g03503(new_n3878, new_n3513, new_n3880);
xnor_4 g03504(new_n3510, new_n3509, new_n3881);
xor_4  g03505(new_n3875, new_n3874, new_n3882);
nor_5  g03506(new_n3882, new_n3881, new_n3883);
xnor_4 g03507(new_n3508, new_n3507, new_n3884);
xor_4  g03508(new_n3872, new_n3870, new_n3885);
and_5  g03509(new_n3885, new_n3884, new_n3886);
xnor_4 g03510(new_n3885, new_n3884, new_n3887);
xor_4  g03511(new_n3506, new_n3501, new_n3888);
xor_4  g03512(new_n3866, new_n3846, new_n3889);
nor_5  g03513(new_n3889, new_n3888, new_n3890);
xor_4  g03514(new_n3864, new_n3852, new_n3891);
and_5  g03515(n7862, n1798, new_n3892);
nor_5  g03516(new_n3892, new_n3460, new_n3893);
nor_5  g03517(new_n3893, new_n3502, new_n3894);
or_5   g03518(new_n3892, new_n3460, new_n3895);
nor_5  g03519(new_n3895, new_n3459, new_n3896);
nor_5  g03520(new_n3896, new_n3894, new_n3897);
nor_5  g03521(new_n3897, new_n3891, new_n3898);
xnor_4 g03522(new_n3897, new_n3891, new_n3899);
xnor_4 g03523(new_n3859, new_n3597, new_n3900);
and_5  g03524(new_n3900, new_n3892, new_n3901);
xor_4  g03525(new_n3504, new_n3503, new_n3902);
nor_5  g03526(new_n3902, new_n3901, new_n3903);
xnor_4 g03527(new_n3862, new_n3860, new_n3904);
xor_4  g03528(new_n3902, new_n3901, new_n3905);
and_5  g03529(new_n3905, new_n3904, new_n3906);
nor_5  g03530(new_n3906, new_n3903, new_n3907);
nor_5  g03531(new_n3907, new_n3899, new_n3908);
nor_5  g03532(new_n3908, new_n3898, new_n3909);
xnor_4 g03533(new_n3889, new_n3888, new_n3910);
nor_5  g03534(new_n3910, new_n3909, new_n3911);
nor_5  g03535(new_n3911, new_n3890, new_n3912);
nor_5  g03536(new_n3912, new_n3887, new_n3913);
or_5   g03537(new_n3913, new_n3886, new_n3914);
xnor_4 g03538(new_n3882, new_n3881, new_n3915);
nor_5  g03539(new_n3915, new_n3914, new_n3916);
nor_5  g03540(new_n3916, new_n3883, new_n3917);
nor_5  g03541(new_n3917, new_n3880, new_n3918);
nor_5  g03542(new_n3918, new_n3879, new_n3919);
nor_5  g03543(new_n3591, new_n3566, new_n3920);
nor_5  g03544(new_n3607, new_n3592, new_n3921);
nor_5  g03545(new_n3921, new_n3920, new_n3922);
nand_5 g03546(n7862, n753, new_n3923);
nor_5  g03547(new_n3682, new_n3679, new_n3924);
nor_5  g03548(new_n3692, new_n3683, new_n3925);
nor_5  g03549(new_n3925, new_n3924, new_n3926);
xnor_4 g03550(new_n3926, new_n3923, new_n3927);
and_5  g03551(new_n3685, new_n3684, new_n3928);
nor_5  g03552(new_n3691, new_n3686, new_n3929);
nor_5  g03553(new_n3929, new_n3928, new_n3930);
and_5  g03554(n3146, n1067, new_n3931);
and_5  g03555(n2551, n137, new_n3932_1);
xnor_4 g03556(new_n3932_1, new_n3931, new_n3933);
and_5  g03557(n12826, n5283, new_n3934);
and_5  g03558(n8665, n6797, new_n3935);
xnor_4 g03559(new_n3935, new_n3934, new_n3936);
xnor_4 g03560(new_n3936, new_n3933, new_n3937);
xnor_4 g03561(new_n3937, new_n3930, new_n3938);
and_5  g03562(new_n3755, new_n3754_1, new_n3939);
nor_5  g03563(new_n3761, new_n3756, new_n3940);
nor_5  g03564(new_n3940, new_n3939, new_n3941);
nor_5  g03565(new_n3768, new_n3767, new_n3942);
nor_5  g03566(new_n3769, new_n3766, new_n3943);
nor_5  g03567(new_n3943, new_n3942, new_n3944);
and_5  g03568(n8384, n1510, new_n3945);
and_5  g03569(n5198, n2749, new_n3946);
xor_4  g03570(new_n3946, new_n3945, new_n3947);
xnor_4 g03571(new_n3947, new_n3944, new_n3948);
xnor_4 g03572(new_n3948, new_n3941, new_n3949);
xnor_4 g03573(new_n3949, new_n3938, new_n3950);
xnor_4 g03574(new_n3950, new_n3927, new_n3951);
xnor_4 g03575(new_n3951, new_n3922, new_n3952);
nor_5  g03576(new_n3493, new_n3492, new_n3953);
nor_5  g03577(new_n3495, new_n3490, new_n3954);
nor_5  g03578(new_n3954, new_n3953, new_n3955);
nor_5  g03579(new_n3696, new_n3695, new_n3956);
nor_5  g03580(new_n3698, new_n3693, new_n3957);
nor_5  g03581(new_n3957, new_n3956, new_n3958);
xnor_4 g03582(new_n3958, new_n3955, new_n3959);
and_5  g03583(n12511, n7236, new_n3960);
and_5  g03584(n6826, n1798, new_n3961);
xnor_4 g03585(new_n3961, new_n3960, new_n3962);
nor_5  g03586(new_n3689, new_n3688, new_n3963);
nor_5  g03587(new_n3690, new_n3687, new_n3964);
nor_5  g03588(new_n3964, new_n3963, new_n3965);
nor_5  g03589(new_n3759, new_n3758, new_n3966);
nor_5  g03590(new_n3760, new_n3757, new_n3967);
nor_5  g03591(new_n3967, new_n3966, new_n3968);
xnor_4 g03592(new_n3968, new_n3965, new_n3969);
xnor_4 g03593(new_n3969, new_n3962, new_n3970);
nand_5 g03594(n6358, n159, new_n3971);
nor_5  g03595(new_n3678, new_n3675, new_n3972);
or_5   g03596(new_n3972, new_n3676, new_n3973);
nand_5 g03597(n11478, n4094, new_n3974);
nor_5  g03598(new_n3974, new_n3973, new_n3975);
or_5   g03599(new_n3974, new_n3609, new_n3976);
and_5  g03600(new_n3976, new_n3973, new_n3977);
nor_5  g03601(new_n3977, new_n3975, new_n3978);
xnor_4 g03602(new_n3978, new_n3971, new_n3979);
xnor_4 g03603(new_n3979, new_n3970, new_n3980);
xnor_4 g03604(new_n3980, new_n3959, new_n3981);
xnor_4 g03605(new_n3981, new_n3952, new_n3982);
nor_5  g03606(new_n3775, new_n3774, new_n3983);
nor_5  g03607(new_n3777, new_n3772, new_n3984);
nor_5  g03608(new_n3984, new_n3983, new_n3985);
and_5  g03609(n5645, n4938, new_n3986_1);
and_5  g03610(n10898, n7646, new_n3987);
xor_4  g03611(new_n3987, new_n3986_1, new_n3988);
xnor_4 g03612(new_n3988, new_n3985, new_n3989);
xnor_4 g03613(new_n3989, new_n3982, new_n3990);
nor_5  g03614(new_n3795, new_n3701, new_n3991);
nor_5  g03615(new_n3836, new_n3796, new_n3992_1);
nor_5  g03616(new_n3992_1, new_n3991, new_n3993);
nand_5 g03617(n11922, n6294, new_n3994);
nor_5  g03618(new_n3699, new_n3674, new_n3995);
nor_5  g03619(new_n3700, new_n3673, new_n3996);
nor_5  g03620(new_n3996, new_n3995, new_n3997);
xnor_4 g03621(new_n3997, new_n3994, new_n3998);
nor_5  g03622(new_n3496, new_n3471, new_n3999);
nor_5  g03623(new_n3512, new_n3497, new_n4000);
nor_5  g03624(new_n4000, new_n3999, new_n4001);
nor_5  g03625(new_n3588, new_n3587, new_n4002);
nor_5  g03626(new_n3590, new_n3585, new_n4003);
nor_5  g03627(new_n4003, new_n4002, new_n4004);
nor_5  g03628(new_n3574, new_n3569, new_n4005_1);
nor_5  g03629(new_n3584, new_n3575, new_n4006);
nor_5  g03630(new_n4006, new_n4005_1, new_n4007);
and_5  g03631(new_n3581, new_n3580, new_n4008);
nor_5  g03632(new_n3581, new_n3580, new_n4009);
nor_5  g03633(new_n4009, new_n3579, new_n4010);
nor_5  g03634(new_n4010, new_n4008, new_n4011);
and_5  g03635(n4203, n3022, new_n4012);
and_5  g03636(n11023, n4187, new_n4013);
xnor_4 g03637(new_n4013, new_n4012, new_n4014);
xnor_4 g03638(new_n4014, new_n4011, new_n4015);
and_5  g03639(n7456, n5240, new_n4016);
and_5  g03640(n12753, n9640, new_n4017);
xnor_4 g03641(new_n4017, new_n4016, new_n4018);
and_5  g03642(n9583, n1333, new_n4019);
and_5  g03643(n12591, n11821, new_n4020);
xnor_4 g03644(new_n4020, new_n4019, new_n4021);
xor_4  g03645(new_n4021, new_n4018, new_n4022);
xnor_4 g03646(new_n4022, new_n4015, new_n4023);
xnor_4 g03647(new_n4023, new_n4007, new_n4024);
nor_5  g03648(new_n3479, new_n3474, new_n4025);
nor_5  g03649(new_n3489, new_n3480, new_n4026);
nor_5  g03650(new_n4026, new_n4025, new_n4027);
and_5  g03651(n9080, n3932, new_n4028);
and_5  g03652(n10174, n6703, new_n4029);
and_5  g03653(n6877, n2278, new_n4030);
xnor_4 g03654(new_n4030, new_n4029, new_n4031);
xnor_4 g03655(new_n4031, new_n4028, new_n4032);
xnor_4 g03656(new_n4032, new_n4027, new_n4033);
xnor_4 g03657(new_n4033, new_n4024, new_n4034);
xnor_4 g03658(new_n4034, new_n4004, new_n4035);
xnor_4 g03659(new_n4035, new_n4001, new_n4036);
xnor_4 g03660(new_n4036, new_n3998, new_n4037);
xnor_4 g03661(new_n4037, new_n3993, new_n4038);
xnor_4 g03662(new_n4038, new_n3990, new_n4039);
xnor_4 g03663(new_n4039, new_n3919, new_n4040);
nor_5  g03664(new_n3770, new_n3765, new_n4041);
nor_5  g03665(new_n3771, new_n3762, new_n4042);
nor_5  g03666(new_n4042, new_n4041, new_n4043);
and_5  g03667(new_n3482, new_n3481, new_n4044);
nor_5  g03668(new_n3488, new_n3483, new_n4045);
nor_5  g03669(new_n4045, new_n4044, new_n4046);
and_5  g03670(new_n3572, new_n3571, new_n4047);
nor_5  g03671(new_n3572, new_n3571, new_n4048);
nor_5  g03672(new_n4048, new_n3570, new_n4049);
or_5   g03673(new_n4049, new_n4047, new_n4050);
xnor_4 g03674(new_n4050, new_n4046, new_n4051);
nor_5  g03675(new_n3477, new_n3476, new_n4052);
nor_5  g03676(new_n3478, new_n3475, new_n4053);
nor_5  g03677(new_n4053, new_n4052, new_n4054);
and_5  g03678(new_n3486, new_n3485, new_n4055);
nor_5  g03679(new_n3486, new_n3485, new_n4056);
nor_5  g03680(new_n4056, new_n3484, new_n4057);
nor_5  g03681(new_n4057, new_n4055, new_n4058);
and_5  g03682(n10278, n2464, new_n4059);
and_5  g03683(n11757, n11662, new_n4060);
xnor_4 g03684(new_n4060, new_n4059, new_n4061);
and_5  g03685(n10327, n3172, new_n4062);
and_5  g03686(n11423, n9400, new_n4063);
xnor_4 g03687(new_n4063, new_n4062, new_n4064);
xor_4  g03688(new_n4064, new_n4061, new_n4065);
xnor_4 g03689(new_n4065, new_n4058, new_n4066);
xnor_4 g03690(new_n4066, new_n4054, new_n4067);
xnor_4 g03691(new_n4067, new_n4051, new_n4068);
xnor_4 g03692(new_n4068, new_n4043, new_n4069);
and_5  g03693(n3754, n1471, new_n4070);
and_5  g03694(n11311, n10451, new_n4071);
xnor_4 g03695(new_n4071, new_n4070, new_n4072);
and_5  g03696(new_n3577, new_n3576, new_n4073);
nor_5  g03697(new_n3583, new_n3578, new_n4074);
nor_5  g03698(new_n4074, new_n4073, new_n4075);
and_5  g03699(n11876, n4722, new_n4076);
and_5  g03700(n10685, n4805, new_n4077);
and_5  g03701(n12247, n3992, new_n4078);
xnor_4 g03702(new_n4078, new_n4077, new_n4079);
xnor_4 g03703(new_n4079, new_n4076, new_n4080);
xnor_4 g03704(new_n4080, new_n4075, new_n4081);
xnor_4 g03705(new_n4081, new_n4072, new_n4082);
xnor_4 g03706(new_n4082, new_n4069, new_n4083);
nor_5  g03707(new_n3778, new_n3753, new_n4084);
nor_5  g03708(new_n3794, new_n3779, new_n4085);
or_5   g03709(new_n4085, new_n4084, new_n4086_1);
nor_5  g03710(new_n3837, new_n3608, new_n4087);
nor_5  g03711(new_n3877, new_n3838, new_n4088_1);
nor_5  g03712(new_n4088_1, new_n4087, new_n4089);
xnor_4 g03713(new_n4089, new_n4086_1, new_n4090);
xnor_4 g03714(new_n4090, new_n4083, new_n4091);
xnor_4 g03715(new_n4091, new_n4040, n1269);
and_5  g03716(n10223, n4312, new_n4093);
nand_5 g03717(n12705, n7265, new_n4094_1);
and_5  g03718(n4312, n2879, new_n4095);
xor_4  g03719(new_n4094_1, new_n888, new_n4096);
nor_5  g03720(new_n4096, new_n4095, new_n4097);
nor_5  g03721(new_n4097, new_n4094_1, new_n4098);
nor_5  g03722(new_n4098, new_n4093, new_n4099);
or_5   g03723(new_n4098, new_n894, new_n4100);
and_5  g03724(new_n4100, new_n4093, new_n4101);
or_5   g03725(new_n4101, new_n4099, new_n4102);
and_5  g03726(n12025, n7265, new_n4103);
and_5  g03727(n12705, n2879, new_n4104);
xnor_4 g03728(new_n4104, new_n4103, new_n4105);
xnor_4 g03729(new_n4105, new_n4102, new_n4106);
and_5  g03730(n9195, n5964, new_n4107);
and_5  g03731(n4634, n1097, new_n4108);
xnor_4 g03732(new_n4108, new_n4107, new_n4109);
xnor_4 g03733(new_n4109, new_n4106, new_n4110);
nand_5 g03734(n5964, n4634, new_n4111);
nor_5  g03735(new_n896, new_n895, new_n4112);
and_5  g03736(new_n896, new_n895, new_n4113);
nor_5  g03737(new_n4113, new_n894, new_n4114);
or_5   g03738(new_n4114, new_n4112, new_n4115);
nor_5  g03739(new_n4115, new_n4111, new_n4116);
xor_4  g03740(new_n4096, new_n4095, new_n4117);
xnor_4 g03741(new_n4115, new_n4111, new_n4118);
nor_5  g03742(new_n4118, new_n4117, new_n4119);
nor_5  g03743(new_n4119, new_n4116, new_n4120);
xnor_4 g03744(new_n4120, new_n4110, new_n4121);
and_5  g03745(n9195, n5305, new_n4122);
nor_5  g03746(new_n892, new_n883, new_n4123);
nor_5  g03747(new_n898, new_n893, new_n4124);
or_5   g03748(new_n4124, new_n4123, new_n4125);
nor_5  g03749(new_n4125, new_n4122, new_n4126);
xor_4  g03750(new_n4118, new_n4117, new_n4127);
xnor_4 g03751(new_n4125, new_n4122, new_n4128);
nor_5  g03752(new_n4128, new_n4127, new_n4129);
or_5   g03753(new_n4129, new_n4126, new_n4130);
or_5   g03754(new_n4130, new_n4121, new_n4131);
nor_5  g03755(new_n4105, new_n4102, new_n4132);
or_5   g03756(new_n4132, new_n4101, new_n4133);
and_5  g03757(n5964, n2253, new_n4134);
and_5  g03758(n9195, n1097, new_n4135);
and_5  g03759(n5305, n3865, new_n4136);
xnor_4 g03760(new_n4136, new_n4135, new_n4137);
xnor_4 g03761(new_n4137, new_n4134, new_n4138);
xnor_4 g03762(new_n4138, new_n4133, new_n4139);
and_5  g03763(new_n4104, new_n4103, new_n4140);
and_5  g03764(n4634, n4312, new_n4141_1);
xnor_4 g03765(new_n4141_1, new_n4140, new_n4142);
and_5  g03766(n12025, n2879, new_n4143);
and_5  g03767(n11257, n7265, new_n4144);
and_5  g03768(n12705, n10223, new_n4145);
xnor_4 g03769(new_n4145, new_n4144, new_n4146);
xor_4  g03770(new_n4146, new_n4143, new_n4147);
xor_4  g03771(new_n4147, new_n4142, new_n4148);
xor_4  g03772(new_n4148, new_n4139, new_n4149);
nor_5  g03773(new_n4109, new_n4106, new_n4150);
nand_5 g03774(new_n4108, new_n4107, new_n4151);
or_5   g03775(new_n4120, new_n4110, new_n4152);
xor_4  g03776(new_n4152, new_n4151, new_n4153);
nor_5  g03777(new_n4153, new_n4150, new_n4154);
xnor_4 g03778(new_n4154, new_n4149, new_n4155_1);
xnor_4 g03779(new_n4155_1, new_n4131, new_n4156);
nand_5 g03780(n5305, n2253, new_n4157);
xnor_4 g03781(new_n4130, new_n4121, new_n4158);
nor_5  g03782(new_n4158, new_n4157, new_n4159_1);
or_5   g03783(new_n904, new_n899, new_n4160);
xor_4  g03784(new_n4128, new_n4127, new_n4161);
or_5   g03785(new_n4161, new_n4160, new_n4162);
xnor_4 g03786(new_n4158, new_n4157, new_n4163);
nor_5  g03787(new_n4163, new_n4162, new_n4164);
nor_5  g03788(new_n4164, new_n4159_1, new_n4165);
xor_4  g03789(new_n4165, new_n4156, new_n4166);
xor_4  g03790(new_n4163, new_n4162, new_n4167);
or_5   g03791(new_n996_1, new_n995, new_n4168);
nand_5 g03792(n12145, n8759, new_n4169);
nor_5  g03793(new_n988, new_n985, new_n4170);
nor_5  g03794(new_n994, new_n989, new_n4171);
nor_5  g03795(new_n4171, new_n4170, new_n4172);
xnor_4 g03796(new_n4172, new_n4169, new_n4173);
nand_5 g03797(n6776, n2522, new_n4174);
nor_5  g03798(new_n992_1, new_n991, new_n4175);
and_5  g03799(new_n992_1, new_n991, new_n4176);
nor_5  g03800(new_n4176, new_n990, new_n4177);
or_5   g03801(new_n4177, new_n4175, new_n4178);
xnor_4 g03802(new_n4178, new_n4174, new_n4179);
and_5  g03803(n7436, n2024, new_n4180);
nand_5 g03804(n12299, n9189, new_n4181);
nand_5 g03805(n8276, n7946, new_n4182);
xnor_4 g03806(new_n4182, new_n4181, new_n4183);
xor_4  g03807(new_n4183, new_n4180, new_n4184);
xnor_4 g03808(new_n4184, new_n4179, new_n4185);
xnor_4 g03809(new_n4185, new_n4173, new_n4186);
or_5   g03810(new_n4186, new_n4168, new_n4187_1);
nand_5 g03811(n12221, n8759, new_n4188);
nor_5  g03812(new_n4178, new_n4174, new_n4189_1);
nor_5  g03813(new_n4184, new_n4179, new_n4190_1);
nor_5  g03814(new_n4190_1, new_n4189_1, new_n4191);
and_5  g03815(n12145, n6776, new_n4192);
and_5  g03816(n12299, n2522, new_n4193);
xnor_4 g03817(new_n4193, new_n4192, new_n4194);
xnor_4 g03818(new_n4194, new_n4191, new_n4195);
and_5  g03819(n9189, n7436, new_n4196);
nor_5  g03820(new_n4183, new_n4180, new_n4197);
nor_5  g03821(new_n4197, new_n4182, new_n4198);
nor_5  g03822(new_n4198, new_n4196, new_n4199);
or_5   g03823(new_n4198, new_n990, new_n4200);
and_5  g03824(new_n4200, new_n4196, new_n4201);
or_5   g03825(new_n4201, new_n4199, new_n4202);
and_5  g03826(n8276, n2024, new_n4203_1);
and_5  g03827(n9241, n7946, new_n4204);
xnor_4 g03828(new_n4204, new_n4203_1, new_n4205);
xnor_4 g03829(new_n4205, new_n4202, new_n4206);
xnor_4 g03830(new_n4206, new_n4195, new_n4207);
nor_5  g03831(new_n4172, new_n4169, new_n4208);
nor_5  g03832(new_n4185, new_n4173, new_n4209);
nor_5  g03833(new_n4209, new_n4208, new_n4210);
xnor_4 g03834(new_n4210, new_n4207, new_n4211);
xnor_4 g03835(new_n4211, new_n4188, new_n4212);
xnor_4 g03836(new_n4212, new_n4187_1, new_n4213);
xnor_4 g03837(new_n4186, new_n4168, new_n4214);
or_5   g03838(new_n1014, new_n1012, new_n4215);
nand_5 g03839(n6016, n5331, new_n4216);
and_5  g03840(n8476, n521, new_n4217);
nor_5  g03841(new_n1009, new_n1008, new_n4218);
nor_5  g03842(new_n1010, new_n1007, new_n4219);
nor_5  g03843(new_n4219, new_n4218, new_n4220);
xnor_4 g03844(new_n4220, new_n4217, new_n4221);
and_5  g03845(n12648, n2498, new_n4222);
and_5  g03846(n10545, n2558, new_n4223);
xnor_4 g03847(new_n4223, new_n963, new_n4224);
xor_4  g03848(new_n4224, new_n4222, new_n4225);
xnor_4 g03849(new_n4225, new_n4221, new_n4226_1);
xnor_4 g03850(new_n4226_1, new_n4216, new_n4227);
nor_5  g03851(new_n1005, new_n1002, new_n4228);
nor_5  g03852(new_n1011, new_n1006, new_n4229);
nor_5  g03853(new_n4229, new_n4228, new_n4230_1);
xnor_4 g03854(new_n4230_1, new_n4227, new_n4231);
xor_4  g03855(new_n4231, new_n4215, new_n4232);
or_5   g03856(new_n1026, new_n1025, new_n4233);
nand_5 g03857(n7965, n7270, new_n4234);
and_5  g03858(n7388, n806, new_n4235);
nor_5  g03859(new_n1022, new_n1021, new_n4236);
nor_5  g03860(new_n1023, new_n1020_1, new_n4237);
nor_5  g03861(new_n4237, new_n4236, new_n4238);
xnor_4 g03862(new_n4238, new_n4235, new_n4239);
and_5  g03863(n9111, n2393, new_n4240);
and_5  g03864(n9763, n5860, new_n4241);
xnor_4 g03865(new_n4241, new_n946, new_n4242);
xor_4  g03866(new_n4242, new_n4240, new_n4243);
xnor_4 g03867(new_n4243, new_n4239, new_n4244);
xnor_4 g03868(new_n4244, new_n4234, new_n4245);
nor_5  g03869(new_n1018, new_n1016, new_n4246);
nor_5  g03870(new_n1024, new_n1019, new_n4247);
nor_5  g03871(new_n4247, new_n4246, new_n4248);
xnor_4 g03872(new_n4248, new_n4245, new_n4249);
xor_4  g03873(new_n4249, new_n4233, new_n4250);
xnor_4 g03874(new_n4250, new_n4232, new_n4251);
nor_5  g03875(new_n1027, new_n1015, new_n4252);
nor_5  g03876(new_n1031, new_n1028, new_n4253);
nor_5  g03877(new_n4253, new_n4252, new_n4254);
xor_4  g03878(new_n4254, new_n4251, new_n4255);
nor_5  g03879(new_n4255, new_n4214, new_n4256);
nor_5  g03880(new_n1000, new_n997, new_n4257);
nor_5  g03881(new_n1032, new_n1001, new_n4258);
nor_5  g03882(new_n4258, new_n4257, new_n4259);
xnor_4 g03883(new_n4255, new_n4214, new_n4260);
nor_5  g03884(new_n4260, new_n4259, new_n4261);
nor_5  g03885(new_n4261, new_n4256, new_n4262);
xnor_4 g03886(new_n4262, new_n4213, new_n4263);
or_5   g03887(new_n4231, new_n4215, new_n4264);
and_5  g03888(n5798, n5331, new_n4265);
nand_5 g03889(n12648, n5579, new_n4266);
and_5  g03890(n10545, n2498, new_n4267);
and_5  g03891(n7690, n2558, new_n4268);
xnor_4 g03892(new_n4268, new_n4267, new_n4269);
xnor_4 g03893(new_n4269, new_n4266, new_n4270);
nor_5  g03894(new_n4223, new_n963, new_n4271);
and_5  g03895(new_n4223, new_n963, new_n4272);
nor_5  g03896(new_n4272, new_n4222, new_n4273);
or_5   g03897(new_n4273, new_n4271, new_n4274);
xnor_4 g03898(new_n4274, new_n4270, new_n4275);
and_5  g03899(n8476, n6016, new_n4276);
and_5  g03900(n2530, n521, new_n4277);
xnor_4 g03901(new_n4277, new_n4276, new_n4278);
xnor_4 g03902(new_n4278, new_n4275, new_n4279);
and_5  g03903(new_n4220, new_n4217, new_n4280);
nor_5  g03904(new_n4225, new_n4221, new_n4281);
nor_5  g03905(new_n4281, new_n4280, new_n4282);
xnor_4 g03906(new_n4282, new_n4279, new_n4283);
nor_5  g03907(new_n4226_1, new_n4216, new_n4284);
nor_5  g03908(new_n4230_1, new_n4227, new_n4285);
nor_5  g03909(new_n4285, new_n4284, new_n4286);
xor_4  g03910(new_n4286, new_n4283, new_n4287);
xnor_4 g03911(new_n4287, new_n4265, new_n4288);
xor_4  g03912(new_n4288, new_n4264, new_n4289);
nor_5  g03913(new_n4249, new_n4233, new_n4290);
and_5  g03914(n7965, n5153, new_n4291);
nand_5 g03915(n3342, n2393, new_n4292);
and_5  g03916(n9763, n3986, new_n4293);
and_5  g03917(n9111, n5860, new_n4294);
xnor_4 g03918(new_n4294, new_n4293, new_n4295);
xnor_4 g03919(new_n4295, new_n4292, new_n4296);
nor_5  g03920(new_n4241, new_n946, new_n4297);
and_5  g03921(new_n4241, new_n946, new_n4298);
nor_5  g03922(new_n4298, new_n4240, new_n4299);
or_5   g03923(new_n4299, new_n4297, new_n4300_1);
xnor_4 g03924(new_n4300_1, new_n4296, new_n4301);
and_5  g03925(n7388, n7270, new_n4302);
and_5  g03926(n11892, n806, new_n4303);
xnor_4 g03927(new_n4303, new_n4302, new_n4304);
xnor_4 g03928(new_n4304, new_n4301, new_n4305);
and_5  g03929(new_n4238, new_n4235, new_n4306);
nor_5  g03930(new_n4243, new_n4239, new_n4307);
nor_5  g03931(new_n4307, new_n4306, new_n4308);
xnor_4 g03932(new_n4308, new_n4305, new_n4309);
nor_5  g03933(new_n4244, new_n4234, new_n4310);
nor_5  g03934(new_n4248, new_n4245, new_n4311);
nor_5  g03935(new_n4311, new_n4310, new_n4312_1);
xor_4  g03936(new_n4312_1, new_n4309, new_n4313);
xnor_4 g03937(new_n4313, new_n4291, new_n4314);
xnor_4 g03938(new_n4314, new_n4290, new_n4315);
xnor_4 g03939(new_n4315, new_n4289, new_n4316);
nor_5  g03940(new_n4250, new_n4232, new_n4317);
nor_5  g03941(new_n4254, new_n4251, new_n4318);
nor_5  g03942(new_n4318, new_n4317, new_n4319);
xor_4  g03943(new_n4319, new_n4316, new_n4320);
xor_4  g03944(new_n4320, new_n4263, new_n4321);
nor_5  g03945(new_n4321, new_n4167, new_n4322);
xnor_4 g03946(new_n4321, new_n4167, new_n4323);
xor_4  g03947(new_n4161, new_n4160, new_n4324);
xor_4  g03948(new_n4260, new_n4259, new_n4325);
nor_5  g03949(new_n4325, new_n4324, new_n4326_1);
nor_5  g03950(new_n983, new_n905, new_n4327);
nor_5  g03951(new_n1033, new_n984, new_n4328);
nor_5  g03952(new_n4328, new_n4327, new_n4329);
xor_4  g03953(new_n4325, new_n4324, new_n4330);
and_5  g03954(new_n4330, new_n4329, new_n4331);
nor_5  g03955(new_n4331, new_n4326_1, new_n4332);
nor_5  g03956(new_n4332, new_n4323, new_n4333_1);
nor_5  g03957(new_n4333_1, new_n4322, new_n4334);
xnor_4 g03958(new_n4334, new_n4166, new_n4335);
nor_5  g03959(new_n4211, new_n4188, new_n4336);
nor_5  g03960(new_n4212, new_n4187_1, new_n4337);
nor_5  g03961(new_n4337, new_n4336, new_n4338);
or_5   g03962(new_n4210, new_n4207, new_n4339);
nor_5  g03963(new_n4205, new_n4202, new_n4340);
or_5   g03964(new_n4340, new_n4201, new_n4341);
and_5  g03965(n12221, n6776, new_n4342);
and_5  g03966(n12299, n12145, new_n4343);
and_5  g03967(n10217, n8759, new_n4344);
xnor_4 g03968(new_n4344, new_n4343, new_n4345);
xnor_4 g03969(new_n4345, new_n4342, new_n4346);
xnor_4 g03970(new_n4346, new_n4341, new_n4347);
and_5  g03971(new_n4204, new_n4203_1, new_n4348);
and_5  g03972(n7436, n2522, new_n4349);
xnor_4 g03973(new_n4349, new_n4348, new_n4350);
nand_5 g03974(n9241, n2024, new_n4351);
and_5  g03975(n10510, n7946, new_n4352);
and_5  g03976(n9189, n8276, new_n4353);
xnor_4 g03977(new_n4353, new_n4352, new_n4354);
xnor_4 g03978(new_n4354, new_n4351, new_n4355);
xor_4  g03979(new_n4355, new_n4350, new_n4356);
xor_4  g03980(new_n4356, new_n4347, new_n4357);
nor_5  g03981(new_n4194, new_n4191, new_n4358);
nand_5 g03982(new_n4193, new_n4192, new_n4359);
or_5   g03983(new_n4206, new_n4195, new_n4360);
xor_4  g03984(new_n4360, new_n4359, new_n4361);
nor_5  g03985(new_n4361, new_n4358, new_n4362);
xnor_4 g03986(new_n4362, new_n4357, new_n4363);
xnor_4 g03987(new_n4363, new_n4339, new_n4364);
xnor_4 g03988(new_n4364, new_n4338, new_n4365);
nor_5  g03989(new_n4262, new_n4213, new_n4366);
nor_5  g03990(new_n4320, new_n4263, new_n4367);
nor_5  g03991(new_n4367, new_n4366, new_n4368);
xnor_4 g03992(new_n4368, new_n4365, new_n4369);
or_5   g03993(new_n4286, new_n4283, new_n4370_1);
and_5  g03994(n8476, n5798, new_n4371);
nand_5 g03995(n6016, n2530, new_n4372);
nand_5 g03996(n5331, n2347, new_n4373);
xnor_4 g03997(new_n4373, new_n4372, new_n4374);
xnor_4 g03998(new_n4374, new_n4371, new_n4375);
nor_5  g03999(new_n4269, new_n4266, new_n4376);
nor_5  g04000(new_n4274, new_n4270, new_n4377);
or_5   g04001(new_n4377, new_n4376, new_n4378_1);
xnor_4 g04002(new_n4378_1, new_n4375, new_n4379);
and_5  g04003(new_n4268, new_n4267, new_n4380);
and_5  g04004(n12648, n521, new_n4381);
xnor_4 g04005(new_n4381, new_n4380, new_n4382);
and_5  g04006(n7690, n2498, new_n4383);
and_5  g04007(n10545, n5579, new_n4384);
and_5  g04008(n3616, n2558, new_n4385);
xnor_4 g04009(new_n4385, new_n4384, new_n4386);
xor_4  g04010(new_n4386, new_n4383, new_n4387);
xor_4  g04011(new_n4387, new_n4382, new_n4388);
xor_4  g04012(new_n4388, new_n4379, new_n4389);
nor_5  g04013(new_n4278, new_n4275, new_n4390);
nand_5 g04014(new_n4277, new_n4276, new_n4391);
or_5   g04015(new_n4282, new_n4279, new_n4392);
xor_4  g04016(new_n4392, new_n4391, new_n4393);
nor_5  g04017(new_n4393, new_n4390, new_n4394);
xnor_4 g04018(new_n4394, new_n4389, new_n4395);
xnor_4 g04019(new_n4395, new_n4370_1, new_n4396);
and_5  g04020(new_n4287, new_n4265, new_n4397_1);
nor_5  g04021(new_n4288, new_n4264, new_n4398);
nor_5  g04022(new_n4398, new_n4397_1, new_n4399);
xor_4  g04023(new_n4399, new_n4396, new_n4400);
nor_5  g04024(new_n4312_1, new_n4309, new_n4401);
nor_5  g04025(new_n4295, new_n4292, new_n4402);
nor_5  g04026(new_n4300_1, new_n4296, new_n4403);
or_5   g04027(new_n4403, new_n4402, new_n4404);
and_5  g04028(n7388, n5153, new_n4405);
and_5  g04029(n11892, n7270, new_n4406);
and_5  g04030(n7965, n2507, new_n4407);
xnor_4 g04031(new_n4407, new_n4406, new_n4408);
xnor_4 g04032(new_n4408, new_n4405, new_n4409);
xnor_4 g04033(new_n4409, new_n4404, new_n4410);
and_5  g04034(new_n4294, new_n4293, new_n4411);
and_5  g04035(n2393, n806, new_n4412);
xnor_4 g04036(new_n4412, new_n4411, new_n4413);
and_5  g04037(n9111, n3986, new_n4414);
and_5  g04038(n5860, n3342, new_n4415);
and_5  g04039(n9763, n5857, new_n4416);
xnor_4 g04040(new_n4416, new_n4415, new_n4417);
xor_4  g04041(new_n4417, new_n4414, new_n4418);
xor_4  g04042(new_n4418, new_n4413, new_n4419);
xor_4  g04043(new_n4419, new_n4410, new_n4420);
nor_5  g04044(new_n4304, new_n4301, new_n4421);
nand_5 g04045(new_n4303, new_n4302, new_n4422);
or_5   g04046(new_n4308, new_n4305, new_n4423);
xor_4  g04047(new_n4423, new_n4422, new_n4424);
nor_5  g04048(new_n4424, new_n4421, new_n4425);
xor_4  g04049(new_n4425, new_n4420, new_n4426);
xnor_4 g04050(new_n4426, new_n4401, new_n4427);
nor_5  g04051(new_n4313, new_n4291, new_n4428);
nor_5  g04052(new_n4314, new_n4290, new_n4429);
or_5   g04053(new_n4429, new_n4428, new_n4430);
xor_4  g04054(new_n4430, new_n4427, new_n4431);
xnor_4 g04055(new_n4431, new_n4400, new_n4432);
nor_5  g04056(new_n4315, new_n4289, new_n4433);
nor_5  g04057(new_n4319, new_n4316, new_n4434);
nor_5  g04058(new_n4434, new_n4433, new_n4435);
xor_4  g04059(new_n4435, new_n4432, new_n4436_1);
xor_4  g04060(new_n4436_1, new_n4369, new_n4437);
xnor_4 g04061(new_n4437, new_n4335, n1523);
nand_5 g04062(n6687, n4634, new_n4439);
and_5  g04063(n10223, n4189, new_n4440);
and_5  g04064(new_n4440, new_n3410, new_n4441);
and_5  g04065(n10223, n6687, new_n4442);
and_5  g04066(n7265, n4189, new_n4443);
nor_5  g04067(new_n4443, new_n4442, new_n4444);
nand_5 g04068(n2879, n2564, new_n4445);
nor_5  g04069(new_n4445, new_n4444, new_n4446);
nor_5  g04070(new_n4446, new_n4441, new_n4447);
xnor_4 g04071(new_n4447, new_n4439, new_n4448);
and_5  g04072(n4189, n2879, new_n4449);
and_5  g04073(n10223, n2564, new_n4450);
and_5  g04074(n7265, n6770, new_n4451);
xnor_4 g04075(new_n4451, new_n4450, new_n4452);
xor_4  g04076(new_n4452, new_n4449, new_n4453);
xnor_4 g04077(new_n4453, new_n4448, new_n4454);
nor_5  g04078(new_n4444, new_n4441, new_n4455);
and_5  g04079(n7265, n2564, new_n4456);
and_5  g04080(n6687, n2879, new_n4457);
nand_5 g04081(new_n4457, new_n4456, new_n4458);
or_5   g04082(new_n4458, new_n4455, new_n4459);
or_5   g04083(new_n4459, new_n4454, new_n4460);
nand_5 g04084(n9195, n6687, new_n4461);
nand_5 g04085(n4634, n2564, new_n4462);
and_5  g04086(n6770, n2879, new_n4463);
and_5  g04087(n9920, n7265, new_n4464);
xnor_4 g04088(new_n4464, new_n4440, new_n4465);
xor_4  g04089(new_n4465, new_n4463, new_n4466);
xnor_4 g04090(new_n4466, new_n4462, new_n4467);
nor_5  g04091(new_n4451, new_n4450, new_n4468);
nor_5  g04092(new_n4452, new_n4449, new_n4469);
or_5   g04093(new_n4469, new_n4468, new_n4470);
xnor_4 g04094(new_n4470, new_n4467, new_n4471);
xnor_4 g04095(new_n4471, new_n4461, new_n4472);
nor_5  g04096(new_n4447, new_n4439, new_n4473);
nor_5  g04097(new_n4453, new_n4448, new_n4474);
nor_5  g04098(new_n4474, new_n4473, new_n4475);
xnor_4 g04099(new_n4475, new_n4472, new_n4476);
xor_4  g04100(new_n4476, new_n4460, new_n4477);
nand_5 g04101(n8336, n2522, new_n4478);
and_5  g04102(n9189, n8336, new_n4479);
and_5  g04103(n7946, n6986, new_n4480);
nor_5  g04104(new_n4480, new_n4479, new_n4481);
and_5  g04105(n9189, n6986, new_n4482);
and_5  g04106(new_n4482, new_n3411, new_n4483);
and_5  g04107(n10928, n2024, new_n4484);
nor_5  g04108(new_n4484, new_n4483, new_n4485);
or_5   g04109(new_n4485, new_n4481, new_n4486);
xnor_4 g04110(new_n4486, new_n4478, new_n4487);
and_5  g04111(n6986, n2024, new_n4488);
and_5  g04112(n10928, n9189, new_n4489);
and_5  g04113(n7946, n2226, new_n4490);
xnor_4 g04114(new_n4490, new_n4489, new_n4491);
xor_4  g04115(new_n4491, new_n4488, new_n4492);
xnor_4 g04116(new_n4492, new_n4487, new_n4493);
nand_5 g04117(n10928, n2024, new_n4494);
or_5   g04118(new_n4494, new_n3411, new_n4495);
or_5   g04119(new_n4483, new_n4481, new_n4496);
and_5  g04120(new_n4496, new_n4495, new_n4497);
nand_5 g04121(new_n4497, new_n4484, new_n4498);
or_5   g04122(new_n4498, new_n4493, new_n4499_1);
nand_5 g04123(n12145, n8336, new_n4500);
nand_5 g04124(n10928, n2522, new_n4501);
nor_5  g04125(new_n4490, new_n4489, new_n4502);
and_5  g04126(new_n4490, new_n4489, new_n4503);
nor_5  g04127(new_n4503, new_n4488, new_n4504);
or_5   g04128(new_n4504, new_n4502, new_n4505);
xnor_4 g04129(new_n4505, new_n4501, new_n4506);
and_5  g04130(n2226, n2024, new_n4507);
and_5  g04131(n7946, n1094, new_n4508);
xnor_4 g04132(new_n4508, new_n4482, new_n4509);
xor_4  g04133(new_n4509, new_n4507, new_n4510);
xnor_4 g04134(new_n4510, new_n4506, new_n4511);
xnor_4 g04135(new_n4511, new_n4500, new_n4512);
nor_5  g04136(new_n4486, new_n4478, new_n4513);
nor_5  g04137(new_n4492, new_n4487, new_n4514);
nor_5  g04138(new_n4514, new_n4513, new_n4515);
xnor_4 g04139(new_n4515, new_n4512, new_n4516_1);
xnor_4 g04140(new_n4516_1, new_n4499_1, new_n4517);
xnor_4 g04141(new_n4498, new_n4493, new_n4518);
nand_5 g04142(n12069, n521, new_n4519);
and_5  g04143(n7891, n5579, new_n4520);
and_5  g04144(new_n4520, new_n3413, new_n4521);
and_5  g04145(n12069, n5579, new_n4522);
and_5  g04146(n7891, n2558, new_n4523);
nor_5  g04147(new_n4523, new_n4522, new_n4524);
nand_5 g04148(n12391, n2498, new_n4525);
nor_5  g04149(new_n4525, new_n4524, new_n4526);
nor_5  g04150(new_n4526, new_n4521, new_n4527);
xnor_4 g04151(new_n4527, new_n4519, new_n4528);
and_5  g04152(n7891, n2498, new_n4529);
and_5  g04153(n12391, n5579, new_n4530);
and_5  g04154(n7160, n2558, new_n4531);
xnor_4 g04155(new_n4531, new_n4530, new_n4532);
xor_4  g04156(new_n4532, new_n4529, new_n4533);
xnor_4 g04157(new_n4533, new_n4528, new_n4534);
nor_5  g04158(new_n4524, new_n4521, new_n4535);
and_5  g04159(n12391, n2558, new_n4536);
and_5  g04160(n12069, n2498, new_n4537);
nand_5 g04161(new_n4537, new_n4536, new_n4538);
or_5   g04162(new_n4538, new_n4535, new_n4539);
xor_4  g04163(new_n4539, new_n4534, new_n4540);
nand_5 g04164(n11222, n806, new_n4541);
and_5  g04165(n11222, n3342, new_n4542);
and_5  g04166(n9763, n5314, new_n4543);
nor_5  g04167(new_n4543, new_n4542, new_n4544);
and_5  g04168(n5314, n3342, new_n4545);
and_5  g04169(new_n4545, new_n3412, new_n4546);
and_5  g04170(n11153, n9111, new_n4547);
nor_5  g04171(new_n4547, new_n4546, new_n4548);
or_5   g04172(new_n4548, new_n4544, new_n4549);
xor_4  g04173(new_n4549, new_n4541, new_n4550);
and_5  g04174(n9111, n5314, new_n4551);
and_5  g04175(n11153, n3342, new_n4552);
and_5  g04176(n9763, n996, new_n4553_1);
xnor_4 g04177(new_n4553_1, new_n4552, new_n4554);
xnor_4 g04178(new_n4554, new_n4551, new_n4555);
xnor_4 g04179(new_n4555, new_n4550, new_n4556);
nand_5 g04180(n11153, n9111, new_n4557);
or_5   g04181(new_n4557, new_n3412, new_n4558);
and_5  g04182(new_n4558, new_n4544, new_n4559);
nor_5  g04183(new_n4559, new_n4546, new_n4560);
or_5   g04184(new_n4560, new_n4557, new_n4561);
xor_4  g04185(new_n4561, new_n4556, new_n4562);
xnor_4 g04186(new_n4562, new_n4540, new_n4563);
or_5   g04187(new_n4558, new_n4544, new_n4564);
and_5  g04188(new_n4564, new_n4560, new_n4565);
and_5  g04189(new_n3413, new_n3412, new_n4566);
xor_4  g04190(new_n4537, new_n4536, new_n4567);
nor_5  g04191(new_n4567, new_n4566, new_n4568);
xnor_4 g04192(new_n4567, new_n4566, new_n4569);
and_5  g04193(n11153, n9763, new_n4570);
and_5  g04194(n11222, n9111, new_n4571);
xor_4  g04195(new_n4571, new_n4570, new_n4572);
nor_5  g04196(new_n4572, new_n4569, new_n4573);
nor_5  g04197(new_n4573, new_n4568, new_n4574);
nor_5  g04198(new_n4574, new_n4565, new_n4575);
xnor_4 g04199(new_n4574, new_n4565, new_n4576);
nor_5  g04200(new_n4525, new_n3413, new_n4577);
nor_5  g04201(new_n4577, new_n4535, new_n4578);
or_5   g04202(new_n4525, new_n3413, new_n4579);
nor_5  g04203(new_n4579, new_n4524, new_n4580);
nor_5  g04204(new_n4580, new_n4578, new_n4581);
nor_5  g04205(new_n4581, new_n4576, new_n4582);
nor_5  g04206(new_n4582, new_n4575, new_n4583);
xor_4  g04207(new_n4583, new_n4563, new_n4584);
nor_5  g04208(new_n4584, new_n4518, new_n4585);
xnor_4 g04209(new_n4584, new_n4518, new_n4586);
nor_5  g04210(new_n4495, new_n4481, new_n4587);
or_5   g04211(new_n4587, new_n4497, new_n4588);
xor_4  g04212(new_n4581, new_n4576, new_n4589);
nor_5  g04213(new_n4589, new_n4588, new_n4590);
xnor_4 g04214(new_n4589, new_n4588, new_n4591);
xor_4  g04215(new_n4572, new_n4569, new_n4592);
and_5  g04216(n10928, n7946, new_n4593);
and_5  g04217(n8336, n2024, new_n4594);
xnor_4 g04218(new_n4594, new_n4593, new_n4595);
nor_5  g04219(new_n4595, new_n4592, new_n4596);
nand_5 g04220(n8336, n7946, new_n4597);
or_5   g04221(new_n3414, new_n4597, new_n4598);
xnor_4 g04222(new_n4595, new_n4592, new_n4599);
nor_5  g04223(new_n4599, new_n4598, new_n4600);
nor_5  g04224(new_n4600, new_n4596, new_n4601);
nor_5  g04225(new_n4601, new_n4591, new_n4602);
nor_5  g04226(new_n4602, new_n4590, new_n4603);
nor_5  g04227(new_n4603, new_n4586, new_n4604);
nor_5  g04228(new_n4604, new_n4585, new_n4605);
xnor_4 g04229(new_n4605, new_n4517, new_n4606);
or_5   g04230(new_n4539, new_n4534, new_n4607);
nand_5 g04231(n12069, n6016, new_n4608);
nand_5 g04232(n12391, n521, new_n4609);
nor_5  g04233(new_n4531, new_n4530, new_n4610);
and_5  g04234(new_n4531, new_n4530, new_n4611);
nor_5  g04235(new_n4611, new_n4529, new_n4612);
or_5   g04236(new_n4612, new_n4610, new_n4613);
xnor_4 g04237(new_n4613, new_n4609, new_n4614);
and_5  g04238(n7160, n2498, new_n4615);
nand_5 g04239(n4828, n2558, new_n4616);
xor_4  g04240(new_n4616, new_n4520, new_n4617);
xor_4  g04241(new_n4617, new_n4615, new_n4618);
xnor_4 g04242(new_n4618, new_n4614, new_n4619);
xnor_4 g04243(new_n4619, new_n4608, new_n4620);
nor_5  g04244(new_n4527, new_n4519, new_n4621);
nor_5  g04245(new_n4533, new_n4528, new_n4622);
nor_5  g04246(new_n4622, new_n4621, new_n4623);
xnor_4 g04247(new_n4623, new_n4620, new_n4624);
xor_4  g04248(new_n4624, new_n4607, new_n4625);
or_5   g04249(new_n4561, new_n4556, new_n4626);
nand_5 g04250(n11222, n7270, new_n4627);
nand_5 g04251(n11153, n806, new_n4628);
nor_5  g04252(new_n4553_1, new_n4552, new_n4629);
and_5  g04253(new_n4553_1, new_n4552, new_n4630);
nor_5  g04254(new_n4630, new_n4551, new_n4631);
or_5   g04255(new_n4631, new_n4629, new_n4632);
xnor_4 g04256(new_n4632, new_n4628, new_n4633);
and_5  g04257(n9111, n996, new_n4634_1);
and_5  g04258(n9763, n5767, new_n4635);
xnor_4 g04259(new_n4635, new_n4545, new_n4636);
xor_4  g04260(new_n4636, new_n4634_1, new_n4637);
xnor_4 g04261(new_n4637, new_n4633, new_n4638);
xnor_4 g04262(new_n4638, new_n4627, new_n4639);
nor_5  g04263(new_n4549, new_n4541, new_n4640);
and_5  g04264(new_n4555, new_n4550, new_n4641);
nor_5  g04265(new_n4641, new_n4640, new_n4642);
xnor_4 g04266(new_n4642, new_n4639, new_n4643);
xor_4  g04267(new_n4643, new_n4626, new_n4644);
xnor_4 g04268(new_n4644, new_n4625, new_n4645);
nor_5  g04269(new_n4562, new_n4540, new_n4646);
nor_5  g04270(new_n4583, new_n4563, new_n4647);
nor_5  g04271(new_n4647, new_n4646, new_n4648);
xor_4  g04272(new_n4648, new_n4645, new_n4649);
xor_4  g04273(new_n4649, new_n4606, new_n4650);
xnor_4 g04274(new_n4650, new_n4477, new_n4651);
xor_4  g04275(new_n4459, new_n4454, new_n4652);
xor_4  g04276(new_n4603, new_n4586, new_n4653);
nor_5  g04277(new_n4653, new_n4652, new_n4654);
xor_4  g04278(new_n4601, new_n4591, new_n4655);
nor_5  g04279(new_n4445, new_n3410, new_n4656);
nor_5  g04280(new_n4656, new_n4455, new_n4657);
or_5   g04281(new_n4445, new_n3410, new_n4658);
nor_5  g04282(new_n4658, new_n4444, new_n4659);
nor_5  g04283(new_n4659, new_n4657, new_n4660);
nor_5  g04284(new_n4660, new_n4655, new_n4661);
xnor_4 g04285(new_n4660, new_n4655, new_n4662);
and_5  g04286(new_n3415, new_n3410, new_n4663);
xor_4  g04287(new_n4457, new_n4456, new_n4664);
nor_5  g04288(new_n4664, new_n4663, new_n4665);
xnor_4 g04289(new_n4599, new_n4598, new_n4666);
xor_4  g04290(new_n4664, new_n4663, new_n4667);
and_5  g04291(new_n4667, new_n4666, new_n4668);
nor_5  g04292(new_n4668, new_n4665, new_n4669);
nor_5  g04293(new_n4669, new_n4662, new_n4670);
nor_5  g04294(new_n4670, new_n4661, new_n4671);
xnor_4 g04295(new_n4653, new_n4652, new_n4672);
nor_5  g04296(new_n4672, new_n4671, new_n4673);
nor_5  g04297(new_n4673, new_n4654, new_n4674);
xnor_4 g04298(new_n4674, new_n4651, n1658);
nand_5 g04299(n7862, n4634, new_n4676);
and_5  g04300(n10223, n7862, new_n4677);
and_5  g04301(n7265, n3172, new_n4678);
nor_5  g04302(new_n4678, new_n4677, new_n4679);
and_5  g04303(n7862, n7265, new_n4680);
and_5  g04304(n10223, n3172, new_n4681);
and_5  g04305(new_n4681, new_n4680, new_n4682);
and_5  g04306(n2879, n1333, new_n4683);
nor_5  g04307(new_n4683, new_n4682, new_n4684);
or_5   g04308(new_n4684, new_n4679, new_n4685);
xnor_4 g04309(new_n4685, new_n4676, new_n4686_1);
and_5  g04310(n3172, n2879, new_n4687);
and_5  g04311(n10223, n1333, new_n4688);
and_5  g04312(n11757, n7265, new_n4689_1);
xnor_4 g04313(new_n4689_1, new_n4688, new_n4690);
xor_4  g04314(new_n4690, new_n4687, new_n4691);
xnor_4 g04315(new_n4691, new_n4686_1, new_n4692);
nand_5 g04316(n2879, n1333, new_n4693);
or_5   g04317(new_n4693, new_n4680, new_n4694);
and_5  g04318(new_n4694, new_n4679, new_n4695);
nor_5  g04319(new_n4695, new_n4682, new_n4696);
or_5   g04320(new_n4696, new_n4693, new_n4697);
xor_4  g04321(new_n4697, new_n4692, new_n4698);
nand_5 g04322(n6877, n2522, new_n4699);
and_5  g04323(n2464, n2024, new_n4700);
and_5  g04324(n9400, n9189, new_n4701);
and_5  g04325(n11311, n7946, new_n4702);
xnor_4 g04326(new_n4702, new_n4701, new_n4703);
xor_4  g04327(new_n4703, new_n4700, new_n4704);
xnor_4 g04328(new_n4704, new_n4699, new_n4705);
and_5  g04329(n9189, n6877, new_n4706);
and_5  g04330(n7946, n2464, new_n4707);
nor_5  g04331(new_n4707, new_n4706, new_n4708);
and_5  g04332(n7946, n6877, new_n4709);
and_5  g04333(n9189, n2464, new_n4710);
and_5  g04334(new_n4710, new_n4709, new_n4711);
and_5  g04335(n9400, n2024, new_n4712);
nor_5  g04336(new_n4712, new_n4711, new_n4713);
or_5   g04337(new_n4713, new_n4708, new_n4714);
xnor_4 g04338(new_n4714, new_n4705, new_n4715);
nand_5 g04339(n9400, n2024, new_n4716);
or_5   g04340(new_n4716, new_n4709, new_n4717);
or_5   g04341(new_n4711, new_n4708, new_n4718);
nand_5 g04342(new_n4718, new_n4717, new_n4719);
or_5   g04343(new_n4719, new_n4716, new_n4720);
xnor_4 g04344(new_n4720, new_n4715, new_n4721);
or_5   g04345(new_n4717, new_n4708, new_n4722_1);
and_5  g04346(new_n4722_1, new_n4719, new_n4723);
nand_5 g04347(n7946, n6877, new_n4724);
and_5  g04348(n4805, n2558, new_n4725);
and_5  g04349(n9763, n7236, new_n4726);
xnor_4 g04350(new_n4726, new_n4725, new_n4727);
nor_5  g04351(new_n4727, new_n4724, new_n4728);
and_5  g04352(n9400, n7946, new_n4729);
and_5  g04353(n6877, n2024, new_n4730);
xor_4  g04354(new_n4730, new_n4729, new_n4731);
and_5  g04355(new_n4731, new_n4728, new_n4732);
and_5  g04356(new_n4726, new_n4725, new_n4733_1);
and_5  g04357(n9111, n7236, new_n4734);
and_5  g04358(n9763, n3992, new_n4735);
xor_4  g04359(new_n4735, new_n4734, new_n4736);
xnor_4 g04360(new_n4736, new_n4733_1, new_n4737);
and_5  g04361(n4805, n2498, new_n4738);
and_5  g04362(n11478, n2558, new_n4739);
xor_4  g04363(new_n4739, new_n4738, new_n4740);
xor_4  g04364(new_n4740, new_n4737, new_n4741);
xnor_4 g04365(new_n4731, new_n4728, new_n4742);
nor_5  g04366(new_n4742, new_n4741, new_n4743);
or_5   g04367(new_n4743, new_n4732, new_n4744);
nor_5  g04368(new_n4744, new_n4723, new_n4745);
nor_5  g04369(new_n4736, new_n4733_1, new_n4746);
nor_5  g04370(new_n4740, new_n4737, new_n4747);
nor_5  g04371(new_n4747, new_n4746, new_n4748);
nand_5 g04372(n11478, n2498, new_n4749);
or_5   g04373(new_n4749, new_n4725, new_n4750);
and_5  g04374(n5283, n2558, new_n4751);
and_5  g04375(n5579, n4805, new_n4752);
xnor_4 g04376(new_n4752, new_n4751, new_n4753);
nand_5 g04377(new_n4753, new_n4750, new_n4754);
nor_5  g04378(new_n4752, new_n4751, new_n4755);
or_5   g04379(new_n4755, new_n4750, new_n4756);
and_5  g04380(new_n4756, new_n4754, new_n4757_1);
xnor_4 g04381(new_n4757_1, new_n4748, new_n4758);
nand_5 g04382(n9111, n3992, new_n4759);
nor_5  g04383(new_n4759, new_n4726, new_n4760);
and_5  g04384(n9763, n8384, new_n4761);
and_5  g04385(n7236, n3342, new_n4762);
nor_5  g04386(new_n4762, new_n4761, new_n4763);
and_5  g04387(new_n4763, new_n4760, new_n4764);
xnor_4 g04388(new_n4762, new_n4761, new_n4765);
nor_5  g04389(new_n4765, new_n4760, new_n4766);
or_5   g04390(new_n4766, new_n4764, new_n4767);
xnor_4 g04391(new_n4767, new_n4758, new_n4768);
xnor_4 g04392(new_n4744, new_n4723, new_n4769);
nor_5  g04393(new_n4769, new_n4768, new_n4770);
or_5   g04394(new_n4770, new_n4745, new_n4771);
xnor_4 g04395(new_n4771, new_n4721, new_n4772);
nand_5 g04396(n4805, n521, new_n4773);
nand_5 g04397(new_n4752, new_n4751, new_n4774);
and_5  g04398(new_n4774, new_n4749, new_n4775);
or_5   g04399(new_n4775, new_n4755, new_n4776);
xnor_4 g04400(new_n4776, new_n4773, new_n4777);
and_5  g04401(n5283, n2498, new_n4778);
and_5  g04402(n2558, n137, new_n4779);
and_5  g04403(n11478, n5579, new_n4780);
xnor_4 g04404(new_n4780, new_n4779, new_n4781);
xor_4  g04405(new_n4781, new_n4778, new_n4782);
xnor_4 g04406(new_n4782, new_n4777, new_n4783);
or_5   g04407(new_n4754, new_n4749, new_n4784);
xor_4  g04408(new_n4784, new_n4783, new_n4785);
nand_5 g04409(n7236, n806, new_n4786);
and_5  g04410(new_n4762, new_n4761, new_n4787);
nor_5  g04411(new_n4763, new_n4759, new_n4788);
nor_5  g04412(new_n4788, new_n4787, new_n4789);
xor_4  g04413(new_n4789, new_n4786, new_n4790);
and_5  g04414(n9111, n8384, new_n4791);
and_5  g04415(n9763, n6358, new_n4792);
and_5  g04416(n3992, n3342, new_n4793);
xnor_4 g04417(new_n4793, new_n4792, new_n4794);
xnor_4 g04418(new_n4794, new_n4791, new_n4795);
xnor_4 g04419(new_n4795, new_n4790, new_n4796);
and_5  g04420(new_n4735, new_n4734, new_n4797);
nand_5 g04421(new_n4765, new_n4797, new_n4798);
xor_4  g04422(new_n4798, new_n4796, new_n4799);
xnor_4 g04423(new_n4799, new_n4785, new_n4800);
nor_5  g04424(new_n4757_1, new_n4748, new_n4801);
nor_5  g04425(new_n4767, new_n4758, new_n4802);
nor_5  g04426(new_n4802, new_n4801, new_n4803);
xor_4  g04427(new_n4803, new_n4800, new_n4804);
xor_4  g04428(new_n4804, new_n4772, new_n4805_1);
xnor_4 g04429(new_n4805_1, new_n4698, new_n4806);
or_5   g04430(new_n4694, new_n4679, new_n4807);
nand_5 g04431(new_n4807, new_n4696, new_n4808);
xor_4  g04432(new_n4769, new_n4768, new_n4809);
nor_5  g04433(new_n4809, new_n4808, new_n4810);
xnor_4 g04434(new_n4727, new_n4709, new_n4811);
and_5  g04435(new_n4811, new_n4680, new_n4812);
and_5  g04436(n7265, n1333, new_n4813);
and_5  g04437(n7862, n2879, new_n4814);
xor_4  g04438(new_n4814, new_n4813, new_n4815);
nor_5  g04439(new_n4815, new_n4812, new_n4816);
xnor_4 g04440(new_n4742, new_n4741, new_n4817_1);
xor_4  g04441(new_n4815, new_n4812, new_n4818);
and_5  g04442(new_n4818, new_n4817_1, new_n4819);
or_5   g04443(new_n4819, new_n4816, new_n4820);
xnor_4 g04444(new_n4809, new_n4808, new_n4821);
nor_5  g04445(new_n4821, new_n4820, new_n4822);
or_5   g04446(new_n4822, new_n4810, new_n4823);
xnor_4 g04447(new_n4823, new_n4806, n1847);
nand_5 g04448(n5305, n1798, new_n4825);
nand_5 g04449(n8759, n6703, new_n4826_1);
and_5  g04450(n5645, n5331, new_n4827);
and_5  g04451(n11876, n7965, new_n4828_1);
xnor_4 g04452(new_n4828_1, new_n4827, new_n4829);
xnor_4 g04453(new_n4829, new_n4826_1, new_n4830);
nor_5  g04454(new_n4830, new_n4825, new_n4831);
and_5  g04455(n5305, n3932, new_n4832);
and_5  g04456(n5964, n1798, new_n4833);
xor_4  g04457(new_n4833, new_n4832, new_n4834);
xnor_4 g04458(new_n4834, new_n4831, new_n4835);
nor_5  g04459(new_n4829, new_n4826_1, new_n4836);
and_5  g04460(n9640, n8759, new_n4837);
and_5  g04461(n6776, n6703, new_n4838);
xor_4  g04462(new_n4838, new_n4837, new_n4839);
xnor_4 g04463(new_n4839, new_n4836, new_n4840);
and_5  g04464(new_n4828_1, new_n4827, new_n4841);
and_5  g04465(n10898, n7965, new_n4842);
and_5  g04466(n11876, n7388, new_n4843);
xor_4  g04467(new_n4843, new_n4842, new_n4844);
xnor_4 g04468(new_n4844, new_n4841, new_n4845);
and_5  g04469(n5331, n1067, new_n4846);
and_5  g04470(n8476, n5645, new_n4847);
xnor_4 g04471(new_n4847, new_n4846, new_n4848);
xnor_4 g04472(new_n4848, new_n4845, new_n4849);
xnor_4 g04473(new_n4849, new_n4840, new_n4850);
xor_4  g04474(new_n4850, new_n4835, n2096);
xor_4  g04475(new_n2907, new_n2906, n2131);
and_5  g04476(n7456, n2564, new_n4853);
nor_5  g04477(new_n3030, new_n3029, new_n4854);
and_5  g04478(new_n3030, new_n3029, new_n4855);
nor_5  g04479(new_n4855, new_n3028, new_n4856);
nor_5  g04480(new_n4856, new_n4854, new_n4857);
and_5  g04481(new_n4857, new_n4853, new_n4858);
xnor_4 g04482(new_n4857, new_n4853, new_n4859);
and_5  g04483(n6770, n3932, new_n4860);
and_5  g04484(n9920, n1798, new_n4861);
xnor_4 g04485(new_n4861, new_n3022_1, new_n4862);
xor_4  g04486(new_n4862, new_n4860, new_n4863);
nor_5  g04487(new_n4863, new_n4859, new_n4864);
nor_5  g04488(new_n4864, new_n4858, new_n4865);
and_5  g04489(n11662, n2564, new_n4866);
and_5  g04490(n7456, n4189, new_n4867);
xnor_4 g04491(new_n4867, new_n4866, new_n4868);
xnor_4 g04492(new_n4868, new_n4865, new_n4869);
nand_5 g04493(n12591, n6770, new_n4870);
and_5  g04494(n3627, n1798, new_n4871);
and_5  g04495(n9920, n3932, new_n4872);
xnor_4 g04496(new_n4872, new_n4871, new_n4873);
xnor_4 g04497(new_n4873, new_n4870, new_n4874);
nor_5  g04498(new_n4861, new_n3022_1, new_n4875);
and_5  g04499(new_n4861, new_n3022_1, new_n4876);
nor_5  g04500(new_n4876, new_n4860, new_n4877);
or_5   g04501(new_n4877, new_n4875, new_n4878);
xnor_4 g04502(new_n4878, new_n4874, new_n4879);
xnor_4 g04503(new_n4879, new_n4869, new_n4880);
and_5  g04504(n11662, n6687, new_n4881);
nor_5  g04505(new_n3026, new_n3017, new_n4882);
nor_5  g04506(new_n3032, new_n3027, new_n4883);
or_5   g04507(new_n4883, new_n4882, new_n4884);
nor_5  g04508(new_n4884, new_n4881, new_n4885);
xor_4  g04509(new_n4863, new_n4859, new_n4886);
xnor_4 g04510(new_n4884, new_n4881, new_n4887);
nor_5  g04511(new_n4887, new_n4886, new_n4888);
or_5   g04512(new_n4888, new_n4885, new_n4889);
or_5   g04513(new_n4889, new_n4880, new_n4890);
nor_5  g04514(new_n4873, new_n4870, new_n4891);
nor_5  g04515(new_n4878, new_n4874, new_n4892);
or_5   g04516(new_n4892, new_n4891, new_n4893);
and_5  g04517(n10327, n2564, new_n4894);
and_5  g04518(n11662, n4189, new_n4895);
and_5  g04519(n9583, n6687, new_n4896);
xnor_4 g04520(new_n4896, new_n4895, new_n4897);
xnor_4 g04521(new_n4897, new_n4894, new_n4898);
xnor_4 g04522(new_n4898, new_n4893, new_n4899);
and_5  g04523(new_n4872, new_n4871, new_n4900);
and_5  g04524(n7456, n6770, new_n4901);
xnor_4 g04525(new_n4901, new_n4900, new_n4902);
nand_5 g04526(n3932, n3627, new_n4903_1);
and_5  g04527(n12591, n9920, new_n4904);
and_5  g04528(n4516, n1798, new_n4905);
xnor_4 g04529(new_n4905, new_n4904, new_n4906);
xnor_4 g04530(new_n4906, new_n4903_1, new_n4907);
xor_4  g04531(new_n4907, new_n4902, new_n4908);
xor_4  g04532(new_n4908, new_n4899, new_n4909);
nor_5  g04533(new_n4868, new_n4865, new_n4910);
nand_5 g04534(new_n4867, new_n4866, new_n4911);
or_5   g04535(new_n4879, new_n4869, new_n4912);
xor_4  g04536(new_n4912, new_n4911, new_n4913);
nor_5  g04537(new_n4913, new_n4910, new_n4914);
xnor_4 g04538(new_n4914, new_n4909, new_n4915);
xnor_4 g04539(new_n4915, new_n4890, new_n4916);
and_5  g04540(n10327, n6687, new_n4917);
xor_4  g04541(new_n4889, new_n4880, new_n4918);
and_5  g04542(new_n4918, new_n4917, new_n4919);
or_5   g04543(new_n3038, new_n3033, new_n4920);
xor_4  g04544(new_n4887, new_n4886, new_n4921_1);
or_5   g04545(new_n4921_1, new_n4920, new_n4922);
xnor_4 g04546(new_n4918, new_n4917, new_n4923);
nor_5  g04547(new_n4923, new_n4922, new_n4924);
nor_5  g04548(new_n4924, new_n4919, new_n4925);
xor_4  g04549(new_n4925, new_n4916, new_n4926);
nand_5 g04550(n3022, n2226, new_n4927);
and_5  g04551(n9640, n1094, new_n4928_1);
and_5  g04552(n10678, n6703, new_n4929);
xnor_4 g04553(new_n4929, new_n4928_1, new_n4930);
xnor_4 g04554(new_n4930, new_n4927, new_n4931);
and_5  g04555(n6703, n1094, new_n4932);
nor_5  g04556(new_n4932, new_n3069, new_n4933);
nand_5 g04557(new_n4932, new_n3069, new_n4934);
nand_5 g04558(n9640, n2226, new_n4935);
and_5  g04559(new_n4935, new_n4934, new_n4936);
or_5   g04560(new_n4936, new_n4933, new_n4937);
xnor_4 g04561(new_n4937, new_n4931, new_n4938_1);
and_5  g04562(n10928, n10451, new_n4939);
and_5  g04563(n11023, n6986, new_n4940);
xnor_4 g04564(new_n4940, new_n4939, new_n4941);
xnor_4 g04565(new_n4941, new_n4938_1, new_n4942);
nand_5 g04566(n11023, n10928, new_n4943);
nor_5  g04567(new_n3153, new_n3152, new_n4944);
and_5  g04568(new_n3153, new_n3152, new_n4945);
nor_5  g04569(new_n4945, new_n3151, new_n4946);
or_5   g04570(new_n4946, new_n4944, new_n4947);
nor_5  g04571(new_n4947, new_n4943, new_n4948);
xnor_4 g04572(new_n4947, new_n4943, new_n4949);
xnor_4 g04573(new_n4932, new_n3069, new_n4950);
xnor_4 g04574(new_n4950, new_n4935, new_n4951);
nor_5  g04575(new_n4951, new_n4949, new_n4952);
nor_5  g04576(new_n4952, new_n4948, new_n4953);
xnor_4 g04577(new_n4953, new_n4942, new_n4954);
nand_5 g04578(n10451, n8336, new_n4955);
xnor_4 g04579(new_n4951, new_n4949, new_n4956);
nor_5  g04580(new_n4956, new_n4955, new_n4957);
nor_5  g04581(new_n3149, new_n3146_1, new_n4958);
nor_5  g04582(new_n3155, new_n3150, new_n4959);
nor_5  g04583(new_n4959, new_n4958, new_n4960);
xnor_4 g04584(new_n4956, new_n4955, new_n4961);
nor_5  g04585(new_n4961, new_n4960, new_n4962);
nor_5  g04586(new_n4962, new_n4957, new_n4963);
or_5   g04587(new_n4963, new_n4954, new_n4964);
nor_5  g04588(new_n4930, new_n4927, new_n4965);
nor_5  g04589(new_n4937, new_n4931, new_n4966);
or_5   g04590(new_n4966, new_n4965, new_n4967);
and_5  g04591(n10928, n10278, new_n4968);
and_5  g04592(n10451, n6986, new_n4969);
and_5  g04593(n11423, n8336, new_n4970_1);
xnor_4 g04594(new_n4970_1, new_n4969, new_n4971_1);
xnor_4 g04595(new_n4971_1, new_n4968, new_n4972);
xnor_4 g04596(new_n4972, new_n4967, new_n4973);
and_5  g04597(new_n4929, new_n4928_1, new_n4974);
and_5  g04598(n11023, n2226, new_n4975);
xnor_4 g04599(new_n4975, new_n4974, new_n4976);
and_5  g04600(n10678, n9640, new_n4977);
and_5  g04601(n3022, n1094, new_n4978);
and_5  g04602(n7320, n6703, new_n4979);
xnor_4 g04603(new_n4979, new_n4978, new_n4980);
xor_4  g04604(new_n4980, new_n4977, new_n4981);
xor_4  g04605(new_n4981, new_n4976, new_n4982);
xor_4  g04606(new_n4982, new_n4973, new_n4983);
nor_5  g04607(new_n4941, new_n4938_1, new_n4984);
nand_5 g04608(new_n4940, new_n4939, new_n4985);
or_5   g04609(new_n4953, new_n4942, new_n4986);
xor_4  g04610(new_n4986, new_n4985, new_n4987);
nor_5  g04611(new_n4987, new_n4984, new_n4988);
xnor_4 g04612(new_n4988, new_n4983, new_n4989);
xnor_4 g04613(new_n4989, new_n4964, new_n4990);
and_5  g04614(n10278, n8336, new_n4991);
xor_4  g04615(new_n4963, new_n4954, new_n4992);
nor_5  g04616(new_n4992, new_n4991, new_n4993);
or_5   g04617(new_n3157, new_n3156, new_n4994);
xnor_4 g04618(new_n4961, new_n4960, new_n4995);
nor_5  g04619(new_n4995, new_n4994, new_n4996);
xnor_4 g04620(new_n4992, new_n4991, new_n4997);
nor_5  g04621(new_n4997, new_n4996, new_n4998);
or_5   g04622(new_n4998, new_n4993, new_n4999);
xnor_4 g04623(new_n4999, new_n4990, new_n5000);
nand_5 g04624(n8665, n7160, new_n5001);
and_5  g04625(n4828, n1067, new_n5002);
and_5  g04626(n5645, n2515, new_n5003);
xnor_4 g04627(new_n5003, new_n5002, new_n5004);
xnor_4 g04628(new_n5004, new_n5001, new_n5005);
and_5  g04629(n5645, n4828, new_n5006);
and_5  g04630(n8665, n7891, new_n5007);
nor_5  g04631(new_n5007, new_n5006, new_n5008);
and_5  g04632(n7160, n1067, new_n5009);
xnor_4 g04633(new_n5007, new_n5006, new_n5010);
nor_5  g04634(new_n5010, new_n5009, new_n5011);
or_5   g04635(new_n5011, new_n5008, new_n5012);
xnor_4 g04636(new_n5012, new_n5005, new_n5013);
and_5  g04637(n12391, n2551, new_n5014);
and_5  g04638(n11922, n7891, new_n5015);
xnor_4 g04639(new_n5015, new_n5014, new_n5016);
xnor_4 g04640(new_n5016, new_n5013, new_n5017);
and_5  g04641(n12391, n11922, new_n5018);
nor_5  g04642(new_n3123, new_n3122, new_n5019);
nor_5  g04643(new_n3124_1, new_n3121, new_n5020);
nor_5  g04644(new_n5020, new_n5019, new_n5021);
and_5  g04645(new_n5021, new_n5018, new_n5022);
xor_4  g04646(new_n5010, new_n5009, new_n5023);
xnor_4 g04647(new_n5021, new_n5018, new_n5024);
nor_5  g04648(new_n5024, new_n5023, new_n5025);
nor_5  g04649(new_n5025, new_n5022, new_n5026);
xnor_4 g04650(new_n5026, new_n5017, new_n5027);
and_5  g04651(n12069, n2551, new_n5028);
xor_4  g04652(new_n5024, new_n5023, new_n5029);
and_5  g04653(new_n5029, new_n5028, new_n5030_1);
nor_5  g04654(new_n5029, new_n5028, new_n5031);
nor_5  g04655(new_n3119, new_n3116, new_n5032);
nor_5  g04656(new_n3125, new_n3120, new_n5033);
nor_5  g04657(new_n5033, new_n5032, new_n5034_1);
nor_5  g04658(new_n5034_1, new_n5031, new_n5035);
nor_5  g04659(new_n5035, new_n5030_1, new_n5036);
nor_5  g04660(new_n5036, new_n5027, new_n5037);
nor_5  g04661(new_n5004, new_n5001, new_n5038);
nor_5  g04662(new_n5012, new_n5005, new_n5039);
or_5   g04663(new_n5039, new_n5038, new_n5040);
and_5  g04664(n12826, n12391, new_n5041);
and_5  g04665(n7891, n2551, new_n5042);
and_5  g04666(n12069, n4094, new_n5043);
xnor_4 g04667(new_n5043, new_n5042, new_n5044);
xnor_4 g04668(new_n5044, new_n5041, new_n5045);
xnor_4 g04669(new_n5045, new_n5040, new_n5046);
and_5  g04670(new_n5003, new_n5002, new_n5047);
and_5  g04671(n11922, n7160, new_n5048);
xnor_4 g04672(new_n5048, new_n5047, new_n5049);
nand_5 g04673(n2515, n1067, new_n5050);
and_5  g04674(n8665, n4828, new_n5051);
and_5  g04675(n5645, n1199, new_n5052);
xnor_4 g04676(new_n5052, new_n5051, new_n5053);
xnor_4 g04677(new_n5053, new_n5050, new_n5054);
xor_4  g04678(new_n5054, new_n5049, new_n5055);
xor_4  g04679(new_n5055, new_n5046, new_n5056);
nor_5  g04680(new_n5016, new_n5013, new_n5057);
nand_5 g04681(new_n5015, new_n5014, new_n5058);
or_5   g04682(new_n5026, new_n5017, new_n5059);
xor_4  g04683(new_n5059, new_n5058, new_n5060);
nor_5  g04684(new_n5060, new_n5057, new_n5061);
xor_4  g04685(new_n5061, new_n5056, new_n5062);
xnor_4 g04686(new_n5062, new_n5037, new_n5063);
and_5  g04687(n12826, n12069, new_n5064);
xor_4  g04688(new_n5036, new_n5027, new_n5065);
nor_5  g04689(new_n5065, new_n5064, new_n5066);
or_5   g04690(new_n3126, new_n3115, new_n5067);
xnor_4 g04691(new_n5029, new_n5028, new_n5068);
xnor_4 g04692(new_n5068, new_n5034_1, new_n5069_1);
nor_5  g04693(new_n5069_1, new_n5067, new_n5070);
xnor_4 g04694(new_n5065, new_n5064, new_n5071);
nor_5  g04695(new_n5071, new_n5070, new_n5072);
or_5   g04696(new_n5072, new_n5066, new_n5073);
xor_4  g04697(new_n5073, new_n5063, new_n5074);
nand_5 g04698(n3754, n996, new_n5075);
and_5  g04699(n10898, n5767, new_n5076);
and_5  g04700(n11876, n5319, new_n5077);
xnor_4 g04701(new_n5077, new_n5076, new_n5078);
xnor_4 g04702(new_n5078, new_n5075, new_n5079);
and_5  g04703(n10898, n996, new_n5080);
nor_5  g04704(new_n5080, new_n3092, new_n5081);
and_5  g04705(n11876, n5767, new_n5082);
xnor_4 g04706(new_n5080, new_n3092, new_n5083);
nor_5  g04707(new_n5083, new_n5082, new_n5084);
or_5   g04708(new_n5084, new_n5081, new_n5085);
xnor_4 g04709(new_n5085, new_n5079, new_n5086);
and_5  g04710(n11153, n159, new_n5087);
and_5  g04711(n5314, n2749, new_n5088);
xnor_4 g04712(new_n5088, new_n5087, new_n5089);
xnor_4 g04713(new_n5089, new_n5086, new_n5090);
and_5  g04714(n11153, n2749, new_n5091);
nor_5  g04715(new_n3135, new_n3134, new_n5092);
nor_5  g04716(new_n3136, new_n3133, new_n5093);
nor_5  g04717(new_n5093, new_n5092, new_n5094_1);
and_5  g04718(new_n5094_1, new_n5091, new_n5095);
xnor_4 g04719(new_n5094_1, new_n5091, new_n5096);
xor_4  g04720(new_n5083, new_n5082, new_n5097);
nor_5  g04721(new_n5097, new_n5096, new_n5098);
nor_5  g04722(new_n5098, new_n5095, new_n5099);
xnor_4 g04723(new_n5099, new_n5090, new_n5100);
and_5  g04724(n11222, n159, new_n5101);
xor_4  g04725(new_n5097, new_n5096, new_n5102);
and_5  g04726(new_n5102, new_n5101, new_n5103);
nor_5  g04727(new_n5102, new_n5101, new_n5104);
and_5  g04728(new_n3131, new_n3128, new_n5105_1);
nor_5  g04729(new_n3137, new_n3132, new_n5106);
nor_5  g04730(new_n5106, new_n5105_1, new_n5107);
nor_5  g04731(new_n5107, new_n5104, new_n5108);
nor_5  g04732(new_n5108, new_n5103, new_n5109);
or_5   g04733(new_n5109, new_n5100, new_n5110);
nor_5  g04734(new_n5089, new_n5086, new_n5111);
nand_5 g04735(new_n5088, new_n5087, new_n5112);
or_5   g04736(new_n5099, new_n5090, new_n5113);
xor_4  g04737(new_n5113, new_n5112, new_n5114);
nor_5  g04738(new_n5114, new_n5111, new_n5115);
nor_5  g04739(new_n5078, new_n5075, new_n5116);
nor_5  g04740(new_n5085, new_n5079, new_n5117);
nor_5  g04741(new_n5117, new_n5116, new_n5118);
and_5  g04742(n11153, n1510, new_n5119);
and_5  g04743(n5314, n159, new_n5120);
and_5  g04744(n12247, n11222, new_n5121);
xnor_4 g04745(new_n5121, new_n5120, new_n5122);
xor_4  g04746(new_n5122, new_n5119, new_n5123);
xnor_4 g04747(new_n5123, new_n5118, new_n5124);
and_5  g04748(new_n5077, new_n5076, new_n5125);
and_5  g04749(n2749, n996, new_n5126);
xnor_4 g04750(new_n5126, new_n5125, new_n5127);
and_5  g04751(n10898, n5319, new_n5128);
and_5  g04752(n11876, n9457, new_n5129);
and_5  g04753(n5767, n3754, new_n5130);
xnor_4 g04754(new_n5130, new_n5129, new_n5131);
xor_4  g04755(new_n5131, new_n5128, new_n5132_1);
xnor_4 g04756(new_n5132_1, new_n5127, new_n5133);
xnor_4 g04757(new_n5133, new_n5124, new_n5134);
xnor_4 g04758(new_n5134, new_n5115, new_n5135);
xnor_4 g04759(new_n5135, new_n5110, new_n5136);
and_5  g04760(n11222, n1510, new_n5137);
xor_4  g04761(new_n5109, new_n5100, new_n5138);
nor_5  g04762(new_n5138, new_n5137, new_n5139);
or_5   g04763(new_n3139, new_n3138, new_n5140);
xnor_4 g04764(new_n5102, new_n5101, new_n5141);
xnor_4 g04765(new_n5141, new_n5107, new_n5142);
nor_5  g04766(new_n5142, new_n5140, new_n5143);
xnor_4 g04767(new_n5138, new_n5137, new_n5144);
nor_5  g04768(new_n5144, new_n5143, new_n5145);
or_5   g04769(new_n5145, new_n5139, new_n5146);
xor_4  g04770(new_n5146, new_n5136, new_n5147);
xor_4  g04771(new_n5144, new_n5143, new_n5148);
xor_4  g04772(new_n5071, new_n5070, new_n5149);
nor_5  g04773(new_n5149, new_n5148, new_n5150);
nand_5 g04774(new_n5149, new_n5148, new_n5151);
xor_4  g04775(new_n5069_1, new_n5067, new_n5152);
nor_5  g04776(new_n3140, new_n3127, new_n5153_1);
nor_5  g04777(new_n3144, new_n3141, new_n5154);
nor_5  g04778(new_n5154, new_n5153_1, new_n5155);
nor_5  g04779(new_n5155, new_n5152, new_n5156);
xor_4  g04780(new_n5142, new_n5140, new_n5157);
xnor_4 g04781(new_n5155, new_n5152, new_n5158);
nor_5  g04782(new_n5158, new_n5157, new_n5159);
nor_5  g04783(new_n5159, new_n5156, new_n5160);
and_5  g04784(new_n5160, new_n5151, new_n5161);
or_5   g04785(new_n5161, new_n5150, new_n5162);
xnor_4 g04786(new_n5162, new_n5147, new_n5163);
xor_4  g04787(new_n5163, new_n5074, new_n5164);
xnor_4 g04788(new_n5164, new_n5000, new_n5165);
xor_4  g04789(new_n4997, new_n4996, new_n5166);
xnor_4 g04790(new_n4995, new_n4994, new_n5167);
xor_4  g04791(new_n5158, new_n5157, new_n5168);
nor_5  g04792(new_n5168, new_n5167, new_n5169);
or_5   g04793(new_n3160, new_n3159, new_n5170);
nor_5  g04794(new_n5170, new_n3158, new_n5171);
nor_5  g04795(new_n3162, new_n3145, new_n5172);
nor_5  g04796(new_n5172, new_n5171, new_n5173);
xnor_4 g04797(new_n5168, new_n5167, new_n5174);
nor_5  g04798(new_n5174, new_n5173, new_n5175);
nor_5  g04799(new_n5175, new_n5169, new_n5176);
nor_5  g04800(new_n5176, new_n5166, new_n5177);
xnor_4 g04801(new_n5176, new_n5166, new_n5178);
xor_4  g04802(new_n5149, new_n5148, new_n5179);
xnor_4 g04803(new_n5179, new_n5160, new_n5180);
nor_5  g04804(new_n5180, new_n5178, new_n5181);
nor_5  g04805(new_n5181, new_n5177, new_n5182);
xor_4  g04806(new_n5182, new_n5165, new_n5183);
xor_4  g04807(new_n5183, new_n4926, new_n5184);
xor_4  g04808(new_n4923, new_n4922, new_n5185);
xor_4  g04809(new_n5180, new_n5178, new_n5186);
and_5  g04810(new_n5186, new_n5185, new_n5187);
nor_5  g04811(new_n5186, new_n5185, new_n5188);
xor_4  g04812(new_n4921_1, new_n4920, new_n5189);
xor_4  g04813(new_n5174, new_n5173, new_n5190);
nor_5  g04814(new_n5190, new_n5189, new_n5191_1);
nor_5  g04815(new_n3113, new_n3039, new_n5192);
nor_5  g04816(new_n3163, new_n3114, new_n5193);
nor_5  g04817(new_n5193, new_n5192, new_n5194);
xor_4  g04818(new_n5190, new_n5189, new_n5195);
and_5  g04819(new_n5195, new_n5194, new_n5196);
or_5   g04820(new_n5196, new_n5191_1, new_n5197);
nor_5  g04821(new_n5197, new_n5188, new_n5198_1);
nor_5  g04822(new_n5198_1, new_n5187, new_n5199);
xnor_4 g04823(new_n5199, new_n5184, n2301);
xor_4  g04824(new_n3111, new_n3110, n2316);
nand_5 g04825(n4634, n1333, new_n5202);
nor_5  g04826(new_n4689_1, new_n4688, new_n5203);
and_5  g04827(new_n4689_1, new_n4688, new_n5204);
nor_5  g04828(new_n5204, new_n4687, new_n5205);
or_5   g04829(new_n5205, new_n5203, new_n5206);
nor_5  g04830(new_n5206, new_n5202, new_n5207);
xnor_4 g04831(new_n5206, new_n5202, new_n5208);
and_5  g04832(n11757, n2879, new_n5209);
and_5  g04833(n7265, n5240, new_n5210);
xnor_4 g04834(new_n5210, new_n4681, new_n5211);
xor_4  g04835(new_n5211, new_n5209, new_n5212_1);
nor_5  g04836(new_n5212_1, new_n5208, new_n5213);
nor_5  g04837(new_n5213, new_n5207, new_n5214);
and_5  g04838(n4634, n3172, new_n5215);
and_5  g04839(n9195, n1333, new_n5216);
xnor_4 g04840(new_n5216, new_n5215, new_n5217);
xnor_4 g04841(new_n5217, new_n5214, new_n5218);
and_5  g04842(n11757, n10223, new_n5219);
and_5  g04843(n5240, n2879, new_n5220);
and_5  g04844(n11821, n7265, new_n5221);
xor_4  g04845(new_n5221, new_n5220, new_n5222);
xnor_4 g04846(new_n5222, new_n5219, new_n5223);
nor_5  g04847(new_n5210, new_n4681, new_n5224);
and_5  g04848(new_n5210, new_n4681, new_n5225);
nor_5  g04849(new_n5225, new_n5209, new_n5226);
nor_5  g04850(new_n5226, new_n5224, new_n5227);
xor_4  g04851(new_n5227, new_n5223, new_n5228);
xnor_4 g04852(new_n5228, new_n5218, new_n5229);
nand_5 g04853(n9195, n7862, new_n5230);
xnor_4 g04854(new_n5212_1, new_n5208, new_n5231);
nor_5  g04855(new_n5231, new_n5230, new_n5232);
nor_5  g04856(new_n4685, new_n4676, new_n5233);
nor_5  g04857(new_n4691, new_n4686_1, new_n5234);
nor_5  g04858(new_n5234, new_n5233, new_n5235);
xnor_4 g04859(new_n5231, new_n5230, new_n5236);
nor_5  g04860(new_n5236, new_n5235, new_n5237);
nor_5  g04861(new_n5237, new_n5232, new_n5238);
or_5   g04862(new_n5238, new_n5229, new_n5239);
nor_5  g04863(new_n5222, new_n5219, new_n5240_1);
nor_5  g04864(new_n5227, new_n5223, new_n5241);
nor_5  g04865(new_n5241, new_n5240_1, new_n5242);
nand_5 g04866(n2253, n1333, new_n5243);
and_5  g04867(n9195, n3172, new_n5244);
and_5  g04868(n7862, n3865, new_n5245);
xnor_4 g04869(new_n5245, new_n5244, new_n5246);
xor_4  g04870(new_n5246, new_n5243, new_n5247);
xnor_4 g04871(new_n5247, new_n5242, new_n5248);
and_5  g04872(new_n5221, new_n5220, new_n5249);
and_5  g04873(n11757, n4634, new_n5250);
xnor_4 g04874(new_n5250, new_n5249, new_n5251);
and_5  g04875(n11821, n2879, new_n5252);
and_5  g04876(n10223, n5240, new_n5253);
and_5  g04877(n9080, n7265, new_n5254);
xnor_4 g04878(new_n5254, new_n5253, new_n5255);
xnor_4 g04879(new_n5255, new_n5252, new_n5256);
xnor_4 g04880(new_n5256, new_n5251, new_n5257_1);
xor_4  g04881(new_n5257_1, new_n5248, new_n5258);
nor_5  g04882(new_n5217, new_n5214, new_n5259);
nand_5 g04883(new_n5216, new_n5215, new_n5260);
or_5   g04884(new_n5228, new_n5218, new_n5261);
xor_4  g04885(new_n5261, new_n5260, new_n5262);
nor_5  g04886(new_n5262, new_n5259, new_n5263);
xnor_4 g04887(new_n5263, new_n5258, new_n5264);
xnor_4 g04888(new_n5264, new_n5239, new_n5265);
nand_5 g04889(n7862, n2253, new_n5266);
xnor_4 g04890(new_n5238, new_n5229, new_n5267);
nor_5  g04891(new_n5267, new_n5266, new_n5268);
or_5   g04892(new_n4697, new_n4692, new_n5269);
xnor_4 g04893(new_n5236, new_n5235, new_n5270);
or_5   g04894(new_n5270, new_n5269, new_n5271);
xnor_4 g04895(new_n5267, new_n5266, new_n5272);
nor_5  g04896(new_n5272, new_n5271, new_n5273);
nor_5  g04897(new_n5273, new_n5268, new_n5274);
xor_4  g04898(new_n5274, new_n5265, new_n5275);
xor_4  g04899(new_n5272, new_n5271, new_n5276);
xnor_4 g04900(new_n5270, new_n5269, new_n5277);
or_5   g04901(new_n4720, new_n4715, new_n5278);
nand_5 g04902(n12145, n6877, new_n5279);
and_5  g04903(n9400, n2522, new_n5280);
and_5  g04904(n11311, n2024, new_n5281);
and_5  g04905(n7946, n4187, new_n5282);
xnor_4 g04906(new_n5282, new_n4710, new_n5283_1);
xnor_4 g04907(new_n5283_1, new_n5281, new_n5284);
xnor_4 g04908(new_n5284, new_n5280, new_n5285);
nor_5  g04909(new_n4702, new_n4701, new_n5286);
nor_5  g04910(new_n4703, new_n4700, new_n5287);
nor_5  g04911(new_n5287, new_n5286, new_n5288);
xor_4  g04912(new_n5288, new_n5285, new_n5289);
xnor_4 g04913(new_n5289, new_n5279, new_n5290);
nor_5  g04914(new_n4704, new_n4699, new_n5291);
nor_5  g04915(new_n4714, new_n4705, new_n5292);
nor_5  g04916(new_n5292, new_n5291, new_n5293);
xnor_4 g04917(new_n5293, new_n5290, new_n5294);
xor_4  g04918(new_n5294, new_n5278, new_n5295);
nor_5  g04919(new_n4771, new_n4721, new_n5296);
nor_5  g04920(new_n4804, new_n4772, new_n5297);
or_5   g04921(new_n5297, new_n5296, new_n5298);
xnor_4 g04922(new_n5298, new_n5295, new_n5299);
or_5   g04923(new_n4784, new_n4783, new_n5300);
and_5  g04924(n11478, n521, new_n5301);
nor_5  g04925(new_n4780, new_n4779, new_n5302);
and_5  g04926(new_n4780, new_n4779, new_n5303);
nor_5  g04927(new_n5303, new_n4778, new_n5304);
nor_5  g04928(new_n5304, new_n5302, new_n5305_1);
xnor_4 g04929(new_n5305_1, new_n5301, new_n5306);
and_5  g04930(n2498, n137, new_n5307);
and_5  g04931(n5579, n5283, new_n5308);
and_5  g04932(n6294, n2558, new_n5309);
xnor_4 g04933(new_n5309, new_n5308, new_n5310);
xor_4  g04934(new_n5310, new_n5307, new_n5311);
xor_4  g04935(new_n5311, new_n5306, new_n5312);
and_5  g04936(n6016, n4805, new_n5313);
nor_5  g04937(new_n4776, new_n4773, new_n5314_1);
nor_5  g04938(new_n4782, new_n4777, new_n5315);
or_5   g04939(new_n5315, new_n5314_1, new_n5316);
xnor_4 g04940(new_n5316, new_n5313, new_n5317);
xor_4  g04941(new_n5317, new_n5312, new_n5318);
xor_4  g04942(new_n5318, new_n5300, new_n5319_1);
or_5   g04943(new_n4798, new_n4796, new_n5320_1);
and_5  g04944(n7270, n7236, new_n5321);
nor_5  g04945(new_n4789, new_n4786, new_n5322);
and_5  g04946(new_n4795, new_n4790, new_n5323);
or_5   g04947(new_n5323, new_n5322, new_n5324);
xnor_4 g04948(new_n5324, new_n5321, new_n5325);
nand_5 g04949(n3992, n806, new_n5326);
nor_5  g04950(new_n4793, new_n4792, new_n5327);
and_5  g04951(new_n4793, new_n4792, new_n5328);
nor_5  g04952(new_n5328, new_n4791, new_n5329);
or_5   g04953(new_n5329, new_n5327, new_n5330);
xnor_4 g04954(new_n5330, new_n5326, new_n5331_1);
and_5  g04955(n9111, n6358, new_n5332);
and_5  g04956(n8384, n3342, new_n5333);
and_5  g04957(n9763, n5198, new_n5334);
xnor_4 g04958(new_n5334, new_n5333, new_n5335);
xor_4  g04959(new_n5335, new_n5332, new_n5336);
xor_4  g04960(new_n5336, new_n5331_1, new_n5337);
xor_4  g04961(new_n5337, new_n5325, new_n5338);
xor_4  g04962(new_n5338, new_n5320_1, new_n5339);
xnor_4 g04963(new_n5339, new_n5319_1, new_n5340);
nor_5  g04964(new_n4799, new_n4785, new_n5341);
nor_5  g04965(new_n4803, new_n4800, new_n5342);
nor_5  g04966(new_n5342, new_n5341, new_n5343);
xnor_4 g04967(new_n5343, new_n5340, new_n5344);
xor_4  g04968(new_n5344, new_n5299, new_n5345);
and_5  g04969(new_n5345, new_n5277, new_n5346);
xnor_4 g04970(new_n5345, new_n5277, new_n5347);
nor_5  g04971(new_n4805_1, new_n4698, new_n5348);
and_5  g04972(new_n4805_1, new_n4698, new_n5349);
nor_5  g04973(new_n4823, new_n5349, new_n5350);
nor_5  g04974(new_n5350, new_n5348, new_n5351);
nor_5  g04975(new_n5351, new_n5347, new_n5352);
nor_5  g04976(new_n5352, new_n5346, new_n5353);
nor_5  g04977(new_n5353, new_n5276, new_n5354);
nor_5  g04978(new_n5298, new_n5295, new_n5355);
nor_5  g04979(new_n5344, new_n5299, new_n5356);
or_5   g04980(new_n5356, new_n5355, new_n5357);
or_5   g04981(new_n5294, new_n5278, new_n5358);
nand_5 g04982(n12221, n6877, new_n5359);
nor_5  g04983(new_n5289, new_n5279, new_n5360);
nor_5  g04984(new_n5293, new_n5290, new_n5361);
nor_5  g04985(new_n5361, new_n5360, new_n5362);
nor_5  g04986(new_n5284, new_n5280, new_n5363);
nor_5  g04987(new_n5288, new_n5285, new_n5364);
or_5   g04988(new_n5364, new_n5363, new_n5365);
and_5  g04989(n11311, n9189, new_n5366);
and_5  g04990(n7946, n4203, new_n5367);
and_5  g04991(n4187, n2024, new_n5368);
xor_4  g04992(new_n5368, new_n5367, new_n5369);
xnor_4 g04993(new_n5369, new_n5366, new_n5370);
nor_5  g04994(new_n5282, new_n4710, new_n5371);
and_5  g04995(new_n5282, new_n4710, new_n5372);
nor_5  g04996(new_n5372, new_n5281, new_n5373);
nor_5  g04997(new_n5373, new_n5371, new_n5374);
xnor_4 g04998(new_n5374, new_n5370, new_n5375);
and_5  g04999(n12145, n9400, new_n5376);
and_5  g05000(n2522, n2464, new_n5377);
xor_4  g05001(new_n5377, new_n5376, new_n5378);
xnor_4 g05002(new_n5378, new_n5375, new_n5379);
xnor_4 g05003(new_n5379, new_n5365, new_n5380);
xnor_4 g05004(new_n5380, new_n5362, new_n5381);
xnor_4 g05005(new_n5381, new_n5359, new_n5382);
xnor_4 g05006(new_n5382, new_n5358, new_n5383);
xnor_4 g05007(new_n5383, new_n5357, new_n5384);
nor_5  g05008(new_n5338, new_n5320_1, new_n5385);
and_5  g05009(n7236, n5153, new_n5386);
nand_5 g05010(n6358, n3342, new_n5387);
and_5  g05011(n9111, n5198, new_n5388);
and_5  g05012(n9763, n1471, new_n5389);
xnor_4 g05013(new_n5389, new_n5388, new_n5390);
xnor_4 g05014(new_n5390, new_n5387, new_n5391);
nor_5  g05015(new_n5334, new_n5333, new_n5392);
nor_5  g05016(new_n5335, new_n5332, new_n5393);
or_5   g05017(new_n5393, new_n5392, new_n5394);
xnor_4 g05018(new_n5394, new_n5391, new_n5395);
and_5  g05019(n7270, n3992, new_n5396);
and_5  g05020(n8384, n806, new_n5397);
xnor_4 g05021(new_n5397, new_n5396, new_n5398);
xnor_4 g05022(new_n5398, new_n5395, new_n5399);
nor_5  g05023(new_n5330, new_n5326, new_n5400);
nor_5  g05024(new_n5336, new_n5331_1, new_n5401);
nor_5  g05025(new_n5401, new_n5400, new_n5402);
xnor_4 g05026(new_n5402, new_n5399, new_n5403);
nor_5  g05027(new_n5324, new_n5321, new_n5404);
nor_5  g05028(new_n5337, new_n5325, new_n5405);
or_5   g05029(new_n5405, new_n5404, new_n5406);
xor_4  g05030(new_n5406, new_n5403, new_n5407);
xnor_4 g05031(new_n5407, new_n5386, new_n5408);
xnor_4 g05032(new_n5408, new_n5385, new_n5409);
or_5   g05033(new_n5318, new_n5300, new_n5410);
and_5  g05034(n5798, n4805, new_n5411_1);
nand_5 g05035(n5579, n137, new_n5412);
and_5  g05036(n6797, n2558, new_n5413);
and_5  g05037(n6294, n2498, new_n5414);
xnor_4 g05038(new_n5414, new_n5413, new_n5415);
xnor_4 g05039(new_n5415, new_n5412, new_n5416);
nor_5  g05040(new_n5309, new_n5308, new_n5417);
and_5  g05041(new_n5309, new_n5308, new_n5418);
nor_5  g05042(new_n5418, new_n5307, new_n5419);
or_5   g05043(new_n5419, new_n5417, new_n5420);
xnor_4 g05044(new_n5420, new_n5416, new_n5421);
and_5  g05045(n11478, n6016, new_n5422);
and_5  g05046(n5283, n521, new_n5423);
xnor_4 g05047(new_n5423, new_n5422, new_n5424);
xnor_4 g05048(new_n5424, new_n5421, new_n5425);
and_5  g05049(new_n5305_1, new_n5301, new_n5426);
nor_5  g05050(new_n5311, new_n5306, new_n5427);
nor_5  g05051(new_n5427, new_n5426, new_n5428);
xnor_4 g05052(new_n5428, new_n5425, new_n5429);
nor_5  g05053(new_n5316, new_n5313, new_n5430);
nor_5  g05054(new_n5317, new_n5312, new_n5431);
or_5   g05055(new_n5431, new_n5430, new_n5432);
xor_4  g05056(new_n5432, new_n5429, new_n5433);
xor_4  g05057(new_n5433, new_n5411_1, new_n5434);
xnor_4 g05058(new_n5434, new_n5410, new_n5435_1);
xnor_4 g05059(new_n5435_1, new_n5409, new_n5436);
nor_5  g05060(new_n5339, new_n5319_1, new_n5437);
nor_5  g05061(new_n5343, new_n5340, new_n5438);
nor_5  g05062(new_n5438, new_n5437, new_n5439);
xor_4  g05063(new_n5439, new_n5436, new_n5440);
xnor_4 g05064(new_n5440, new_n5384, new_n5441);
xor_4  g05065(new_n5353, new_n5276, new_n5442);
and_5  g05066(new_n5442, new_n5441, new_n5443);
nor_5  g05067(new_n5443, new_n5354, new_n5444);
nor_5  g05068(new_n5444, new_n5275, new_n5445);
xnor_4 g05069(new_n5444, new_n5275, new_n5446);
or_5   g05070(new_n5380, new_n5362, new_n5447);
nor_5  g05071(new_n5369, new_n5366, new_n5448);
nor_5  g05072(new_n5374, new_n5370, new_n5449);
nor_5  g05073(new_n5449, new_n5448, new_n5450);
and_5  g05074(n12221, n9400, new_n5451);
and_5  g05075(n12145, n2464, new_n5452);
and_5  g05076(n10217, n6877, new_n5453);
xnor_4 g05077(new_n5453, new_n5452, new_n5454);
xnor_4 g05078(new_n5454, new_n5451, new_n5455);
xnor_4 g05079(new_n5455, new_n5450, new_n5456);
and_5  g05080(new_n5368, new_n5367, new_n5457);
and_5  g05081(n11311, n2522, new_n5458);
xnor_4 g05082(new_n5458, new_n5457, new_n5459);
nand_5 g05083(n4203, n2024, new_n5460);
and_5  g05084(n9189, n4187, new_n5461);
and_5  g05085(n12753, n7946, new_n5462);
xnor_4 g05086(new_n5462, new_n5461, new_n5463);
xnor_4 g05087(new_n5463, new_n5460, new_n5464);
xor_4  g05088(new_n5464, new_n5459, new_n5465);
xor_4  g05089(new_n5465, new_n5456, new_n5466);
and_5  g05090(new_n5378, new_n5375, new_n5467);
nand_5 g05091(new_n5377, new_n5376, new_n5468);
nor_5  g05092(new_n5378, new_n5375, new_n5469);
or_5   g05093(new_n5469, new_n5365, new_n5470);
xor_4  g05094(new_n5470, new_n5468, new_n5471);
nor_5  g05095(new_n5471, new_n5467, new_n5472);
xnor_4 g05096(new_n5472, new_n5466, new_n5473);
xnor_4 g05097(new_n5473, new_n5447, new_n5474);
nor_5  g05098(new_n5381, new_n5359, new_n5475);
nor_5  g05099(new_n5382, new_n5358, new_n5476);
nor_5  g05100(new_n5476, new_n5475, new_n5477);
xnor_4 g05101(new_n5477, new_n5474, new_n5478);
or_5   g05102(new_n5432, new_n5429, new_n5479);
and_5  g05103(n4805, n2347, new_n5480);
and_5  g05104(n6016, n5283, new_n5481);
and_5  g05105(n11478, n5798, new_n5482);
xnor_4 g05106(new_n5482, new_n5481, new_n5483);
xnor_4 g05107(new_n5483, new_n5480, new_n5484);
nor_5  g05108(new_n5415, new_n5412, new_n5485);
nor_5  g05109(new_n5420, new_n5416, new_n5486);
or_5   g05110(new_n5486, new_n5485, new_n5487);
xnor_4 g05111(new_n5487, new_n5484, new_n5488);
and_5  g05112(new_n5414, new_n5413, new_n5489);
and_5  g05113(n521, n137, new_n5490);
xnor_4 g05114(new_n5490, new_n5489, new_n5491);
and_5  g05115(n6797, n2498, new_n5492);
and_5  g05116(n6294, n5579, new_n5493);
and_5  g05117(n3146, n2558, new_n5494);
xnor_4 g05118(new_n5494, new_n5493, new_n5495);
xor_4  g05119(new_n5495, new_n5492, new_n5496);
xor_4  g05120(new_n5496, new_n5491, new_n5497);
xor_4  g05121(new_n5497, new_n5488, new_n5498);
nor_5  g05122(new_n5424, new_n5421, new_n5499);
nand_5 g05123(new_n5423, new_n5422, new_n5500);
or_5   g05124(new_n5428, new_n5425, new_n5501);
xor_4  g05125(new_n5501, new_n5500, new_n5502);
nor_5  g05126(new_n5502, new_n5499, new_n5503);
xnor_4 g05127(new_n5503, new_n5498, new_n5504);
xnor_4 g05128(new_n5504, new_n5479, new_n5505);
and_5  g05129(new_n5433, new_n5411_1, new_n5506);
nor_5  g05130(new_n5433, new_n5411_1, new_n5507);
nor_5  g05131(new_n5507, new_n5410, new_n5508);
nor_5  g05132(new_n5508, new_n5506, new_n5509);
xor_4  g05133(new_n5509, new_n5505, new_n5510);
nor_5  g05134(new_n5406, new_n5403, new_n5511);
nor_5  g05135(new_n5398, new_n5395, new_n5512);
nand_5 g05136(new_n5397, new_n5396, new_n5513);
or_5   g05137(new_n5402, new_n5399, new_n5514);
xor_4  g05138(new_n5514, new_n5513, new_n5515);
nor_5  g05139(new_n5515, new_n5512, new_n5516);
and_5  g05140(new_n5389, new_n5388, new_n5517);
and_5  g05141(n6358, n806, new_n5518);
xnor_4 g05142(new_n5518, new_n5517, new_n5519);
nand_5 g05143(n9111, n1471, new_n5520);
and_5  g05144(n5198, n3342, new_n5521);
and_5  g05145(n9763, n7646, new_n5522);
xnor_4 g05146(new_n5522, new_n5521, new_n5523);
xnor_4 g05147(new_n5523, new_n5520, new_n5524);
xor_4  g05148(new_n5524, new_n5519, new_n5525);
nor_5  g05149(new_n5390, new_n5387, new_n5526);
nor_5  g05150(new_n5394, new_n5391, new_n5527);
or_5   g05151(new_n5527, new_n5526, new_n5528);
and_5  g05152(n5153, n3992, new_n5529);
and_5  g05153(n8384, n7270, new_n5530);
and_5  g05154(n7236, n2507, new_n5531);
xnor_4 g05155(new_n5531, new_n5530, new_n5532);
xnor_4 g05156(new_n5532, new_n5529, new_n5533);
xnor_4 g05157(new_n5533, new_n5528, new_n5534);
xor_4  g05158(new_n5534, new_n5525, new_n5535);
xor_4  g05159(new_n5535, new_n5516, new_n5536);
xnor_4 g05160(new_n5536, new_n5511, new_n5537);
nor_5  g05161(new_n5407, new_n5386, new_n5538);
and_5  g05162(new_n5407, new_n5386, new_n5539);
nor_5  g05163(new_n5539, new_n5385, new_n5540);
or_5   g05164(new_n5540, new_n5538, new_n5541);
xor_4  g05165(new_n5541, new_n5537, new_n5542);
xnor_4 g05166(new_n5542, new_n5510, new_n5543);
nor_5  g05167(new_n5435_1, new_n5409, new_n5544);
nor_5  g05168(new_n5439, new_n5436, new_n5545);
nor_5  g05169(new_n5545, new_n5544, new_n5546);
xor_4  g05170(new_n5546, new_n5543, new_n5547);
xnor_4 g05171(new_n5547, new_n5478, new_n5548);
nor_5  g05172(new_n5383, new_n5357, new_n5549);
nor_5  g05173(new_n5440, new_n5384, new_n5550);
nor_5  g05174(new_n5550, new_n5549, new_n5551);
xor_4  g05175(new_n5551, new_n5548, new_n5552);
nor_5  g05176(new_n5552, new_n5446, new_n5553);
nor_5  g05177(new_n5553, new_n5445, new_n5554);
nor_5  g05178(new_n5547, new_n5478, new_n5555);
nor_5  g05179(new_n5551, new_n5548, new_n5556);
nor_5  g05180(new_n5556, new_n5555, new_n5557);
and_5  g05181(n4805, n1576, new_n5558);
nor_5  g05182(new_n5501, new_n5500, new_n5559);
nor_5  g05183(new_n5503, new_n5498, new_n5560);
nor_5  g05184(new_n5560, new_n5559, new_n5561);
xnor_4 g05185(new_n5561, new_n5558, new_n5562);
xnor_4 g05186(new_n5562, new_n5557, new_n5563);
nor_5  g05187(new_n5473, new_n5447, new_n5564);
nor_5  g05188(new_n5477, new_n5474, new_n5565);
or_5   g05189(new_n5565, new_n5564, new_n5566);
and_5  g05190(new_n5536, new_n5511, new_n5567);
nor_5  g05191(new_n5541, new_n5537, new_n5568);
nor_5  g05192(new_n5568, new_n5567, new_n5569);
nor_5  g05193(new_n5455, new_n5450, new_n5570);
nor_5  g05194(new_n5465, new_n5456, new_n5571);
nor_5  g05195(new_n5571, new_n5570, new_n5572);
and_5  g05196(n9189, n4203, new_n5573);
and_5  g05197(n4187, n2522, new_n5574);
xnor_4 g05198(new_n5574, new_n5573, new_n5575);
and_5  g05199(n9763, n4722, new_n5576);
and_5  g05200(n10217, n9400, new_n5577);
xnor_4 g05201(new_n5577, new_n5576, new_n5578);
xnor_4 g05202(new_n5578, new_n5575, new_n5579_1);
nand_5 g05203(n9111, n7646, new_n5580);
and_5  g05204(n12221, n2464, new_n5581);
and_5  g05205(n12145, n11311, new_n5582);
xnor_4 g05206(new_n5582, new_n5581, new_n5583);
xnor_4 g05207(new_n5583, new_n5580, new_n5584);
xnor_4 g05208(new_n5584, new_n5579_1, new_n5585);
xnor_4 g05209(new_n5585, new_n5572, new_n5586);
xnor_4 g05210(new_n5586, new_n5569, new_n5587);
xnor_4 g05211(new_n5587, new_n5566, new_n5588);
nor_5  g05212(new_n5470, new_n5468, new_n5589);
nor_5  g05213(new_n5472, new_n5466, new_n5590);
or_5   g05214(new_n5590, new_n5589, new_n5591);
nor_5  g05215(new_n5514, new_n5513, new_n5592);
nor_5  g05216(new_n5535, new_n5516, new_n5593);
nor_5  g05217(new_n5593, new_n5592, new_n5594);
xnor_4 g05218(new_n5594, new_n5591, new_n5595);
and_5  g05219(n11821, n10223, new_n5596);
and_5  g05220(n9080, n2879, new_n5597);
xnor_4 g05221(new_n5597, new_n5596, new_n5598);
and_5  g05222(n11757, n9195, new_n5599);
and_5  g05223(n7862, n2512, new_n5600);
xnor_4 g05224(new_n5600, new_n5599, new_n5601);
xor_4  g05225(new_n5601, new_n5598, new_n5602);
and_5  g05226(new_n5245, new_n5244, new_n5603);
nor_5  g05227(new_n5245, new_n5244, new_n5604);
nor_5  g05228(new_n5604, new_n5243, new_n5605);
nor_5  g05229(new_n5605, new_n5603, new_n5606);
xnor_4 g05230(new_n5606, new_n5602, new_n5607);
and_5  g05231(n12753, n2024, new_n5608);
and_5  g05232(n3865, n1333, new_n5609);
and_5  g05233(n5240, n4634, new_n5610);
xnor_4 g05234(new_n5610, new_n5609, new_n5611);
xnor_4 g05235(new_n5611, new_n5608, new_n5612);
xnor_4 g05236(new_n5612, new_n5607, new_n5613);
xnor_4 g05237(new_n5613, new_n5595, new_n5614);
nor_5  g05238(new_n5261, new_n5260, new_n5615);
nor_5  g05239(new_n5263, new_n5258, new_n5616);
nor_5  g05240(new_n5616, new_n5615, new_n5617);
nor_5  g05241(new_n5247, new_n5242, new_n5618);
nor_5  g05242(new_n5257_1, new_n5248, new_n5619);
nor_5  g05243(new_n5619, new_n5618, new_n5620);
and_5  g05244(new_n5458, new_n5457, new_n5621);
nor_5  g05245(new_n5464, new_n5459, new_n5622);
nor_5  g05246(new_n5622, new_n5621, new_n5623);
and_5  g05247(n8384, n5153, new_n5624);
and_5  g05248(n7270, n6358, new_n5625);
xnor_4 g05249(new_n5625, new_n5624, new_n5626);
and_5  g05250(new_n5462, new_n5461, new_n5627);
nor_5  g05251(new_n5462, new_n5461, new_n5628);
nor_5  g05252(new_n5628, new_n5460, new_n5629);
nor_5  g05253(new_n5629, new_n5627, new_n5630);
xnor_4 g05254(new_n5630, new_n5626, new_n5631);
xnor_4 g05255(new_n5631, new_n5623, new_n5632);
xnor_4 g05256(new_n5632, new_n5620, new_n5633);
and_5  g05257(n5198, n806, new_n5634);
and_5  g05258(n3992, n2507, new_n5635);
xnor_4 g05259(new_n5635, new_n5634, new_n5636);
and_5  g05260(n7823, n6877, new_n5637);
and_5  g05261(n3342, n1471, new_n5638);
xnor_4 g05262(new_n5638, new_n5637, new_n5639);
xor_4  g05263(new_n5639, new_n5636, new_n5640);
and_5  g05264(new_n5522, new_n5521, new_n5641_1);
nor_5  g05265(new_n5522, new_n5521, new_n5642);
nor_5  g05266(new_n5642, new_n5520, new_n5643);
nor_5  g05267(new_n5643, new_n5641_1, new_n5644);
xnor_4 g05268(new_n5644, new_n5640, new_n5645_1);
xnor_4 g05269(new_n5645_1, new_n5633, new_n5646);
nor_5  g05270(new_n5533, new_n5528, new_n5647);
nor_5  g05271(new_n5534, new_n5525, new_n5648);
nor_5  g05272(new_n5648, new_n5647, new_n5649);
nor_5  g05273(new_n5453, new_n5452, new_n5650);
nor_5  g05274(new_n5454, new_n5451, new_n5651);
nor_5  g05275(new_n5651, new_n5650, new_n5652);
and_5  g05276(n7236, n6431, new_n5653);
and_5  g05277(n10174, n7946, new_n5654);
xor_4  g05278(new_n5654, new_n5653, new_n5655);
xnor_4 g05279(new_n5655, new_n5652, new_n5656);
xnor_4 g05280(new_n5656, new_n5649, new_n5657);
xnor_4 g05281(new_n5657, new_n5646, new_n5658);
xnor_4 g05282(new_n5658, new_n5617, new_n5659);
xnor_4 g05283(new_n5659, new_n5614, new_n5660);
xnor_4 g05284(new_n5660, new_n5588, new_n5661);
nor_5  g05285(new_n5542, new_n5510, new_n5662);
nor_5  g05286(new_n5546, new_n5543, new_n5663);
nor_5  g05287(new_n5663, new_n5662, new_n5664);
nor_5  g05288(new_n5264, new_n5239, new_n5665);
nor_5  g05289(new_n5274, new_n5265, new_n5666);
nor_5  g05290(new_n5666, new_n5665, new_n5667);
nor_5  g05291(new_n5504, new_n5479, new_n5668);
nor_5  g05292(new_n5509, new_n5505, new_n5669);
nor_5  g05293(new_n5669, new_n5668, new_n5670_1);
and_5  g05294(new_n5518, new_n5517, new_n5671);
nor_5  g05295(new_n5524, new_n5519, new_n5672);
nor_5  g05296(new_n5672, new_n5671, new_n5673);
and_5  g05297(new_n5490, new_n5489, new_n5674);
nor_5  g05298(new_n5496, new_n5491, new_n5675);
nor_5  g05299(new_n5675, new_n5674, new_n5676);
xor_4  g05300(new_n5676, new_n5673, new_n5677);
nor_5  g05301(new_n5250, new_n5249, new_n5678);
nor_5  g05302(new_n5256, new_n5251, new_n5679);
nor_5  g05303(new_n5679, new_n5678, new_n5680);
and_5  g05304(n3172, n2253, new_n5681);
and_5  g05305(n6797, n5579, new_n5682);
and_5  g05306(n5798, n5283, new_n5683);
xnor_4 g05307(new_n5683, new_n5682, new_n5684);
xnor_4 g05308(new_n5684, new_n5681, new_n5685);
xnor_4 g05309(new_n5685, new_n5680, new_n5686);
nor_5  g05310(new_n5482, new_n5481, new_n5687);
nor_5  g05311(new_n5483, new_n5480, new_n5688);
nor_5  g05312(new_n5688, new_n5687, new_n5689);
nor_5  g05313(new_n5494, new_n5493, new_n5690);
nor_5  g05314(new_n5495, new_n5492, new_n5691);
nor_5  g05315(new_n5691, new_n5690, new_n5692);
xnor_4 g05316(new_n5692, new_n5689, new_n5693_1);
and_5  g05317(n11478, n2347, new_n5694_1);
and_5  g05318(n3146, n2498, new_n5695);
xnor_4 g05319(new_n5695, new_n5694_1, new_n5696);
xnor_4 g05320(new_n5696, new_n5693_1, new_n5697);
xnor_4 g05321(new_n5697, new_n5686, new_n5698);
xnor_4 g05322(new_n5698, new_n5677, new_n5699);
nor_5  g05323(new_n5487, new_n5484, new_n5700);
nor_5  g05324(new_n5497, new_n5488, new_n5701);
nor_5  g05325(new_n5701, new_n5700, new_n5702);
nor_5  g05326(new_n5254, new_n5253, new_n5703);
nor_5  g05327(new_n5255, new_n5252, new_n5704);
nor_5  g05328(new_n5704, new_n5703, new_n5705);
and_5  g05329(n6016, n137, new_n5706);
and_5  g05330(n7265, n6826, new_n5707);
and_5  g05331(n6294, n521, new_n5708);
xnor_4 g05332(new_n5708, new_n5707, new_n5709);
xnor_4 g05333(new_n5709, new_n5706, new_n5710);
xnor_4 g05334(new_n5710, new_n5705, new_n5711);
and_5  g05335(n4938, n2558, new_n5712);
nor_5  g05336(new_n5531, new_n5530, new_n5713);
nor_5  g05337(new_n5532, new_n5529, new_n5714);
nor_5  g05338(new_n5714, new_n5713, new_n5715);
xnor_4 g05339(new_n5715, new_n5712, new_n5716);
xnor_4 g05340(new_n5716, new_n5711, new_n5717);
xnor_4 g05341(new_n5717, new_n5702, new_n5718);
xnor_4 g05342(new_n5718, new_n5699, new_n5719);
xnor_4 g05343(new_n5719, new_n5670_1, new_n5720);
xnor_4 g05344(new_n5720, new_n5667, new_n5721);
xnor_4 g05345(new_n5721, new_n5664, new_n5722);
xnor_4 g05346(new_n5722, new_n5661, new_n5723);
xnor_4 g05347(new_n5723, new_n5563, new_n5724);
xnor_4 g05348(new_n5724, new_n5554, n2383);
xnor_4 g05349(new_n4669, new_n4662, n2425);
xor_4  g05350(new_n2347_1, new_n2310, n2431);
xnor_4 g05351(new_n1670, new_n1669, n2434);
xnor_4 g05352(new_n3905, new_n3904, n2581);
xor_4  g05353(new_n5186, new_n5185, new_n5730);
xnor_4 g05354(new_n5730, new_n5197, n2624);
and_5  g05355(n11917, n6770, new_n5732);
and_5  g05356(n9920, n4921, new_n5733);
and_5  g05357(n9956, n3627, new_n5734);
xor_4  g05358(new_n5734, new_n5733, new_n5735);
xnor_4 g05359(new_n5735, new_n5732, new_n5736);
nor_5  g05360(new_n3200, new_n3170, new_n5737);
nor_5  g05361(new_n3201, new_n3199, new_n5738);
nor_5  g05362(new_n5738, new_n5737, new_n5739);
xor_4  g05363(new_n5739, new_n5736, new_n5740);
and_5  g05364(n2577, n2564, new_n5741);
and_5  g05365(n4189, n3842, new_n5742);
xnor_4 g05366(new_n5742, new_n5741, new_n5743);
xnor_4 g05367(new_n5743, new_n5740, new_n5744);
nor_5  g05368(new_n3197, new_n3193, new_n5745);
nor_5  g05369(new_n3202, new_n3198, new_n5746);
nor_5  g05370(new_n5746, new_n5745, new_n5747);
xnor_4 g05371(new_n5747, new_n5744, new_n5748);
nor_5  g05372(new_n3191, new_n3188, new_n5749);
nor_5  g05373(new_n3203, new_n3192, new_n5750);
nor_5  g05374(new_n5750, new_n5749, new_n5751);
nor_5  g05375(new_n5751, new_n5748, new_n5752);
and_5  g05376(new_n5734, new_n5733, new_n5753);
and_5  g05377(n6770, n3842, new_n5754);
xnor_4 g05378(new_n5754, new_n5753, new_n5755);
and_5  g05379(n4921, n3627, new_n5756);
and_5  g05380(n11917, n9920, new_n5757);
and_5  g05381(n9956, n4516, new_n5758);
xnor_4 g05382(new_n5758, new_n5757, new_n5759);
xnor_4 g05383(new_n5759, new_n5756, new_n5760_1);
xor_4  g05384(new_n5760_1, new_n5755, new_n5761);
nor_5  g05385(new_n5735, new_n5732, new_n5762);
nor_5  g05386(new_n5739, new_n5736, new_n5763);
or_5   g05387(new_n5763, new_n5762, new_n5764);
and_5  g05388(n9637, n2564, new_n5765);
and_5  g05389(n4189, n2577, new_n5766);
and_5  g05390(n6687, n1835, new_n5767_1);
xnor_4 g05391(new_n5767_1, new_n5766, new_n5768);
xor_4  g05392(new_n5768, new_n5765, new_n5769);
xnor_4 g05393(new_n5769, new_n5764, new_n5770);
xnor_4 g05394(new_n5770, new_n5761, new_n5771);
nor_5  g05395(new_n5743, new_n5740, new_n5772);
nand_5 g05396(new_n5742, new_n5741, new_n5773);
or_5   g05397(new_n5747, new_n5744, new_n5774);
xor_4  g05398(new_n5774, new_n5773, new_n5775);
nor_5  g05399(new_n5775, new_n5772, new_n5776);
xor_4  g05400(new_n5776, new_n5771, new_n5777);
xnor_4 g05401(new_n5777, new_n5752, new_n5778);
nand_5 g05402(n9637, n6687, new_n5779);
xnor_4 g05403(new_n5751, new_n5748, new_n5780);
nor_5  g05404(new_n5780, new_n5779, new_n5781);
or_5   g05405(new_n3204, new_n3187, new_n5782);
xnor_4 g05406(new_n5780, new_n5779, new_n5783);
nor_5  g05407(new_n5783, new_n5782, new_n5784);
nor_5  g05408(new_n5784, new_n5781, new_n5785);
xnor_4 g05409(new_n5785, new_n5778, new_n5786);
and_5  g05410(n6126, n2226, new_n5787);
and_5  g05411(n3602, n1094, new_n5788);
and_5  g05412(n10678, n3719, new_n5789);
xor_4  g05413(new_n5789, new_n5788, new_n5790);
xnor_4 g05414(new_n5790, new_n5787, new_n5791);
nor_5  g05415(new_n3355, new_n3212, new_n5792);
nor_5  g05416(new_n3356, new_n3354, new_n5793);
nor_5  g05417(new_n5793, new_n5792, new_n5794);
xor_4  g05418(new_n5794, new_n5791, new_n5795);
and_5  g05419(n10928, n10439, new_n5796);
and_5  g05420(n8595, n6986, new_n5797);
xnor_4 g05421(new_n5797, new_n5796, new_n5798_1);
xnor_4 g05422(new_n5798_1, new_n5795, new_n5799);
nor_5  g05423(new_n3352, new_n3348, new_n5800);
nor_5  g05424(new_n3357, new_n3353, new_n5801);
nor_5  g05425(new_n5801, new_n5800, new_n5802);
xnor_4 g05426(new_n5802, new_n5799, new_n5803);
nor_5  g05427(new_n3346, new_n3343, new_n5804);
nor_5  g05428(new_n3358, new_n3347, new_n5805);
nor_5  g05429(new_n5805, new_n5804, new_n5806);
or_5   g05430(new_n5806, new_n5803, new_n5807);
nor_5  g05431(new_n5790, new_n5787, new_n5808);
nor_5  g05432(new_n5794, new_n5791, new_n5809);
nor_5  g05433(new_n5809, new_n5808, new_n5810);
and_5  g05434(n10928, n8065, new_n5811);
and_5  g05435(n10439, n6986, new_n5812);
and_5  g05436(n10391, n8336, new_n5813);
xnor_4 g05437(new_n5813, new_n5812, new_n5814_1);
xnor_4 g05438(new_n5814_1, new_n5811, new_n5815);
xnor_4 g05439(new_n5815, new_n5810, new_n5816);
and_5  g05440(new_n5789, new_n5788, new_n5817);
and_5  g05441(n8595, n2226, new_n5818);
xnor_4 g05442(new_n5818, new_n5817, new_n5819);
and_5  g05443(n10678, n3602, new_n5820);
and_5  g05444(n6126, n1094, new_n5821);
and_5  g05445(n7320, n3719, new_n5822);
xnor_4 g05446(new_n5822, new_n5821, new_n5823);
xor_4  g05447(new_n5823, new_n5820, new_n5824);
xor_4  g05448(new_n5824, new_n5819, new_n5825);
xor_4  g05449(new_n5825, new_n5816, new_n5826);
nor_5  g05450(new_n5798_1, new_n5795, new_n5827);
nand_5 g05451(new_n5797, new_n5796, new_n5828);
or_5   g05452(new_n5802, new_n5799, new_n5829);
xor_4  g05453(new_n5829, new_n5828, new_n5830);
nor_5  g05454(new_n5830, new_n5827, new_n5831);
xnor_4 g05455(new_n5831, new_n5826, new_n5832);
xnor_4 g05456(new_n5832, new_n5807, new_n5833);
and_5  g05457(n8336, n8065, new_n5834);
xor_4  g05458(new_n5806, new_n5803, new_n5835);
nor_5  g05459(new_n5835, new_n5834, new_n5836);
nor_5  g05460(new_n3359, new_n3342_1, new_n5837);
xnor_4 g05461(new_n5835, new_n5834, new_n5838);
nor_5  g05462(new_n5838, new_n5837, new_n5839);
or_5   g05463(new_n5839, new_n5836, new_n5840);
xor_4  g05464(new_n5840, new_n5833, new_n5841);
nand_5 g05465(n7160, n4826, new_n5842);
and_5  g05466(n7733, n4828, new_n5843);
and_5  g05467(n12925, n2515, new_n5844);
xnor_4 g05468(new_n5844, new_n5843, new_n5845);
xnor_4 g05469(new_n5845, new_n5842, new_n5846);
nor_5  g05470(new_n3389, new_n3235, new_n5847);
nor_5  g05471(new_n3390, new_n3388, new_n5848);
or_5   g05472(new_n5848, new_n5847, new_n5849);
xnor_4 g05473(new_n5849, new_n5846, new_n5850);
and_5  g05474(n12391, n4970, new_n5851);
and_5  g05475(n7891, n7610, new_n5852);
xnor_4 g05476(new_n5852, new_n5851, new_n5853);
xnor_4 g05477(new_n5853, new_n5850, new_n5854);
and_5  g05478(new_n3386, new_n3383, new_n5855);
nor_5  g05479(new_n3391, new_n3387, new_n5856);
nor_5  g05480(new_n5856, new_n5855, new_n5857_1);
xnor_4 g05481(new_n5857_1, new_n5854, new_n5858);
nor_5  g05482(new_n3392, new_n3382, new_n5859);
nor_5  g05483(new_n3396, new_n3393, new_n5860_1);
nor_5  g05484(new_n5860_1, new_n5859, new_n5861);
or_5   g05485(new_n5861, new_n5858, new_n5862);
nor_5  g05486(new_n5845, new_n5842, new_n5863);
nor_5  g05487(new_n5849, new_n5846, new_n5864);
or_5   g05488(new_n5864, new_n5863, new_n5865);
and_5  g05489(n12391, n503, new_n5866);
and_5  g05490(n7891, n4970, new_n5867);
and_5  g05491(n12069, n10965, new_n5868);
xnor_4 g05492(new_n5868, new_n5867, new_n5869);
xnor_4 g05493(new_n5869, new_n5866, new_n5870);
xnor_4 g05494(new_n5870, new_n5865, new_n5871);
and_5  g05495(new_n5844, new_n5843, new_n5872);
and_5  g05496(n7610, n7160, new_n5873);
xnor_4 g05497(new_n5873, new_n5872, new_n5874);
and_5  g05498(n7733, n2515, new_n5875);
and_5  g05499(n4828, n4826, new_n5876);
and_5  g05500(n12925, n1199, new_n5877);
xnor_4 g05501(new_n5877, new_n5876, new_n5878);
xor_4  g05502(new_n5878, new_n5875, new_n5879);
xor_4  g05503(new_n5879, new_n5874, new_n5880);
xor_4  g05504(new_n5880, new_n5871, new_n5881);
nor_5  g05505(new_n5853, new_n5850, new_n5882);
nand_5 g05506(new_n5852, new_n5851, new_n5883);
or_5   g05507(new_n5857_1, new_n5854, new_n5884);
xor_4  g05508(new_n5884, new_n5883, new_n5885);
nor_5  g05509(new_n5885, new_n5882, new_n5886);
xnor_4 g05510(new_n5886, new_n5881, new_n5887);
xnor_4 g05511(new_n5887, new_n5862, new_n5888);
nand_5 g05512(n12069, n503, new_n5889);
xnor_4 g05513(new_n5861, new_n5858, new_n5890);
nor_5  g05514(new_n5890, new_n5889, new_n5891);
or_5   g05515(new_n3397, new_n3381, new_n5892);
xnor_4 g05516(new_n5890, new_n5889, new_n5893);
nor_5  g05517(new_n5893, new_n5892, new_n5894);
nor_5  g05518(new_n5894, new_n5891, new_n5895);
xor_4  g05519(new_n5895, new_n5888, new_n5896);
and_5  g05520(n11222, n6359, new_n5897);
nand_5 g05521(n4086, n996, new_n5898);
and_5  g05522(n5767, n405, new_n5899);
and_5  g05523(n8433, n5319, new_n5900);
xnor_4 g05524(new_n5900, new_n5899, new_n5901);
xnor_4 g05525(new_n5901, new_n5898, new_n5902);
nor_5  g05526(new_n3366, new_n3365, new_n5903);
and_5  g05527(new_n3366, new_n3365, new_n5904);
nor_5  g05528(new_n5904, new_n3364, new_n5905);
or_5   g05529(new_n5905, new_n5903, new_n5906);
xnor_4 g05530(new_n5906, new_n5902, new_n5907);
and_5  g05531(n11153, n6611, new_n5908);
and_5  g05532(n5314, n217, new_n5909);
xnor_4 g05533(new_n5909, new_n5908, new_n5910);
xnor_4 g05534(new_n5910, new_n5907, new_n5911);
nor_5  g05535(new_n3368, new_n3363, new_n5912);
nor_5  g05536(new_n3373, new_n3369, new_n5913);
nor_5  g05537(new_n5913, new_n5912, new_n5914);
xnor_4 g05538(new_n5914, new_n5911, new_n5915);
and_5  g05539(new_n3374, new_n3362, new_n5916);
nor_5  g05540(new_n3378, new_n3375, new_n5917);
nor_5  g05541(new_n5917, new_n5916, new_n5918);
xor_4  g05542(new_n5918, new_n5915, new_n5919);
and_5  g05543(new_n5919, new_n5897, new_n5920);
or_5   g05544(new_n3379, new_n3361, new_n5921);
xnor_4 g05545(new_n5919, new_n5897, new_n5922);
nor_5  g05546(new_n5922, new_n5921, new_n5923);
nor_5  g05547(new_n5923, new_n5920, new_n5924);
or_5   g05548(new_n5918, new_n5915, new_n5925);
and_5  g05549(new_n5900, new_n5899, new_n5926);
and_5  g05550(n996, n217, new_n5927);
xnor_4 g05551(new_n5927, new_n5926, new_n5928);
and_5  g05552(n5319, n405, new_n5929);
and_5  g05553(n5767, n4086, new_n5930);
and_5  g05554(n9457, n8433, new_n5931);
xnor_4 g05555(new_n5931, new_n5930, new_n5932);
xor_4  g05556(new_n5932, new_n5929, new_n5933);
xor_4  g05557(new_n5933, new_n5928, new_n5934_1);
and_5  g05558(n11153, n6359, new_n5935);
nand_5 g05559(n6611, n5314, new_n5936);
nand_5 g05560(n11296, n11222, new_n5937);
xnor_4 g05561(new_n5937, new_n5936, new_n5938);
xnor_4 g05562(new_n5938, new_n5935, new_n5939);
nor_5  g05563(new_n5901, new_n5898, new_n5940);
nor_5  g05564(new_n5906, new_n5902, new_n5941);
or_5   g05565(new_n5941, new_n5940, new_n5942);
xnor_4 g05566(new_n5942, new_n5939, new_n5943);
xor_4  g05567(new_n5943, new_n5934_1, new_n5944);
nor_5  g05568(new_n5910, new_n5907, new_n5945);
nand_5 g05569(new_n5909, new_n5908, new_n5946);
or_5   g05570(new_n5914, new_n5911, new_n5947);
xor_4  g05571(new_n5947, new_n5946, new_n5948);
nor_5  g05572(new_n5948, new_n5945, new_n5949);
xnor_4 g05573(new_n5949, new_n5944, new_n5950);
xnor_4 g05574(new_n5950, new_n5925, new_n5951);
xor_4  g05575(new_n5951, new_n5924, new_n5952);
xnor_4 g05576(new_n5952, new_n5896, new_n5953);
xor_4  g05577(new_n5893, new_n5892, new_n5954);
xor_4  g05578(new_n5922, new_n5921, new_n5955);
nor_5  g05579(new_n5955, new_n5954, new_n5956);
nor_5  g05580(new_n3401, new_n3398, new_n5957);
nor_5  g05581(new_n3402, new_n3380, new_n5958);
nor_5  g05582(new_n5958, new_n5957, new_n5959);
xnor_4 g05583(new_n5955, new_n5954, new_n5960);
nor_5  g05584(new_n5960, new_n5959, new_n5961);
nor_5  g05585(new_n5961, new_n5956, new_n5962);
xnor_4 g05586(new_n5962, new_n5953, new_n5963);
xnor_4 g05587(new_n5963, new_n5841, new_n5964_1);
xnor_4 g05588(new_n5838, new_n5837, new_n5965);
xnor_4 g05589(new_n5960, new_n5959, new_n5966);
nor_5  g05590(new_n5966, new_n5965, new_n5967);
xnor_4 g05591(new_n5966, new_n5965, new_n5968);
nor_5  g05592(new_n3403, new_n3360, new_n5969);
nor_5  g05593(new_n3407, new_n3404, new_n5970);
or_5   g05594(new_n5970, new_n5969, new_n5971);
nor_5  g05595(new_n5971, new_n5968, new_n5972);
nor_5  g05596(new_n5972, new_n5967, new_n5973);
xor_4  g05597(new_n5973, new_n5964_1, new_n5974);
nor_5  g05598(new_n5974, new_n5786, new_n5975);
xor_4  g05599(new_n5783, new_n5782, new_n5976);
and_5  g05600(new_n3340, new_n3205, new_n5977);
nor_5  g05601(new_n3408, new_n3341, new_n5978);
or_5   g05602(new_n5978, new_n5977, new_n5979);
nor_5  g05603(new_n5979, new_n5976, new_n5980);
xor_4  g05604(new_n5971, new_n5968, new_n5981);
xor_4  g05605(new_n5979, new_n5976, new_n5982);
and_5  g05606(new_n5982, new_n5981, new_n5983);
or_5   g05607(new_n5983, new_n5980, new_n5984);
xnor_4 g05608(new_n5974, new_n5786, new_n5985);
nor_5  g05609(new_n5985, new_n5984, new_n5986);
nor_5  g05610(new_n5986, new_n5975, new_n5987);
nor_5  g05611(new_n5884, new_n5883, new_n5988);
nor_5  g05612(new_n5886, new_n5881, new_n5989);
nor_5  g05613(new_n5989, new_n5988, new_n5990);
and_5  g05614(new_n5873, new_n5872, new_n5991);
nor_5  g05615(new_n5879, new_n5874, new_n5992);
nor_5  g05616(new_n5992, new_n5991, new_n5993);
nor_5  g05617(new_n5767_1, new_n5766, new_n5994);
nor_5  g05618(new_n5768, new_n5765, new_n5995);
nor_5  g05619(new_n5995, new_n5994, new_n5996);
and_5  g05620(n6770, n2577, new_n5997);
xnor_4 g05621(new_n5997, new_n5996, new_n5998);
and_5  g05622(n9637, n4189, new_n5999);
and_5  g05623(n11917, n3627, new_n6000);
xnor_4 g05624(new_n6000, new_n5999, new_n6001);
xnor_4 g05625(new_n6001, new_n5998, new_n6002);
nor_5  g05626(new_n5868, new_n5867, new_n6003);
nor_5  g05627(new_n5869, new_n5866, new_n6004);
or_5   g05628(new_n6004, new_n6003, new_n6005);
nor_5  g05629(new_n5754, new_n5753, new_n6006);
nor_5  g05630(new_n5760_1, new_n5755, new_n6007);
nor_5  g05631(new_n6007, new_n6006, new_n6008);
xnor_4 g05632(new_n6008, new_n6005, new_n6009);
xnor_4 g05633(new_n6009, new_n6002, new_n6010);
xnor_4 g05634(new_n6010, new_n5993, new_n6011);
nor_5  g05635(new_n5870, new_n5865, new_n6012);
nor_5  g05636(new_n5880, new_n5871, new_n6013);
nor_5  g05637(new_n6013, new_n6012, new_n6014);
nor_5  g05638(new_n5822, new_n5821, new_n6015);
nor_5  g05639(new_n5823, new_n5820, new_n6016_1);
nor_5  g05640(new_n6016_1, new_n6015, new_n6017);
and_5  g05641(n7523, n3719, new_n6018);
and_5  g05642(n11222, n1357, new_n6019);
xnor_4 g05643(new_n6019, new_n6018, new_n6020);
and_5  g05644(n8336, n4190, new_n6021);
and_5  g05645(n7320, n3602, new_n6022);
xnor_4 g05646(new_n6022, new_n6021, new_n6023);
xor_4  g05647(new_n6023, new_n6020, new_n6024);
xnor_4 g05648(new_n6024, new_n6017, new_n6025);
xnor_4 g05649(new_n6025, new_n6014, new_n6026);
xnor_4 g05650(new_n6026, new_n6011, new_n6027);
nor_5  g05651(new_n5774, new_n5773, new_n6028);
nor_5  g05652(new_n5776, new_n5771, new_n6029);
nor_5  g05653(new_n6029, new_n6028, new_n6030);
nor_5  g05654(new_n5829, new_n5828, new_n6031);
nor_5  g05655(new_n5831, new_n5826, new_n6032);
nor_5  g05656(new_n6032, new_n6031, new_n6033);
xnor_4 g05657(new_n6033, new_n6030, new_n6034);
xnor_4 g05658(new_n6034, new_n6027, new_n6035);
xnor_4 g05659(new_n6035, new_n5990, new_n6036);
nor_5  g05660(new_n5832, new_n5807, new_n6037);
nor_5  g05661(new_n5840, new_n5833, new_n6038_1);
nor_5  g05662(new_n6038_1, new_n6037, new_n6039);
nor_5  g05663(new_n5813, new_n5812, new_n6040);
nor_5  g05664(new_n5814_1, new_n5811, new_n6041);
nor_5  g05665(new_n6041, new_n6040, new_n6042);
and_5  g05666(n5319, n4086, new_n6043);
and_5  g05667(n10928, n10391, new_n6044);
xor_4  g05668(new_n6044, new_n6043, new_n6045);
xnor_4 g05669(new_n6045, new_n6042, new_n6046);
xnor_4 g05670(new_n6046, new_n6039, new_n6047);
xnor_4 g05671(new_n6047, new_n6036, new_n6048);
nor_5  g05672(new_n5887, new_n5862, new_n6049);
nor_5  g05673(new_n5895, new_n5888, new_n6050);
or_5   g05674(new_n6050, new_n6049, new_n6051);
nor_5  g05675(new_n5950, new_n5925, new_n6052);
nor_5  g05676(new_n5951, new_n5924, new_n6053);
nor_5  g05677(new_n6053, new_n6052, new_n6054);
xnor_4 g05678(new_n6054, new_n6051, new_n6055);
xnor_4 g05679(new_n6055, new_n6048, new_n6056);
and_5  g05680(n4826, n2515, new_n6057);
and_5  g05681(n12925, n6578, new_n6058);
xnor_4 g05682(new_n6058, new_n6057, new_n6059);
and_5  g05683(n6359, n5314, new_n6060);
and_5  g05684(n12069, n7546, new_n6061);
xnor_4 g05685(new_n6061, new_n6060, new_n6062);
xor_4  g05686(new_n6062, new_n6059, new_n6063);
nor_5  g05687(new_n5931, new_n5930, new_n6064);
nor_5  g05688(new_n5932, new_n5929, new_n6065);
or_5   g05689(new_n6065, new_n6064, new_n6066);
nor_5  g05690(new_n5938, new_n5935, new_n6067);
or_5   g05691(new_n6067, new_n5936, new_n6068);
nand_5 g05692(n11296, n11153, new_n6069);
nor_5  g05693(new_n6069, new_n6068, new_n6070);
or_5   g05694(new_n6069, new_n5897, new_n6071);
and_5  g05695(new_n6071, new_n6068, new_n6072);
nor_5  g05696(new_n6072, new_n6070, new_n6073);
xnor_4 g05697(new_n6073, new_n6066, new_n6074);
xnor_4 g05698(new_n6074, new_n6063, new_n6075);
xnor_4 g05699(new_n6075, new_n6056, new_n6076);
nor_5  g05700(new_n5963, new_n5841, new_n6077);
nor_5  g05701(new_n5973, new_n5964_1, new_n6078);
nor_5  g05702(new_n6078, new_n6077, new_n6079);
nor_5  g05703(new_n5952, new_n5896, new_n6080);
nor_5  g05704(new_n5962, new_n5953, new_n6081);
nor_5  g05705(new_n6081, new_n6080, new_n6082);
and_5  g05706(new_n5777, new_n5752, new_n6083);
nor_5  g05707(new_n5785, new_n5778, new_n6084);
nor_5  g05708(new_n6084, new_n6083, new_n6085);
nor_5  g05709(new_n5947, new_n5946, new_n6086);
nor_5  g05710(new_n5949, new_n5944, new_n6087);
nor_5  g05711(new_n6087, new_n6086, new_n6088);
nor_5  g05712(new_n5769, new_n5764, new_n6089_1);
nor_5  g05713(new_n5770, new_n5761, new_n6090);
nor_5  g05714(new_n6090, new_n6089_1, new_n6091);
nor_5  g05715(new_n5815, new_n5810, new_n6092);
nor_5  g05716(new_n5825, new_n5816, new_n6093);
nor_5  g05717(new_n6093, new_n6092, new_n6094);
xnor_4 g05718(new_n6094, new_n6091, new_n6095);
and_5  g05719(new_n5927, new_n5926, new_n6096);
nor_5  g05720(new_n5933, new_n5928, new_n6097);
nor_5  g05721(new_n6097, new_n6096, new_n6098);
and_5  g05722(n8595, n1094, new_n6099);
and_5  g05723(n2564, n1835, new_n6100);
xnor_4 g05724(new_n6100, new_n6099, new_n6101);
xnor_4 g05725(new_n6101, new_n6098, new_n6102);
nor_5  g05726(new_n5877, new_n5876, new_n6103);
nor_5  g05727(new_n5878, new_n5875, new_n6104);
nor_5  g05728(new_n6104, new_n6103, new_n6105);
nand_5 g05729(n12391, n10965, new_n6106);
and_5  g05730(n7891, n503, new_n6107);
and_5  g05731(n9457, n405, new_n6108);
xnor_4 g05732(new_n6108, new_n6107, new_n6109);
xnor_4 g05733(new_n6109, new_n6106, new_n6110);
xnor_4 g05734(new_n6110, new_n6105, new_n6111);
and_5  g05735(n8065, n6986, new_n6112);
and_5  g05736(n10439, n2226, new_n6113);
xnor_4 g05737(new_n6113, new_n6112, new_n6114);
xnor_4 g05738(new_n6114, new_n6111, new_n6115);
xnor_4 g05739(new_n6115, new_n6102, new_n6116);
nor_5  g05740(new_n5758, new_n5757, new_n6117);
nor_5  g05741(new_n5759, new_n5756, new_n6118);
nor_5  g05742(new_n6118, new_n6117, new_n6119);
and_5  g05743(n11536, n6687, new_n6120);
and_5  g05744(n6611, n996, new_n6121);
xnor_4 g05745(new_n6121, new_n6120, new_n6122);
and_5  g05746(n4921, n4516, new_n6123);
and_5  g05747(n9920, n3842, new_n6124);
xnor_4 g05748(new_n6124, new_n6123, new_n6125);
xnor_4 g05749(new_n6125, new_n6122, new_n6126_1);
xnor_4 g05750(new_n6126_1, new_n6119, new_n6127);
nand_5 g05751(n9956, n2087, new_n6128);
and_5  g05752(n7733, n1199, new_n6129);
and_5  g05753(n5767, n217, new_n6130);
xnor_4 g05754(new_n6130, new_n6129, new_n6131);
and_5  g05755(n7160, n4970, new_n6132);
and_5  g05756(n7610, n4828, new_n6133);
xnor_4 g05757(new_n6133, new_n6132, new_n6134);
xnor_4 g05758(new_n6134, new_n6131, new_n6135);
xnor_4 g05759(new_n6135, new_n6128, new_n6136);
xnor_4 g05760(new_n6136, new_n6127, new_n6137);
and_5  g05761(new_n5818, new_n5817, new_n6138);
nor_5  g05762(new_n5824, new_n5819, new_n6139);
nor_5  g05763(new_n6139, new_n6138, new_n6140);
and_5  g05764(n8433, n4817, new_n6141);
and_5  g05765(n10678, n6126, new_n6142);
xnor_4 g05766(new_n6142, new_n6141, new_n6143);
xnor_4 g05767(new_n6143, new_n6140, new_n6144);
xnor_4 g05768(new_n6144, new_n6137, new_n6145);
xnor_4 g05769(new_n6145, new_n6116, new_n6146);
xnor_4 g05770(new_n6146, new_n6095, new_n6147);
xnor_4 g05771(new_n6147, new_n6088, new_n6148);
xnor_4 g05772(new_n6148, new_n6085, new_n6149);
xnor_4 g05773(new_n6149, new_n6082, new_n6150);
nor_5  g05774(new_n5942, new_n5939, new_n6151);
nor_5  g05775(new_n5943, new_n5934_1, new_n6152);
nor_5  g05776(new_n6152, new_n6151, new_n6153);
xnor_4 g05777(new_n6153, new_n6150, new_n6154);
xnor_4 g05778(new_n6154, new_n6079, new_n6155);
xnor_4 g05779(new_n6155, new_n6076, new_n6156);
xnor_4 g05780(new_n6156, new_n5987, n2679);
nor_5  g05781(new_n4476, new_n4460, new_n6158);
and_5  g05782(n6687, n2253, new_n6159);
nand_5 g05783(n10223, n6770, new_n6160);
and_5  g05784(n9920, n2879, new_n6161);
and_5  g05785(n7265, n3627, new_n6162);
xnor_4 g05786(new_n6162, new_n6161, new_n6163);
xnor_4 g05787(new_n6163, new_n6160, new_n6164);
nor_5  g05788(new_n4464, new_n4440, new_n6165);
nor_5  g05789(new_n4465, new_n4463, new_n6166);
or_5   g05790(new_n6166, new_n6165, new_n6167);
xnor_4 g05791(new_n6167, new_n6164, new_n6168);
and_5  g05792(n9195, n2564, new_n6169);
and_5  g05793(n4634, n4189, new_n6170);
xnor_4 g05794(new_n6170, new_n6169, new_n6171);
xnor_4 g05795(new_n6171, new_n6168, new_n6172);
nor_5  g05796(new_n4466, new_n4462, new_n6173);
nor_5  g05797(new_n4470, new_n4467, new_n6174);
nor_5  g05798(new_n6174, new_n6173, new_n6175);
xnor_4 g05799(new_n6175, new_n6172, new_n6176);
nor_5  g05800(new_n4471, new_n4461, new_n6177);
nor_5  g05801(new_n4475, new_n4472, new_n6178);
nor_5  g05802(new_n6178, new_n6177, new_n6179);
xor_4  g05803(new_n6179, new_n6176, new_n6180);
xnor_4 g05804(new_n6180, new_n6159, new_n6181);
xnor_4 g05805(new_n6181, new_n6158, new_n6182);
nor_5  g05806(new_n4650, new_n4477, new_n6183);
nor_5  g05807(new_n4674, new_n4651, new_n6184);
nor_5  g05808(new_n6184, new_n6183, new_n6185);
xnor_4 g05809(new_n6185, new_n6182, new_n6186);
or_5   g05810(new_n4516_1, new_n4499_1, new_n6187);
nand_5 g05811(n12221, n8336, new_n6188);
nand_5 g05812(n9189, n2226, new_n6189);
and_5  g05813(n2024, n1094, new_n6190);
and_5  g05814(n10678, n7946, new_n6191);
xnor_4 g05815(new_n6191, new_n6190, new_n6192_1);
xnor_4 g05816(new_n6192_1, new_n6189, new_n6193);
nor_5  g05817(new_n4508, new_n4482, new_n6194);
nor_5  g05818(new_n4509, new_n4507, new_n6195);
or_5   g05819(new_n6195, new_n6194, new_n6196);
xnor_4 g05820(new_n6196, new_n6193, new_n6197);
and_5  g05821(n12145, n10928, new_n6198);
and_5  g05822(n6986, n2522, new_n6199);
xnor_4 g05823(new_n6199, new_n6198, new_n6200);
xnor_4 g05824(new_n6200, new_n6197, new_n6201);
nor_5  g05825(new_n4505, new_n4501, new_n6202);
nor_5  g05826(new_n4510, new_n4506, new_n6203);
nor_5  g05827(new_n6203, new_n6202, new_n6204);
xnor_4 g05828(new_n6204, new_n6201, new_n6205);
nor_5  g05829(new_n4511, new_n4500, new_n6206);
nor_5  g05830(new_n4515, new_n4512, new_n6207);
nor_5  g05831(new_n6207, new_n6206, new_n6208);
xnor_4 g05832(new_n6208, new_n6205, new_n6209);
xnor_4 g05833(new_n6209, new_n6188, new_n6210);
xnor_4 g05834(new_n6210, new_n6187, new_n6211);
nor_5  g05835(new_n4605, new_n4517, new_n6212);
nor_5  g05836(new_n4649, new_n4606, new_n6213);
nor_5  g05837(new_n6213, new_n6212, new_n6214);
xnor_4 g05838(new_n6214, new_n6211, new_n6215);
or_5   g05839(new_n4624, new_n4607, new_n6216);
nand_5 g05840(n12069, n5798, new_n6217);
and_5  g05841(n7160, n5579, new_n6218);
nor_5  g05842(new_n4617, new_n4615, new_n6219);
nor_5  g05843(new_n6219, new_n4616, new_n6220);
nor_5  g05844(new_n6220, new_n6218, new_n6221);
or_5   g05845(new_n6220, new_n4529, new_n6222);
and_5  g05846(new_n6222, new_n6218, new_n6223);
or_5   g05847(new_n6223, new_n6221, new_n6224);
and_5  g05848(n4828, n2498, new_n6225);
and_5  g05849(n2558, n2515, new_n6226);
xnor_4 g05850(new_n6226, new_n6225, new_n6227);
xnor_4 g05851(new_n6227, new_n6224, new_n6228);
and_5  g05852(n12391, n6016, new_n6229);
and_5  g05853(n7891, n521, new_n6230);
xnor_4 g05854(new_n6230, new_n6229, new_n6231);
xnor_4 g05855(new_n6231, new_n6228, new_n6232);
nor_5  g05856(new_n4613, new_n4609, new_n6233);
nor_5  g05857(new_n4618, new_n4614, new_n6234);
nor_5  g05858(new_n6234, new_n6233, new_n6235);
xnor_4 g05859(new_n6235, new_n6232, new_n6236);
nor_5  g05860(new_n4619, new_n4608, new_n6237);
nor_5  g05861(new_n4623, new_n4620, new_n6238);
nor_5  g05862(new_n6238, new_n6237, new_n6239);
xnor_4 g05863(new_n6239, new_n6236, new_n6240);
xnor_4 g05864(new_n6240, new_n6217, new_n6241);
xnor_4 g05865(new_n6241, new_n6216, new_n6242);
nor_5  g05866(new_n4643, new_n4626, new_n6243);
and_5  g05867(n11222, n5153, new_n6244);
nand_5 g05868(n3342, n996, new_n6245);
and_5  g05869(n9111, n5767, new_n6246);
and_5  g05870(n9763, n5319, new_n6247);
xnor_4 g05871(new_n6247, new_n6246, new_n6248);
xnor_4 g05872(new_n6248, new_n6245, new_n6249);
nor_5  g05873(new_n4635, new_n4545, new_n6250);
and_5  g05874(new_n4635, new_n4545, new_n6251);
nor_5  g05875(new_n6251, new_n4634_1, new_n6252);
or_5   g05876(new_n6252, new_n6250, new_n6253);
xnor_4 g05877(new_n6253, new_n6249, new_n6254_1);
and_5  g05878(n11153, n7270, new_n6255);
and_5  g05879(n5314, n806, new_n6256);
xnor_4 g05880(new_n6256, new_n6255, new_n6257);
xnor_4 g05881(new_n6257, new_n6254_1, new_n6258);
nor_5  g05882(new_n4632, new_n4628, new_n6259);
nor_5  g05883(new_n4637, new_n4633, new_n6260);
nor_5  g05884(new_n6260, new_n6259, new_n6261);
xnor_4 g05885(new_n6261, new_n6258, new_n6262);
nor_5  g05886(new_n4638, new_n4627, new_n6263);
nor_5  g05887(new_n4642, new_n4639, new_n6264);
nor_5  g05888(new_n6264, new_n6263, new_n6265);
xor_4  g05889(new_n6265, new_n6262, new_n6266);
xnor_4 g05890(new_n6266, new_n6244, new_n6267);
xor_4  g05891(new_n6267, new_n6243, new_n6268);
xnor_4 g05892(new_n6268, new_n6242, new_n6269);
nor_5  g05893(new_n4644, new_n4625, new_n6270);
nor_5  g05894(new_n4648, new_n4645, new_n6271);
or_5   g05895(new_n6271, new_n6270, new_n6272);
xnor_4 g05896(new_n6272, new_n6269, new_n6273_1);
xnor_4 g05897(new_n6273_1, new_n6215, new_n6274);
xor_4  g05898(new_n6274, new_n6186, n2708);
xnor_4 g05899(new_n762, new_n761, n2818);
xnor_4 g05900(new_n1672, new_n1650, n2902);
and_5  g05901(n11407, n5305, new_n6278);
and_5  g05902(n12709, n8759, new_n6279);
and_5  g05903(n12489, n5331, new_n6280);
and_5  g05904(n10990, n7965, new_n6281);
xnor_4 g05905(new_n6281, new_n6280, new_n6282);
xnor_4 g05906(new_n6282, new_n6279, new_n6283);
xor_4  g05907(new_n6283, new_n6278, n3071);
xnor_4 g05908(new_n2340, new_n2339, n3124);
and_5  g05909(new_n6283, new_n6278, new_n6286);
and_5  g05910(n11407, n5964, new_n6287);
and_5  g05911(n5305, n5212, new_n6288);
xor_4  g05912(new_n6288, new_n6287, new_n6289);
nor_5  g05913(new_n6289, new_n6286, new_n6290);
nand_5 g05914(n12709, n8759, new_n6291);
nor_5  g05915(new_n6282, new_n6291, new_n6292);
and_5  g05916(n11728, n8759, new_n6293);
and_5  g05917(n12709, n6776, new_n6294_1);
xor_4  g05918(new_n6294_1, new_n6293, new_n6295);
xnor_4 g05919(new_n6295, new_n6292, new_n6296);
and_5  g05920(new_n6281, new_n6280, new_n6297);
and_5  g05921(n7159, n5331, new_n6298);
and_5  g05922(n12489, n8476, new_n6299);
xor_4  g05923(new_n6299, new_n6298, new_n6300);
xnor_4 g05924(new_n6300, new_n6297, new_n6301);
and_5  g05925(n7965, n5760, new_n6302);
and_5  g05926(n10990, n7388, new_n6303);
xor_4  g05927(new_n6303, new_n6302, new_n6304);
xor_4  g05928(new_n6304, new_n6301, new_n6305);
xnor_4 g05929(new_n6305, new_n6296, new_n6306);
xor_4  g05930(new_n6289, new_n6286, new_n6307);
and_5  g05931(new_n6307, new_n6306, new_n6308);
nor_5  g05932(new_n6308, new_n6290, new_n6309);
nand_5 g05933(n5964, n5212, new_n6310);
nor_5  g05934(new_n6310, new_n6278, new_n6311);
and_5  g05935(n11407, n1097, new_n6312);
and_5  g05936(n11877, n5305, new_n6313);
xor_4  g05937(new_n6313, new_n6312, new_n6314);
or_5   g05938(new_n6314, new_n6311, new_n6315);
or_5   g05939(new_n6310, new_n6278, new_n6316);
nor_5  g05940(new_n6313, new_n6312, new_n6317);
or_5   g05941(new_n6317, new_n6316, new_n6318);
and_5  g05942(new_n6318, new_n6315, new_n6319);
xnor_4 g05943(new_n6319, new_n6309, new_n6320);
and_5  g05944(new_n6295, new_n6292, new_n6321);
nor_5  g05945(new_n6305, new_n6296, new_n6322);
nor_5  g05946(new_n6322, new_n6321, new_n6323);
nand_5 g05947(n11728, n6776, new_n6324);
or_5   g05948(new_n6324, new_n6279, new_n6325);
and_5  g05949(n12709, n12299, new_n6326);
and_5  g05950(n8759, n6429, new_n6327);
xnor_4 g05951(new_n6327, new_n6326, new_n6328);
nand_5 g05952(new_n6328, new_n6325, new_n6329);
nor_5  g05953(new_n6327, new_n6326, new_n6330);
or_5   g05954(new_n6330, new_n6325, new_n6331);
nand_5 g05955(new_n6331, new_n6329, new_n6332);
xnor_4 g05956(new_n6332, new_n6323, new_n6333);
nand_5 g05957(n8476, n7159, new_n6334);
or_5   g05958(new_n6334, new_n6280, new_n6335);
and_5  g05959(n12489, n2530, new_n6336);
and_5  g05960(n12777, n5331, new_n6337);
nor_5  g05961(new_n6337, new_n6336, new_n6338);
and_5  g05962(n12777, n2530, new_n6339);
and_5  g05963(new_n6339, new_n6280, new_n6340);
or_5   g05964(new_n6340, new_n6338, new_n6341);
nand_5 g05965(new_n6341, new_n6335, new_n6342);
or_5   g05966(new_n6338, new_n6335, new_n6343);
and_5  g05967(new_n6343, new_n6342, new_n6344);
nand_5 g05968(n7388, n5760, new_n6345);
nor_5  g05969(new_n6345, new_n6281, new_n6346);
and_5  g05970(n11892, n10990, new_n6347);
and_5  g05971(n7965, n1478, new_n6348);
xor_4  g05972(new_n6348, new_n6347, new_n6349);
or_5   g05973(new_n6349, new_n6346, new_n6350);
or_5   g05974(new_n6345, new_n6281, new_n6351);
nor_5  g05975(new_n6348, new_n6347, new_n6352);
or_5   g05976(new_n6352, new_n6351, new_n6353);
and_5  g05977(new_n6353, new_n6350, new_n6354);
xnor_4 g05978(new_n6354, new_n6344, new_n6355);
nor_5  g05979(new_n6300, new_n6297, new_n6356);
nor_5  g05980(new_n6304, new_n6301, new_n6357);
or_5   g05981(new_n6357, new_n6356, new_n6358_1);
xnor_4 g05982(new_n6358_1, new_n6355, new_n6359_1);
xnor_4 g05983(new_n6359_1, new_n6333, new_n6360);
xor_4  g05984(new_n6360, new_n6320, n3214);
xnor_4 g05985(new_n4330, new_n4329, n3230);
xor_4  g05986(new_n3917, new_n3880, n3272);
and_5  g05987(n5964, n4370, new_n6364);
and_5  g05988(n11407, n4312, new_n6365);
and_5  g05989(n11877, n5964, new_n6366);
nor_5  g05990(new_n6366, new_n6365, new_n6367);
nand_5 g05991(new_n6366, new_n6365, new_n6368);
nand_5 g05992(n5212, n1097, new_n6369);
and_5  g05993(new_n6369, new_n6368, new_n6370);
nor_5  g05994(new_n6370, new_n6367, new_n6371);
and_5  g05995(new_n6371, new_n6364, new_n6372);
xnor_4 g05996(new_n6371, new_n6364, new_n6373);
and_5  g05997(n5212, n4312, new_n6374);
and_5  g05998(n11877, n1097, new_n6375);
and_5  g05999(n12705, n11407, new_n6376);
xnor_4 g06000(new_n6376, new_n6375, new_n6377);
xor_4  g06001(new_n6377, new_n6374, new_n6378);
nor_5  g06002(new_n6378, new_n6373, new_n6379);
nor_5  g06003(new_n6379, new_n6372, new_n6380);
and_5  g06004(n5964, n5320, new_n6381);
and_5  g06005(n4370, n1097, new_n6382);
xnor_4 g06006(new_n6382, new_n6381, new_n6383);
xnor_4 g06007(new_n6383, new_n6380, new_n6384);
and_5  g06008(n11877, n4312, new_n6385);
and_5  g06009(n12705, n5212, new_n6386);
and_5  g06010(n12025, n11407, new_n6387);
xor_4  g06011(new_n6387, new_n6386, new_n6388);
xnor_4 g06012(new_n6388, new_n6385, new_n6389);
nor_5  g06013(new_n6376, new_n6375, new_n6390);
and_5  g06014(new_n6376, new_n6375, new_n6391);
nor_5  g06015(new_n6391, new_n6374, new_n6392);
nor_5  g06016(new_n6392, new_n6390, new_n6393);
xor_4  g06017(new_n6393, new_n6389, new_n6394);
xnor_4 g06018(new_n6394, new_n6384, new_n6395);
and_5  g06019(n5320, n5305, new_n6396);
xor_4  g06020(new_n6378, new_n6373, new_n6397);
nor_5  g06021(new_n6397, new_n6396, new_n6398);
xnor_4 g06022(new_n6397, new_n6396, new_n6399);
nand_5 g06023(n5305, n4370, new_n6400);
nand_5 g06024(new_n6313, new_n6312, new_n6401);
and_5  g06025(new_n6401, new_n6310, new_n6402);
or_5   g06026(new_n6402, new_n6317, new_n6403);
nor_5  g06027(new_n6403, new_n6400, new_n6404);
xnor_4 g06028(new_n6403, new_n6400, new_n6405);
xnor_4 g06029(new_n6366, new_n6365, new_n6406);
xnor_4 g06030(new_n6406, new_n6369, new_n6407);
nor_5  g06031(new_n6407, new_n6405, new_n6408);
or_5   g06032(new_n6408, new_n6404, new_n6409);
nor_5  g06033(new_n6409, new_n6399, new_n6410);
or_5   g06034(new_n6410, new_n6398, new_n6411);
nor_5  g06035(new_n6411, new_n6395, new_n6412);
nor_5  g06036(new_n6388, new_n6385, new_n6413);
nor_5  g06037(new_n6393, new_n6389, new_n6414);
nor_5  g06038(new_n6414, new_n6413, new_n6415);
and_5  g06039(n12000, n5964, new_n6416);
and_5  g06040(n5320, n1097, new_n6417);
and_5  g06041(n9725, n5305, new_n6418);
xnor_4 g06042(new_n6418, new_n6417, new_n6419);
xnor_4 g06043(new_n6419, new_n6416, new_n6420);
xnor_4 g06044(new_n6420, new_n6415, new_n6421);
and_5  g06045(new_n6387, new_n6386, new_n6422);
and_5  g06046(n4370, n4312, new_n6423);
xnor_4 g06047(new_n6423, new_n6422, new_n6424);
and_5  g06048(n12025, n5212, new_n6425);
and_5  g06049(n12705, n11877, new_n6426);
and_5  g06050(n11407, n11257, new_n6427);
xnor_4 g06051(new_n6427, new_n6426, new_n6428);
xnor_4 g06052(new_n6428, new_n6425, new_n6429_1);
xnor_4 g06053(new_n6429_1, new_n6424, new_n6430);
xor_4  g06054(new_n6430, new_n6421, new_n6431_1);
nor_5  g06055(new_n6383, new_n6380, new_n6432);
nand_5 g06056(new_n6382, new_n6381, new_n6433);
or_5   g06057(new_n6394, new_n6384, new_n6434);
xor_4  g06058(new_n6434, new_n6433, new_n6435);
nor_5  g06059(new_n6435, new_n6432, new_n6436);
xor_4  g06060(new_n6436, new_n6431_1, new_n6437);
xnor_4 g06061(new_n6437, new_n6412, new_n6438);
and_5  g06062(n12000, n5305, new_n6439);
xor_4  g06063(new_n6411, new_n6395, new_n6440);
and_5  g06064(new_n6440, new_n6439, new_n6441_1);
xnor_4 g06065(new_n6407, new_n6405, new_n6442);
or_5   g06066(new_n6315, new_n6310, new_n6443);
or_5   g06067(new_n6443, new_n6442, new_n6444);
xor_4  g06068(new_n6409, new_n6399, new_n6445_1);
or_5   g06069(new_n6445_1, new_n6444, new_n6446);
xnor_4 g06070(new_n6440, new_n6439, new_n6447);
nor_5  g06071(new_n6447, new_n6446, new_n6448);
nor_5  g06072(new_n6448, new_n6441_1, new_n6449);
xnor_4 g06073(new_n6449, new_n6438, new_n6450);
and_5  g06074(n8759, n8717, new_n6451);
and_5  g06075(n7436, n6429, new_n6452);
and_5  g06076(n12709, n9241, new_n6453);
and_5  g06077(n11728, n8276, new_n6454);
xor_4  g06078(new_n6454, new_n6453, new_n6455);
xnor_4 g06079(new_n6455, new_n6452, new_n6456);
and_5  g06080(n12299, n6429, new_n6457);
and_5  g06081(n12709, n8276, new_n6458);
nor_5  g06082(new_n6458, new_n6457, new_n6459);
nand_5 g06083(new_n6458, new_n6457, new_n6460);
nand_5 g06084(n11728, n7436, new_n6461);
and_5  g06085(new_n6461, new_n6460, new_n6462);
nor_5  g06086(new_n6462, new_n6459, new_n6463);
xor_4  g06087(new_n6463, new_n6456, new_n6464);
and_5  g06088(n6776, n2433, new_n6465);
and_5  g06089(n12299, n8819, new_n6466);
xnor_4 g06090(new_n6466, new_n6465, new_n6467);
xnor_4 g06091(new_n6467, new_n6464, new_n6468);
nand_5 g06092(n8819, n6776, new_n6469);
and_5  g06093(n12709, n7436, new_n6470);
and_5  g06094(n6776, n6429, new_n6471);
nor_5  g06095(new_n6471, new_n6470, new_n6472);
nand_5 g06096(new_n6471, new_n6470, new_n6473);
nand_5 g06097(n12299, n11728, new_n6474);
and_5  g06098(new_n6474, new_n6473, new_n6475);
or_5   g06099(new_n6475, new_n6472, new_n6476);
nor_5  g06100(new_n6476, new_n6469, new_n6477);
xnor_4 g06101(new_n6476, new_n6469, new_n6478);
xnor_4 g06102(new_n6458, new_n6457, new_n6479);
xnor_4 g06103(new_n6479, new_n6461, new_n6480);
nor_5  g06104(new_n6480, new_n6478, new_n6481);
nor_5  g06105(new_n6481, new_n6477, new_n6482);
xnor_4 g06106(new_n6482, new_n6468, new_n6483);
and_5  g06107(n8759, n2433, new_n6484);
xor_4  g06108(new_n6480, new_n6478, new_n6485);
nor_5  g06109(new_n6485, new_n6484, new_n6486);
xnor_4 g06110(new_n6485, new_n6484, new_n6487);
nand_5 g06111(n8819, n8759, new_n6488);
nand_5 g06112(new_n6327, new_n6326, new_n6489);
and_5  g06113(new_n6489, new_n6324, new_n6490);
or_5   g06114(new_n6490, new_n6330, new_n6491);
nor_5  g06115(new_n6491, new_n6488, new_n6492);
xnor_4 g06116(new_n6491, new_n6488, new_n6493);
xnor_4 g06117(new_n6471, new_n6470, new_n6494);
xnor_4 g06118(new_n6494, new_n6474, new_n6495);
nor_5  g06119(new_n6495, new_n6493, new_n6496);
or_5   g06120(new_n6496, new_n6492, new_n6497);
nor_5  g06121(new_n6497, new_n6487, new_n6498);
or_5   g06122(new_n6498, new_n6486, new_n6499);
xor_4  g06123(new_n6499, new_n6483, new_n6500);
and_5  g06124(new_n6500, new_n6451, new_n6501);
xnor_4 g06125(new_n6495, new_n6493, new_n6502);
or_5   g06126(new_n6329, new_n6324, new_n6503);
or_5   g06127(new_n6503, new_n6502, new_n6504);
xor_4  g06128(new_n6497, new_n6487, new_n6505);
or_5   g06129(new_n6505, new_n6504, new_n6506);
xnor_4 g06130(new_n6500, new_n6451, new_n6507);
nor_5  g06131(new_n6507, new_n6506, new_n6508);
nor_5  g06132(new_n6508, new_n6501, new_n6509);
or_5   g06133(new_n6499, new_n6483, new_n6510);
nor_5  g06134(new_n6455, new_n6452, new_n6511);
nor_5  g06135(new_n6463, new_n6456, new_n6512);
nor_5  g06136(new_n6512, new_n6511, new_n6513);
nand_5 g06137(n8717, n6776, new_n6514);
and_5  g06138(n12299, n2433, new_n6515);
and_5  g06139(n8759, n7730, new_n6516);
xnor_4 g06140(new_n6516, new_n6515, new_n6517);
xor_4  g06141(new_n6517, new_n6514, new_n6518);
xnor_4 g06142(new_n6518, new_n6513, new_n6519);
and_5  g06143(new_n6454, new_n6453, new_n6520);
and_5  g06144(n8819, n7436, new_n6521);
xnor_4 g06145(new_n6521, new_n6520, new_n6522);
and_5  g06146(n11728, n9241, new_n6523);
and_5  g06147(n8276, n6429, new_n6524);
and_5  g06148(n12709, n10510, new_n6525);
xnor_4 g06149(new_n6525, new_n6524, new_n6526);
xor_4  g06150(new_n6526, new_n6523, new_n6527);
xor_4  g06151(new_n6527, new_n6522, new_n6528);
xor_4  g06152(new_n6528, new_n6519, new_n6529);
nor_5  g06153(new_n6467, new_n6464, new_n6530);
nand_5 g06154(new_n6466, new_n6465, new_n6531);
or_5   g06155(new_n6482, new_n6468, new_n6532);
xor_4  g06156(new_n6532, new_n6531, new_n6533);
nor_5  g06157(new_n6533, new_n6530, new_n6534);
xnor_4 g06158(new_n6534, new_n6529, new_n6535);
xnor_4 g06159(new_n6535, new_n6510, new_n6536);
xor_4  g06160(new_n6536, new_n6509, new_n6537);
nand_5 g06161(n2393, n1478, new_n6538);
and_5  g06162(n5860, n5760, new_n6539);
and_5  g06163(n10990, n3986, new_n6540);
xnor_4 g06164(new_n6540, new_n6539, new_n6541);
xnor_4 g06165(new_n6541, new_n6538, new_n6542);
and_5  g06166(n11892, n1478, new_n6543);
and_5  g06167(n10990, n5860, new_n6544);
nor_5  g06168(new_n6544, new_n6543, new_n6545);
nand_5 g06169(new_n6544, new_n6543, new_n6546);
nand_5 g06170(n5760, n2393, new_n6547);
and_5  g06171(new_n6547, new_n6546, new_n6548);
or_5   g06172(new_n6548, new_n6545, new_n6549);
xnor_4 g06173(new_n6549, new_n6542, new_n6550);
and_5  g06174(n12947, n7388, new_n6551);
and_5  g06175(n11892, n11791, new_n6552);
xnor_4 g06176(new_n6552, new_n6551, new_n6553);
xnor_4 g06177(new_n6553, new_n6550, new_n6554);
nand_5 g06178(n11791, n7388, new_n6555);
and_5  g06179(n10990, n2393, new_n6556);
and_5  g06180(n7388, n1478, new_n6557);
nor_5  g06181(new_n6557, new_n6556, new_n6558);
nand_5 g06182(new_n6557, new_n6556, new_n6559);
nand_5 g06183(n11892, n5760, new_n6560);
and_5  g06184(new_n6560, new_n6559, new_n6561);
or_5   g06185(new_n6561, new_n6558, new_n6562);
nor_5  g06186(new_n6562, new_n6555, new_n6563);
xnor_4 g06187(new_n6562, new_n6555, new_n6564);
xnor_4 g06188(new_n6544, new_n6543, new_n6565);
xnor_4 g06189(new_n6565, new_n6547, new_n6566);
nor_5  g06190(new_n6566, new_n6564, new_n6567);
nor_5  g06191(new_n6567, new_n6563, new_n6568);
xnor_4 g06192(new_n6568, new_n6554, new_n6569);
and_5  g06193(n12947, n7965, new_n6570);
nand_5 g06194(n11791, n7965, new_n6571);
nand_5 g06195(new_n6348, new_n6347, new_n6572);
and_5  g06196(new_n6572, new_n6345, new_n6573);
or_5   g06197(new_n6573, new_n6352, new_n6574);
nor_5  g06198(new_n6574, new_n6571, new_n6575);
xnor_4 g06199(new_n6574, new_n6571, new_n6576);
xnor_4 g06200(new_n6557, new_n6556, new_n6577);
xnor_4 g06201(new_n6577, new_n6560, new_n6578_1);
nor_5  g06202(new_n6578_1, new_n6576, new_n6579);
or_5   g06203(new_n6579, new_n6575, new_n6580);
nor_5  g06204(new_n6580, new_n6570, new_n6581);
xor_4  g06205(new_n6566, new_n6564, new_n6582);
xnor_4 g06206(new_n6580, new_n6570, new_n6583);
nor_5  g06207(new_n6583, new_n6582, new_n6584);
or_5   g06208(new_n6584, new_n6581, new_n6585);
or_5   g06209(new_n6585, new_n6569, new_n6586);
and_5  g06210(new_n6540, new_n6539, new_n6587);
and_5  g06211(n11791, n2393, new_n6588);
xnor_4 g06212(new_n6588, new_n6587, new_n6589);
nand_5 g06213(n5760, n3986, new_n6590);
and_5  g06214(n5860, n1478, new_n6591);
and_5  g06215(n10990, n5857, new_n6592);
xnor_4 g06216(new_n6592, new_n6591, new_n6593);
xnor_4 g06217(new_n6593, new_n6590, new_n6594);
xor_4  g06218(new_n6594, new_n6589, new_n6595);
and_5  g06219(n7388, n6441, new_n6596);
nand_5 g06220(n12947, n11892, new_n6597);
nand_5 g06221(n11999, n7965, new_n6598);
xnor_4 g06222(new_n6598, new_n6597, new_n6599);
xnor_4 g06223(new_n6599, new_n6596, new_n6600);
nor_5  g06224(new_n6541, new_n6538, new_n6601);
nor_5  g06225(new_n6549, new_n6542, new_n6602);
or_5   g06226(new_n6602, new_n6601, new_n6603);
xnor_4 g06227(new_n6603, new_n6600, new_n6604_1);
xor_4  g06228(new_n6604_1, new_n6595, new_n6605);
nor_5  g06229(new_n6553, new_n6550, new_n6606);
nand_5 g06230(new_n6552, new_n6551, new_n6607);
or_5   g06231(new_n6568, new_n6554, new_n6608);
xor_4  g06232(new_n6608, new_n6607, new_n6609);
nor_5  g06233(new_n6609, new_n6606, new_n6610);
xnor_4 g06234(new_n6610, new_n6605, new_n6611_1);
xnor_4 g06235(new_n6611_1, new_n6586, new_n6612);
and_5  g06236(n7965, n6441, new_n6613);
xor_4  g06237(new_n6585, new_n6569, new_n6614);
and_5  g06238(new_n6614, new_n6613, new_n6615);
nor_5  g06239(new_n6614, new_n6613, new_n6616);
xnor_4 g06240(new_n6578_1, new_n6576, new_n6617);
or_5   g06241(new_n6350, new_n6345, new_n6618);
or_5   g06242(new_n6618, new_n6617, new_n6619);
xor_4  g06243(new_n6583, new_n6582, new_n6620);
or_5   g06244(new_n6620, new_n6619, new_n6621);
nor_5  g06245(new_n6621, new_n6616, new_n6622);
nor_5  g06246(new_n6622, new_n6615, new_n6623);
xor_4  g06247(new_n6623, new_n6612, new_n6624);
nand_5 g06248(n12777, n12648, new_n6625);
and_5  g06249(n10545, n7159, new_n6626);
and_5  g06250(n12489, n7690, new_n6627);
xnor_4 g06251(new_n6627, new_n6626, new_n6628);
xnor_4 g06252(new_n6628, new_n6625, new_n6629);
and_5  g06253(n12489, n10545, new_n6630);
nor_5  g06254(new_n6630, new_n6339, new_n6631);
nand_5 g06255(new_n6630, new_n6339, new_n6632);
nand_5 g06256(n12648, n7159, new_n6633);
and_5  g06257(new_n6633, new_n6632, new_n6634);
or_5   g06258(new_n6634, new_n6631, new_n6635);
xnor_4 g06259(new_n6635, new_n6629, new_n6636);
and_5  g06260(n6254, n2530, new_n6637);
and_5  g06261(n11967, n8476, new_n6638);
xnor_4 g06262(new_n6638, new_n6637, new_n6639);
xnor_4 g06263(new_n6639, new_n6636, new_n6640);
nand_5 g06264(n8476, n6254, new_n6641);
and_5  g06265(n12648, n12489, new_n6642);
and_5  g06266(n12777, n8476, new_n6643);
nor_5  g06267(new_n6643, new_n6642, new_n6644);
nand_5 g06268(new_n6643, new_n6642, new_n6645_1);
nand_5 g06269(n7159, n2530, new_n6646);
and_5  g06270(new_n6646, new_n6645_1, new_n6647);
or_5   g06271(new_n6647, new_n6644, new_n6648);
nor_5  g06272(new_n6648, new_n6641, new_n6649);
xnor_4 g06273(new_n6648, new_n6641, new_n6650);
xnor_4 g06274(new_n6630, new_n6339, new_n6651);
xnor_4 g06275(new_n6651, new_n6633, new_n6652);
nor_5  g06276(new_n6652, new_n6650, new_n6653);
nor_5  g06277(new_n6653, new_n6649, new_n6654);
xnor_4 g06278(new_n6654, new_n6640, new_n6655);
and_5  g06279(n11967, n5331, new_n6656);
xor_4  g06280(new_n6652, new_n6650, new_n6657);
nor_5  g06281(new_n6657, new_n6656, new_n6658);
xnor_4 g06282(new_n6657, new_n6656, new_n6659);
nand_5 g06283(n6254, n5331, new_n6660);
and_5  g06284(n8476, n7159, new_n6661);
nor_5  g06285(new_n6340, new_n6661, new_n6662);
or_5   g06286(new_n6662, new_n6338, new_n6663);
nor_5  g06287(new_n6663, new_n6660, new_n6664);
xnor_4 g06288(new_n6663, new_n6660, new_n6665);
xnor_4 g06289(new_n6643, new_n6642, new_n6666);
xnor_4 g06290(new_n6666, new_n6646, new_n6667);
nor_5  g06291(new_n6667, new_n6665, new_n6668);
or_5   g06292(new_n6668, new_n6664, new_n6669);
nor_5  g06293(new_n6669, new_n6659, new_n6670);
or_5   g06294(new_n6670, new_n6658, new_n6671);
or_5   g06295(new_n6671, new_n6655, new_n6672);
and_5  g06296(n5331, n1353, new_n6673);
and_5  g06297(n11967, n2530, new_n6674);
and_5  g06298(n8476, n447, new_n6675);
xnor_4 g06299(new_n6675, new_n6674, new_n6676);
xnor_4 g06300(new_n6676, new_n6673, new_n6677);
nor_5  g06301(new_n6628, new_n6625, new_n6678);
nor_5  g06302(new_n6635, new_n6629, new_n6679);
or_5   g06303(new_n6679, new_n6678, new_n6680);
xnor_4 g06304(new_n6680, new_n6677, new_n6681);
and_5  g06305(new_n6627, new_n6626, new_n6682);
and_5  g06306(n12648, n6254, new_n6683);
xnor_4 g06307(new_n6683, new_n6682, new_n6684);
and_5  g06308(n7690, n7159, new_n6685);
and_5  g06309(n12777, n10545, new_n6686);
and_5  g06310(n12489, n3616, new_n6687_1);
xnor_4 g06311(new_n6687_1, new_n6686, new_n6688);
xor_4  g06312(new_n6688, new_n6685, new_n6689_1);
xor_4  g06313(new_n6689_1, new_n6684, new_n6690);
xor_4  g06314(new_n6690, new_n6681, new_n6691);
nor_5  g06315(new_n6639, new_n6636, new_n6692);
nand_5 g06316(new_n6638, new_n6637, new_n6693);
or_5   g06317(new_n6654, new_n6640, new_n6694);
xor_4  g06318(new_n6694, new_n6693, new_n6695);
nor_5  g06319(new_n6695, new_n6692, new_n6696);
xnor_4 g06320(new_n6696, new_n6691, new_n6697);
xnor_4 g06321(new_n6697, new_n6672, new_n6698);
and_5  g06322(n5331, n447, new_n6699);
xor_4  g06323(new_n6671, new_n6655, new_n6700);
and_5  g06324(new_n6700, new_n6699, new_n6701);
nor_5  g06325(new_n6700, new_n6699, new_n6702);
xnor_4 g06326(new_n6667, new_n6665, new_n6703_1);
or_5   g06327(new_n6342, new_n6334, new_n6704);
or_5   g06328(new_n6704, new_n6703_1, new_n6705);
xor_4  g06329(new_n6669, new_n6659, new_n6706);
or_5   g06330(new_n6706, new_n6705, new_n6707);
nor_5  g06331(new_n6707, new_n6702, new_n6708);
nor_5  g06332(new_n6708, new_n6701, new_n6709);
xor_4  g06333(new_n6709, new_n6698, new_n6710);
xnor_4 g06334(new_n6710, new_n6624, new_n6711);
xor_4  g06335(new_n6614, new_n6613, new_n6712);
xnor_4 g06336(new_n6712, new_n6621, new_n6713);
xor_4  g06337(new_n6700, new_n6699, new_n6714);
xnor_4 g06338(new_n6714, new_n6707, new_n6715);
nor_5  g06339(new_n6715, new_n6713, new_n6716);
xor_4  g06340(new_n6706, new_n6705, new_n6717);
xor_4  g06341(new_n6620, new_n6619, new_n6718);
nor_5  g06342(new_n6718, new_n6717, new_n6719);
xnor_4 g06343(new_n6718, new_n6717, new_n6720);
xnor_4 g06344(new_n6704, new_n6703_1, new_n6721);
xnor_4 g06345(new_n6618, new_n6617, new_n6722);
nor_5  g06346(new_n6722, new_n6721, new_n6723);
and_5  g06347(new_n6354, new_n6344, new_n6724);
nor_5  g06348(new_n6358_1, new_n6355, new_n6725);
nor_5  g06349(new_n6725, new_n6724, new_n6726);
xnor_4 g06350(new_n6722, new_n6721, new_n6727);
nor_5  g06351(new_n6727, new_n6726, new_n6728);
or_5   g06352(new_n6728, new_n6723, new_n6729);
nor_5  g06353(new_n6729, new_n6720, new_n6730);
nor_5  g06354(new_n6730, new_n6719, new_n6731);
xnor_4 g06355(new_n6715, new_n6713, new_n6732);
nor_5  g06356(new_n6732, new_n6731, new_n6733);
nor_5  g06357(new_n6733, new_n6716, new_n6734);
xnor_4 g06358(new_n6734, new_n6711, new_n6735);
xnor_4 g06359(new_n6735, new_n6537, new_n6736);
xor_4  g06360(new_n6507, new_n6506, new_n6737);
xnor_4 g06361(new_n6732, new_n6731, new_n6738);
nor_5  g06362(new_n6738, new_n6737, new_n6739);
xnor_4 g06363(new_n6738, new_n6737, new_n6740);
xnor_4 g06364(new_n6505, new_n6504, new_n6741);
xor_4  g06365(new_n6729, new_n6720, new_n6742_1);
nor_5  g06366(new_n6742_1, new_n6741, new_n6743);
xnor_4 g06367(new_n6503, new_n6502, new_n6744);
xnor_4 g06368(new_n6727, new_n6726, new_n6745);
nor_5  g06369(new_n6745, new_n6744, new_n6746);
xnor_4 g06370(new_n6745, new_n6744, new_n6747);
nor_5  g06371(new_n6332, new_n6323, new_n6748);
nor_5  g06372(new_n6359_1, new_n6333, new_n6749);
nor_5  g06373(new_n6749, new_n6748, new_n6750);
nor_5  g06374(new_n6750, new_n6747, new_n6751);
nor_5  g06375(new_n6751, new_n6746, new_n6752);
xnor_4 g06376(new_n6742_1, new_n6741, new_n6753);
nor_5  g06377(new_n6753, new_n6752, new_n6754);
or_5   g06378(new_n6754, new_n6743, new_n6755);
nor_5  g06379(new_n6755, new_n6740, new_n6756);
nor_5  g06380(new_n6756, new_n6739, new_n6757);
xor_4  g06381(new_n6757, new_n6736, new_n6758);
nor_5  g06382(new_n6758, new_n6450, new_n6759);
xnor_4 g06383(new_n6758, new_n6450, new_n6760);
xnor_4 g06384(new_n6447, new_n6446, new_n6761);
xor_4  g06385(new_n6755, new_n6740, new_n6762);
and_5  g06386(new_n6762, new_n6761, new_n6763);
xnor_4 g06387(new_n6762, new_n6761, new_n6764);
xor_4  g06388(new_n6445_1, new_n6444, new_n6765);
xor_4  g06389(new_n6753, new_n6752, new_n6766);
nor_5  g06390(new_n6766, new_n6765, new_n6767);
xnor_4 g06391(new_n6766, new_n6765, new_n6768);
xor_4  g06392(new_n6443, new_n6442, new_n6769);
xor_4  g06393(new_n6750, new_n6747, new_n6770_1);
nor_5  g06394(new_n6770_1, new_n6769, new_n6771);
and_5  g06395(new_n6319, new_n6309, new_n6772);
nor_5  g06396(new_n6360, new_n6320, new_n6773);
nor_5  g06397(new_n6773, new_n6772, new_n6774);
xor_4  g06398(new_n6770_1, new_n6769, new_n6775);
and_5  g06399(new_n6775, new_n6774, new_n6776_1);
nor_5  g06400(new_n6776_1, new_n6771, new_n6777);
nor_5  g06401(new_n6777, new_n6768, new_n6778);
nor_5  g06402(new_n6778, new_n6767, new_n6779);
nor_5  g06403(new_n6779, new_n6764, new_n6780);
or_5   g06404(new_n6780, new_n6763, new_n6781);
nor_5  g06405(new_n6781, new_n6760, new_n6782);
nor_5  g06406(new_n6782, new_n6759, new_n6783);
nor_5  g06407(new_n6735, new_n6537, new_n6784);
nor_5  g06408(new_n6757, new_n6736, new_n6785);
nor_5  g06409(new_n6785, new_n6784, new_n6786);
and_5  g06410(new_n6437, new_n6412, new_n6787);
nor_5  g06411(new_n6449, new_n6438, new_n6788);
nor_5  g06412(new_n6788, new_n6787, new_n6789);
nor_5  g06413(new_n6427, new_n6426, new_n6790);
nor_5  g06414(new_n6428, new_n6425, new_n6791);
or_5   g06415(new_n6791, new_n6790, new_n6792);
nor_5  g06416(new_n6418, new_n6417, new_n6793);
nor_5  g06417(new_n6419, new_n6416, new_n6794);
nor_5  g06418(new_n6794, new_n6793, new_n6795);
and_5  g06419(n9725, n5964, new_n6796);
xnor_4 g06420(new_n6796, new_n6795, new_n6797_1);
xnor_4 g06421(new_n6797_1, new_n6792, new_n6798);
xnor_4 g06422(new_n6798, new_n6789, new_n6799);
nor_5  g06423(new_n6535, new_n6510, new_n6800);
nor_5  g06424(new_n6536, new_n6509, new_n6801);
nor_5  g06425(new_n6801, new_n6800, new_n6802);
nor_5  g06426(new_n6697, new_n6672, new_n6803);
nor_5  g06427(new_n6709, new_n6698, new_n6804);
nor_5  g06428(new_n6804, new_n6803, new_n6805);
xnor_4 g06429(new_n6805, new_n6802, new_n6806_1);
nor_5  g06430(new_n6611_1, new_n6586, new_n6807);
nor_5  g06431(new_n6623, new_n6612, new_n6808);
nor_5  g06432(new_n6808, new_n6807, new_n6809_1);
nor_5  g06433(new_n6680, new_n6677, new_n6810);
nor_5  g06434(new_n6690, new_n6681, new_n6811);
nor_5  g06435(new_n6811, new_n6810, new_n6812);
and_5  g06436(new_n6516, new_n6515, new_n6813);
nor_5  g06437(new_n6516, new_n6515, new_n6814);
nor_5  g06438(new_n6814, new_n6514, new_n6815);
nor_5  g06439(new_n6815, new_n6813, new_n6816);
and_5  g06440(n3986, n1478, new_n6817);
and_5  g06441(n9241, n6429, new_n6818);
and_5  g06442(n10022, n7965, new_n6819);
xnor_4 g06443(new_n6819, new_n6818, new_n6820);
xnor_4 g06444(new_n6820, new_n6817, new_n6821);
xnor_4 g06445(new_n6821, new_n6816, new_n6822_1);
xnor_4 g06446(new_n6822_1, new_n6812, new_n6823);
nor_5  g06447(new_n6687_1, new_n6686, new_n6824);
nor_5  g06448(new_n6688, new_n6685, new_n6825);
nor_5  g06449(new_n6825, new_n6824, new_n6826_1);
nor_5  g06450(new_n6599, new_n6596, new_n6827);
or_5   g06451(new_n6827, new_n6597, new_n6828);
nand_5 g06452(n11999, n7388, new_n6829);
nor_5  g06453(new_n6829, new_n6828, new_n6830);
or_5   g06454(new_n6829, new_n6613, new_n6831);
and_5  g06455(new_n6831, new_n6828, new_n6832);
nor_5  g06456(new_n6832, new_n6830, new_n6833);
xnor_4 g06457(new_n6833, new_n6826_1, new_n6834);
and_5  g06458(new_n6683, new_n6682, new_n6835);
nor_5  g06459(new_n6689_1, new_n6684, new_n6836);
nor_5  g06460(new_n6836, new_n6835, new_n6837);
and_5  g06461(new_n6592, new_n6591, new_n6838);
nor_5  g06462(new_n6592, new_n6591, new_n6839);
nor_5  g06463(new_n6839, new_n6590, new_n6840);
nor_5  g06464(new_n6840, new_n6838, new_n6841);
nand_5 g06465(n2530, n447, new_n6842);
and_5  g06466(n12777, n7690, new_n6843);
and_5  g06467(n8476, n1353, new_n6844);
xnor_4 g06468(new_n6844, new_n6843, new_n6845);
xnor_4 g06469(new_n6845, new_n6842, new_n6846);
xnor_4 g06470(new_n6846, new_n6841, new_n6847);
xnor_4 g06471(new_n6847, new_n6837, new_n6848);
xnor_4 g06472(new_n6848, new_n6834, new_n6849);
and_5  g06473(n8759, n1198, new_n6850);
and_5  g06474(n11728, n10510, new_n6851);
xnor_4 g06475(new_n6851, new_n6850, new_n6852);
and_5  g06476(n12489, n4499, new_n6853);
and_5  g06477(n10545, n6254, new_n6854);
xnor_4 g06478(new_n6854, new_n6853, new_n6855);
and_5  g06479(n5331, n4436, new_n6856);
and_5  g06480(n12947, n2393, new_n6857);
xnor_4 g06481(new_n6857, new_n6856, new_n6858);
xnor_4 g06482(new_n6858, new_n6855, new_n6859);
xnor_4 g06483(new_n6859, new_n6852, new_n6860_1);
and_5  g06484(n12648, n11967, new_n6861);
and_5  g06485(n7159, n3616, new_n6862);
and_5  g06486(n12709, n10644, new_n6863);
xnor_4 g06487(new_n6863, new_n6862, new_n6864);
xnor_4 g06488(new_n6864, new_n6861, new_n6865);
and_5  g06489(n8819, n8276, new_n6866);
and_5  g06490(n7730, n6776, new_n6867);
xnor_4 g06491(new_n6867, new_n6866, new_n6868);
xnor_4 g06492(new_n6868, new_n6865, new_n6869);
xnor_4 g06493(new_n6869, new_n6860_1, new_n6870);
xnor_4 g06494(new_n6870, new_n6849, new_n6871);
xnor_4 g06495(new_n6871, new_n6823, new_n6872);
nor_5  g06496(new_n6608, new_n6607, new_n6873);
nor_5  g06497(new_n6610, new_n6605, new_n6874);
nor_5  g06498(new_n6874, new_n6873, new_n6875);
and_5  g06499(n12705, n4370, new_n6876);
nor_5  g06500(new_n6420, new_n6415, new_n6877_1);
nor_5  g06501(new_n6430, new_n6421, new_n6878);
nor_5  g06502(new_n6878, new_n6877_1, new_n6879);
nor_5  g06503(new_n6603, new_n6600, new_n6880);
nor_5  g06504(new_n6604_1, new_n6595, new_n6881);
nor_5  g06505(new_n6881, new_n6880, new_n6882);
xnor_4 g06506(new_n6882, new_n6879, new_n6883);
xnor_4 g06507(new_n6883, new_n6876, new_n6884);
xnor_4 g06508(new_n6884, new_n6875, new_n6885);
xnor_4 g06509(new_n6885, new_n6872, new_n6886);
xnor_4 g06510(new_n6886, new_n6809_1, new_n6887);
xnor_4 g06511(new_n6887, new_n6806_1, new_n6888);
xnor_4 g06512(new_n6888, new_n6799, new_n6889);
nor_5  g06513(new_n6710, new_n6624, new_n6890);
nor_5  g06514(new_n6734, new_n6711, new_n6891);
nor_5  g06515(new_n6891, new_n6890, new_n6892);
nor_5  g06516(new_n6532, new_n6531, new_n6893);
nor_5  g06517(new_n6534, new_n6529, new_n6894);
nor_5  g06518(new_n6894, new_n6893, new_n6895);
and_5  g06519(n11407, n10547, new_n6896);
and_5  g06520(n5320, n4312, new_n6897);
xnor_4 g06521(new_n6897, new_n6896, new_n6898);
and_5  g06522(n12299, n8717, new_n6899);
and_5  g06523(n5857, n5760, new_n6900);
xnor_4 g06524(new_n6900, new_n6899, new_n6901);
and_5  g06525(n12025, n11877, new_n6902);
and_5  g06526(n12000, n1097, new_n6903);
xnor_4 g06527(new_n6903, new_n6902, new_n6904);
xnor_4 g06528(new_n6904, new_n6901, new_n6905);
xnor_4 g06529(new_n6905, new_n6898, new_n6906);
nor_5  g06530(new_n6525, new_n6524, new_n6907);
nor_5  g06531(new_n6526, new_n6523, new_n6908);
nor_5  g06532(new_n6908, new_n6907, new_n6909);
nand_5 g06533(n10990, n45, new_n6910);
xnor_4 g06534(new_n6910, new_n6909, new_n6911);
xnor_4 g06535(new_n6911, new_n6906, new_n6912);
and_5  g06536(new_n6521, new_n6520, new_n6913);
nor_5  g06537(new_n6527, new_n6522, new_n6914);
nor_5  g06538(new_n6914, new_n6913, new_n6915);
nand_5 g06539(n7436, n2433, new_n6916);
xnor_4 g06540(new_n6916, new_n6915, new_n6917);
xnor_4 g06541(new_n6917, new_n6912, new_n6918);
nor_5  g06542(new_n6675, new_n6674, new_n6919);
nor_5  g06543(new_n6676, new_n6673, new_n6920);
or_5   g06544(new_n6920, new_n6919, new_n6921);
nor_5  g06545(new_n6518, new_n6513, new_n6922);
nor_5  g06546(new_n6528, new_n6519, new_n6923);
nor_5  g06547(new_n6923, new_n6922, new_n6924);
xnor_4 g06548(new_n6924, new_n6921, new_n6925);
xnor_4 g06549(new_n6925, new_n6918, new_n6926);
xnor_4 g06550(new_n6926, new_n6895, new_n6927);
nor_5  g06551(new_n6694, new_n6693, new_n6928);
nor_5  g06552(new_n6696, new_n6691, new_n6929);
nor_5  g06553(new_n6929, new_n6928, new_n6930);
and_5  g06554(new_n6588, new_n6587, new_n6931);
nor_5  g06555(new_n6594, new_n6589, new_n6932);
nor_5  g06556(new_n6932, new_n6931, new_n6933);
and_5  g06557(n11892, n6441, new_n6934);
and_5  g06558(n11791, n5860, new_n6935);
xnor_4 g06559(new_n6935, new_n6934, new_n6936);
and_5  g06560(n11257, n5212, new_n6937);
and_5  g06561(n6604, n5305, new_n6938);
xnor_4 g06562(new_n6938, new_n6937, new_n6939);
xor_4  g06563(new_n6939, new_n6936, new_n6940);
xnor_4 g06564(new_n6940, new_n6933, new_n6941);
xnor_4 g06565(new_n6941, new_n6930, new_n6942);
xnor_4 g06566(new_n6942, new_n6927, new_n6943);
nor_5  g06567(new_n6423, new_n6422, new_n6944);
nor_5  g06568(new_n6429_1, new_n6424, new_n6945);
or_5   g06569(new_n6945, new_n6944, new_n6946);
nor_5  g06570(new_n6434, new_n6433, new_n6947);
nor_5  g06571(new_n6436, new_n6431_1, new_n6948);
nor_5  g06572(new_n6948, new_n6947, new_n6949);
xnor_4 g06573(new_n6949, new_n6946, new_n6950);
xnor_4 g06574(new_n6950, new_n6943, new_n6951);
xnor_4 g06575(new_n6951, new_n6892, new_n6952);
xnor_4 g06576(new_n6952, new_n6889, new_n6953);
xnor_4 g06577(new_n6953, new_n6786, new_n6954);
xnor_4 g06578(new_n6954, new_n6783, n3287);
xnor_4 g06579(new_n6779, new_n6764, n3339);
xnor_4 g06580(new_n3108, new_n3107, n3456);
and_5  g06581(n6687, n4005, new_n6958);
and_5  g06582(n12720, n6770, new_n6959);
and_5  g06583(n9920, n2509, new_n6960);
and_5  g06584(n6038, n3627, new_n6961);
xor_4  g06585(new_n6961, new_n6960, new_n6962);
xnor_4 g06586(new_n6962, new_n6959, new_n6963);
and_5  g06587(n9920, n6038, new_n6964);
and_5  g06588(n12720, n4189, new_n6965);
nor_5  g06589(new_n6965, new_n6964, new_n6966);
and_5  g06590(n6770, n2509, new_n6967);
xnor_4 g06591(new_n6965, new_n6964, new_n6968);
nor_5  g06592(new_n6968, new_n6967, new_n6969);
nor_5  g06593(new_n6969, new_n6966, new_n6970);
xor_4  g06594(new_n6970, new_n6963, new_n6971);
and_5  g06595(n2564, n2508, new_n6972);
and_5  g06596(n6770, n6038, new_n6973);
and_5  g06597(n4189, n2509, new_n6974);
nor_5  g06598(new_n6974, new_n6973, new_n6975);
and_5  g06599(n12720, n2564, new_n6976);
xnor_4 g06600(new_n6974, new_n6973, new_n6977);
nor_5  g06601(new_n6977, new_n6976, new_n6978);
nor_5  g06602(new_n6978, new_n6975, new_n6979);
and_5  g06603(new_n6979, new_n6972, new_n6980);
xor_4  g06604(new_n6968, new_n6967, new_n6981);
xnor_4 g06605(new_n6979, new_n6972, new_n6982);
nor_5  g06606(new_n6982, new_n6981, new_n6983);
nor_5  g06607(new_n6983, new_n6980, new_n6984);
and_5  g06608(n2585, n2564, new_n6985);
and_5  g06609(n4189, n2508, new_n6986_1);
xnor_4 g06610(new_n6986_1, new_n6985, new_n6987);
xnor_4 g06611(new_n6987, new_n6984, new_n6988);
xnor_4 g06612(new_n6988, new_n6971, new_n6989);
and_5  g06613(n6687, n2585, new_n6990);
nand_5 g06614(n6687, n2508, new_n6991);
and_5  g06615(new_n6965, new_n377, new_n6992);
and_5  g06616(n6038, n4189, new_n6993);
and_5  g06617(n12720, n6687, new_n6994);
nor_5  g06618(new_n6994, new_n6993, new_n6995);
nand_5 g06619(n2564, n2509, new_n6996);
nor_5  g06620(new_n6996, new_n6995, new_n6997);
nor_5  g06621(new_n6997, new_n6992, new_n6998);
nor_5  g06622(new_n6998, new_n6991, new_n6999);
xnor_4 g06623(new_n6998, new_n6991, new_n7000);
xor_4  g06624(new_n6977, new_n6976, new_n7001);
nor_5  g06625(new_n7001, new_n7000, new_n7002);
or_5   g06626(new_n7002, new_n6999, new_n7003);
nor_5  g06627(new_n7003, new_n6990, new_n7004);
xor_4  g06628(new_n6982, new_n6981, new_n7005);
xnor_4 g06629(new_n7003, new_n6990, new_n7006);
nor_5  g06630(new_n7006, new_n7005, new_n7007);
or_5   g06631(new_n7007, new_n7004, new_n7008);
xor_4  g06632(new_n7008, new_n6989, new_n7009);
and_5  g06633(new_n7009, new_n6958, new_n7010);
xnor_4 g06634(new_n7001, new_n7000, new_n7011);
nor_5  g06635(new_n6995, new_n6992, new_n7012);
and_5  g06636(n6687, n2509, new_n7013);
and_5  g06637(n6038, n2564, new_n7014);
nand_5 g06638(new_n7014, new_n7013, new_n7015);
or_5   g06639(new_n7015, new_n7012, new_n7016);
or_5   g06640(new_n7016, new_n7011, new_n7017);
xor_4  g06641(new_n7006, new_n7005, new_n7018);
or_5   g06642(new_n7018, new_n7017, new_n7019);
xnor_4 g06643(new_n7009, new_n6958, new_n7020);
nor_5  g06644(new_n7020, new_n7019, new_n7021);
nor_5  g06645(new_n7021, new_n7010, new_n7022);
or_5   g06646(new_n7008, new_n6989, new_n7023);
nor_5  g06647(new_n6962, new_n6959, new_n7024);
nor_5  g06648(new_n6970, new_n6963, new_n7025);
nor_5  g06649(new_n7025, new_n7024, new_n7026);
and_5  g06650(n4005, n2564, new_n7027);
and_5  g06651(n4189, n2585, new_n7028);
and_5  g06652(n12706, n6687, new_n7029);
xnor_4 g06653(new_n7029, new_n7028, new_n7030);
xnor_4 g06654(new_n7030, new_n7027, new_n7031);
xnor_4 g06655(new_n7031, new_n7026, new_n7032);
and_5  g06656(new_n6961, new_n6960, new_n7033);
and_5  g06657(n6770, n2508, new_n7034);
xnor_4 g06658(new_n7034, new_n7033, new_n7035);
nand_5 g06659(n3627, n2509, new_n7036);
and_5  g06660(n12720, n9920, new_n7037);
and_5  g06661(n6038, n4516, new_n7038);
xnor_4 g06662(new_n7038, new_n7037, new_n7039);
xor_4  g06663(new_n7039, new_n7036, new_n7040);
xnor_4 g06664(new_n7040, new_n7035, new_n7041);
xor_4  g06665(new_n7041, new_n7032, new_n7042);
nor_5  g06666(new_n6987, new_n6984, new_n7043);
nand_5 g06667(new_n6986_1, new_n6985, new_n7044);
or_5   g06668(new_n6988, new_n6971, new_n7045);
xor_4  g06669(new_n7045, new_n7044, new_n7046);
nor_5  g06670(new_n7046, new_n7043, new_n7047);
xnor_4 g06671(new_n7047, new_n7042, new_n7048);
xnor_4 g06672(new_n7048, new_n7023, new_n7049);
xnor_4 g06673(new_n7049, new_n7022, new_n7050);
nand_5 g06674(n8336, n5105, new_n7051);
nand_5 g06675(n10928, n7500, new_n7052);
and_5  g06676(n8336, n1209, new_n7053);
and_5  g06677(n7354, n6986, new_n7054);
nor_5  g06678(new_n7054, new_n7053, new_n7055);
nor_5  g06679(new_n7055, new_n7052, new_n7056);
and_5  g06680(new_n7054, new_n7053, new_n7057);
nor_5  g06681(new_n7057, new_n7056, new_n7058);
xnor_4 g06682(new_n7058, new_n7051, new_n7059);
and_5  g06683(n7500, n6986, new_n7060);
and_5  g06684(n7354, n2226, new_n7061);
and_5  g06685(n10928, n1209, new_n7062);
xnor_4 g06686(new_n7062, new_n7061, new_n7063);
xor_4  g06687(new_n7063, new_n7060, new_n7064);
xnor_4 g06688(new_n7064, new_n7059, new_n7065);
xnor_4 g06689(new_n7054, new_n7053, new_n7066);
and_5  g06690(n10928, n7354, new_n7067);
and_5  g06691(n8336, n7500, new_n7068);
and_5  g06692(new_n7068, new_n7067, new_n7069);
nand_5 g06693(new_n7069, new_n7066, new_n7070);
or_5   g06694(new_n7070, new_n7065, new_n7071);
and_5  g06695(n8336, n4141, new_n7072);
nor_5  g06696(new_n7058, new_n7051, new_n7073);
nor_5  g06697(new_n7064, new_n7059, new_n7074);
or_5   g06698(new_n7074, new_n7073, new_n7075);
xnor_4 g06699(new_n7075, new_n7072, new_n7076);
nand_5 g06700(n10928, n5105, new_n7077);
nor_5  g06701(new_n7062, new_n7061, new_n7078);
and_5  g06702(new_n7062, new_n7061, new_n7079);
nor_5  g06703(new_n7079, new_n7060, new_n7080);
or_5   g06704(new_n7080, new_n7078, new_n7081);
xnor_4 g06705(new_n7081, new_n7077, new_n7082);
and_5  g06706(n6986, n1209, new_n7083);
and_5  g06707(n7354, n1094, new_n7084);
and_5  g06708(n7500, n2226, new_n7085);
xnor_4 g06709(new_n7085, new_n7084, new_n7086);
xor_4  g06710(new_n7086, new_n7083, new_n7087);
xor_4  g06711(new_n7087, new_n7082, new_n7088);
xor_4  g06712(new_n7088, new_n7076, new_n7089);
nor_5  g06713(new_n7089, new_n7071, new_n7090);
and_5  g06714(n8336, n4928, new_n7091);
and_5  g06715(n2226, n1209, new_n7092);
nor_5  g06716(new_n7085, new_n7084, new_n7093);
nor_5  g06717(new_n7086, new_n7083, new_n7094);
nor_5  g06718(new_n7094, new_n7093, new_n7095);
xnor_4 g06719(new_n7095, new_n7092, new_n7096);
and_5  g06720(n7500, n1094, new_n7097);
and_5  g06721(n10678, n7354, new_n7098);
xnor_4 g06722(new_n7098, new_n7097, new_n7099);
xor_4  g06723(new_n7099, new_n7096, new_n7100);
and_5  g06724(n10928, n4141, new_n7101);
and_5  g06725(n6986, n5105, new_n7102);
xor_4  g06726(new_n7102, new_n7101, new_n7103);
xnor_4 g06727(new_n7103, new_n7100, new_n7104);
nor_5  g06728(new_n7081, new_n7077, new_n7105);
nor_5  g06729(new_n7087, new_n7082, new_n7106);
nor_5  g06730(new_n7106, new_n7105, new_n7107);
xnor_4 g06731(new_n7107, new_n7104, new_n7108);
nor_5  g06732(new_n7075, new_n7072, new_n7109);
nor_5  g06733(new_n7088, new_n7076, new_n7110);
or_5   g06734(new_n7110, new_n7109, new_n7111);
xor_4  g06735(new_n7111, new_n7108, new_n7112);
xnor_4 g06736(new_n7112, new_n7091, new_n7113);
xor_4  g06737(new_n7113, new_n7090, new_n7114);
nand_5 g06738(n11222, n7294, new_n7115);
and_5  g06739(n11222, n1980, new_n7116);
and_5  g06740(n8028, n5314, new_n7117);
and_5  g06741(new_n7117, new_n7116, new_n7118);
nor_5  g06742(new_n7117, new_n7116, new_n7119);
nand_5 g06743(n11153, n10848, new_n7120);
nor_5  g06744(new_n7120, new_n7119, new_n7121);
nor_5  g06745(new_n7121, new_n7118, new_n7122);
xor_4  g06746(new_n7122, new_n7115, new_n7123);
and_5  g06747(n10848, n5314, new_n7124);
and_5  g06748(n8028, n996, new_n7125);
and_5  g06749(n11153, n1980, new_n7126);
xnor_4 g06750(new_n7126, new_n7125, new_n7127);
xnor_4 g06751(new_n7127, new_n7124, new_n7128);
xnor_4 g06752(new_n7128, new_n7123, new_n7129);
xor_4  g06753(new_n7117, new_n7116, new_n7130);
and_5  g06754(n11153, n8028, new_n7131);
and_5  g06755(n11222, n10848, new_n7132);
nand_5 g06756(new_n7132, new_n7131, new_n7133);
or_5   g06757(new_n7133, new_n7130, new_n7134);
or_5   g06758(new_n7134, new_n7129, new_n7135);
nor_5  g06759(new_n7122, new_n7115, new_n7136);
and_5  g06760(new_n7128, new_n7123, new_n7137);
or_5   g06761(new_n7137, new_n7136, new_n7138);
and_5  g06762(n12704, n11222, new_n7139);
and_5  g06763(n11153, n7294, new_n7140);
nor_5  g06764(new_n7126, new_n7125, new_n7141);
and_5  g06765(new_n7126, new_n7125, new_n7142);
nor_5  g06766(new_n7142, new_n7124, new_n7143);
nor_5  g06767(new_n7143, new_n7141, new_n7144);
xnor_4 g06768(new_n7144, new_n7140, new_n7145);
and_5  g06769(n10848, n996, new_n7146);
and_5  g06770(n5314, n1980, new_n7147);
and_5  g06771(n8028, n5767, new_n7148);
xnor_4 g06772(new_n7148, new_n7147, new_n7149);
xor_4  g06773(new_n7149, new_n7146, new_n7150);
xor_4  g06774(new_n7150, new_n7145, new_n7151);
xnor_4 g06775(new_n7151, new_n7139, new_n7152);
xor_4  g06776(new_n7152, new_n7138, new_n7153);
or_5   g06777(new_n7153, new_n7135, new_n7154);
and_5  g06778(n11222, n5814, new_n7155);
nand_5 g06779(n1980, n996, new_n7156);
and_5  g06780(n8028, n5319, new_n7157);
and_5  g06781(n10848, n5767, new_n7158);
xnor_4 g06782(new_n7158, new_n7157, new_n7159_1);
xnor_4 g06783(new_n7159_1, new_n7156, new_n7160_1);
nor_5  g06784(new_n7148, new_n7147, new_n7161);
and_5  g06785(new_n7148, new_n7147, new_n7162);
nor_5  g06786(new_n7162, new_n7146, new_n7163);
or_5   g06787(new_n7163, new_n7161, new_n7164);
xnor_4 g06788(new_n7164, new_n7160_1, new_n7165);
and_5  g06789(n12704, n11153, new_n7166);
and_5  g06790(n7294, n5314, new_n7167);
xnor_4 g06791(new_n7167, new_n7166, new_n7168);
xnor_4 g06792(new_n7168, new_n7165, new_n7169);
and_5  g06793(new_n7144, new_n7140, new_n7170);
nor_5  g06794(new_n7150, new_n7145, new_n7171);
nor_5  g06795(new_n7171, new_n7170, new_n7172);
xnor_4 g06796(new_n7172, new_n7169, new_n7173);
nor_5  g06797(new_n7151, new_n7139, new_n7174);
nor_5  g06798(new_n7152, new_n7138, new_n7175);
or_5   g06799(new_n7175, new_n7174, new_n7176);
xor_4  g06800(new_n7176, new_n7173, new_n7177);
xnor_4 g06801(new_n7177, new_n7155, new_n7178);
xor_4  g06802(new_n7178, new_n7154, new_n7179);
nand_5 g06803(n12069, n2802, new_n7180);
and_5  g06804(n7891, n1564, new_n7181);
and_5  g06805(n12069, n533, new_n7182);
nor_5  g06806(new_n7182, new_n7181, new_n7183);
nand_5 g06807(n12391, n1512, new_n7184);
or_5   g06808(new_n7184, new_n7183, new_n7185);
nand_5 g06809(new_n7182, new_n7181, new_n7186);
and_5  g06810(new_n7186, new_n7185, new_n7187);
xnor_4 g06811(new_n7187, new_n7180, new_n7188);
and_5  g06812(n7891, n1512, new_n7189);
and_5  g06813(n7160, n1564, new_n7190);
and_5  g06814(n12391, n533, new_n7191);
xnor_4 g06815(new_n7191, new_n7190, new_n7192);
xor_4  g06816(new_n7192, new_n7189, new_n7193_1);
xnor_4 g06817(new_n7193_1, new_n7188, new_n7194);
xor_4  g06818(new_n7182, new_n7181, new_n7195);
and_5  g06819(n12391, n1564, new_n7196);
and_5  g06820(n12069, n1512, new_n7197);
nand_5 g06821(new_n7197, new_n7196, new_n7198);
or_5   g06822(new_n7198, new_n7195, new_n7199);
or_5   g06823(new_n7199, new_n7194, new_n7200);
and_5  g06824(n12069, n6806, new_n7201);
and_5  g06825(n12391, n2802, new_n7202);
nor_5  g06826(new_n7191, new_n7190, new_n7203);
nor_5  g06827(new_n7192, new_n7189, new_n7204);
nor_5  g06828(new_n7204, new_n7203, new_n7205);
xnor_4 g06829(new_n7205, new_n7202, new_n7206);
and_5  g06830(n7891, n533, new_n7207);
and_5  g06831(n4828, n1564, new_n7208);
and_5  g06832(n7160, n1512, new_n7209);
xnor_4 g06833(new_n7209, new_n7208, new_n7210);
xor_4  g06834(new_n7210, new_n7207, new_n7211);
xor_4  g06835(new_n7211, new_n7206, new_n7212);
xnor_4 g06836(new_n7212, new_n7201, new_n7213);
nor_5  g06837(new_n7187, new_n7180, new_n7214);
nor_5  g06838(new_n7193_1, new_n7188, new_n7215);
or_5   g06839(new_n7215, new_n7214, new_n7216);
xor_4  g06840(new_n7216, new_n7213, new_n7217);
or_5   g06841(new_n7217, new_n7200, new_n7218);
and_5  g06842(n12069, n5069, new_n7219);
nand_5 g06843(n7160, n533, new_n7220);
and_5  g06844(n2515, n1564, new_n7221);
and_5  g06845(n4828, n1512, new_n7222);
xnor_4 g06846(new_n7222, new_n7221, new_n7223);
xnor_4 g06847(new_n7223, new_n7220, new_n7224);
nor_5  g06848(new_n7209, new_n7208, new_n7225);
nor_5  g06849(new_n7210, new_n7207, new_n7226);
or_5   g06850(new_n7226, new_n7225, new_n7227);
xnor_4 g06851(new_n7227, new_n7224, new_n7228);
and_5  g06852(n7891, n2802, new_n7229);
and_5  g06853(n12391, n6806, new_n7230);
xnor_4 g06854(new_n7230, new_n7229, new_n7231);
xnor_4 g06855(new_n7231, new_n7228, new_n7232);
and_5  g06856(new_n7205, new_n7202, new_n7233);
nor_5  g06857(new_n7211, new_n7206, new_n7234);
nor_5  g06858(new_n7234, new_n7233, new_n7235);
xnor_4 g06859(new_n7235, new_n7232, new_n7236_1);
nor_5  g06860(new_n7212, new_n7201, new_n7237);
nor_5  g06861(new_n7216, new_n7213, new_n7238);
or_5   g06862(new_n7238, new_n7237, new_n7239);
xor_4  g06863(new_n7239, new_n7236_1, new_n7240);
xor_4  g06864(new_n7240, new_n7219, new_n7241);
xnor_4 g06865(new_n7241, new_n7218, new_n7242);
xnor_4 g06866(new_n7242, new_n7179, new_n7243);
xor_4  g06867(new_n7153, new_n7135, new_n7244);
xor_4  g06868(new_n7199, new_n7194, new_n7245);
xor_4  g06869(new_n7134, new_n7129, new_n7246);
nor_5  g06870(new_n7246, new_n7245, new_n7247);
nor_5  g06871(new_n7184, new_n380, new_n7248);
nor_5  g06872(new_n7248, new_n7195, new_n7249);
nor_5  g06873(new_n7185, new_n380, new_n7250);
or_5   g06874(new_n7250, new_n7249, new_n7251);
nor_5  g06875(new_n7120, new_n379, new_n7252);
nor_5  g06876(new_n7252, new_n7130, new_n7253);
or_5   g06877(new_n7120, new_n379, new_n7254);
nor_5  g06878(new_n7254, new_n7119, new_n7255);
or_5   g06879(new_n7255, new_n7253, new_n7256);
nor_5  g06880(new_n7256, new_n7251, new_n7257);
and_5  g06881(new_n380, new_n379, new_n7258);
xor_4  g06882(new_n7132, new_n7131, new_n7259);
nor_5  g06883(new_n7259, new_n7258, new_n7260);
xnor_4 g06884(new_n7259, new_n7258, new_n7261);
xor_4  g06885(new_n7197, new_n7196, new_n7262);
nor_5  g06886(new_n7262, new_n7261, new_n7263);
nor_5  g06887(new_n7263, new_n7260, new_n7264);
xor_4  g06888(new_n7256, new_n7251, new_n7265_1);
and_5  g06889(new_n7265_1, new_n7264, new_n7266);
or_5   g06890(new_n7266, new_n7257, new_n7267);
xnor_4 g06891(new_n7246, new_n7245, new_n7268);
nor_5  g06892(new_n7268, new_n7267, new_n7269);
nor_5  g06893(new_n7269, new_n7247, new_n7270_1);
nor_5  g06894(new_n7270_1, new_n7244, new_n7271);
xor_4  g06895(new_n7217, new_n7200, new_n7272);
xnor_4 g06896(new_n7270_1, new_n7244, new_n7273);
nor_5  g06897(new_n7273, new_n7272, new_n7274);
nor_5  g06898(new_n7274, new_n7271, new_n7275);
xor_4  g06899(new_n7275, new_n7243, new_n7276);
nor_5  g06900(new_n7276, new_n7114, new_n7277);
xnor_4 g06901(new_n7276, new_n7114, new_n7278);
xnor_4 g06902(new_n7089, new_n7071, new_n7279);
xor_4  g06903(new_n7273, new_n7272, new_n7280);
nor_5  g06904(new_n7280, new_n7279, new_n7281);
xnor_4 g06905(new_n7280, new_n7279, new_n7282);
xnor_4 g06906(new_n7070, new_n7065, new_n7283);
xor_4  g06907(new_n7268, new_n7267, new_n7284);
nor_5  g06908(new_n7284, new_n7283, new_n7285);
xnor_4 g06909(new_n7284, new_n7283, new_n7286);
xor_4  g06910(new_n7265_1, new_n7264, new_n7287);
nor_5  g06911(new_n7052, new_n378, new_n7288);
and_5  g06912(new_n7288, new_n7055, new_n7289);
nor_5  g06913(new_n7288, new_n7066, new_n7290);
or_5   g06914(new_n7290, new_n7289, new_n7291);
nor_5  g06915(new_n7291, new_n7287, new_n7292);
xor_4  g06916(new_n7291, new_n7287, new_n7293);
xor_4  g06917(new_n7262, new_n7261, new_n7294_1);
xnor_4 g06918(new_n7068, new_n7067, new_n7295);
nor_5  g06919(new_n7295, new_n7294_1, new_n7296);
nand_5 g06920(n8336, n7354, new_n7297);
or_5   g06921(new_n381_1, new_n7297, new_n7298);
xnor_4 g06922(new_n7295, new_n7294_1, new_n7299);
nor_5  g06923(new_n7299, new_n7298, new_n7300);
nor_5  g06924(new_n7300, new_n7296, new_n7301);
and_5  g06925(new_n7301, new_n7293, new_n7302);
or_5   g06926(new_n7302, new_n7292, new_n7303);
nor_5  g06927(new_n7303, new_n7286, new_n7304);
nor_5  g06928(new_n7304, new_n7285, new_n7305);
nor_5  g06929(new_n7305, new_n7282, new_n7306);
nor_5  g06930(new_n7306, new_n7281, new_n7307);
nor_5  g06931(new_n7307, new_n7278, new_n7308);
or_5   g06932(new_n7308, new_n7277, new_n7309);
or_5   g06933(new_n7111, new_n7108, new_n7310);
and_5  g06934(new_n7095, new_n7092, new_n7311);
nor_5  g06935(new_n7099, new_n7096, new_n7312);
or_5   g06936(new_n7312, new_n7311, new_n7313);
and_5  g06937(n10928, n4928, new_n7314);
and_5  g06938(n6986, n4141, new_n7315);
and_5  g06939(n8336, n8236, new_n7316);
xnor_4 g06940(new_n7316, new_n7315, new_n7317);
xnor_4 g06941(new_n7317, new_n7314, new_n7318);
xnor_4 g06942(new_n7318, new_n7313, new_n7319);
and_5  g06943(new_n7098, new_n7097, new_n7320_1);
and_5  g06944(n5105, n2226, new_n7321);
xnor_4 g06945(new_n7321, new_n7320_1, new_n7322);
and_5  g06946(n10678, n7500, new_n7323);
and_5  g06947(n7354, n7320, new_n7324);
and_5  g06948(n1209, n1094, new_n7325);
xnor_4 g06949(new_n7325, new_n7324, new_n7326);
xor_4  g06950(new_n7326, new_n7323, new_n7327);
xor_4  g06951(new_n7327, new_n7322, new_n7328);
xor_4  g06952(new_n7328, new_n7319, new_n7329);
and_5  g06953(new_n7103, new_n7100, new_n7330);
nand_5 g06954(new_n7102, new_n7101, new_n7331);
or_5   g06955(new_n7107, new_n7104, new_n7332);
xor_4  g06956(new_n7332, new_n7331, new_n7333);
nor_5  g06957(new_n7333, new_n7330, new_n7334);
xnor_4 g06958(new_n7334, new_n7329, new_n7335);
xnor_4 g06959(new_n7335, new_n7310, new_n7336);
nor_5  g06960(new_n7112, new_n7091, new_n7337);
nor_5  g06961(new_n7113, new_n7090, new_n7338);
or_5   g06962(new_n7338, new_n7337, new_n7339);
xor_4  g06963(new_n7339, new_n7336, new_n7340);
or_5   g06964(new_n7176, new_n7173, new_n7341);
nor_5  g06965(new_n7159_1, new_n7156, new_n7342);
nor_5  g06966(new_n7164, new_n7160_1, new_n7343);
or_5   g06967(new_n7343, new_n7342, new_n7344);
and_5  g06968(n11153, n5814, new_n7345);
and_5  g06969(n12704, n5314, new_n7346);
and_5  g06970(n11222, n4903, new_n7347);
xnor_4 g06971(new_n7347, new_n7346, new_n7348);
xnor_4 g06972(new_n7348, new_n7345, new_n7349);
xnor_4 g06973(new_n7349, new_n7344, new_n7350);
and_5  g06974(new_n7158, new_n7157, new_n7351);
and_5  g06975(n7294, n996, new_n7352);
xnor_4 g06976(new_n7352, new_n7351, new_n7353);
and_5  g06977(n10848, n5319, new_n7354_1);
and_5  g06978(n5767, n1980, new_n7355);
and_5  g06979(n9457, n8028, new_n7356);
xnor_4 g06980(new_n7356, new_n7355, new_n7357);
xor_4  g06981(new_n7357, new_n7354_1, new_n7358);
xor_4  g06982(new_n7358, new_n7353, new_n7359);
xor_4  g06983(new_n7359, new_n7350, new_n7360);
nor_5  g06984(new_n7168, new_n7165, new_n7361);
nand_5 g06985(new_n7167, new_n7166, new_n7362);
or_5   g06986(new_n7172, new_n7169, new_n7363);
xor_4  g06987(new_n7363, new_n7362, new_n7364);
nor_5  g06988(new_n7364, new_n7361, new_n7365);
xnor_4 g06989(new_n7365, new_n7360, new_n7366);
xnor_4 g06990(new_n7366, new_n7341, new_n7367);
and_5  g06991(new_n7177, new_n7155, new_n7368);
nor_5  g06992(new_n7178, new_n7154, new_n7369);
nor_5  g06993(new_n7369, new_n7368, new_n7370);
xor_4  g06994(new_n7370, new_n7367, new_n7371);
or_5   g06995(new_n7239, new_n7236_1, new_n7372);
nor_5  g06996(new_n7231, new_n7228, new_n7373);
nand_5 g06997(new_n7230, new_n7229, new_n7374);
or_5   g06998(new_n7235, new_n7232, new_n7375);
xor_4  g06999(new_n7375, new_n7374, new_n7376);
nor_5  g07000(new_n7376, new_n7373, new_n7377);
and_5  g07001(new_n7222, new_n7221, new_n7378);
and_5  g07002(n7160, n2802, new_n7379);
xnor_4 g07003(new_n7379, new_n7378, new_n7380);
nand_5 g07004(n2515, n1512, new_n7381);
and_5  g07005(n1564, n1199, new_n7382);
and_5  g07006(n4828, n533, new_n7383);
xnor_4 g07007(new_n7383, new_n7382, new_n7384);
xnor_4 g07008(new_n7384, new_n7381, new_n7385);
xor_4  g07009(new_n7385, new_n7380, new_n7386);
nor_5  g07010(new_n7223, new_n7220, new_n7387);
nor_5  g07011(new_n7227, new_n7224, new_n7388_1);
or_5   g07012(new_n7388_1, new_n7387, new_n7389);
and_5  g07013(n12391, n5069, new_n7390);
and_5  g07014(n7891, n6806, new_n7391);
and_5  g07015(n12069, n12044, new_n7392);
xnor_4 g07016(new_n7392, new_n7391, new_n7393);
xnor_4 g07017(new_n7393, new_n7390, new_n7394);
xnor_4 g07018(new_n7394, new_n7389, new_n7395);
xor_4  g07019(new_n7395, new_n7386, new_n7396);
xnor_4 g07020(new_n7396, new_n7377, new_n7397);
xnor_4 g07021(new_n7397, new_n7372, new_n7398);
and_5  g07022(new_n7240, new_n7219, new_n7399);
nor_5  g07023(new_n7240, new_n7219, new_n7400);
nor_5  g07024(new_n7400, new_n7218, new_n7401);
nor_5  g07025(new_n7401, new_n7399, new_n7402);
xor_4  g07026(new_n7402, new_n7398, new_n7403);
nor_5  g07027(new_n7242, new_n7179, new_n7404);
nor_5  g07028(new_n7275, new_n7243, new_n7405);
nor_5  g07029(new_n7405, new_n7404, new_n7406);
xnor_4 g07030(new_n7406, new_n7403, new_n7407);
xnor_4 g07031(new_n7407, new_n7371, new_n7408);
xnor_4 g07032(new_n7408, new_n7340, new_n7409);
xor_4  g07033(new_n7409, new_n7309, new_n7410);
and_5  g07034(new_n7410, new_n7050, new_n7411);
xor_4  g07035(new_n7020, new_n7019, new_n7412);
xor_4  g07036(new_n7018, new_n7017, new_n7413);
xor_4  g07037(new_n7305, new_n7282, new_n7414);
nor_5  g07038(new_n7414, new_n7413, new_n7415);
xor_4  g07039(new_n7016, new_n7011, new_n7416);
xor_4  g07040(new_n7303, new_n7286, new_n7417);
nor_5  g07041(new_n7417, new_n7416, new_n7418);
xnor_4 g07042(new_n7417, new_n7416, new_n7419);
xnor_4 g07043(new_n7301, new_n7293, new_n7420);
nor_5  g07044(new_n6996, new_n377, new_n7421);
nor_5  g07045(new_n7421, new_n7012, new_n7422);
or_5   g07046(new_n6996, new_n377, new_n7423);
nor_5  g07047(new_n7423, new_n6995, new_n7424);
nor_5  g07048(new_n7424, new_n7422, new_n7425);
nor_5  g07049(new_n7425, new_n7420, new_n7426);
xnor_4 g07050(new_n7425, new_n7420, new_n7427);
and_5  g07051(new_n382, new_n377, new_n7428);
xor_4  g07052(new_n7014, new_n7013, new_n7429);
nor_5  g07053(new_n7429, new_n7428, new_n7430);
xnor_4 g07054(new_n7299, new_n7298, new_n7431);
xor_4  g07055(new_n7429, new_n7428, new_n7432);
and_5  g07056(new_n7432, new_n7431, new_n7433);
nor_5  g07057(new_n7433, new_n7430, new_n7434);
nor_5  g07058(new_n7434, new_n7427, new_n7435);
nor_5  g07059(new_n7435, new_n7426, new_n7436_1);
nor_5  g07060(new_n7436_1, new_n7419, new_n7437);
or_5   g07061(new_n7437, new_n7418, new_n7438);
xor_4  g07062(new_n7414, new_n7413, new_n7439);
and_5  g07063(new_n7439, new_n7438, new_n7440);
nor_5  g07064(new_n7440, new_n7415, new_n7441);
nor_5  g07065(new_n7441, new_n7412, new_n7442);
xnor_4 g07066(new_n7307, new_n7278, new_n7443);
xor_4  g07067(new_n7441, new_n7412, new_n7444);
and_5  g07068(new_n7444, new_n7443, new_n7445);
nor_5  g07069(new_n7445, new_n7442, new_n7446);
xnor_4 g07070(new_n7410, new_n7050, new_n7447);
nor_5  g07071(new_n7447, new_n7446, new_n7448);
nor_5  g07072(new_n7448, new_n7411, new_n7449);
nor_5  g07073(new_n7406, new_n7403, new_n7450);
nor_5  g07074(new_n7407, new_n7371, new_n7451);
nor_5  g07075(new_n7451, new_n7450, new_n7452);
nor_5  g07076(new_n7408, new_n7340, new_n7453);
nor_5  g07077(new_n7409, new_n7309, new_n7454);
nor_5  g07078(new_n7454, new_n7453, new_n7455);
xnor_4 g07079(new_n7455, new_n7452, new_n7456_1);
nor_5  g07080(new_n7335, new_n7310, new_n7457);
nor_5  g07081(new_n7339, new_n7336, new_n7458);
nor_5  g07082(new_n7458, new_n7457, new_n7459);
nor_5  g07083(new_n7375, new_n7374, new_n7460);
nor_5  g07084(new_n7396, new_n7377, new_n7461);
nor_5  g07085(new_n7461, new_n7460, new_n7462);
and_5  g07086(new_n7352, new_n7351, new_n7463);
nor_5  g07087(new_n7358, new_n7353, new_n7464);
nor_5  g07088(new_n7464, new_n7463, new_n7465);
and_5  g07089(new_n7383, new_n7382, new_n7466);
nor_5  g07090(new_n7383, new_n7382, new_n7467);
nor_5  g07091(new_n7467, new_n7381, new_n7468);
or_5   g07092(new_n7468, new_n7466, new_n7469);
xnor_4 g07093(new_n7469, new_n7465, new_n7470);
and_5  g07094(n8028, n4817, new_n7471);
and_5  g07095(n7523, n7354, new_n7472);
xor_4  g07096(new_n7472, new_n7471, new_n7473);
and_5  g07097(n10848, n9457, new_n7474);
and_5  g07098(n11222, n1906, new_n7475);
xnor_4 g07099(new_n7475, new_n7474, new_n7476);
and_5  g07100(n6986, n4928, new_n7477);
and_5  g07101(n4141, n2226, new_n7478);
xnor_4 g07102(new_n7478, new_n7477, new_n7479);
xnor_4 g07103(new_n7479, new_n7476, new_n7480);
xnor_4 g07104(new_n7480, new_n7473, new_n7481);
and_5  g07105(new_n7038, new_n7037, new_n7482);
nor_5  g07106(new_n7038, new_n7037, new_n7483);
nor_5  g07107(new_n7483, new_n7036, new_n7484);
nor_5  g07108(new_n7484, new_n7482, new_n7485);
nand_5 g07109(n4516, n2509, new_n7486);
and_5  g07110(n12704, n996, new_n7487);
and_5  g07111(n12720, n3627, new_n7488);
xnor_4 g07112(new_n7488, new_n7487, new_n7489);
xnor_4 g07113(new_n7489, new_n7486, new_n7490);
xnor_4 g07114(new_n7490, new_n7485, new_n7491);
xnor_4 g07115(new_n7491, new_n7481, new_n7492);
nand_5 g07116(n2515, n533, new_n7493);
and_5  g07117(n1512, n1199, new_n7494);
and_5  g07118(n12391, n12044, new_n7495);
xnor_4 g07119(new_n7495, new_n7494, new_n7496);
xnor_4 g07120(new_n7496, new_n7493, new_n7497);
xnor_4 g07121(new_n7497, new_n7492, new_n7498);
xnor_4 g07122(new_n7498, new_n7470, new_n7499);
nor_5  g07123(new_n7349, new_n7344, new_n7500_1);
nor_5  g07124(new_n7359, new_n7350, new_n7501);
nor_5  g07125(new_n7501, new_n7500_1, new_n7502);
nor_5  g07126(new_n7356, new_n7355, new_n7503);
nor_5  g07127(new_n7357, new_n7354_1, new_n7504);
nor_5  g07128(new_n7504, new_n7503, new_n7505);
and_5  g07129(n12069, n5694, new_n7506);
and_5  g07130(n11153, n4903, new_n7507);
xnor_4 g07131(new_n7507, new_n7506, new_n7508);
and_5  g07132(n7294, n5767, new_n7509);
and_5  g07133(n8336, n783, new_n7510);
xnor_4 g07134(new_n7510, new_n7509, new_n7511);
xnor_4 g07135(new_n7511, new_n7508, new_n7512);
xnor_4 g07136(new_n7512, new_n7505, new_n7513);
and_5  g07137(n4189, n4005, new_n7514);
and_5  g07138(n5814, n5314, new_n7515);
xnor_4 g07139(new_n7515, new_n7514, new_n7516);
xnor_4 g07140(new_n7516, new_n7513, new_n7517);
xnor_4 g07141(new_n7517, new_n7502, new_n7518);
xnor_4 g07142(new_n7518, new_n7499, new_n7519);
xnor_4 g07143(new_n7519, new_n7462, new_n7520);
xnor_4 g07144(new_n7520, new_n7459, new_n7521);
nor_5  g07145(new_n7397, new_n7372, new_n7522);
nor_5  g07146(new_n7402, new_n7398, new_n7523_1);
or_5   g07147(new_n7523_1, new_n7522, new_n7524);
nor_5  g07148(new_n7366, new_n7341, new_n7525);
nor_5  g07149(new_n7370, new_n7367, new_n7526);
nor_5  g07150(new_n7526, new_n7525, new_n7527);
nor_5  g07151(new_n7031, new_n7026, new_n7528);
nor_5  g07152(new_n7041, new_n7032, new_n7529);
nor_5  g07153(new_n7529, new_n7528, new_n7530);
nor_5  g07154(new_n7029, new_n7028, new_n7531);
nor_5  g07155(new_n7030, new_n7027, new_n7532);
nor_5  g07156(new_n7532, new_n7531, new_n7533);
xnor_4 g07157(new_n7533, new_n7530, new_n7534);
nor_5  g07158(new_n7347, new_n7346, new_n7535);
nor_5  g07159(new_n7348, new_n7345, new_n7536);
nor_5  g07160(new_n7536, new_n7535, new_n7537);
nor_5  g07161(new_n7392, new_n7391, new_n7538);
nor_5  g07162(new_n7393, new_n7390, new_n7539);
nor_5  g07163(new_n7539, new_n7538, new_n7540);
xnor_4 g07164(new_n7540, new_n7537, new_n7541);
xnor_4 g07165(new_n7541, new_n7534, new_n7542);
xnor_4 g07166(new_n7542, new_n7527, new_n7543);
nor_5  g07167(new_n7048, new_n7023, new_n7544);
nor_5  g07168(new_n7049, new_n7022, new_n7545);
nor_5  g07169(new_n7545, new_n7544, new_n7546_1);
nor_5  g07170(new_n7394, new_n7389, new_n7547);
nor_5  g07171(new_n7395, new_n7386, new_n7548);
nor_5  g07172(new_n7548, new_n7547, new_n7549);
nand_5 g07173(n6578, n1564, new_n7550);
xnor_4 g07174(new_n7550, new_n7549, new_n7551);
xnor_4 g07175(new_n7551, new_n7546_1, new_n7552);
xnor_4 g07176(new_n7552, new_n7543, new_n7553);
nor_5  g07177(new_n7363, new_n7362, new_n7554);
nor_5  g07178(new_n7365, new_n7360, new_n7555);
nor_5  g07179(new_n7555, new_n7554, new_n7556);
and_5  g07180(new_n7321, new_n7320_1, new_n7557);
nor_5  g07181(new_n7327, new_n7322, new_n7558);
nor_5  g07182(new_n7558, new_n7557, new_n7559);
nor_5  g07183(new_n7316, new_n7315, new_n7560);
nor_5  g07184(new_n7317, new_n7314, new_n7561);
nor_5  g07185(new_n7561, new_n7560, new_n7562);
and_5  g07186(n5319, n1980, new_n7563);
and_5  g07187(n9920, n2508, new_n7564);
and_5  g07188(n10678, n1209, new_n7565);
xnor_4 g07189(new_n7565, new_n7564, new_n7566);
xnor_4 g07190(new_n7566, new_n7563, new_n7567);
xnor_4 g07191(new_n7567, new_n7562, new_n7568_1);
xnor_4 g07192(new_n7568_1, new_n7559, new_n7569);
xnor_4 g07193(new_n7569, new_n7556, new_n7570);
nor_5  g07194(new_n7318, new_n7313, new_n7571);
nor_5  g07195(new_n7328, new_n7319, new_n7572);
nor_5  g07196(new_n7572, new_n7571, new_n7573);
nor_5  g07197(new_n7325, new_n7324, new_n7574);
nor_5  g07198(new_n7326, new_n7323, new_n7575);
nor_5  g07199(new_n7575, new_n7574, new_n7576);
and_5  g07200(n4828, n2802, new_n7577);
and_5  g07201(n10928, n8236, new_n7578);
and_5  g07202(n5105, n1094, new_n7579);
xnor_4 g07203(new_n7579, new_n7578, new_n7580);
xnor_4 g07204(new_n7580, new_n7577, new_n7581);
xnor_4 g07205(new_n7581, new_n7576, new_n7582);
xnor_4 g07206(new_n7582, new_n7573, new_n7583);
xnor_4 g07207(new_n7583, new_n7570, new_n7584);
and_5  g07208(new_n7379, new_n7378, new_n7585);
nor_5  g07209(new_n7385, new_n7380, new_n7586);
nor_5  g07210(new_n7586, new_n7585, new_n7587);
and_5  g07211(n7891, n5069, new_n7588);
and_5  g07212(n6038, n2087, new_n7589);
xor_4  g07213(new_n7589, new_n7588, new_n7590);
xnor_4 g07214(new_n7590, new_n7587, new_n7591);
and_5  g07215(n7160, n6806, new_n7592);
and_5  g07216(n6687, n615, new_n7593);
xor_4  g07217(new_n7593, new_n7592, new_n7594);
xnor_4 g07218(new_n7594, new_n7591, new_n7595);
xnor_4 g07219(new_n7595, new_n7584, new_n7596);
nor_5  g07220(new_n7045, new_n7044, new_n7597);
nor_5  g07221(new_n7047, new_n7042, new_n7598);
or_5   g07222(new_n7598, new_n7597, new_n7599);
nor_5  g07223(new_n7332, new_n7331, new_n7600);
nor_5  g07224(new_n7334, new_n7329, new_n7601);
nor_5  g07225(new_n7601, new_n7600, new_n7602);
nor_5  g07226(new_n7034, new_n7033, new_n7603);
nor_5  g07227(new_n7040, new_n7035, new_n7604);
nor_5  g07228(new_n7604, new_n7603, new_n7605);
and_5  g07229(n7500, n7320, new_n7606);
and_5  g07230(n12706, n2564, new_n7607);
and_5  g07231(n6770, n2585, new_n7608);
xnor_4 g07232(new_n7608, new_n7607, new_n7609);
xnor_4 g07233(new_n7609, new_n7606, new_n7610_1);
xnor_4 g07234(new_n7610_1, new_n7605, new_n7611);
xnor_4 g07235(new_n7611, new_n7602, new_n7612);
xnor_4 g07236(new_n7612, new_n7599, new_n7613);
xnor_4 g07237(new_n7613, new_n7596, new_n7614);
xnor_4 g07238(new_n7614, new_n7553, new_n7615);
xnor_4 g07239(new_n7615, new_n7524, new_n7616);
xnor_4 g07240(new_n7616, new_n7521, new_n7617);
xnor_4 g07241(new_n7617, new_n7456_1, new_n7618);
xnor_4 g07242(new_n7618, new_n7449, n3654);
xnor_4 g07243(new_n7444, new_n7443, n3661);
nand_5 g07244(n7456, n5305, new_n7621);
nand_5 g07245(n5964, n3932, new_n7622);
and_5  g07246(n1798, n1097, new_n7623);
and_5  g07247(n12591, n5305, new_n7624);
nor_5  g07248(new_n7624, new_n7623, new_n7625);
nor_5  g07249(new_n7625, new_n7622, new_n7626);
and_5  g07250(new_n7624, new_n7623, new_n7627);
nor_5  g07251(new_n7627, new_n7626, new_n7628);
xnor_4 g07252(new_n7628, new_n7621, new_n7629);
and_5  g07253(n3932, n1097, new_n7630);
and_5  g07254(n4312, n1798, new_n7631);
and_5  g07255(n12591, n5964, new_n7632);
xnor_4 g07256(new_n7632, new_n7631, new_n7633);
xor_4  g07257(new_n7633, new_n7630, new_n7634);
xnor_4 g07258(new_n7634, new_n7629, new_n7635);
and_5  g07259(new_n4833, new_n4832, new_n7636);
xnor_4 g07260(new_n7624, new_n7623, new_n7637);
nand_5 g07261(new_n7637, new_n7636, new_n7638);
or_5   g07262(new_n7638, new_n7635, new_n7639);
nand_5 g07263(n11662, n5305, new_n7640);
nand_5 g07264(n7456, n5964, new_n7641);
and_5  g07265(n4312, n3932, new_n7642);
and_5  g07266(n12591, n1097, new_n7643);
and_5  g07267(n12705, n1798, new_n7644);
xnor_4 g07268(new_n7644, new_n7643, new_n7645);
xor_4  g07269(new_n7645, new_n7642, new_n7646_1);
xnor_4 g07270(new_n7646_1, new_n7641, new_n7647);
nor_5  g07271(new_n7632, new_n7631, new_n7648);
nor_5  g07272(new_n7633, new_n7630, new_n7649);
or_5   g07273(new_n7649, new_n7648, new_n7650);
xnor_4 g07274(new_n7650, new_n7647, new_n7651);
xnor_4 g07275(new_n7651, new_n7640, new_n7652);
nor_5  g07276(new_n7628, new_n7621, new_n7653);
nor_5  g07277(new_n7634, new_n7629, new_n7654);
nor_5  g07278(new_n7654, new_n7653, new_n7655);
xnor_4 g07279(new_n7655, new_n7652, new_n7656);
xnor_4 g07280(new_n7656, new_n7639, new_n7657);
xnor_4 g07281(new_n7638, new_n7635, new_n7658);
nand_5 g07282(n11023, n8759, new_n7659);
and_5  g07283(n8759, n3022, new_n7660);
and_5  g07284(n12299, n6703, new_n7661);
nor_5  g07285(new_n7661, new_n7660, new_n7662);
and_5  g07286(n8759, n6703, new_n7663);
and_5  g07287(n12299, n3022, new_n7664);
and_5  g07288(new_n7664, new_n7663, new_n7665);
and_5  g07289(n9640, n6776, new_n7666);
nor_5  g07290(new_n7666, new_n7665, new_n7667);
or_5   g07291(new_n7667, new_n7662, new_n7668);
xnor_4 g07292(new_n7668, new_n7659, new_n7669);
and_5  g07293(n12299, n9640, new_n7670);
and_5  g07294(n6776, n3022, new_n7671);
and_5  g07295(n7436, n6703, new_n7672);
xnor_4 g07296(new_n7672, new_n7671, new_n7673);
xor_4  g07297(new_n7673, new_n7670, new_n7674);
xnor_4 g07298(new_n7674, new_n7669, new_n7675);
nand_5 g07299(n9640, n6776, new_n7676_1);
or_5   g07300(new_n7676_1, new_n7663, new_n7677);
or_5   g07301(new_n7665, new_n7662, new_n7678);
nand_5 g07302(new_n7678, new_n7677, new_n7679);
or_5   g07303(new_n7679, new_n7676_1, new_n7680);
xor_4  g07304(new_n7680, new_n7675, new_n7681);
nand_5 g07305(n11922, n5331, new_n7682);
and_5  g07306(n2530, n1067, new_n7683);
and_5  g07307(n8665, n8476, new_n7684);
and_5  g07308(n12648, n5645, new_n7685);
xnor_4 g07309(new_n7685, new_n7684, new_n7686);
xor_4  g07310(new_n7686, new_n7683, new_n7687);
xnor_4 g07311(new_n7687, new_n7682, new_n7688);
and_5  g07312(n8665, n5331, new_n7689);
and_5  g07313(n5645, n2530, new_n7690_1);
nor_5  g07314(new_n7690_1, new_n7689, new_n7691);
and_5  g07315(n8476, n1067, new_n7692);
and_5  g07316(n8665, n2530, new_n7693);
and_5  g07317(new_n7693, new_n4827, new_n7694);
nor_5  g07318(new_n7694, new_n7692, new_n7695);
or_5   g07319(new_n7695, new_n7691, new_n7696);
xnor_4 g07320(new_n7696, new_n7688, new_n7697);
nand_5 g07321(new_n4847, new_n4846, new_n7698);
nor_5  g07322(new_n7694, new_n7691, new_n7699);
or_5   g07323(new_n7699, new_n7698, new_n7700);
xor_4  g07324(new_n7700, new_n7697, new_n7701);
and_5  g07325(n7965, n2749, new_n7702);
and_5  g07326(n7965, n3754, new_n7703);
and_5  g07327(n11892, n11876, new_n7704);
nor_5  g07328(new_n7704, new_n7703, new_n7705);
and_5  g07329(n11892, n3754, new_n7706);
and_5  g07330(new_n7706, new_n4828_1, new_n7707);
and_5  g07331(n10898, n7388, new_n7708);
nor_5  g07332(new_n7708, new_n7707, new_n7709);
nor_5  g07333(new_n7709, new_n7705, new_n7710);
xnor_4 g07334(new_n7710, new_n7702, new_n7711);
and_5  g07335(n11892, n10898, new_n7712);
and_5  g07336(n7388, n3754, new_n7713);
and_5  g07337(n11876, n2393, new_n7714);
xnor_4 g07338(new_n7714, new_n7713, new_n7715);
xor_4  g07339(new_n7715, new_n7712, new_n7716);
xnor_4 g07340(new_n7716, new_n7711, new_n7717);
nand_5 g07341(n10898, n7388, new_n7718);
or_5   g07342(new_n7718, new_n4828_1, new_n7719);
or_5   g07343(new_n7707, new_n7705, new_n7720);
and_5  g07344(new_n7720, new_n7719, new_n7721);
nand_5 g07345(new_n7721, new_n7708, new_n7722);
xor_4  g07346(new_n7722, new_n7717, new_n7723);
xnor_4 g07347(new_n7723, new_n7701, new_n7724);
nor_5  g07348(new_n7719, new_n7705, new_n7725);
nor_5  g07349(new_n7725, new_n7721, new_n7726);
and_5  g07350(new_n4844, new_n4841, new_n7727);
nor_5  g07351(new_n4848, new_n4845, new_n7728);
or_5   g07352(new_n7728, new_n7727, new_n7729);
nor_5  g07353(new_n7729, new_n7726, new_n7730_1);
xnor_4 g07354(new_n7729, new_n7726, new_n7731);
or_5   g07355(new_n7690_1, new_n7689, new_n7732);
nand_5 g07356(n8476, n1067, new_n7733_1);
or_5   g07357(new_n7733_1, new_n4827, new_n7734);
nor_5  g07358(new_n7734, new_n7732, new_n7735);
and_5  g07359(new_n7734, new_n7699, new_n7736);
or_5   g07360(new_n7736, new_n7735, new_n7737);
nor_5  g07361(new_n7737, new_n7731, new_n7738);
nor_5  g07362(new_n7738, new_n7730_1, new_n7739);
xnor_4 g07363(new_n7739, new_n7724, new_n7740);
xnor_4 g07364(new_n7740, new_n7681, new_n7741);
or_5   g07365(new_n7677, new_n7662, new_n7742);
and_5  g07366(new_n7742, new_n7679, new_n7743);
and_5  g07367(new_n4839, new_n4836, new_n7744);
nor_5  g07368(new_n4849, new_n4840, new_n7745);
or_5   g07369(new_n7745, new_n7744, new_n7746);
nor_5  g07370(new_n7746, new_n7743, new_n7747);
xnor_4 g07371(new_n7737, new_n7731, new_n7748);
xnor_4 g07372(new_n7746, new_n7743, new_n7749);
nor_5  g07373(new_n7749, new_n7748, new_n7750);
nor_5  g07374(new_n7750, new_n7747, new_n7751);
xor_4  g07375(new_n7751, new_n7741, new_n7752);
nor_5  g07376(new_n7752, new_n7658, new_n7753);
xnor_4 g07377(new_n7752, new_n7658, new_n7754);
xnor_4 g07378(new_n7749, new_n7748, new_n7755);
and_5  g07379(n5305, n1798, new_n7756);
nor_5  g07380(new_n7622, new_n7756, new_n7757);
and_5  g07381(new_n7757, new_n7625, new_n7758);
nor_5  g07382(new_n7757, new_n7637, new_n7759);
or_5   g07383(new_n7759, new_n7758, new_n7760);
nor_5  g07384(new_n7760, new_n7755, new_n7761);
and_5  g07385(new_n4834, new_n4831, new_n7762);
nor_5  g07386(new_n4850, new_n4835, new_n7763);
nor_5  g07387(new_n7763, new_n7762, new_n7764);
xor_4  g07388(new_n7760, new_n7755, new_n7765);
and_5  g07389(new_n7765, new_n7764, new_n7766);
or_5   g07390(new_n7766, new_n7761, new_n7767);
nor_5  g07391(new_n7767, new_n7754, new_n7768);
nor_5  g07392(new_n7768, new_n7753, new_n7769);
xnor_4 g07393(new_n7769, new_n7657, new_n7770);
or_5   g07394(new_n7680, new_n7675, new_n7771);
nand_5 g07395(n10451, n8759, new_n7772);
nand_5 g07396(n11023, n6776, new_n7773);
nor_5  g07397(new_n7672, new_n7671, new_n7774);
and_5  g07398(new_n7672, new_n7671, new_n7775);
nor_5  g07399(new_n7775, new_n7670, new_n7776);
or_5   g07400(new_n7776, new_n7774, new_n7777);
xnor_4 g07401(new_n7777, new_n7773, new_n7778);
and_5  g07402(n9640, n7436, new_n7779);
and_5  g07403(n8276, n6703, new_n7780);
xnor_4 g07404(new_n7780, new_n7664, new_n7781);
xor_4  g07405(new_n7781, new_n7779, new_n7782);
xnor_4 g07406(new_n7782, new_n7778, new_n7783);
xnor_4 g07407(new_n7783, new_n7772, new_n7784);
nor_5  g07408(new_n7668, new_n7659, new_n7785);
nor_5  g07409(new_n7674, new_n7669, new_n7786);
nor_5  g07410(new_n7786, new_n7785, new_n7787);
xnor_4 g07411(new_n7787, new_n7784, new_n7788);
xnor_4 g07412(new_n7788, new_n7771, new_n7789);
or_5   g07413(new_n7722, new_n7717, new_n7790);
nand_5 g07414(n7965, n159, new_n7791);
and_5  g07415(new_n7710, new_n7702, new_n7792);
nor_5  g07416(new_n7716, new_n7711, new_n7793);
nor_5  g07417(new_n7793, new_n7792, new_n7794);
xnor_4 g07418(new_n7794, new_n7791, new_n7795);
and_5  g07419(n7388, n2749, new_n7796);
nor_5  g07420(new_n7714, new_n7713, new_n7797);
nor_5  g07421(new_n7715, new_n7712, new_n7798);
nor_5  g07422(new_n7798, new_n7797, new_n7799);
xnor_4 g07423(new_n7799, new_n7796, new_n7800);
and_5  g07424(n11876, n5860, new_n7801);
and_5  g07425(n10898, n2393, new_n7802);
xnor_4 g07426(new_n7802, new_n7801, new_n7803);
xor_4  g07427(new_n7803, new_n7706, new_n7804);
xnor_4 g07428(new_n7804, new_n7800, new_n7805);
xnor_4 g07429(new_n7805, new_n7795, new_n7806);
xor_4  g07430(new_n7806, new_n7790, new_n7807);
or_5   g07431(new_n7700, new_n7697, new_n7808);
nand_5 g07432(n5331, n2551, new_n7809);
nand_5 g07433(n11922, n8476, new_n7810);
nor_5  g07434(new_n7685, new_n7684, new_n7811);
and_5  g07435(new_n7685, new_n7684, new_n7812);
nor_5  g07436(new_n7812, new_n7683, new_n7813);
or_5   g07437(new_n7813, new_n7811, new_n7814);
xnor_4 g07438(new_n7814, new_n7810, new_n7815);
and_5  g07439(n12648, n1067, new_n7816);
and_5  g07440(n10545, n5645, new_n7817);
xnor_4 g07441(new_n7817, new_n7693, new_n7818);
xor_4  g07442(new_n7818, new_n7816, new_n7819);
xnor_4 g07443(new_n7819, new_n7815, new_n7820);
xnor_4 g07444(new_n7820, new_n7809, new_n7821);
nor_5  g07445(new_n7687, new_n7682, new_n7822);
nor_5  g07446(new_n7696, new_n7688, new_n7823_1);
nor_5  g07447(new_n7823_1, new_n7822, new_n7824);
xnor_4 g07448(new_n7824, new_n7821, new_n7825);
xor_4  g07449(new_n7825, new_n7808, new_n7826);
xnor_4 g07450(new_n7826, new_n7807, new_n7827);
nor_5  g07451(new_n7723, new_n7701, new_n7828);
nor_5  g07452(new_n7739, new_n7724, new_n7829);
nor_5  g07453(new_n7829, new_n7828, new_n7830);
xor_4  g07454(new_n7830, new_n7827, new_n7831);
xnor_4 g07455(new_n7831, new_n7789, new_n7832);
nor_5  g07456(new_n7740, new_n7681, new_n7833);
nor_5  g07457(new_n7751, new_n7741, new_n7834);
or_5   g07458(new_n7834, new_n7833, new_n7835);
xnor_4 g07459(new_n7835, new_n7832, new_n7836);
xor_4  g07460(new_n7836, new_n7770, n3677);
xnor_4 g07461(new_n6775, new_n6774, n3849);
xor_4  g07462(new_n4821, new_n4820, n4088);
xor_4  g07463(new_n971, new_n887, n4155);
xor_4  g07464(new_n2345, new_n2344, n4159);
xor_4  g07465(new_n4811, new_n4680, n4226);
and_5  g07466(n12591, n4312, new_n7843);
nor_5  g07467(new_n7644, new_n7643, new_n7844);
nor_5  g07468(new_n7645, new_n7642, new_n7845);
nor_5  g07469(new_n7845, new_n7844, new_n7846);
xnor_4 g07470(new_n7846, new_n7843, new_n7847);
and_5  g07471(n12705, n3932, new_n7848);
and_5  g07472(n12025, n1798, new_n7849);
xor_4  g07473(new_n7849, new_n7848, new_n7850);
xor_4  g07474(new_n7850, new_n7847, new_n7851);
and_5  g07475(n11662, n5964, new_n7852);
and_5  g07476(n7456, n1097, new_n7853);
xnor_4 g07477(new_n7853, new_n7852, new_n7854);
xnor_4 g07478(new_n7854, new_n7851, new_n7855);
nor_5  g07479(new_n7646_1, new_n7641, new_n7856);
nor_5  g07480(new_n7650, new_n7647, new_n7857);
nor_5  g07481(new_n7857, new_n7856, new_n7858);
xnor_4 g07482(new_n7858, new_n7855, new_n7859);
nor_5  g07483(new_n7651, new_n7640, new_n7860);
nor_5  g07484(new_n7655, new_n7652, new_n7861);
nor_5  g07485(new_n7861, new_n7860, new_n7862_1);
or_5   g07486(new_n7862_1, new_n7859, new_n7863);
nor_5  g07487(new_n7846, new_n7843, new_n7864);
nor_5  g07488(new_n7850, new_n7847, new_n7865);
nor_5  g07489(new_n7865, new_n7864, new_n7866);
and_5  g07490(n10327, n5964, new_n7867);
and_5  g07491(n11662, n1097, new_n7868);
and_5  g07492(n9583, n5305, new_n7869);
xnor_4 g07493(new_n7869, new_n7868, new_n7870);
xnor_4 g07494(new_n7870, new_n7867, new_n7871);
xnor_4 g07495(new_n7871, new_n7866, new_n7872);
and_5  g07496(new_n7849, new_n7848, new_n7873);
and_5  g07497(n7456, n4312, new_n7874);
xnor_4 g07498(new_n7874, new_n7873, new_n7875);
and_5  g07499(n12025, n3932, new_n7876);
and_5  g07500(n12705, n12591, new_n7877);
and_5  g07501(n11257, n1798, new_n7878);
xnor_4 g07502(new_n7878, new_n7877, new_n7879);
xnor_4 g07503(new_n7879, new_n7876, new_n7880);
xnor_4 g07504(new_n7880, new_n7875, new_n7881);
xor_4  g07505(new_n7881, new_n7872, new_n7882);
nor_5  g07506(new_n7854, new_n7851, new_n7883);
nand_5 g07507(new_n7853, new_n7852, new_n7884);
or_5   g07508(new_n7858, new_n7855, new_n7885);
xor_4  g07509(new_n7885, new_n7884, new_n7886);
nor_5  g07510(new_n7886, new_n7883, new_n7887);
xnor_4 g07511(new_n7887, new_n7882, new_n7888);
xnor_4 g07512(new_n7888, new_n7863, new_n7889);
and_5  g07513(n10327, n5305, new_n7890);
xor_4  g07514(new_n7862_1, new_n7859, new_n7891_1);
nor_5  g07515(new_n7891_1, new_n7890, new_n7892);
nor_5  g07516(new_n7656, new_n7639, new_n7893);
xnor_4 g07517(new_n7891_1, new_n7890, new_n7894);
nor_5  g07518(new_n7894, new_n7893, new_n7895);
or_5   g07519(new_n7895, new_n7892, new_n7896);
xnor_4 g07520(new_n7896, new_n7889, new_n7897);
nor_5  g07521(new_n7777, new_n7773, new_n7898);
nor_5  g07522(new_n7782, new_n7778, new_n7899);
nor_5  g07523(new_n7899, new_n7898, new_n7900);
and_5  g07524(n10451, n6776, new_n7901);
and_5  g07525(n12299, n11023, new_n7902);
xnor_4 g07526(new_n7902, new_n7901, new_n7903);
xnor_4 g07527(new_n7903, new_n7900, new_n7904);
and_5  g07528(n7436, n3022, new_n7905);
and_5  g07529(n9640, n8276, new_n7906);
and_5  g07530(n9241, n6703, new_n7907);
xor_4  g07531(new_n7907, new_n7906, new_n7908);
xnor_4 g07532(new_n7908, new_n7905, new_n7909);
nor_5  g07533(new_n7780, new_n7664, new_n7910);
and_5  g07534(new_n7780, new_n7664, new_n7911);
nor_5  g07535(new_n7911, new_n7779, new_n7912);
nor_5  g07536(new_n7912, new_n7910, new_n7913);
xor_4  g07537(new_n7913, new_n7909, new_n7914);
xnor_4 g07538(new_n7914, new_n7904, new_n7915);
nor_5  g07539(new_n7783, new_n7772, new_n7916);
nor_5  g07540(new_n7787, new_n7784, new_n7917);
nor_5  g07541(new_n7917, new_n7916, new_n7918);
or_5   g07542(new_n7918, new_n7915, new_n7919);
nor_5  g07543(new_n7908, new_n7905, new_n7920);
nor_5  g07544(new_n7913, new_n7909, new_n7921);
nor_5  g07545(new_n7921, new_n7920, new_n7922);
and_5  g07546(n10278, n6776, new_n7923);
and_5  g07547(n12299, n10451, new_n7924);
and_5  g07548(n11423, n8759, new_n7925);
xnor_4 g07549(new_n7925, new_n7924, new_n7926);
xnor_4 g07550(new_n7926, new_n7923, new_n7927);
xnor_4 g07551(new_n7927, new_n7922, new_n7928);
and_5  g07552(new_n7907, new_n7906, new_n7929);
and_5  g07553(n11023, n7436, new_n7930);
xnor_4 g07554(new_n7930, new_n7929, new_n7931);
and_5  g07555(n9640, n9241, new_n7932);
and_5  g07556(n8276, n3022, new_n7933);
and_5  g07557(n10510, n6703, new_n7934);
xnor_4 g07558(new_n7934, new_n7933, new_n7935);
xor_4  g07559(new_n7935, new_n7932, new_n7936);
xor_4  g07560(new_n7936, new_n7931, new_n7937);
xor_4  g07561(new_n7937, new_n7928, new_n7938);
nor_5  g07562(new_n7903, new_n7900, new_n7939);
nand_5 g07563(new_n7902, new_n7901, new_n7940);
or_5   g07564(new_n7914, new_n7904, new_n7941);
xor_4  g07565(new_n7941, new_n7940, new_n7942);
nor_5  g07566(new_n7942, new_n7939, new_n7943);
xnor_4 g07567(new_n7943, new_n7938, new_n7944);
xnor_4 g07568(new_n7944, new_n7919, new_n7945);
nand_5 g07569(n10278, n8759, new_n7946_1);
xnor_4 g07570(new_n7918, new_n7915, new_n7947);
nor_5  g07571(new_n7947, new_n7946_1, new_n7948);
or_5   g07572(new_n7788, new_n7771, new_n7949);
xnor_4 g07573(new_n7947, new_n7946_1, new_n7950);
nor_5  g07574(new_n7950, new_n7949, new_n7951);
nor_5  g07575(new_n7951, new_n7948, new_n7952);
xor_4  g07576(new_n7952, new_n7945, new_n7953);
nand_5 g07577(n12648, n8665, new_n7954);
and_5  g07578(n10545, n1067, new_n7955);
and_5  g07579(n7690, n5645, new_n7956);
xnor_4 g07580(new_n7956, new_n7955, new_n7957);
xnor_4 g07581(new_n7957, new_n7954, new_n7958);
nor_5  g07582(new_n7817, new_n7693, new_n7959);
and_5  g07583(new_n7817, new_n7693, new_n7960);
nor_5  g07584(new_n7960, new_n7816, new_n7961);
or_5   g07585(new_n7961, new_n7959, new_n7962);
xnor_4 g07586(new_n7962, new_n7958, new_n7963);
and_5  g07587(n8476, n2551, new_n7964);
and_5  g07588(n11922, n2530, new_n7965_1);
xnor_4 g07589(new_n7965_1, new_n7964, new_n7966_1);
xnor_4 g07590(new_n7966_1, new_n7963, new_n7967);
nor_5  g07591(new_n7814, new_n7810, new_n7968);
nor_5  g07592(new_n7819, new_n7815, new_n7969);
nor_5  g07593(new_n7969, new_n7968, new_n7970);
xnor_4 g07594(new_n7970, new_n7967, new_n7971);
nor_5  g07595(new_n7820, new_n7809, new_n7972);
nor_5  g07596(new_n7824, new_n7821, new_n7973);
nor_5  g07597(new_n7973, new_n7972, new_n7974);
or_5   g07598(new_n7974, new_n7971, new_n7975);
and_5  g07599(new_n7956, new_n7955, new_n7976);
and_5  g07600(n12648, n11922, new_n7977);
xnor_4 g07601(new_n7977, new_n7976, new_n7978);
and_5  g07602(n7690, n1067, new_n7979);
and_5  g07603(n10545, n8665, new_n7980);
and_5  g07604(n5645, n3616, new_n7981_1);
xnor_4 g07605(new_n7981_1, new_n7980, new_n7982);
xor_4  g07606(new_n7982, new_n7979, new_n7983);
xor_4  g07607(new_n7983, new_n7978, new_n7984);
nor_5  g07608(new_n7957, new_n7954, new_n7985);
nor_5  g07609(new_n7962, new_n7958, new_n7986);
or_5   g07610(new_n7986, new_n7985, new_n7987);
and_5  g07611(n12826, n8476, new_n7988);
and_5  g07612(n2551, n2530, new_n7989);
and_5  g07613(n5331, n4094, new_n7990);
xnor_4 g07614(new_n7990, new_n7989, new_n7991);
xnor_4 g07615(new_n7991, new_n7988, new_n7992);
xnor_4 g07616(new_n7992, new_n7987, new_n7993);
xor_4  g07617(new_n7993, new_n7984, new_n7994);
nor_5  g07618(new_n7966_1, new_n7963, new_n7995);
nand_5 g07619(new_n7965_1, new_n7964, new_n7996);
or_5   g07620(new_n7970, new_n7967, new_n7997);
xor_4  g07621(new_n7997, new_n7996, new_n7998);
nor_5  g07622(new_n7998, new_n7995, new_n7999);
xnor_4 g07623(new_n7999, new_n7994, new_n8000);
xnor_4 g07624(new_n8000, new_n7975, new_n8001);
and_5  g07625(n12826, n5331, new_n8002);
xor_4  g07626(new_n7974, new_n7971, new_n8003);
nor_5  g07627(new_n8003, new_n8002, new_n8004);
nor_5  g07628(new_n7825, new_n7808, new_n8005);
xnor_4 g07629(new_n8003, new_n8002, new_n8006);
nor_5  g07630(new_n8006, new_n8005, new_n8007);
or_5   g07631(new_n8007, new_n8004, new_n8008);
xor_4  g07632(new_n8008, new_n8001, new_n8009);
and_5  g07633(n7965, n1510, new_n8010);
and_5  g07634(new_n7799, new_n7796, new_n8011);
nor_5  g07635(new_n7804, new_n7800, new_n8012);
or_5   g07636(new_n8012, new_n8011, new_n8013);
and_5  g07637(n7388, n159, new_n8014);
and_5  g07638(n11892, n2749, new_n8015);
xor_4  g07639(new_n8015, new_n8014, new_n8016);
xnor_4 g07640(new_n8016, new_n8013, new_n8017);
nand_5 g07641(n3754, n2393, new_n8018);
and_5  g07642(n10898, n5860, new_n8019);
and_5  g07643(n11876, n3986, new_n8020);
xnor_4 g07644(new_n8020, new_n8019, new_n8021);
xnor_4 g07645(new_n8021, new_n8018, new_n8022);
nor_5  g07646(new_n7802, new_n7801, new_n8023);
nor_5  g07647(new_n7803, new_n7706, new_n8024);
or_5   g07648(new_n8024, new_n8023, new_n8025);
xor_4  g07649(new_n8025, new_n8022, new_n8026);
xor_4  g07650(new_n8026, new_n8017, new_n8027);
nor_5  g07651(new_n7794, new_n7791, new_n8028_1);
nor_5  g07652(new_n7805, new_n7795, new_n8029);
nor_5  g07653(new_n8029, new_n8028_1, new_n8030);
xor_4  g07654(new_n8030, new_n8027, new_n8031);
and_5  g07655(new_n8031, new_n8010, new_n8032);
or_5   g07656(new_n7806, new_n7790, new_n8033);
xnor_4 g07657(new_n8031, new_n8010, new_n8034);
nor_5  g07658(new_n8034, new_n8033, new_n8035);
nor_5  g07659(new_n8035, new_n8032, new_n8036);
or_5   g07660(new_n8030, new_n8027, new_n8037);
nand_5 g07661(new_n8015, new_n8014, new_n8038);
nor_5  g07662(new_n8016, new_n8013, new_n8039);
nor_5  g07663(new_n8026, new_n8017, new_n8040);
or_5   g07664(new_n8040, new_n8039, new_n8041);
xnor_4 g07665(new_n8041, new_n8038, new_n8042);
and_5  g07666(n7388, n1510, new_n8043);
nand_5 g07667(n11892, n159, new_n8044);
nand_5 g07668(n12247, n7965, new_n8045);
xnor_4 g07669(new_n8045, new_n8044, new_n8046);
xnor_4 g07670(new_n8046, new_n8043, new_n8047);
nor_5  g07671(new_n8021, new_n8018, new_n8048);
nor_5  g07672(new_n8025, new_n8022, new_n8049);
or_5   g07673(new_n8049, new_n8048, new_n8050);
xnor_4 g07674(new_n8050, new_n8047, new_n8051);
and_5  g07675(new_n8020, new_n8019, new_n8052);
and_5  g07676(n2749, n2393, new_n8053);
xnor_4 g07677(new_n8053, new_n8052, new_n8054);
and_5  g07678(n10898, n3986, new_n8055);
and_5  g07679(n11876, n5857, new_n8056);
and_5  g07680(n5860, n3754, new_n8057);
xnor_4 g07681(new_n8057, new_n8056, new_n8058);
xor_4  g07682(new_n8058, new_n8055, new_n8059);
xor_4  g07683(new_n8059, new_n8054, new_n8060);
xor_4  g07684(new_n8060, new_n8051, new_n8061);
xnor_4 g07685(new_n8061, new_n8042, new_n8062);
xnor_4 g07686(new_n8062, new_n8037, new_n8063);
xor_4  g07687(new_n8063, new_n8036, new_n8064);
xnor_4 g07688(new_n8064, new_n8009, new_n8065_1);
xor_4  g07689(new_n8034, new_n8033, new_n8066);
xnor_4 g07690(new_n8006, new_n8005, new_n8067);
nor_5  g07691(new_n8067, new_n8066, new_n8068);
nor_5  g07692(new_n7826, new_n7807, new_n8069);
nor_5  g07693(new_n7830, new_n7827, new_n8070);
nor_5  g07694(new_n8070, new_n8069, new_n8071);
xnor_4 g07695(new_n8067, new_n8066, new_n8072);
nor_5  g07696(new_n8072, new_n8071, new_n8073);
nor_5  g07697(new_n8073, new_n8068, new_n8074);
xnor_4 g07698(new_n8074, new_n8065_1, new_n8075);
xnor_4 g07699(new_n8075, new_n7953, new_n8076);
xor_4  g07700(new_n7950, new_n7949, new_n8077);
xnor_4 g07701(new_n8072, new_n8071, new_n8078);
nor_5  g07702(new_n8078, new_n8077, new_n8079);
nor_5  g07703(new_n7831, new_n7789, new_n8080);
nor_5  g07704(new_n7835, new_n7832, new_n8081);
or_5   g07705(new_n8081, new_n8080, new_n8082);
xnor_4 g07706(new_n8078, new_n8077, new_n8083);
nor_5  g07707(new_n8083, new_n8082, new_n8084);
nor_5  g07708(new_n8084, new_n8079, new_n8085);
xor_4  g07709(new_n8085, new_n8076, new_n8086);
and_5  g07710(new_n8086, new_n7897, new_n8087);
xnor_4 g07711(new_n8086, new_n7897, new_n8088);
xnor_4 g07712(new_n7894, new_n7893, new_n8089);
xnor_4 g07713(new_n8083, new_n8082, new_n8090);
nor_5  g07714(new_n8090, new_n8089, new_n8091);
xor_4  g07715(new_n8090, new_n8089, new_n8092);
nor_5  g07716(new_n7769, new_n7657, new_n8093);
nor_5  g07717(new_n7836, new_n7770, new_n8094);
nor_5  g07718(new_n8094, new_n8093, new_n8095);
and_5  g07719(new_n8095, new_n8092, new_n8096);
nor_5  g07720(new_n8096, new_n8091, new_n8097);
nor_5  g07721(new_n8097, new_n8088, new_n8098);
nor_5  g07722(new_n8098, new_n8087, new_n8099);
nor_5  g07723(new_n7944, new_n7919, new_n8100_1);
nor_5  g07724(new_n7952, new_n7945, new_n8101);
or_5   g07725(new_n8101, new_n8100_1, new_n8102);
nor_5  g07726(new_n8075, new_n7953, new_n8103);
nor_5  g07727(new_n8085, new_n8076, new_n8104);
nor_5  g07728(new_n8104, new_n8103, new_n8105);
nor_5  g07729(new_n7874, new_n7873, new_n8106);
nor_5  g07730(new_n7880, new_n7875, new_n8107);
nor_5  g07731(new_n8107, new_n8106, new_n8108);
and_5  g07732(n11662, n4312, new_n8109);
xnor_4 g07733(new_n8109, new_n8108, new_n8110);
and_5  g07734(new_n7930, new_n7929, new_n8111);
nor_5  g07735(new_n7936, new_n7931, new_n8112);
nor_5  g07736(new_n8112, new_n8111, new_n8113);
and_5  g07737(n12299, n10278, new_n8114);
xnor_4 g07738(new_n8114, new_n8113, new_n8115);
nor_5  g07739(new_n7925, new_n7924, new_n8116);
nor_5  g07740(new_n7926, new_n7923, new_n8117);
nor_5  g07741(new_n8117, new_n8116, new_n8118);
and_5  g07742(n10451, n7436, new_n8119);
and_5  g07743(n9241, n3022, new_n8120);
xnor_4 g07744(new_n8120, new_n8119, new_n8121);
and_5  g07745(n11257, n3932, new_n8122);
and_5  g07746(n10327, n1097, new_n8123);
xnor_4 g07747(new_n8123, new_n8122, new_n8124);
xor_4  g07748(new_n8124, new_n8121, new_n8125);
xnor_4 g07749(new_n8125, new_n8118, new_n8126);
nor_5  g07750(new_n8057, new_n8056, new_n8127);
nor_5  g07751(new_n8058, new_n8055, new_n8128);
nor_5  g07752(new_n8128, new_n8127, new_n8129);
and_5  g07753(n2393, n159, new_n8130);
and_5  g07754(n5860, n2749, new_n8131);
xor_4  g07755(new_n8131, new_n8130, new_n8132);
xnor_4 g07756(new_n8132, new_n8129, new_n8133);
xnor_4 g07757(new_n8133, new_n8126, new_n8134);
xnor_4 g07758(new_n8134, new_n8115, new_n8135);
xnor_4 g07759(new_n8135, new_n8110, new_n8136);
nor_5  g07760(new_n8000, new_n7975, new_n8137);
nor_5  g07761(new_n8008, new_n8001, new_n8138_1);
nor_5  g07762(new_n8138_1, new_n8137, new_n8139);
xnor_4 g07763(new_n8139, new_n8136, new_n8140);
nor_5  g07764(new_n8041, new_n8038, new_n8141);
nor_5  g07765(new_n8061, new_n8042, new_n8142);
nor_5  g07766(new_n8142, new_n8141, new_n8143);
nor_5  g07767(new_n8046, new_n8043, new_n8144);
or_5   g07768(new_n8144, new_n8044, new_n8145);
nand_5 g07769(n12247, n7388, new_n8146);
nor_5  g07770(new_n8146, new_n8145, new_n8147);
or_5   g07771(new_n8146, new_n8010, new_n8148);
and_5  g07772(new_n8148, new_n8145, new_n8149);
nor_5  g07773(new_n8149, new_n8147, new_n8150);
and_5  g07774(n10898, n5857, new_n8151);
and_5  g07775(n12591, n12025, new_n8152);
and_5  g07776(n11876, n45, new_n8153);
xnor_4 g07777(new_n8153, new_n8152, new_n8154);
xnor_4 g07778(new_n8154, new_n8151, new_n8155);
xnor_4 g07779(new_n8155, new_n8150, new_n8156);
xnor_4 g07780(new_n8156, new_n8143, new_n8157);
nor_5  g07781(new_n7934, new_n7933, new_n8158);
nor_5  g07782(new_n7935, new_n7932, new_n8159);
nor_5  g07783(new_n8159, new_n8158, new_n8160);
and_5  g07784(n12705, n7456, new_n8161);
and_5  g07785(n11023, n8276, new_n8162);
xor_4  g07786(new_n8162, new_n8161, new_n8163);
xnor_4 g07787(new_n8163, new_n8160, new_n8164);
and_5  g07788(n9583, n5964, new_n8165);
and_5  g07789(n12511, n7965, new_n8166);
xnor_4 g07790(new_n8166, new_n8165, new_n8167);
xnor_4 g07791(new_n8167, new_n8164, new_n8168);
nor_5  g07792(new_n7941, new_n7940, new_n8169);
nor_5  g07793(new_n7943, new_n7938, new_n8170);
nor_5  g07794(new_n8170, new_n8169, new_n8171);
nor_5  g07795(new_n7927, new_n7922, new_n8172);
nor_5  g07796(new_n7937, new_n7928, new_n8173);
or_5   g07797(new_n8173, new_n8172, new_n8174);
xnor_4 g07798(new_n8174, new_n8171, new_n8175);
xnor_4 g07799(new_n8175, new_n8168, new_n8176);
xnor_4 g07800(new_n8176, new_n8157, new_n8177);
nor_5  g07801(new_n8062, new_n8037, new_n8178);
nor_5  g07802(new_n8063, new_n8036, new_n8179);
nor_5  g07803(new_n8179, new_n8178, new_n8180);
nor_5  g07804(new_n7997, new_n7996, new_n8181);
nor_5  g07805(new_n7999, new_n7994, new_n8182);
nor_5  g07806(new_n8182, new_n8181, new_n8183);
nor_5  g07807(new_n7871, new_n7866, new_n8184);
nor_5  g07808(new_n7881, new_n7872, new_n8185);
or_5   g07809(new_n8185, new_n8184, new_n8186);
xnor_4 g07810(new_n8186, new_n8183, new_n8187);
and_5  g07811(n3986, n3754, new_n8188);
and_5  g07812(n11423, n6776, new_n8189);
xnor_4 g07813(new_n8189, new_n8188, new_n8190);
and_5  g07814(n8759, n2278, new_n8191);
and_5  g07815(n10510, n9640, new_n8192);
xnor_4 g07816(new_n8192, new_n8191, new_n8193);
xnor_4 g07817(new_n8193, new_n8190, new_n8194);
and_5  g07818(n8476, n4094, new_n8195);
and_5  g07819(n5305, n753, new_n8196);
xnor_4 g07820(new_n8196, new_n8195, new_n8197);
and_5  g07821(n3616, n1067, new_n8198);
and_5  g07822(n10644, n6703, new_n8199);
xnor_4 g07823(new_n8199, new_n8198, new_n8200);
xnor_4 g07824(new_n8200, new_n8197, new_n8201);
xnor_4 g07825(new_n8201, new_n8194, new_n8202_1);
nor_5  g07826(new_n7869, new_n7868, new_n8203);
nor_5  g07827(new_n7870, new_n7867, new_n8204);
nor_5  g07828(new_n8204, new_n8203, new_n8205);
nor_5  g07829(new_n7878, new_n7877, new_n8206);
nor_5  g07830(new_n7879, new_n7876, new_n8207);
nor_5  g07831(new_n8207, new_n8206, new_n8208);
xnor_4 g07832(new_n8208, new_n8205, new_n8209);
xnor_4 g07833(new_n8209, new_n8202_1, new_n8210);
xnor_4 g07834(new_n8210, new_n8187, new_n8211);
nor_5  g07835(new_n7885, new_n7884, new_n8212);
nor_5  g07836(new_n7887, new_n7882, new_n8213);
or_5   g07837(new_n8213, new_n8212, new_n8214);
nor_5  g07838(new_n8050, new_n8047, new_n8215);
nor_5  g07839(new_n8060, new_n8051, new_n8216);
nor_5  g07840(new_n8216, new_n8215, new_n8217);
and_5  g07841(new_n8053, new_n8052, new_n8218);
nor_5  g07842(new_n8059, new_n8054, new_n8219);
nor_5  g07843(new_n8219, new_n8218, new_n8220);
nor_5  g07844(new_n7981_1, new_n7980, new_n8221);
nor_5  g07845(new_n7982, new_n7979, new_n8222);
nor_5  g07846(new_n8222, new_n8221, new_n8223);
and_5  g07847(n10547, n1798, new_n8224);
and_5  g07848(n8665, n7690, new_n8225);
xnor_4 g07849(new_n8225, new_n8224, new_n8226);
and_5  g07850(n12826, n2530, new_n8227);
and_5  g07851(n11892, n1510, new_n8228);
xnor_4 g07852(new_n8228, new_n8227, new_n8229);
xor_4  g07853(new_n8229, new_n8226, new_n8230);
xnor_4 g07854(new_n8230, new_n8223, new_n8231);
xnor_4 g07855(new_n8231, new_n8220, new_n8232);
xnor_4 g07856(new_n8232, new_n8217, new_n8233);
nand_5 g07857(n11922, n10545, new_n8234);
nor_5  g07858(new_n7992, new_n7987, new_n8235);
nor_5  g07859(new_n7993, new_n7984, new_n8236_1);
nor_5  g07860(new_n8236_1, new_n8235, new_n8237);
xnor_4 g07861(new_n8237, new_n8234, new_n8238);
and_5  g07862(new_n7977, new_n7976, new_n8239);
nor_5  g07863(new_n7983, new_n7978, new_n8240);
nor_5  g07864(new_n8240, new_n8239, new_n8241);
nor_5  g07865(new_n7990, new_n7989, new_n8242);
nor_5  g07866(new_n7991, new_n7988, new_n8243);
or_5   g07867(new_n8243, new_n8242, new_n8244);
xnor_4 g07868(new_n8244, new_n8241, new_n8245);
nand_5 g07869(n12648, n2551, new_n8246);
and_5  g07870(n10685, n5331, new_n8247);
and_5  g07871(n5645, n4499, new_n8248);
xnor_4 g07872(new_n8248, new_n8247, new_n8249);
xnor_4 g07873(new_n8249, new_n8246, new_n8250);
xnor_4 g07874(new_n8250, new_n8245, new_n8251);
xnor_4 g07875(new_n8251, new_n8238, new_n8252);
xnor_4 g07876(new_n8252, new_n8233, new_n8253);
xnor_4 g07877(new_n8253, new_n8214, new_n8254);
xnor_4 g07878(new_n8254, new_n8211, new_n8255);
xnor_4 g07879(new_n8255, new_n8180, new_n8256);
xnor_4 g07880(new_n8256, new_n8177, new_n8257);
xnor_4 g07881(new_n8257, new_n8140, new_n8258);
nor_5  g07882(new_n7888, new_n7863, new_n8259);
nor_5  g07883(new_n7896, new_n7889, new_n8260);
or_5   g07884(new_n8260, new_n8259, new_n8261);
nor_5  g07885(new_n8064, new_n8009, new_n8262);
nor_5  g07886(new_n8074, new_n8065_1, new_n8263);
nor_5  g07887(new_n8263, new_n8262, new_n8264);
xnor_4 g07888(new_n8264, new_n8261, new_n8265);
xnor_4 g07889(new_n8265, new_n8258, new_n8266);
xnor_4 g07890(new_n8266, new_n8105, new_n8267);
xnor_4 g07891(new_n8267, new_n8102, new_n8268);
xnor_4 g07892(new_n8268, new_n8099, n4230);
xnor_4 g07893(new_n4672, new_n4671, n4300);
xnor_4 g07894(new_n2899, new_n2898, n4326);
or_5   g07895(new_n1062, new_n1056, new_n8272);
nand_5 g07896(n6687, n5320, new_n8273);
nor_5  g07897(new_n1049, new_n1042, new_n8274);
nor_5  g07898(new_n1055, new_n1050, new_n8275);
nor_5  g07899(new_n8275, new_n8274, new_n8276_1);
xnor_4 g07900(new_n8276_1, new_n8273, new_n8277);
and_5  g07901(n4370, n2564, new_n8278);
nor_5  g07902(new_n1053, new_n1052, new_n8279);
nor_5  g07903(new_n1054, new_n1051, new_n8280);
nor_5  g07904(new_n8280, new_n8279, new_n8281);
xnor_4 g07905(new_n8281, new_n8278, new_n8282);
and_5  g07906(n6770, n5212, new_n8283);
and_5  g07907(n11877, n4189, new_n8284);
and_5  g07908(n11407, n9920, new_n8285);
xnor_4 g07909(new_n8285, new_n8284, new_n8286);
xor_4  g07910(new_n8286, new_n8283, new_n8287);
xnor_4 g07911(new_n8287, new_n8282, new_n8288);
xnor_4 g07912(new_n8288, new_n8277, new_n8289);
xnor_4 g07913(new_n8289, new_n8272, new_n8290);
or_5   g07914(new_n1151, new_n1150, new_n8291);
nand_5 g07915(n8336, n2433, new_n8292);
nand_5 g07916(n10928, n8819, new_n8293);
nor_5  g07917(new_n1144, new_n1143, new_n8294);
and_5  g07918(new_n1144, new_n1143, new_n8295);
nor_5  g07919(new_n8295, new_n1142, new_n8296);
or_5   g07920(new_n8296, new_n8294, new_n8297);
xnor_4 g07921(new_n8297, new_n8293, new_n8298);
and_5  g07922(n11728, n2226, new_n8299);
and_5  g07923(n12709, n1094, new_n8300);
xnor_4 g07924(new_n8300, new_n1088, new_n8301);
xor_4  g07925(new_n8301, new_n8299, new_n8302);
xnor_4 g07926(new_n8302, new_n8298, new_n8303_1);
xnor_4 g07927(new_n8303_1, new_n8292, new_n8304);
nor_5  g07928(new_n1146, new_n1141, new_n8305);
nor_5  g07929(new_n1149, new_n1147, new_n8306);
nor_5  g07930(new_n8306, new_n8305, new_n8307);
xnor_4 g07931(new_n8307, new_n8304, new_n8308);
xnor_4 g07932(new_n8308, new_n8291, new_n8309);
nor_5  g07933(new_n1183, new_n1152, new_n8310);
nor_5  g07934(new_n1187, new_n1184, new_n8311);
nor_5  g07935(new_n8311, new_n8310, new_n8312);
xnor_4 g07936(new_n8312, new_n8309, new_n8313);
or_5   g07937(new_n1164, new_n1163, new_n8314);
nand_5 g07938(n12069, n11967, new_n8315);
and_5  g07939(n12391, n6254, new_n8316);
nor_5  g07940(new_n1160, new_n1159, new_n8317);
nor_5  g07941(new_n1161, new_n1158, new_n8318);
nor_5  g07942(new_n8318, new_n8317, new_n8319);
xnor_4 g07943(new_n8319, new_n8316, new_n8320);
and_5  g07944(n7160, n7159, new_n8321);
and_5  g07945(n12777, n7891, new_n8322);
and_5  g07946(n12489, n4828, new_n8323);
xnor_4 g07947(new_n8323, new_n8322, new_n8324);
xor_4  g07948(new_n8324, new_n8321, new_n8325);
xnor_4 g07949(new_n8325, new_n8320, new_n8326);
xnor_4 g07950(new_n8326, new_n8315, new_n8327);
and_5  g07951(new_n1156, new_n1153, new_n8328);
nor_5  g07952(new_n1162, new_n1157, new_n8329);
nor_5  g07953(new_n8329, new_n8328, new_n8330);
xnor_4 g07954(new_n8330, new_n8327, new_n8331);
xnor_4 g07955(new_n8331, new_n8314, new_n8332);
or_5   g07956(new_n1177, new_n1176, new_n8333);
nand_5 g07957(n12947, n11222, new_n8334);
and_5  g07958(n11791, n11153, new_n8335);
nor_5  g07959(new_n1173, new_n1172, new_n8336_1);
nor_5  g07960(new_n1174, new_n1171, new_n8337);
nor_5  g07961(new_n8337, new_n8336_1, new_n8338);
xnor_4 g07962(new_n8338, new_n8335, new_n8339);
and_5  g07963(n5760, n996, new_n8340);
and_5  g07964(n5314, n1478, new_n8341);
and_5  g07965(n10990, n5767, new_n8342);
xnor_4 g07966(new_n8342, new_n8341, new_n8343);
xor_4  g07967(new_n8343, new_n8340, new_n8344);
xnor_4 g07968(new_n8344, new_n8339, new_n8345);
xnor_4 g07969(new_n8345, new_n8334, new_n8346);
and_5  g07970(new_n1169, new_n1166, new_n8347);
nor_5  g07971(new_n1175, new_n1170, new_n8348);
nor_5  g07972(new_n8348, new_n8347, new_n8349);
xnor_4 g07973(new_n8349, new_n8346, new_n8350);
xnor_4 g07974(new_n8350, new_n8333, new_n8351);
nor_5  g07975(new_n1178, new_n1165, new_n8352);
nor_5  g07976(new_n1182, new_n1179, new_n8353);
nor_5  g07977(new_n8353, new_n8352, new_n8354);
xor_4  g07978(new_n8354, new_n8351, new_n8355);
xnor_4 g07979(new_n8355, new_n8332, new_n8356);
xnor_4 g07980(new_n8356, new_n8313, new_n8357);
xnor_4 g07981(new_n8357, new_n8290, new_n8358);
and_5  g07982(new_n1139, new_n1063, new_n8359);
nor_5  g07983(new_n1188, new_n1140, new_n8360);
nor_5  g07984(new_n8360, new_n8359, new_n8361);
xor_4  g07985(new_n8361, new_n8358, n4333);
and_5  g07986(n11877, n11757, new_n8363);
and_5  g07987(n5240, n5212, new_n8364);
and_5  g07988(n11821, n11407, new_n8365);
xor_4  g07989(new_n8365, new_n8364, new_n8366);
xnor_4 g07990(new_n8366, new_n8363, new_n8367);
and_5  g07991(n11407, n5240, new_n8368);
and_5  g07992(n11877, n3172, new_n8369);
nor_5  g07993(new_n8369, new_n8368, new_n8370);
and_5  g07994(n11757, n5212, new_n8371);
xnor_4 g07995(new_n8369, new_n8368, new_n8372);
nor_5  g07996(new_n8372, new_n8371, new_n8373);
nor_5  g07997(new_n8373, new_n8370, new_n8374);
xnor_4 g07998(new_n8374, new_n8367, new_n8375);
and_5  g07999(n5320, n1333, new_n8376);
and_5  g08000(n4370, n3172, new_n8377);
xor_4  g08001(new_n8377, new_n8376, new_n8378);
xnor_4 g08002(new_n8378, new_n8375, new_n8379);
and_5  g08003(n4370, n1333, new_n8380);
and_5  g08004(n11877, n1333, new_n8381);
and_5  g08005(n11757, n11407, new_n8382);
nor_5  g08006(new_n8382, new_n8381, new_n8383);
and_5  g08007(n5212, n3172, new_n8384_1);
xnor_4 g08008(new_n8382, new_n8381, new_n8385);
nor_5  g08009(new_n8385, new_n8384_1, new_n8386);
nor_5  g08010(new_n8386, new_n8383, new_n8387);
and_5  g08011(new_n8387, new_n8380, new_n8388);
xnor_4 g08012(new_n8387, new_n8380, new_n8389);
xor_4  g08013(new_n8372, new_n8371, new_n8390);
nor_5  g08014(new_n8390, new_n8389, new_n8391);
nor_5  g08015(new_n8391, new_n8388, new_n8392);
xnor_4 g08016(new_n8392, new_n8379, new_n8393);
and_5  g08017(n7862, n5320, new_n8394);
xor_4  g08018(new_n8390, new_n8389, new_n8395);
nor_5  g08019(new_n8395, new_n8394, new_n8396);
xnor_4 g08020(new_n8395, new_n8394, new_n8397);
and_5  g08021(n7862, n4370, new_n8398_1);
and_5  g08022(n11407, n3172, new_n8399);
and_5  g08023(n11877, n7862, new_n8400);
nor_5  g08024(new_n8400, new_n8399, new_n8401);
and_5  g08025(n11407, n7862, new_n8402);
and_5  g08026(new_n8402, new_n8369, new_n8403);
and_5  g08027(n5212, n1333, new_n8404);
nor_5  g08028(new_n8404, new_n8403, new_n8405);
nor_5  g08029(new_n8405, new_n8401, new_n8406);
and_5  g08030(new_n8406, new_n8398_1, new_n8407);
xnor_4 g08031(new_n8406, new_n8398_1, new_n8408);
xor_4  g08032(new_n8385, new_n8384_1, new_n8409);
nor_5  g08033(new_n8409, new_n8408, new_n8410);
or_5   g08034(new_n8410, new_n8407, new_n8411);
nor_5  g08035(new_n8411, new_n8397, new_n8412);
or_5   g08036(new_n8412, new_n8396, new_n8413);
or_5   g08037(new_n8413, new_n8393, new_n8414);
and_5  g08038(new_n8378, new_n8375, new_n8415);
nand_5 g08039(new_n8377, new_n8376, new_n8416);
or_5   g08040(new_n8392, new_n8379, new_n8417);
xor_4  g08041(new_n8417, new_n8416, new_n8418);
nor_5  g08042(new_n8418, new_n8415, new_n8419);
and_5  g08043(new_n8365, new_n8364, new_n8420);
and_5  g08044(n11757, n4370, new_n8421);
xnor_4 g08045(new_n8421, new_n8420, new_n8422);
and_5  g08046(n11821, n5212, new_n8423);
and_5  g08047(n11877, n5240, new_n8424);
and_5  g08048(n11407, n9080, new_n8425);
xnor_4 g08049(new_n8425, new_n8424, new_n8426);
xnor_4 g08050(new_n8426, new_n8423, new_n8427);
xnor_4 g08051(new_n8427, new_n8422, new_n8428);
nor_5  g08052(new_n8366, new_n8363, new_n8429);
nor_5  g08053(new_n8374, new_n8367, new_n8430);
nor_5  g08054(new_n8430, new_n8429, new_n8431);
and_5  g08055(n12000, n1333, new_n8432);
and_5  g08056(n5320, n3172, new_n8433_1);
and_5  g08057(n9725, n7862, new_n8434);
xnor_4 g08058(new_n8434, new_n8433_1, new_n8435);
xnor_4 g08059(new_n8435, new_n8432, new_n8436);
xnor_4 g08060(new_n8436, new_n8431, new_n8437);
xor_4  g08061(new_n8437, new_n8428, new_n8438);
xnor_4 g08062(new_n8438, new_n8419, new_n8439);
xnor_4 g08063(new_n8439, new_n8414, new_n8440);
and_5  g08064(n12000, n7862, new_n8441);
xor_4  g08065(new_n8413, new_n8393, new_n8442);
nor_5  g08066(new_n8442, new_n8441, new_n8443);
xnor_4 g08067(new_n8409, new_n8408, new_n8444);
nor_5  g08068(new_n8403, new_n8401, new_n8445);
and_5  g08069(n11407, n1333, new_n8446);
and_5  g08070(n7862, n5212, new_n8447);
nand_5 g08071(new_n8447, new_n8446, new_n8448);
or_5   g08072(new_n8448, new_n8445, new_n8449);
or_5   g08073(new_n8449, new_n8444, new_n8450);
xor_4  g08074(new_n8411, new_n8397, new_n8451);
nor_5  g08075(new_n8451, new_n8450, new_n8452);
xnor_4 g08076(new_n8442, new_n8441, new_n8453);
nor_5  g08077(new_n8453, new_n8452, new_n8454);
or_5   g08078(new_n8454, new_n8443, new_n8455);
xnor_4 g08079(new_n8455, new_n8440, new_n8456);
nand_5 g08080(n8819, n6877, new_n8457);
and_5  g08081(n12709, n2464, new_n8458);
and_5  g08082(n6877, n6429, new_n8459);
and_5  g08083(new_n8459, new_n8458, new_n8460);
nor_5  g08084(new_n8459, new_n8458, new_n8461);
nand_5 g08085(n11728, n9400, new_n8462);
nor_5  g08086(new_n8462, new_n8461, new_n8463);
nor_5  g08087(new_n8463, new_n8460, new_n8464);
xnor_4 g08088(new_n8464, new_n8457, new_n8465);
and_5  g08089(n11728, n2464, new_n8466);
and_5  g08090(n12709, n11311, new_n8467);
and_5  g08091(n9400, n6429, new_n8468);
xnor_4 g08092(new_n8468, new_n8467, new_n8469);
xor_4  g08093(new_n8469, new_n8466, new_n8470);
xnor_4 g08094(new_n8470, new_n8465, new_n8471);
xor_4  g08095(new_n8459, new_n8458, new_n8472);
and_5  g08096(n12709, n9400, new_n8473);
and_5  g08097(n11728, n6877, new_n8474);
nand_5 g08098(new_n8474, new_n8473, new_n8475);
or_5   g08099(new_n8475, new_n8472, new_n8476_1);
or_5   g08100(new_n8476_1, new_n8471, new_n8477);
nand_5 g08101(n6877, n2433, new_n8478);
nand_5 g08102(n9400, n8819, new_n8479);
nor_5  g08103(new_n8468, new_n8467, new_n8480);
and_5  g08104(new_n8468, new_n8467, new_n8481);
nor_5  g08105(new_n8481, new_n8466, new_n8482);
or_5   g08106(new_n8482, new_n8480, new_n8483);
xnor_4 g08107(new_n8483, new_n8479, new_n8484);
and_5  g08108(n11728, n11311, new_n8485);
and_5  g08109(n6429, n2464, new_n8486);
and_5  g08110(n12709, n4187, new_n8487);
xnor_4 g08111(new_n8487, new_n8486, new_n8488);
xor_4  g08112(new_n8488, new_n8485, new_n8489);
xnor_4 g08113(new_n8489, new_n8484, new_n8490);
xnor_4 g08114(new_n8490, new_n8478, new_n8491);
nor_5  g08115(new_n8464, new_n8457, new_n8492);
nor_5  g08116(new_n8470, new_n8465, new_n8493);
nor_5  g08117(new_n8493, new_n8492, new_n8494);
xnor_4 g08118(new_n8494, new_n8491, new_n8495);
or_5   g08119(new_n8495, new_n8477, new_n8496);
nand_5 g08120(n8717, n6877, new_n8497);
nand_5 g08121(n11311, n6429, new_n8498);
and_5  g08122(n12709, n4203, new_n8499);
and_5  g08123(n11728, n4187, new_n8500);
xnor_4 g08124(new_n8500, new_n8499, new_n8501);
xnor_4 g08125(new_n8501, new_n8498, new_n8502);
nor_5  g08126(new_n8487, new_n8486, new_n8503);
nor_5  g08127(new_n8488, new_n8485, new_n8504);
or_5   g08128(new_n8504, new_n8503, new_n8505);
xnor_4 g08129(new_n8505, new_n8502, new_n8506);
and_5  g08130(n9400, n2433, new_n8507);
and_5  g08131(n8819, n2464, new_n8508);
xnor_4 g08132(new_n8508, new_n8507, new_n8509);
xnor_4 g08133(new_n8509, new_n8506, new_n8510);
nor_5  g08134(new_n8483, new_n8479, new_n8511);
nor_5  g08135(new_n8489, new_n8484, new_n8512);
nor_5  g08136(new_n8512, new_n8511, new_n8513);
xnor_4 g08137(new_n8513, new_n8510, new_n8514);
nor_5  g08138(new_n8490, new_n8478, new_n8515);
nor_5  g08139(new_n8494, new_n8491, new_n8516);
nor_5  g08140(new_n8516, new_n8515, new_n8517);
xnor_4 g08141(new_n8517, new_n8514, new_n8518);
xnor_4 g08142(new_n8518, new_n8497, new_n8519);
xor_4  g08143(new_n8519, new_n8496, new_n8520);
xor_4  g08144(new_n8495, new_n8477, new_n8521);
xnor_4 g08145(new_n8476_1, new_n8471, new_n8522);
and_5  g08146(n12489, n4805, new_n8523);
and_5  g08147(n10990, n7236, new_n8524);
and_5  g08148(new_n8524, new_n8523, new_n8525);
and_5  g08149(n12489, n11478, new_n8526);
and_5  g08150(n7159, n4805, new_n8527);
xor_4  g08151(new_n8527, new_n8526, new_n8528);
nor_5  g08152(new_n8528, new_n8525, new_n8529);
xnor_4 g08153(new_n8528, new_n8525, new_n8530);
and_5  g08154(n10990, n3992, new_n8531);
and_5  g08155(n7236, n5760, new_n8532);
xor_4  g08156(new_n8532, new_n8531, new_n8533);
nor_5  g08157(new_n8533, new_n8530, new_n8534);
nor_5  g08158(new_n8534, new_n8529, new_n8535);
and_5  g08159(n10990, n8384, new_n8536);
and_5  g08160(n7236, n1478, new_n8537);
and_5  g08161(new_n8537, new_n8536, new_n8538);
nand_5 g08162(n5760, n3992, new_n8539);
or_5   g08163(new_n8539, new_n8524, new_n8540);
nor_5  g08164(new_n8537, new_n8536, new_n8541);
and_5  g08165(new_n8541, new_n8540, new_n8542);
nor_5  g08166(new_n8542, new_n8538, new_n8543);
or_5   g08167(new_n8541, new_n8540, new_n8544);
and_5  g08168(new_n8544, new_n8543, new_n8545);
nor_5  g08169(new_n8545, new_n8535, new_n8546);
xnor_4 g08170(new_n8545, new_n8535, new_n8547);
nand_5 g08171(n11478, n7159, new_n8548);
nor_5  g08172(new_n8548, new_n8523, new_n8549);
and_5  g08173(n12489, n5283, new_n8550);
and_5  g08174(n12777, n4805, new_n8551);
xor_4  g08175(new_n8551, new_n8550, new_n8552);
nor_5  g08176(new_n8552, new_n8549, new_n8553);
or_5   g08177(new_n8548, new_n8523, new_n8554);
nor_5  g08178(new_n8551, new_n8550, new_n8555);
nor_5  g08179(new_n8555, new_n8554, new_n8556);
nor_5  g08180(new_n8556, new_n8553, new_n8557);
nor_5  g08181(new_n8557, new_n8547, new_n8558);
nor_5  g08182(new_n8558, new_n8546, new_n8559);
nand_5 g08183(n6254, n4805, new_n8560);
and_5  g08184(new_n8551, new_n8550, new_n8561);
nor_5  g08185(new_n8555, new_n8548, new_n8562);
nor_5  g08186(new_n8562, new_n8561, new_n8563);
xnor_4 g08187(new_n8563, new_n8560, new_n8564);
and_5  g08188(n7159, n5283, new_n8565);
and_5  g08189(n12489, n137, new_n8566);
and_5  g08190(n12777, n11478, new_n8567);
xnor_4 g08191(new_n8567, new_n8566, new_n8568);
xor_4  g08192(new_n8568, new_n8565, new_n8569);
xnor_4 g08193(new_n8569, new_n8564, new_n8570);
nand_5 g08194(new_n8527, new_n8526, new_n8571);
or_5   g08195(new_n8552, new_n8571, new_n8572);
xor_4  g08196(new_n8572, new_n8570, new_n8573);
and_5  g08197(n11791, n7236, new_n8574);
and_5  g08198(n5760, n3992, new_n8575);
nor_5  g08199(new_n8575, new_n8538, new_n8576);
nor_5  g08200(new_n8576, new_n8541, new_n8577);
xnor_4 g08201(new_n8577, new_n8574, new_n8578);
and_5  g08202(n8384, n5760, new_n8579);
and_5  g08203(n10990, n6358, new_n8580);
and_5  g08204(n3992, n1478, new_n8581);
xnor_4 g08205(new_n8581, new_n8580, new_n8582);
xor_4  g08206(new_n8582, new_n8579, new_n8583);
xnor_4 g08207(new_n8583, new_n8578, new_n8584);
or_5   g08208(new_n8543, new_n8539, new_n8585);
xor_4  g08209(new_n8585, new_n8584, new_n8586);
xnor_4 g08210(new_n8586, new_n8573, new_n8587);
xor_4  g08211(new_n8587, new_n8559, new_n8588);
nor_5  g08212(new_n8588, new_n8522, new_n8589);
xnor_4 g08213(new_n8588, new_n8522, new_n8590);
xor_4  g08214(new_n8557, new_n8547, new_n8591);
and_5  g08215(n12709, n6877, new_n8592);
nor_5  g08216(new_n8592, new_n8462, new_n8593);
nor_5  g08217(new_n8593, new_n8472, new_n8594);
or_5   g08218(new_n8592, new_n8462, new_n8595_1);
nor_5  g08219(new_n8595_1, new_n8461, new_n8596);
or_5   g08220(new_n8596, new_n8594, new_n8597);
nor_5  g08221(new_n8597, new_n8591, new_n8598);
xnor_4 g08222(new_n8597, new_n8591, new_n8599);
xor_4  g08223(new_n8533, new_n8530, new_n8600);
xnor_4 g08224(new_n8474, new_n8473, new_n8601);
nor_5  g08225(new_n8601, new_n8600, new_n8602);
nand_5 g08226(n12709, n6877, new_n8603);
xnor_4 g08227(new_n8524, new_n8523, new_n8604);
or_5   g08228(new_n8604, new_n8603, new_n8605);
xnor_4 g08229(new_n8601, new_n8600, new_n8606);
nor_5  g08230(new_n8606, new_n8605, new_n8607);
nor_5  g08231(new_n8607, new_n8602, new_n8608);
nor_5  g08232(new_n8608, new_n8599, new_n8609);
nor_5  g08233(new_n8609, new_n8598, new_n8610);
nor_5  g08234(new_n8610, new_n8590, new_n8611);
or_5   g08235(new_n8611, new_n8589, new_n8612);
nor_5  g08236(new_n8612, new_n8521, new_n8613);
xnor_4 g08237(new_n8612, new_n8521, new_n8614);
or_5   g08238(new_n8572, new_n8570, new_n8615);
and_5  g08239(n7159, n137, new_n8616);
and_5  g08240(n12777, n5283, new_n8617);
and_5  g08241(n12489, n6294, new_n8618);
xnor_4 g08242(new_n8618, new_n8617, new_n8619);
xor_4  g08243(new_n8619, new_n8616, new_n8620);
and_5  g08244(n11478, n6254, new_n8621);
nor_5  g08245(new_n8567, new_n8566, new_n8622);
nor_5  g08246(new_n8568, new_n8565, new_n8623);
nor_5  g08247(new_n8623, new_n8622, new_n8624);
xnor_4 g08248(new_n8624, new_n8621, new_n8625);
xor_4  g08249(new_n8625, new_n8620, new_n8626);
and_5  g08250(n11967, n4805, new_n8627);
nor_5  g08251(new_n8563, new_n8560, new_n8628);
nor_5  g08252(new_n8569, new_n8564, new_n8629);
or_5   g08253(new_n8629, new_n8628, new_n8630);
xnor_4 g08254(new_n8630, new_n8627, new_n8631);
xor_4  g08255(new_n8631, new_n8626, new_n8632);
xor_4  g08256(new_n8632, new_n8615, new_n8633);
or_5   g08257(new_n8585, new_n8584, new_n8634);
and_5  g08258(n6358, n5760, new_n8635);
and_5  g08259(n8384, n1478, new_n8636);
and_5  g08260(n10990, n5198, new_n8637);
xnor_4 g08261(new_n8637, new_n8636, new_n8638);
xor_4  g08262(new_n8638, new_n8635, new_n8639);
and_5  g08263(n11791, n3992, new_n8640);
nor_5  g08264(new_n8581, new_n8580, new_n8641);
nor_5  g08265(new_n8582, new_n8579, new_n8642);
nor_5  g08266(new_n8642, new_n8641, new_n8643);
xnor_4 g08267(new_n8643, new_n8640, new_n8644);
xor_4  g08268(new_n8644, new_n8639, new_n8645);
nand_5 g08269(n12947, n7236, new_n8646);
and_5  g08270(new_n8577, new_n8574, new_n8647);
nor_5  g08271(new_n8583, new_n8578, new_n8648);
nor_5  g08272(new_n8648, new_n8647, new_n8649);
xnor_4 g08273(new_n8649, new_n8646, new_n8650);
xor_4  g08274(new_n8650, new_n8645, new_n8651);
xor_4  g08275(new_n8651, new_n8634, new_n8652);
xnor_4 g08276(new_n8652, new_n8633, new_n8653);
nor_5  g08277(new_n8586, new_n8573, new_n8654);
nor_5  g08278(new_n8587, new_n8559, new_n8655);
or_5   g08279(new_n8655, new_n8654, new_n8656);
xor_4  g08280(new_n8656, new_n8653, new_n8657);
nor_5  g08281(new_n8657, new_n8614, new_n8658);
nor_5  g08282(new_n8658, new_n8613, new_n8659);
nor_5  g08283(new_n8659, new_n8520, new_n8660);
or_5   g08284(new_n8651, new_n8634, new_n8661);
and_5  g08285(n7236, n6441, new_n8662);
and_5  g08286(new_n8643, new_n8640, new_n8663);
nor_5  g08287(new_n8644, new_n8639, new_n8664);
nor_5  g08288(new_n8664, new_n8663, new_n8665_1);
and_5  g08289(n12947, n3992, new_n8666);
and_5  g08290(n11791, n8384, new_n8667);
xnor_4 g08291(new_n8667, new_n8666, new_n8668);
xnor_4 g08292(new_n8668, new_n8665_1, new_n8669);
nand_5 g08293(n6358, n1478, new_n8670);
and_5  g08294(n5760, n5198, new_n8671);
and_5  g08295(n10990, n1471, new_n8672);
xnor_4 g08296(new_n8672, new_n8671, new_n8673);
xnor_4 g08297(new_n8673, new_n8670, new_n8674);
nor_5  g08298(new_n8637, new_n8636, new_n8675);
nor_5  g08299(new_n8638, new_n8635, new_n8676);
or_5   g08300(new_n8676, new_n8675, new_n8677);
xnor_4 g08301(new_n8677, new_n8674, new_n8678);
xnor_4 g08302(new_n8678, new_n8669, new_n8679);
and_5  g08303(new_n8649, new_n8646, new_n8680);
nor_5  g08304(new_n8650, new_n8645, new_n8681);
or_5   g08305(new_n8681, new_n8680, new_n8682);
xor_4  g08306(new_n8682, new_n8679, new_n8683);
xnor_4 g08307(new_n8683, new_n8662, new_n8684);
xor_4  g08308(new_n8684, new_n8661, new_n8685);
or_5   g08309(new_n8632, new_n8615, new_n8686);
and_5  g08310(n4805, n447, new_n8687);
and_5  g08311(new_n8624, new_n8621, new_n8688);
nor_5  g08312(new_n8625, new_n8620, new_n8689);
nor_5  g08313(new_n8689, new_n8688, new_n8690);
and_5  g08314(n11967, n11478, new_n8691);
and_5  g08315(n6254, n5283, new_n8692);
xnor_4 g08316(new_n8692, new_n8691, new_n8693);
xnor_4 g08317(new_n8693, new_n8690, new_n8694);
nand_5 g08318(n12777, n137, new_n8695);
and_5  g08319(n7159, n6294, new_n8696);
and_5  g08320(n12489, n6797, new_n8697);
xnor_4 g08321(new_n8697, new_n8696, new_n8698);
xnor_4 g08322(new_n8698, new_n8695, new_n8699);
nor_5  g08323(new_n8618, new_n8617, new_n8700);
nor_5  g08324(new_n8619, new_n8616, new_n8701);
or_5   g08325(new_n8701, new_n8700, new_n8702);
xnor_4 g08326(new_n8702, new_n8699, new_n8703);
xnor_4 g08327(new_n8703, new_n8694, new_n8704);
nor_5  g08328(new_n8630, new_n8627, new_n8705);
nor_5  g08329(new_n8631, new_n8626, new_n8706);
or_5   g08330(new_n8706, new_n8705, new_n8707);
xor_4  g08331(new_n8707, new_n8704, new_n8708);
xnor_4 g08332(new_n8708, new_n8687, new_n8709);
xor_4  g08333(new_n8709, new_n8686, new_n8710);
and_5  g08334(new_n8652, new_n8633, new_n8711);
nor_5  g08335(new_n8656, new_n8653, new_n8712);
or_5   g08336(new_n8712, new_n8711, new_n8713);
xnor_4 g08337(new_n8713, new_n8710, new_n8714);
xnor_4 g08338(new_n8714, new_n8685, new_n8715);
xnor_4 g08339(new_n8659, new_n8520, new_n8716);
nor_5  g08340(new_n8716, new_n8715, new_n8717_1);
nor_5  g08341(new_n8717_1, new_n8660, new_n8718);
or_5   g08342(new_n8517, new_n8514, new_n8719);
nor_5  g08343(new_n8509, new_n8506, new_n8720);
nand_5 g08344(new_n8508, new_n8507, new_n8721);
or_5   g08345(new_n8513, new_n8510, new_n8722);
xor_4  g08346(new_n8722, new_n8721, new_n8723);
nor_5  g08347(new_n8723, new_n8720, new_n8724);
nor_5  g08348(new_n8501, new_n8498, new_n8725);
nor_5  g08349(new_n8505, new_n8502, new_n8726);
nor_5  g08350(new_n8726, new_n8725, new_n8727);
and_5  g08351(n9400, n8717, new_n8728);
and_5  g08352(n2464, n2433, new_n8729);
and_5  g08353(n7730, n6877, new_n8730);
xnor_4 g08354(new_n8730, new_n8729, new_n8731);
xor_4  g08355(new_n8731, new_n8728, new_n8732);
xnor_4 g08356(new_n8732, new_n8727, new_n8733);
and_5  g08357(new_n8500, new_n8499, new_n8734);
and_5  g08358(n11311, n8819, new_n8735);
xnor_4 g08359(new_n8735, new_n8734, new_n8736);
and_5  g08360(n11728, n4203, new_n8737);
and_5  g08361(n6429, n4187, new_n8738);
and_5  g08362(n12753, n12709, new_n8739);
xnor_4 g08363(new_n8739, new_n8738, new_n8740);
xor_4  g08364(new_n8740, new_n8737, new_n8741);
xnor_4 g08365(new_n8741, new_n8736, new_n8742);
xnor_4 g08366(new_n8742, new_n8733, new_n8743);
xnor_4 g08367(new_n8743, new_n8724, new_n8744);
xnor_4 g08368(new_n8744, new_n8719, new_n8745);
nor_5  g08369(new_n8518, new_n8497, new_n8746);
nor_5  g08370(new_n8519, new_n8496, new_n8747);
nor_5  g08371(new_n8747, new_n8746, new_n8748);
xor_4  g08372(new_n8748, new_n8745, new_n8749);
or_5   g08373(new_n8707, new_n8704, new_n8750);
and_5  g08374(n11478, n447, new_n8751);
nand_5 g08375(n11967, n5283, new_n8752);
nand_5 g08376(n4805, n1353, new_n8753);
xnor_4 g08377(new_n8753, new_n8752, new_n8754);
xnor_4 g08378(new_n8754, new_n8751, new_n8755);
nor_5  g08379(new_n8698, new_n8695, new_n8756);
nor_5  g08380(new_n8702, new_n8699, new_n8757);
or_5   g08381(new_n8757, new_n8756, new_n8758);
xnor_4 g08382(new_n8758, new_n8755, new_n8759_1);
and_5  g08383(new_n8697, new_n8696, new_n8760);
and_5  g08384(n6254, n137, new_n8761);
xnor_4 g08385(new_n8761, new_n8760, new_n8762);
nand_5 g08386(n7159, n6797, new_n8763);
and_5  g08387(n12777, n6294, new_n8764);
and_5  g08388(n12489, n3146, new_n8765);
xnor_4 g08389(new_n8765, new_n8764, new_n8766);
xnor_4 g08390(new_n8766, new_n8763, new_n8767);
xor_4  g08391(new_n8767, new_n8762, new_n8768);
xor_4  g08392(new_n8768, new_n8759_1, new_n8769);
nor_5  g08393(new_n8693, new_n8690, new_n8770);
nand_5 g08394(new_n8692, new_n8691, new_n8771);
or_5   g08395(new_n8703, new_n8694, new_n8772);
xor_4  g08396(new_n8772, new_n8771, new_n8773);
nor_5  g08397(new_n8773, new_n8770, new_n8774);
xnor_4 g08398(new_n8774, new_n8769, new_n8775);
xnor_4 g08399(new_n8775, new_n8750, new_n8776);
and_5  g08400(new_n8708, new_n8687, new_n8777);
nor_5  g08401(new_n8709, new_n8686, new_n8778);
nor_5  g08402(new_n8778, new_n8777, new_n8779);
xnor_4 g08403(new_n8779, new_n8776, new_n8780);
or_5   g08404(new_n8682, new_n8679, new_n8781);
nor_5  g08405(new_n8673, new_n8670, new_n8782);
nor_5  g08406(new_n8677, new_n8674, new_n8783);
or_5   g08407(new_n8783, new_n8782, new_n8784);
and_5  g08408(n6441, n3992, new_n8785);
and_5  g08409(n12947, n8384, new_n8786);
and_5  g08410(n11999, n7236, new_n8787);
xnor_4 g08411(new_n8787, new_n8786, new_n8788);
xnor_4 g08412(new_n8788, new_n8785, new_n8789);
xnor_4 g08413(new_n8789, new_n8784, new_n8790);
and_5  g08414(new_n8672, new_n8671, new_n8791);
and_5  g08415(n11791, n6358, new_n8792);
xnor_4 g08416(new_n8792, new_n8791, new_n8793);
and_5  g08417(n5760, n1471, new_n8794);
and_5  g08418(n5198, n1478, new_n8795);
and_5  g08419(n10990, n7646, new_n8796);
xnor_4 g08420(new_n8796, new_n8795, new_n8797);
xor_4  g08421(new_n8797, new_n8794, new_n8798);
xor_4  g08422(new_n8798, new_n8793, new_n8799);
xor_4  g08423(new_n8799, new_n8790, new_n8800);
nor_5  g08424(new_n8668, new_n8665_1, new_n8801);
nand_5 g08425(new_n8667, new_n8666, new_n8802);
or_5   g08426(new_n8678, new_n8669, new_n8803);
xor_4  g08427(new_n8803, new_n8802, new_n8804);
nor_5  g08428(new_n8804, new_n8801, new_n8805);
xnor_4 g08429(new_n8805, new_n8800, new_n8806);
xnor_4 g08430(new_n8806, new_n8781, new_n8807);
and_5  g08431(new_n8683, new_n8662, new_n8808);
nor_5  g08432(new_n8684, new_n8661, new_n8809);
nor_5  g08433(new_n8809, new_n8808, new_n8810);
xnor_4 g08434(new_n8810, new_n8807, new_n8811);
xnor_4 g08435(new_n8811, new_n8780, new_n8812);
nor_5  g08436(new_n8713, new_n8710, new_n8813);
nor_5  g08437(new_n8714, new_n8685, new_n8814);
or_5   g08438(new_n8814, new_n8813, new_n8815);
xor_4  g08439(new_n8815, new_n8812, new_n8816);
xor_4  g08440(new_n8816, new_n8749, new_n8817);
xnor_4 g08441(new_n8817, new_n8718, new_n8818);
and_5  g08442(new_n8818, new_n8456, new_n8819_1);
xnor_4 g08443(new_n8818, new_n8456, new_n8820);
xnor_4 g08444(new_n8453, new_n8452, new_n8821);
xnor_4 g08445(new_n8451, new_n8450, new_n8822);
xor_4  g08446(new_n8657, new_n8614, new_n8823);
and_5  g08447(new_n8823, new_n8822, new_n8824);
xnor_4 g08448(new_n8823, new_n8822, new_n8825);
xor_4  g08449(new_n8449, new_n8444, new_n8826);
xor_4  g08450(new_n8610, new_n8590, new_n8827);
nor_5  g08451(new_n8827, new_n8826, new_n8828);
xnor_4 g08452(new_n8608, new_n8599, new_n8829);
or_5   g08453(new_n8400, new_n8399, new_n8830);
nand_5 g08454(n5212, n1333, new_n8831);
or_5   g08455(new_n8831, new_n8402, new_n8832);
nor_5  g08456(new_n8832, new_n8830, new_n8833);
and_5  g08457(new_n8832, new_n8445, new_n8834);
nor_5  g08458(new_n8834, new_n8833, new_n8835);
and_5  g08459(new_n8835, new_n8829, new_n8836);
xnor_4 g08460(new_n8835, new_n8829, new_n8837);
xnor_4 g08461(new_n8604, new_n8592, new_n8838);
and_5  g08462(new_n8838, new_n8402, new_n8839);
xor_4  g08463(new_n8447, new_n8446, new_n8840);
nor_5  g08464(new_n8840, new_n8839, new_n8841);
xnor_4 g08465(new_n8606, new_n8605, new_n8842);
xor_4  g08466(new_n8840, new_n8839, new_n8843);
and_5  g08467(new_n8843, new_n8842, new_n8844);
nor_5  g08468(new_n8844, new_n8841, new_n8845);
nor_5  g08469(new_n8845, new_n8837, new_n8846);
nor_5  g08470(new_n8846, new_n8836, new_n8847);
xnor_4 g08471(new_n8827, new_n8826, new_n8848);
nor_5  g08472(new_n8848, new_n8847, new_n8849);
nor_5  g08473(new_n8849, new_n8828, new_n8850);
nor_5  g08474(new_n8850, new_n8825, new_n8851);
nor_5  g08475(new_n8851, new_n8824, new_n8852);
nor_5  g08476(new_n8852, new_n8821, new_n8853);
xor_4  g08477(new_n8716, new_n8715, new_n8854);
xor_4  g08478(new_n8852, new_n8821, new_n8855);
and_5  g08479(new_n8855, new_n8854, new_n8856);
nor_5  g08480(new_n8856, new_n8853, new_n8857);
nor_5  g08481(new_n8857, new_n8820, new_n8858);
nor_5  g08482(new_n8858, new_n8819_1, new_n8859);
and_5  g08483(new_n8816, new_n8749, new_n8860);
or_5   g08484(new_n8816, new_n8749, new_n8861);
and_5  g08485(new_n8861, new_n8718, new_n8862);
nor_5  g08486(new_n8862, new_n8860, new_n8863);
nor_5  g08487(new_n8439, new_n8414, new_n8864);
nor_5  g08488(new_n8455, new_n8440, new_n8865);
nor_5  g08489(new_n8865, new_n8864, new_n8866);
nor_5  g08490(new_n8772, new_n8771, new_n8867);
nor_5  g08491(new_n8774, new_n8769, new_n8868);
or_5   g08492(new_n8868, new_n8867, new_n8869);
nor_5  g08493(new_n8787, new_n8786, new_n8870);
nor_5  g08494(new_n8788, new_n8785, new_n8871);
nor_5  g08495(new_n8871, new_n8870, new_n8872);
and_5  g08496(n4805, n4436, new_n8873);
and_5  g08497(n8384, n6441, new_n8874);
and_5  g08498(n11791, n5198, new_n8875);
xnor_4 g08499(new_n8875, new_n8874, new_n8876);
xnor_4 g08500(new_n8876, new_n8873, new_n8877);
xnor_4 g08501(new_n8877, new_n8872, new_n8878);
and_5  g08502(n7159, n3146, new_n8879);
and_5  g08503(n11967, n137, new_n8880);
xnor_4 g08504(new_n8880, new_n8879, new_n8881);
and_5  g08505(n6294, n6254, new_n8882);
and_5  g08506(n12947, n6358, new_n8883);
xnor_4 g08507(new_n8883, new_n8882, new_n8884);
and_5  g08508(n11407, n6826, new_n8885);
and_5  g08509(n7862, n6604, new_n8886);
xnor_4 g08510(new_n8886, new_n8885, new_n8887);
xnor_4 g08511(new_n8887, new_n8884, new_n8888);
xnor_4 g08512(new_n8888, new_n8881, new_n8889);
xnor_4 g08513(new_n8889, new_n8878, new_n8890);
nand_5 g08514(n6429, n4203, new_n8891);
and_5  g08515(new_n8761, new_n8760, new_n8892);
nor_5  g08516(new_n8767, new_n8762, new_n8893);
nor_5  g08517(new_n8893, new_n8892, new_n8894);
xnor_4 g08518(new_n8894, new_n8891, new_n8895);
xnor_4 g08519(new_n8895, new_n8890, new_n8896);
nor_5  g08520(new_n8758, new_n8755, new_n8897);
nor_5  g08521(new_n8768, new_n8759_1, new_n8898);
nor_5  g08522(new_n8898, new_n8897, new_n8899);
nor_5  g08523(new_n8789, new_n8784, new_n8900);
nor_5  g08524(new_n8799, new_n8790, new_n8901);
nor_5  g08525(new_n8901, new_n8900, new_n8902);
nand_5 g08526(n11478, n1353, new_n8903);
nor_5  g08527(new_n8754, new_n8751, new_n8904);
or_5   g08528(new_n8904, new_n8752, new_n8905);
nor_5  g08529(new_n8905, new_n8903, new_n8906);
or_5   g08530(new_n8903, new_n8687, new_n8907);
and_5  g08531(new_n8907, new_n8905, new_n8908);
nor_5  g08532(new_n8908, new_n8906, new_n8909);
and_5  g08533(new_n8765, new_n8764, new_n8910);
nor_5  g08534(new_n8765, new_n8764, new_n8911);
nor_5  g08535(new_n8911, new_n8763, new_n8912);
nor_5  g08536(new_n8912, new_n8910, new_n8913);
xnor_4 g08537(new_n8913, new_n8909, new_n8914);
xnor_4 g08538(new_n8914, new_n8902, new_n8915);
xnor_4 g08539(new_n8915, new_n8899, new_n8916);
xnor_4 g08540(new_n8916, new_n8896, new_n8917);
nor_5  g08541(new_n8417, new_n8416, new_n8918);
nor_5  g08542(new_n8438, new_n8419, new_n8919);
nor_5  g08543(new_n8919, new_n8918, new_n8920);
nand_5 g08544(n12777, n6797, new_n8921);
xnor_4 g08545(new_n8921, new_n8920, new_n8922);
xnor_4 g08546(new_n8922, new_n8917, new_n8923);
xnor_4 g08547(new_n8923, new_n8869, new_n8924);
xnor_4 g08548(new_n8924, new_n8866, new_n8925);
xnor_4 g08549(new_n8925, new_n8863, new_n8926);
nor_5  g08550(new_n8744, new_n8719, new_n8927);
nor_5  g08551(new_n8748, new_n8745, new_n8928);
nor_5  g08552(new_n8928, new_n8927, new_n8929);
nor_5  g08553(new_n8775, new_n8750, new_n8930);
nor_5  g08554(new_n8779, new_n8776, new_n8931);
nor_5  g08555(new_n8931, new_n8930, new_n8932);
xnor_4 g08556(new_n8932, new_n8929, new_n8933);
nor_5  g08557(new_n8806, new_n8781, new_n8934);
nor_5  g08558(new_n8810, new_n8807, new_n8935);
nor_5  g08559(new_n8935, new_n8934, new_n8936);
nor_5  g08560(new_n8732, new_n8727, new_n8937);
nor_5  g08561(new_n8742, new_n8733, new_n8938);
nor_5  g08562(new_n8938, new_n8937, new_n8939);
nor_5  g08563(new_n8730, new_n8729, new_n8940);
nor_5  g08564(new_n8731, new_n8728, new_n8941);
nor_5  g08565(new_n8941, new_n8940, new_n8942);
and_5  g08566(n5283, n447, new_n8943);
and_5  g08567(n11999, n3992, new_n8944);
xnor_4 g08568(new_n8944, new_n8943, new_n8945);
xnor_4 g08569(new_n8945, new_n8942, new_n8946);
xnor_4 g08570(new_n8946, new_n8939, new_n8947);
and_5  g08571(n7646, n5760, new_n8948);
and_5  g08572(n10990, n4722, new_n8949);
xnor_4 g08573(new_n8949, new_n8948, new_n8950);
xnor_4 g08574(new_n8950, new_n8947, new_n8951);
xnor_4 g08575(new_n8951, new_n8936, new_n8952);
xnor_4 g08576(new_n8952, new_n8933, new_n8953);
nor_5  g08577(new_n8811, new_n8780, new_n8954);
nor_5  g08578(new_n8815, new_n8812, new_n8955);
nor_5  g08579(new_n8955, new_n8954, new_n8956);
nor_5  g08580(new_n8722, new_n8721, new_n8957);
nor_5  g08581(new_n8743, new_n8724, new_n8958);
nor_5  g08582(new_n8958, new_n8957, new_n8959);
nor_5  g08583(new_n8436, new_n8431, new_n8960);
nor_5  g08584(new_n8437, new_n8428, new_n8961);
nor_5  g08585(new_n8961, new_n8960, new_n8962);
nor_5  g08586(new_n8739, new_n8738, new_n8963);
nor_5  g08587(new_n8740, new_n8737, new_n8964);
nor_5  g08588(new_n8964, new_n8963, new_n8965);
nand_5 g08589(n12000, n3172, new_n8966);
and_5  g08590(n9725, n1333, new_n8967);
and_5  g08591(n12709, n10174, new_n8968);
xnor_4 g08592(new_n8968, new_n8967, new_n8969);
xnor_4 g08593(new_n8969, new_n8966, new_n8970);
xnor_4 g08594(new_n8970, new_n8965, new_n8971);
and_5  g08595(new_n8735, new_n8734, new_n8972);
nor_5  g08596(new_n8741, new_n8736, new_n8973);
nor_5  g08597(new_n8973, new_n8972, new_n8974);
nor_5  g08598(new_n8796, new_n8795, new_n8975);
nor_5  g08599(new_n8797, new_n8794, new_n8976);
nor_5  g08600(new_n8976, new_n8975, new_n8977);
and_5  g08601(n6877, n1198, new_n8978);
and_5  g08602(n12753, n11728, new_n8979);
xor_4  g08603(new_n8979, new_n8978, new_n8980);
xnor_4 g08604(new_n8980, new_n8977, new_n8981);
xnor_4 g08605(new_n8981, new_n8974, new_n8982);
xnor_4 g08606(new_n8982, new_n8971, new_n8983);
xnor_4 g08607(new_n8983, new_n8962, new_n8984);
and_5  g08608(n12489, n4938, new_n8985);
nor_5  g08609(new_n8434, new_n8433_1, new_n8986);
nor_5  g08610(new_n8435, new_n8432, new_n8987);
nor_5  g08611(new_n8987, new_n8986, new_n8988);
and_5  g08612(n11757, n5320, new_n8989);
and_5  g08613(n9080, n5212, new_n8990);
xnor_4 g08614(new_n8990, new_n8989, new_n8991);
and_5  g08615(n11877, n11821, new_n8992);
and_5  g08616(n5240, n4370, new_n8993);
xnor_4 g08617(new_n8993, new_n8992, new_n8994);
xor_4  g08618(new_n8994, new_n8991, new_n8995);
xnor_4 g08619(new_n8995, new_n8988, new_n8996);
and_5  g08620(n9400, n7730, new_n8997);
and_5  g08621(n11311, n2433, new_n8998);
xnor_4 g08622(new_n8998, new_n8997, new_n8999);
xnor_4 g08623(new_n8999, new_n8996, new_n9000);
nor_5  g08624(new_n8425, new_n8424, new_n9001);
nor_5  g08625(new_n8426, new_n8423, new_n9002);
or_5   g08626(new_n9002, new_n9001, new_n9003);
nor_5  g08627(new_n8421, new_n8420, new_n9004);
nor_5  g08628(new_n8427, new_n8422, new_n9005);
nor_5  g08629(new_n9005, new_n9004, new_n9006);
xnor_4 g08630(new_n9006, new_n9003, new_n9007);
xnor_4 g08631(new_n9007, new_n9000, new_n9008);
xnor_4 g08632(new_n9008, new_n8985, new_n9009);
xnor_4 g08633(new_n9009, new_n8984, new_n9010);
xnor_4 g08634(new_n9010, new_n8959, new_n9011);
nor_5  g08635(new_n8803, new_n8802, new_n9012);
nor_5  g08636(new_n8805, new_n8800, new_n9013);
nor_5  g08637(new_n9013, new_n9012, new_n9014);
and_5  g08638(n8819, n4187, new_n9015);
and_5  g08639(n1478, n1471, new_n9016);
xnor_4 g08640(new_n9016, new_n9015, new_n9017);
and_5  g08641(n8717, n2464, new_n9018);
and_5  g08642(n10022, n7236, new_n9019);
xnor_4 g08643(new_n9019, new_n9018, new_n9020);
xnor_4 g08644(new_n9020, new_n9017, new_n9021);
and_5  g08645(new_n8792, new_n8791, new_n9022);
nor_5  g08646(new_n8798, new_n8793, new_n9023);
nor_5  g08647(new_n9023, new_n9022, new_n9024);
xnor_4 g08648(new_n9024, new_n9021, new_n9025);
xnor_4 g08649(new_n9025, new_n9014, new_n9026);
xnor_4 g08650(new_n9026, new_n9011, new_n9027);
xnor_4 g08651(new_n9027, new_n8956, new_n9028);
xor_4  g08652(new_n9028, new_n8953, new_n9029);
xnor_4 g08653(new_n9029, new_n8926, new_n9030);
xnor_4 g08654(new_n9030, new_n8859, n4378);
xor_4  g08655(new_n3101, new_n3021, n4397);
xor_4  g08656(new_n3328, new_n3169, n4553);
xor_4  g08657(new_n757, new_n750, n4686);
xnor_4 g08658(new_n7436_1, new_n7419, n4689);
xor_4  g08659(new_n3915, new_n3914, n4733);
xnor_4 g08660(new_n1667, new_n1660, n4757);
xnor_4 g08661(new_n3910, new_n3909, n4971);
xnor_4 g08662(new_n5195, new_n5194, n5030);
xnor_4 g08663(new_n2342, new_n2317, n5034);
xnor_4 g08664(new_n2337, new_n2329, n5094);
and_5  g08665(new_n8281, new_n8278, new_n9042);
nor_5  g08666(new_n8287, new_n8282, new_n9043);
nor_5  g08667(new_n9043, new_n9042, new_n9044);
and_5  g08668(n5320, n2564, new_n9045);
and_5  g08669(n4370, n4189, new_n9046);
xnor_4 g08670(new_n9046, new_n9045, new_n9047);
xnor_4 g08671(new_n9047, new_n9044, new_n9048);
and_5  g08672(n11877, n6770, new_n9049);
nor_5  g08673(new_n8285, new_n8284, new_n9050);
nor_5  g08674(new_n8286, new_n8283, new_n9051);
nor_5  g08675(new_n9051, new_n9050, new_n9052);
xnor_4 g08676(new_n9052, new_n9049, new_n9053);
and_5  g08677(n9920, n5212, new_n9054);
and_5  g08678(n11407, n3627, new_n9055);
xnor_4 g08679(new_n9055, new_n9054, new_n9056);
xnor_4 g08680(new_n9056, new_n9053, new_n9057);
xnor_4 g08681(new_n9057, new_n9048, new_n9058);
nor_5  g08682(new_n8276_1, new_n8273, new_n9059);
nor_5  g08683(new_n8288, new_n8277, new_n9060);
nor_5  g08684(new_n9060, new_n9059, new_n9061);
or_5   g08685(new_n9061, new_n9058, new_n9062);
and_5  g08686(new_n9052, new_n9049, new_n9063);
nor_5  g08687(new_n9056, new_n9053, new_n9064);
or_5   g08688(new_n9064, new_n9063, new_n9065);
nand_5 g08689(n12000, n2564, new_n9066);
and_5  g08690(n5320, n4189, new_n9067);
and_5  g08691(n9725, n6687, new_n9068);
xnor_4 g08692(new_n9068, new_n9067, new_n9069);
xor_4  g08693(new_n9069, new_n9066, new_n9070);
xnor_4 g08694(new_n9070, new_n9065, new_n9071);
and_5  g08695(new_n9055, new_n9054, new_n9072);
and_5  g08696(n6770, n4370, new_n9073);
xnor_4 g08697(new_n9073, new_n9072, new_n9074);
nand_5 g08698(n5212, n3627, new_n9075);
and_5  g08699(n11877, n9920, new_n9076);
and_5  g08700(n11407, n4516, new_n9077);
xnor_4 g08701(new_n9077, new_n9076, new_n9078);
xnor_4 g08702(new_n9078, new_n9075, new_n9079);
xor_4  g08703(new_n9079, new_n9074, new_n9080_1);
xor_4  g08704(new_n9080_1, new_n9071, new_n9081);
nor_5  g08705(new_n9047, new_n9044, new_n9082);
nand_5 g08706(new_n9046, new_n9045, new_n9083);
or_5   g08707(new_n9057, new_n9048, new_n9084);
xor_4  g08708(new_n9084, new_n9083, new_n9085);
nor_5  g08709(new_n9085, new_n9082, new_n9086);
xnor_4 g08710(new_n9086, new_n9081, new_n9087);
xnor_4 g08711(new_n9087, new_n9062, new_n9088);
nand_5 g08712(n12000, n6687, new_n9089);
xnor_4 g08713(new_n9061, new_n9058, new_n9090);
nor_5  g08714(new_n9090, new_n9089, new_n9091);
or_5   g08715(new_n8289, new_n8272, new_n9092);
xnor_4 g08716(new_n9090, new_n9089, new_n9093);
nor_5  g08717(new_n9093, new_n9092, new_n9094);
nor_5  g08718(new_n9094, new_n9091, new_n9095);
xor_4  g08719(new_n9095, new_n9088, new_n9096);
nand_5 g08720(n8717, n8336, new_n9097);
nand_5 g08721(n6429, n2226, new_n9098);
and_5  g08722(n11728, n1094, new_n9099);
and_5  g08723(n12709, n10678, new_n9100);
xnor_4 g08724(new_n9100, new_n9099, new_n9101);
xnor_4 g08725(new_n9101, new_n9098, new_n9102);
nor_5  g08726(new_n8300, new_n1088, new_n9103);
and_5  g08727(new_n8300, new_n1088, new_n9104);
nor_5  g08728(new_n9104, new_n8299, new_n9105);
or_5   g08729(new_n9105, new_n9103, new_n9106);
xnor_4 g08730(new_n9106, new_n9102, new_n9107);
and_5  g08731(n10928, n2433, new_n9108);
and_5  g08732(n8819, n6986, new_n9109);
xnor_4 g08733(new_n9109, new_n9108, new_n9110);
xnor_4 g08734(new_n9110, new_n9107, new_n9111_1);
nor_5  g08735(new_n8297, new_n8293, new_n9112);
nor_5  g08736(new_n8302, new_n8298, new_n9113);
nor_5  g08737(new_n9113, new_n9112, new_n9114);
xnor_4 g08738(new_n9114, new_n9111_1, new_n9115);
nor_5  g08739(new_n8303_1, new_n8292, new_n9116);
nor_5  g08740(new_n8307, new_n8304, new_n9117);
nor_5  g08741(new_n9117, new_n9116, new_n9118);
xnor_4 g08742(new_n9118, new_n9115, new_n9119);
nor_5  g08743(new_n9119, new_n9097, new_n9120);
or_5   g08744(new_n8308, new_n8291, new_n9121);
xnor_4 g08745(new_n9119, new_n9097, new_n9122);
nor_5  g08746(new_n9122, new_n9121, new_n9123);
nor_5  g08747(new_n9123, new_n9120, new_n9124);
or_5   g08748(new_n9118, new_n9115, new_n9125);
nor_5  g08749(new_n9101, new_n9098, new_n9126);
nor_5  g08750(new_n9106, new_n9102, new_n9127);
or_5   g08751(new_n9127, new_n9126, new_n9128);
and_5  g08752(n10928, n8717, new_n9129);
and_5  g08753(n6986, n2433, new_n9130);
and_5  g08754(n8336, n7730, new_n9131);
xnor_4 g08755(new_n9131, new_n9130, new_n9132);
xnor_4 g08756(new_n9132, new_n9129, new_n9133);
xnor_4 g08757(new_n9133, new_n9128, new_n9134);
and_5  g08758(new_n9100, new_n9099, new_n9135);
and_5  g08759(n8819, n2226, new_n9136);
xnor_4 g08760(new_n9136, new_n9135, new_n9137_1);
and_5  g08761(n11728, n10678, new_n9138);
and_5  g08762(n6429, n1094, new_n9139);
and_5  g08763(n12709, n7320, new_n9140);
xnor_4 g08764(new_n9140, new_n9139, new_n9141);
xor_4  g08765(new_n9141, new_n9138, new_n9142);
xor_4  g08766(new_n9142, new_n9137_1, new_n9143);
xor_4  g08767(new_n9143, new_n9134, new_n9144);
nor_5  g08768(new_n9110, new_n9107, new_n9145);
nand_5 g08769(new_n9109, new_n9108, new_n9146);
or_5   g08770(new_n9114, new_n9111_1, new_n9147);
xor_4  g08771(new_n9147, new_n9146, new_n9148);
nor_5  g08772(new_n9148, new_n9145, new_n9149);
xnor_4 g08773(new_n9149, new_n9144, new_n9150);
xnor_4 g08774(new_n9150, new_n9125, new_n9151);
xor_4  g08775(new_n9151, new_n9124, new_n9152);
xor_4  g08776(new_n9122, new_n9121, new_n9153);
nor_5  g08777(new_n8312, new_n8309, new_n9154);
nor_5  g08778(new_n8356, new_n8313, new_n9155);
or_5   g08779(new_n9155, new_n9154, new_n9156);
nor_5  g08780(new_n9156, new_n9153, new_n9157);
or_5   g08781(new_n8350, new_n8333, new_n9158);
nand_5 g08782(n11222, n6441, new_n9159);
and_5  g08783(new_n8338, new_n8335, new_n9160);
nor_5  g08784(new_n8344, new_n8339, new_n9161);
nor_5  g08785(new_n9161, new_n9160, new_n9162);
and_5  g08786(n12947, n11153, new_n9163);
and_5  g08787(n11791, n5314, new_n9164);
xnor_4 g08788(new_n9164, new_n9163, new_n9165);
xnor_4 g08789(new_n9165, new_n9162, new_n9166);
nand_5 g08790(n1478, n996, new_n9167);
and_5  g08791(n10990, n5319, new_n9168);
and_5  g08792(n5767, n5760, new_n9169);
xnor_4 g08793(new_n9169, new_n9168, new_n9170);
xnor_4 g08794(new_n9170, new_n9167, new_n9171);
nor_5  g08795(new_n8342, new_n8341, new_n9172);
and_5  g08796(new_n8342, new_n8341, new_n9173);
nor_5  g08797(new_n9173, new_n8340, new_n9174);
or_5   g08798(new_n9174, new_n9172, new_n9175);
xnor_4 g08799(new_n9175, new_n9171, new_n9176);
xnor_4 g08800(new_n9176, new_n9166, new_n9177);
nor_5  g08801(new_n8345, new_n8334, new_n9178);
nor_5  g08802(new_n8349, new_n8346, new_n9179);
nor_5  g08803(new_n9179, new_n9178, new_n9180);
xnor_4 g08804(new_n9180, new_n9177, new_n9181);
xnor_4 g08805(new_n9181, new_n9159, new_n9182);
xnor_4 g08806(new_n9182, new_n9158, new_n9183);
nor_5  g08807(new_n8331, new_n8314, new_n9184);
and_5  g08808(n12069, n447, new_n9185);
nand_5 g08809(n12777, n7160, new_n9186);
and_5  g08810(n7159, n4828, new_n9187);
and_5  g08811(n12489, n2515, new_n9188);
xnor_4 g08812(new_n9188, new_n9187, new_n9189_1);
xnor_4 g08813(new_n9189_1, new_n9186, new_n9190);
nor_5  g08814(new_n8323, new_n8322, new_n9191);
and_5  g08815(new_n8323, new_n8322, new_n9192);
nor_5  g08816(new_n9192, new_n8321, new_n9193);
or_5   g08817(new_n9193, new_n9191, new_n9194);
xnor_4 g08818(new_n9194, new_n9190, new_n9195_1);
and_5  g08819(n12391, n11967, new_n9196);
and_5  g08820(n7891, n6254, new_n9197);
xnor_4 g08821(new_n9197, new_n9196, new_n9198);
xnor_4 g08822(new_n9198, new_n9195_1, new_n9199);
and_5  g08823(new_n8319, new_n8316, new_n9200);
nor_5  g08824(new_n8325, new_n8320, new_n9201);
nor_5  g08825(new_n9201, new_n9200, new_n9202);
xnor_4 g08826(new_n9202, new_n9199, new_n9203);
nor_5  g08827(new_n8326, new_n8315, new_n9204);
nor_5  g08828(new_n8330, new_n8327, new_n9205);
nor_5  g08829(new_n9205, new_n9204, new_n9206);
xor_4  g08830(new_n9206, new_n9203, new_n9207);
xnor_4 g08831(new_n9207, new_n9185, new_n9208);
xor_4  g08832(new_n9208, new_n9184, new_n9209);
or_5   g08833(new_n8353, new_n8352, new_n9210);
nor_5  g08834(new_n9210, new_n8351, new_n9211);
nor_5  g08835(new_n8355, new_n8332, new_n9212);
nor_5  g08836(new_n9212, new_n9211, new_n9213);
xnor_4 g08837(new_n9213, new_n9209, new_n9214);
xor_4  g08838(new_n9214, new_n9183, new_n9215);
nor_5  g08839(new_n9155, new_n9154, new_n9216);
xor_4  g08840(new_n9216, new_n9153, new_n9217);
nor_5  g08841(new_n9217, new_n9215, new_n9218);
nor_5  g08842(new_n9218, new_n9157, new_n9219);
xnor_4 g08843(new_n9219, new_n9152, new_n9220);
or_5   g08844(new_n9180, new_n9177, new_n9221);
nor_5  g08845(new_n9170, new_n9167, new_n9222);
nor_5  g08846(new_n9175, new_n9171, new_n9223);
or_5   g08847(new_n9223, new_n9222, new_n9224);
and_5  g08848(n11153, n6441, new_n9225);
and_5  g08849(n12947, n5314, new_n9226);
and_5  g08850(n11999, n11222, new_n9227);
xnor_4 g08851(new_n9227, new_n9226, new_n9228);
xnor_4 g08852(new_n9228, new_n9225, new_n9229);
xnor_4 g08853(new_n9229, new_n9224, new_n9230);
and_5  g08854(new_n9169, new_n9168, new_n9231);
and_5  g08855(n11791, n996, new_n9232);
xnor_4 g08856(new_n9232, new_n9231, new_n9233);
and_5  g08857(n5760, n5319, new_n9234);
and_5  g08858(n5767, n1478, new_n9235);
and_5  g08859(n10990, n9457, new_n9236);
xnor_4 g08860(new_n9236, new_n9235, new_n9237);
xor_4  g08861(new_n9237, new_n9234, new_n9238);
xor_4  g08862(new_n9238, new_n9233, new_n9239);
xor_4  g08863(new_n9239, new_n9230, new_n9240);
nor_5  g08864(new_n9165, new_n9162, new_n9241_1);
nand_5 g08865(new_n9164, new_n9163, new_n9242);
or_5   g08866(new_n9176, new_n9166, new_n9243);
xor_4  g08867(new_n9243, new_n9242, new_n9244);
nor_5  g08868(new_n9244, new_n9241_1, new_n9245);
xnor_4 g08869(new_n9245, new_n9240, new_n9246);
xnor_4 g08870(new_n9246, new_n9221, new_n9247);
nor_5  g08871(new_n9181, new_n9159, new_n9248);
nor_5  g08872(new_n9182, new_n9158, new_n9249);
nor_5  g08873(new_n9249, new_n9248, new_n9250);
xnor_4 g08874(new_n9250, new_n9247, new_n9251);
or_5   g08875(new_n9206, new_n9203, new_n9252);
nor_5  g08876(new_n9189_1, new_n9186, new_n9253);
nor_5  g08877(new_n9194, new_n9190, new_n9254);
or_5   g08878(new_n9254, new_n9253, new_n9255);
nand_5 g08879(n12391, n447, new_n9256);
and_5  g08880(n11967, n7891, new_n9257);
and_5  g08881(n12069, n1353, new_n9258);
xnor_4 g08882(new_n9258, new_n9257, new_n9259);
xor_4  g08883(new_n9259, new_n9256, new_n9260);
xnor_4 g08884(new_n9260, new_n9255, new_n9261);
and_5  g08885(new_n9188, new_n9187, new_n9262);
and_5  g08886(n7160, n6254, new_n9263);
xnor_4 g08887(new_n9263, new_n9262, new_n9264);
nand_5 g08888(n7159, n2515, new_n9265);
and_5  g08889(n12777, n4828, new_n9266);
and_5  g08890(n12489, n1199, new_n9267);
xnor_4 g08891(new_n9267, new_n9266, new_n9268);
xnor_4 g08892(new_n9268, new_n9265, new_n9269);
xor_4  g08893(new_n9269, new_n9264, new_n9270);
xor_4  g08894(new_n9270, new_n9261, new_n9271);
nor_5  g08895(new_n9198, new_n9195_1, new_n9272);
nand_5 g08896(new_n9197, new_n9196, new_n9273);
or_5   g08897(new_n9202, new_n9199, new_n9274);
xor_4  g08898(new_n9274, new_n9273, new_n9275);
nor_5  g08899(new_n9275, new_n9272, new_n9276);
xnor_4 g08900(new_n9276, new_n9271, new_n9277);
xnor_4 g08901(new_n9277, new_n9252, new_n9278);
nor_5  g08902(new_n9207, new_n9185, new_n9279);
nor_5  g08903(new_n9208, new_n9184, new_n9280);
or_5   g08904(new_n9280, new_n9279, new_n9281);
xnor_4 g08905(new_n9281, new_n9278, new_n9282);
xnor_4 g08906(new_n9282, new_n9251, new_n9283);
nor_5  g08907(new_n9213, new_n9209, new_n9284);
nor_5  g08908(new_n9214, new_n9183, new_n9285);
nor_5  g08909(new_n9285, new_n9284, new_n9286);
xnor_4 g08910(new_n9286, new_n9283, new_n9287);
xor_4  g08911(new_n9287, new_n9220, new_n9288);
xnor_4 g08912(new_n9288, new_n9096, new_n9289);
xor_4  g08913(new_n9093, new_n9092, new_n9290);
nor_5  g08914(new_n8357, new_n8290, new_n9291);
nor_5  g08915(new_n8361, new_n8358, new_n9292);
or_5   g08916(new_n9292, new_n9291, new_n9293);
nor_5  g08917(new_n9293, new_n9290, new_n9294);
xor_4  g08918(new_n9293, new_n9290, new_n9295);
xor_4  g08919(new_n9217, new_n9215, new_n9296);
and_5  g08920(new_n9296, new_n9295, new_n9297);
nor_5  g08921(new_n9297, new_n9294, new_n9298);
xnor_4 g08922(new_n9298, new_n9289, n5132);
xor_4  g08923(new_n8838, new_n8402, n5191);
and_5  g08924(new_n2911, new_n2614, new_n9301);
nor_5  g08925(new_n2911, new_n2614, new_n9302);
nor_5  g08926(new_n3015, new_n9302, new_n9303);
nor_5  g08927(new_n9303, new_n9301, new_n9304);
nor_5  g08928(new_n3010, new_n2943, new_n9305);
nor_5  g08929(new_n3014, new_n3011, new_n9306);
nor_5  g08930(new_n9306, new_n9305, new_n9307);
nor_5  g08931(new_n2597, new_n2573, new_n9308);
nor_5  g08932(new_n2613, new_n2598, new_n9309);
nor_5  g08933(new_n9309, new_n9308, new_n9310);
nor_5  g08934(new_n2594, new_n2593, new_n9311);
nor_5  g08935(new_n2596, new_n2591, new_n9312);
nor_5  g08936(new_n9312, new_n9311, new_n9313);
and_5  g08937(n11478, n10965, new_n9314);
and_5  g08938(new_n2924, new_n2923, new_n9315);
nor_5  g08939(new_n2930, new_n2925, new_n9316);
nor_5  g08940(new_n9316, new_n9315, new_n9317);
nand_5 g08941(n8433, n4722, new_n9318);
and_5  g08942(n8065, n2464, new_n9319);
and_5  g08943(n7646, n405, new_n9320);
xnor_4 g08944(new_n9320, new_n9319, new_n9321);
xnor_4 g08945(new_n9321, new_n9318, new_n9322);
xnor_4 g08946(new_n9322, new_n9317, new_n9323);
xnor_4 g08947(new_n9323, new_n9314, new_n9324);
xnor_4 g08948(new_n9324, new_n9313, new_n9325);
nor_5  g08949(new_n2983, new_n2980, new_n9326);
nor_5  g08950(new_n2993, new_n2984, new_n9327);
nor_5  g08951(new_n9327, new_n9326, new_n9328);
and_5  g08952(new_n2955, new_n2954, new_n9329);
nor_5  g08953(new_n2961, new_n2956, new_n9330);
nor_5  g08954(new_n9330, new_n9329, new_n9331);
and_5  g08955(new_n2986, new_n2985, new_n9332);
nor_5  g08956(new_n2992, new_n2987, new_n9333);
nor_5  g08957(new_n9333, new_n9332, new_n9334);
xnor_4 g08958(new_n9334, new_n9331, new_n9335);
and_5  g08959(n8384, n6359, new_n9336);
and_5  g08960(n7546, n4805, new_n9337);
xor_4  g08961(new_n9337, new_n9336, new_n9338);
and_5  g08962(n12925, n4938, new_n9339);
and_5  g08963(n11536, n7862, new_n9340);
xnor_4 g08964(new_n9340, new_n9339, new_n9341);
and_5  g08965(new_n2990, new_n2989, new_n9342);
nor_5  g08966(new_n2990, new_n2989, new_n9343);
nor_5  g08967(new_n9343, new_n2988, new_n9344);
nor_5  g08968(new_n9344, new_n9342, new_n9345);
xnor_4 g08969(new_n9345, new_n9341, new_n9346);
xnor_4 g08970(new_n9346, new_n9338, new_n9347);
xnor_4 g08971(new_n9347, new_n9335, new_n9348);
xnor_4 g08972(new_n9348, new_n9328, new_n9349);
nor_5  g08973(new_n2952, new_n2949, new_n9350);
nor_5  g08974(new_n2962, new_n2953, new_n9351);
nor_5  g08975(new_n9351, new_n9350, new_n9352);
nor_5  g08976(new_n2978, new_n2977, new_n9353);
nor_5  g08977(new_n2979, new_n2976, new_n9354);
nor_5  g08978(new_n9354, new_n9353, new_n9355);
and_5  g08979(n9956, n6826, new_n9356);
and_5  g08980(n6797, n4826, new_n9357);
xnor_4 g08981(new_n9357, new_n9356, new_n9358);
and_5  g08982(n7610, n6294, new_n9359);
and_5  g08983(n6611, n6358, new_n9360);
xnor_4 g08984(new_n9360, new_n9359, new_n9361);
xnor_4 g08985(new_n9361, new_n9358, new_n9362);
xnor_4 g08986(new_n9362, new_n9355, new_n9363);
and_5  g08987(n7733, n3146, new_n9364);
nor_5  g08988(new_n2947, new_n2946, new_n9365);
nor_5  g08989(new_n2948, new_n2945, new_n9366);
nor_5  g08990(new_n9366, new_n9365, new_n9367);
xnor_4 g08991(new_n9367, new_n9364, new_n9368);
xnor_4 g08992(new_n9368, new_n9363, new_n9369);
and_5  g08993(n5198, n217, new_n9370);
and_5  g08994(n5283, n503, new_n9371);
xnor_4 g08995(new_n9371, new_n9370, new_n9372);
and_5  g08996(n4970, n137, new_n9373);
and_5  g08997(n11296, n3992, new_n9374);
xnor_4 g08998(new_n9374, new_n9373, new_n9375);
xor_4  g08999(new_n9375, new_n9372, new_n9376);
and_5  g09000(new_n2959, new_n2958, new_n9377);
nor_5  g09001(new_n2959, new_n2958, new_n9378);
nor_5  g09002(new_n9378, new_n2957, new_n9379);
nor_5  g09003(new_n9379, new_n9377, new_n9380);
and_5  g09004(n11311, n10439, new_n9381);
and_5  g09005(n6126, n4203, new_n9382);
xor_4  g09006(new_n9382, new_n9381, new_n9383);
xnor_4 g09007(new_n9383, new_n9380, new_n9384);
xnor_4 g09008(new_n9384, new_n9376, new_n9385);
xnor_4 g09009(new_n9385, new_n9369, new_n9386);
xnor_4 g09010(new_n9386, new_n9352, new_n9387_1);
xnor_4 g09011(new_n9387_1, new_n9349, new_n9388);
nor_5  g09012(new_n2935, new_n2934, new_n9389);
nor_5  g09013(new_n2937, new_n2932, new_n9390);
nor_5  g09014(new_n9390, new_n9389, new_n9391);
nor_5  g09015(new_n2966, new_n2965, new_n9392);
nor_5  g09016(new_n2968, new_n2963, new_n9393);
or_5   g09017(new_n9393, new_n9392, new_n9394);
xnor_4 g09018(new_n9394, new_n9391, new_n9395);
xnor_4 g09019(new_n9395, new_n9388, new_n9396);
xnor_4 g09020(new_n9396, new_n9325, new_n9397);
xnor_4 g09021(new_n9397, new_n9310, new_n9398);
nor_5  g09022(new_n2938, new_n2913, new_n9399);
nor_5  g09023(new_n2942, new_n2939, new_n9400_1);
nor_5  g09024(new_n9400_1, new_n9399, new_n9401);
nor_5  g09025(new_n2921, new_n2918, new_n9402);
nor_5  g09026(new_n2931, new_n2922, new_n9403);
nor_5  g09027(new_n9403, new_n9402, new_n9404);
nand_5 g09028(n4086, n1471, new_n9405);
nand_5 g09029(n10391, n9400, new_n9406);
nor_5  g09030(new_n2917, new_n2914, new_n9407);
or_5   g09031(new_n9407, new_n2915, new_n9408);
nor_5  g09032(new_n9408, new_n9406, new_n9409);
or_5   g09033(new_n9406, new_n2657, new_n9410);
and_5  g09034(new_n9410, new_n9408, new_n9411);
nor_5  g09035(new_n9411, new_n9409, new_n9412);
nand_5 g09036(n11757, n2577, new_n9413);
and_5  g09037(n9637, n3172, new_n9414);
and_5  g09038(n5240, n3842, new_n9415);
xnor_4 g09039(new_n9415, new_n9414, new_n9416);
xnor_4 g09040(new_n9416, new_n9413, new_n9417);
and_5  g09041(new_n2578, new_n2577_1, new_n9418);
nor_5  g09042(new_n2578, new_n2577_1, new_n9419);
nor_5  g09043(new_n9419, new_n2576, new_n9420);
nor_5  g09044(new_n9420, new_n9418, new_n9421);
xnor_4 g09045(new_n9421, new_n9417, new_n9422);
xnor_4 g09046(new_n9422, new_n9412, new_n9423);
xnor_4 g09047(new_n9423, new_n9405, new_n9424);
and_5  g09048(n7236, n1357, new_n9425);
and_5  g09049(new_n2583, new_n2582, new_n9426);
nor_5  g09050(new_n2589, new_n2584, new_n9427);
nor_5  g09051(new_n9427, new_n9426, new_n9428);
xnor_4 g09052(new_n9428, new_n9425, new_n9429);
xnor_4 g09053(new_n9429, new_n9424, new_n9430);
xnor_4 g09054(new_n9430, new_n9404, new_n9431);
and_5  g09055(n1835, n1333, new_n9432);
and_5  g09056(n11917, n11821, new_n9433);
xor_4  g09057(new_n9433, new_n9432, new_n9434);
and_5  g09058(n12753, n3602, new_n9435);
and_5  g09059(n8595, n4187, new_n9436);
xnor_4 g09060(new_n9436, new_n9435, new_n9437);
and_5  g09061(n6877, n4190, new_n9438);
and_5  g09062(n10174, n3719, new_n9439);
xnor_4 g09063(new_n9439, new_n9438, new_n9440);
xnor_4 g09064(new_n9440, new_n9437, new_n9441);
xnor_4 g09065(new_n9441, new_n9434, new_n9442);
nor_5  g09066(new_n2928, new_n2927, new_n9443);
nor_5  g09067(new_n2929, new_n2926, new_n9444);
nor_5  g09068(new_n9444, new_n9443, new_n9445);
nand_5 g09069(n9080, n4921, new_n9446);
xnor_4 g09070(new_n9446, new_n9445, new_n9447);
xnor_4 g09071(new_n9447, new_n9442, new_n9448);
nor_5  g09072(new_n2580, new_n2575, new_n9449);
nor_5  g09073(new_n2590, new_n2581_1, new_n9450);
nor_5  g09074(new_n9450, new_n9449, new_n9451);
xnor_4 g09075(new_n9451, new_n9448, new_n9452);
xnor_4 g09076(new_n9452, new_n9431, new_n9453);
nor_5  g09077(new_n2997, new_n2996, new_n9454);
nor_5  g09078(new_n2999, new_n2994, new_n9455);
nor_5  g09079(new_n9455, new_n9454, new_n9456);
xnor_4 g09080(new_n9456, new_n9453, new_n9457_1);
xnor_4 g09081(new_n9457_1, new_n9401, new_n9458);
nor_5  g09082(new_n2969, new_n2944, new_n9459);
nor_5  g09083(new_n2973, new_n2970, new_n9460);
nor_5  g09084(new_n9460, new_n9459, new_n9461);
xnor_4 g09085(new_n9461, new_n9458, new_n9462);
xnor_4 g09086(new_n9462, new_n9398, new_n9463);
and_5  g09087(new_n3005, new_n2974, new_n9464);
nor_5  g09088(new_n3009, new_n3006, new_n9465);
nor_5  g09089(new_n9465, new_n9464, new_n9466);
nor_5  g09090(new_n3000, new_n2975, new_n9467);
nor_5  g09091(new_n3004, new_n3001, new_n9468);
nor_5  g09092(new_n9468, new_n9467, new_n9469);
nor_5  g09093(new_n2587, new_n2586, new_n9470);
nor_5  g09094(new_n2588, new_n2585_1, new_n9471);
nor_5  g09095(new_n9471, new_n9470, new_n9472);
xnor_4 g09096(new_n9472, new_n9469, new_n9473);
xnor_4 g09097(new_n9473, new_n9466, new_n9474);
xnor_4 g09098(new_n9474, new_n9463, new_n9475);
xnor_4 g09099(new_n9475, new_n9307, new_n9476);
xnor_4 g09100(new_n9476, new_n9304, n5257);
xnor_4 g09101(new_n8845, new_n8837, n5411);
xnor_4 g09102(new_n2901, new_n2893, n5435);
xnor_4 g09103(new_n4830, new_n7756, n5641);
xnor_4 g09104(new_n6777, new_n6768, n5670);
xnor_4 g09105(new_n3912, new_n3887, n5693);
xnor_4 g09106(new_n1137, new_n1127, n5934);
xnor_4 g09107(new_n8848, new_n8847, n6089);
or_5   g09108(new_n6179, new_n6176, new_n9485);
nor_5  g09109(new_n6163, new_n6160, new_n9486);
nor_5  g09110(new_n6167, new_n6164, new_n9487);
or_5   g09111(new_n9487, new_n9486, new_n9488);
nand_5 g09112(n2564, n2253, new_n9489);
and_5  g09113(n9195, n4189, new_n9490);
and_5  g09114(n6687, n3865, new_n9491);
xnor_4 g09115(new_n9491, new_n9490, new_n9492);
xor_4  g09116(new_n9492, new_n9489, new_n9493);
xnor_4 g09117(new_n9493, new_n9488, new_n9494);
and_5  g09118(new_n6162, new_n6161, new_n9495);
and_5  g09119(n6770, n4634, new_n9496);
xnor_4 g09120(new_n9496, new_n9495, new_n9497);
and_5  g09121(n3627, n2879, new_n9498);
and_5  g09122(n10223, n9920, new_n9499);
and_5  g09123(n7265, n4516, new_n9500);
xnor_4 g09124(new_n9500, new_n9499, new_n9501);
xnor_4 g09125(new_n9501, new_n9498, new_n9502);
xnor_4 g09126(new_n9502, new_n9497, new_n9503);
xor_4  g09127(new_n9503, new_n9494, new_n9504);
nor_5  g09128(new_n6171, new_n6168, new_n9505);
nand_5 g09129(new_n6170, new_n6169, new_n9506);
or_5   g09130(new_n6175, new_n6172, new_n9507);
xor_4  g09131(new_n9507, new_n9506, new_n9508);
nor_5  g09132(new_n9508, new_n9505, new_n9509);
xnor_4 g09133(new_n9509, new_n9504, new_n9510);
xnor_4 g09134(new_n9510, new_n9485, new_n9511);
nor_5  g09135(new_n6180, new_n6159, new_n9512);
nor_5  g09136(new_n6181, new_n6158, new_n9513);
or_5   g09137(new_n9513, new_n9512, new_n9514);
xor_4  g09138(new_n9514, new_n9511, new_n9515);
nor_5  g09139(new_n6214, new_n6211, new_n9516);
nor_5  g09140(new_n6273_1, new_n6215, new_n9517);
nor_5  g09141(new_n9517, new_n9516, new_n9518);
nor_5  g09142(new_n6209, new_n6188, new_n9519);
nor_5  g09143(new_n6210, new_n6187, new_n9520);
nor_5  g09144(new_n9520, new_n9519, new_n9521);
or_5   g09145(new_n6208, new_n6205, new_n9522);
nor_5  g09146(new_n6192_1, new_n6189, new_n9523);
nor_5  g09147(new_n6196, new_n6193, new_n9524);
or_5   g09148(new_n9524, new_n9523, new_n9525);
nand_5 g09149(n12221, n10928, new_n9526);
and_5  g09150(n12145, n6986, new_n9527);
and_5  g09151(n10217, n8336, new_n9528);
xnor_4 g09152(new_n9528, new_n9527, new_n9529);
xor_4  g09153(new_n9529, new_n9526, new_n9530);
xnor_4 g09154(new_n9530, new_n9525, new_n9531);
and_5  g09155(new_n6191, new_n6190, new_n9532);
and_5  g09156(n2522, n2226, new_n9533);
xnor_4 g09157(new_n9533, new_n9532, new_n9534);
and_5  g09158(n10678, n2024, new_n9535);
and_5  g09159(n9189, n1094, new_n9536);
and_5  g09160(n7946, n7320, new_n9537);
xnor_4 g09161(new_n9537, new_n9536, new_n9538);
xnor_4 g09162(new_n9538, new_n9535, new_n9539);
xnor_4 g09163(new_n9539, new_n9534, new_n9540);
xor_4  g09164(new_n9540, new_n9531, new_n9541);
nor_5  g09165(new_n6200, new_n6197, new_n9542);
nand_5 g09166(new_n6199, new_n6198, new_n9543);
or_5   g09167(new_n6204, new_n6201, new_n9544);
xor_4  g09168(new_n9544, new_n9543, new_n9545);
nor_5  g09169(new_n9545, new_n9542, new_n9546);
xnor_4 g09170(new_n9546, new_n9541, new_n9547);
xnor_4 g09171(new_n9547, new_n9522, new_n9548);
xor_4  g09172(new_n9548, new_n9521, new_n9549);
or_5   g09173(new_n6239, new_n6236, new_n9550);
and_5  g09174(new_n6226, new_n6225, new_n9551);
and_5  g09175(n7160, n521, new_n9552);
xnor_4 g09176(new_n9552, new_n9551, new_n9553);
nand_5 g09177(n2515, n2498, new_n9554);
and_5  g09178(n2558, n1199, new_n9555);
and_5  g09179(n5579, n4828, new_n9556);
xnor_4 g09180(new_n9556, new_n9555, new_n9557);
xnor_4 g09181(new_n9557, new_n9554, new_n9558);
xnor_4 g09182(new_n9558, new_n9553, new_n9559);
nor_5  g09183(new_n6227, new_n6224, new_n9560);
or_5   g09184(new_n9560, new_n6223, new_n9561);
and_5  g09185(n12391, n5798, new_n9562);
and_5  g09186(n7891, n6016, new_n9563);
and_5  g09187(n12069, n2347, new_n9564);
xnor_4 g09188(new_n9564, new_n9563, new_n9565);
xnor_4 g09189(new_n9565, new_n9562, new_n9566);
xor_4  g09190(new_n9566, new_n9561, new_n9567);
xor_4  g09191(new_n9567, new_n9559, new_n9568);
nor_5  g09192(new_n6231, new_n6228, new_n9569);
nand_5 g09193(new_n6230, new_n6229, new_n9570);
or_5   g09194(new_n6235, new_n6232, new_n9571_1);
xor_4  g09195(new_n9571_1, new_n9570, new_n9572);
nor_5  g09196(new_n9572, new_n9569, new_n9573);
xnor_4 g09197(new_n9573, new_n9568, new_n9574);
xnor_4 g09198(new_n9574, new_n9550, new_n9575);
nor_5  g09199(new_n6240, new_n6217, new_n9576);
nor_5  g09200(new_n6241, new_n6216, new_n9577);
nor_5  g09201(new_n9577, new_n9576, new_n9578_1);
xor_4  g09202(new_n9578_1, new_n9575, new_n9579);
nor_5  g09203(new_n6265, new_n6262, new_n9580);
nor_5  g09204(new_n6248, new_n6245, new_n9581);
nor_5  g09205(new_n6253, new_n6249, new_n9582);
or_5   g09206(new_n9582, new_n9581, new_n9583_1);
and_5  g09207(n11153, n5153, new_n9584);
and_5  g09208(n7270, n5314, new_n9585);
and_5  g09209(n11222, n2507, new_n9586);
xnor_4 g09210(new_n9586, new_n9585, new_n9587);
xnor_4 g09211(new_n9587, new_n9584, new_n9588);
xnor_4 g09212(new_n9588, new_n9583_1, new_n9589);
and_5  g09213(new_n6247, new_n6246, new_n9590);
and_5  g09214(n996, n806, new_n9591);
xnor_4 g09215(new_n9591, new_n9590, new_n9592);
and_5  g09216(n9111, n5319, new_n9593);
and_5  g09217(n5767, n3342, new_n9594);
and_5  g09218(n9763, n9457, new_n9595);
xnor_4 g09219(new_n9595, new_n9594, new_n9596);
xor_4  g09220(new_n9596, new_n9593, new_n9597);
xor_4  g09221(new_n9597, new_n9592, new_n9598);
xor_4  g09222(new_n9598, new_n9589, new_n9599);
nor_5  g09223(new_n6257, new_n6254_1, new_n9600);
nand_5 g09224(new_n6256, new_n6255, new_n9601);
or_5   g09225(new_n6261, new_n6258, new_n9602);
xor_4  g09226(new_n9602, new_n9601, new_n9603);
nor_5  g09227(new_n9603, new_n9600, new_n9604);
xor_4  g09228(new_n9604, new_n9599, new_n9605);
xnor_4 g09229(new_n9605, new_n9580, new_n9606);
nor_5  g09230(new_n6266, new_n6244, new_n9607);
nor_5  g09231(new_n6267, new_n6243, new_n9608);
or_5   g09232(new_n9608, new_n9607, new_n9609);
xor_4  g09233(new_n9609, new_n9606, new_n9610);
xnor_4 g09234(new_n9610, new_n9579, new_n9611);
nor_5  g09235(new_n6268, new_n6242, new_n9612);
nor_5  g09236(new_n6272, new_n6269, new_n9613);
or_5   g09237(new_n9613, new_n9612, new_n9614);
xnor_4 g09238(new_n9614, new_n9611, new_n9615);
xnor_4 g09239(new_n9615, new_n9549, new_n9616);
xor_4  g09240(new_n9616, new_n9518, new_n9617);
nor_5  g09241(new_n9617, new_n9515, new_n9618);
and_5  g09242(new_n6185, new_n6182, new_n9619);
nor_5  g09243(new_n6274, new_n6186, new_n9620);
nor_5  g09244(new_n9620, new_n9619, new_n9621);
xor_4  g09245(new_n9617, new_n9515, new_n9622);
and_5  g09246(new_n9622, new_n9621, new_n9623);
nor_5  g09247(new_n9623, new_n9618, new_n9624);
nor_5  g09248(new_n9615, new_n9549, new_n9625);
or_5   g09249(new_n9517, new_n9516, new_n9626);
nor_5  g09250(new_n9616, new_n9626, new_n9627);
nor_5  g09251(new_n9627, new_n9625, new_n9628);
nor_5  g09252(new_n9610, new_n9579, new_n9629);
nor_5  g09253(new_n9614, new_n9611, new_n9630);
nor_5  g09254(new_n9630, new_n9629, new_n9631);
nor_5  g09255(new_n9544, new_n9543, new_n9632);
nor_5  g09256(new_n9546, new_n9541, new_n9633);
nor_5  g09257(new_n9633, new_n9632, new_n9634);
nor_5  g09258(new_n9493, new_n9488, new_n9635);
nor_5  g09259(new_n9503, new_n9494, new_n9636);
nor_5  g09260(new_n9636, new_n9635, new_n9637_1);
nand_5 g09261(n2522, n1094, new_n9638);
nor_5  g09262(new_n9586, new_n9585, new_n9639);
nor_5  g09263(new_n9587, new_n9584, new_n9640_1);
nor_5  g09264(new_n9640_1, new_n9639, new_n9641);
xnor_4 g09265(new_n9641, new_n9638, new_n9642);
xnor_4 g09266(new_n9642, new_n9637_1, new_n9643);
xnor_4 g09267(new_n9643, new_n9634, new_n9644);
nor_5  g09268(new_n9530, new_n9525, new_n9645);
nor_5  g09269(new_n9540, new_n9531, new_n9646);
nor_5  g09270(new_n9646, new_n9645, new_n9647);
nand_5 g09271(n10678, n9189, new_n9648);
xnor_4 g09272(new_n9648, new_n9647, new_n9649);
nor_5  g09273(new_n9537, new_n9536, new_n9650);
nor_5  g09274(new_n9538, new_n9535, new_n9651);
nor_5  g09275(new_n9651, new_n9650, new_n9652);
and_5  g09276(n7946, n7523, new_n9653);
and_5  g09277(n10223, n3627, new_n9654);
and_5  g09278(n3865, n2564, new_n9655);
xnor_4 g09279(new_n9655, new_n9654, new_n9656);
xnor_4 g09280(new_n9656, new_n9653, new_n9657);
xnor_4 g09281(new_n9657, new_n9652, new_n9658);
and_5  g09282(n12221, n6986, new_n9659);
and_5  g09283(n8336, n7823, new_n9660);
xnor_4 g09284(new_n9660, new_n9659, new_n9661);
xnor_4 g09285(new_n9661, new_n9658, new_n9662);
nor_5  g09286(new_n9500, new_n9499, new_n9663);
nor_5  g09287(new_n9501, new_n9498, new_n9664);
or_5   g09288(new_n9664, new_n9663, new_n9665);
nor_5  g09289(new_n9533, new_n9532, new_n9666);
nor_5  g09290(new_n9539, new_n9534, new_n9667);
nor_5  g09291(new_n9667, new_n9666, new_n9668);
xnor_4 g09292(new_n9668, new_n9665, new_n9669);
nor_5  g09293(new_n9564, new_n9563, new_n9670);
nor_5  g09294(new_n9565, new_n9562, new_n9671);
or_5   g09295(new_n9671, new_n9670, new_n9672);
and_5  g09296(n6687, n2512, new_n9673);
and_5  g09297(new_n9556, new_n9555, new_n9674);
nor_5  g09298(new_n9556, new_n9555, new_n9675);
nor_5  g09299(new_n9675, new_n9554, new_n9676);
nor_5  g09300(new_n9676, new_n9674, new_n9677);
xnor_4 g09301(new_n9677, new_n9673, new_n9678);
xnor_4 g09302(new_n9678, new_n9672, new_n9679);
xnor_4 g09303(new_n9679, new_n9669, new_n9680);
xnor_4 g09304(new_n9680, new_n9662, new_n9681);
and_5  g09305(n11153, n2507, new_n9682);
and_5  g09306(n7270, n996, new_n9683);
xnor_4 g09307(new_n9683, new_n9682, new_n9684);
and_5  g09308(n7160, n6016, new_n9685);
and_5  g09309(n5767, n806, new_n9686);
xnor_4 g09310(new_n9686, new_n9685, new_n9687);
xnor_4 g09311(new_n9687, new_n9684, new_n9688);
and_5  g09312(n4828, n521, new_n9689);
and_5  g09313(n5579, n2515, new_n9690);
xnor_4 g09314(new_n9690, new_n9689, new_n9691);
and_5  g09315(n12069, n1576, new_n9692);
and_5  g09316(n5314, n5153, new_n9693);
xnor_4 g09317(new_n9693, new_n9692, new_n9694);
xnor_4 g09318(new_n9694, new_n9691, new_n9695);
xor_4  g09319(new_n9695, new_n9688, new_n9696);
and_5  g09320(new_n9491, new_n9490, new_n9697);
nor_5  g09321(new_n9491, new_n9490, new_n9698);
nor_5  g09322(new_n9698, new_n9489, new_n9699);
nor_5  g09323(new_n9699, new_n9697, new_n9700);
nand_5 g09324(n4516, n2879, new_n9701);
and_5  g09325(n4189, n2253, new_n9702);
and_5  g09326(n9920, n4634, new_n9703);
xnor_4 g09327(new_n9703, new_n9702, new_n9704);
xnor_4 g09328(new_n9704, new_n9701, new_n9705);
xnor_4 g09329(new_n9705, new_n9700, new_n9706_1);
xnor_4 g09330(new_n9706_1, new_n9696, new_n9707);
nor_5  g09331(new_n9496, new_n9495, new_n9708);
nor_5  g09332(new_n9502, new_n9497, new_n9709);
nor_5  g09333(new_n9709, new_n9708, new_n9710);
and_5  g09334(new_n9591, new_n9590, new_n9711);
nor_5  g09335(new_n9597, new_n9592, new_n9712);
nor_5  g09336(new_n9712, new_n9711, new_n9713);
xnor_4 g09337(new_n9713, new_n9710, new_n9714);
xnor_4 g09338(new_n9714, new_n9707, new_n9715);
xnor_4 g09339(new_n9715, new_n9681, new_n9716);
xnor_4 g09340(new_n9716, new_n9649, new_n9717);
xnor_4 g09341(new_n9717, new_n9644, new_n9718);
nor_5  g09342(new_n9602, new_n9601, new_n9719);
nor_5  g09343(new_n9604, new_n9599, new_n9720);
nor_5  g09344(new_n9720, new_n9719, new_n9721);
and_5  g09345(n12145, n2226, new_n9722);
and_5  g09346(new_n9528, new_n9527, new_n9723);
nor_5  g09347(new_n9528, new_n9527, new_n9724);
nor_5  g09348(new_n9724, new_n9526, new_n9725_1);
nor_5  g09349(new_n9725_1, new_n9723, new_n9726);
and_5  g09350(n9195, n6770, new_n9727);
and_5  g09351(n11222, n6431, new_n9728);
xnor_4 g09352(new_n9728, new_n9727, new_n9729);
and_5  g09353(n10928, n10217, new_n9730);
and_5  g09354(n7320, n2024, new_n9731);
xnor_4 g09355(new_n9731, new_n9730, new_n9732);
xnor_4 g09356(new_n9732, new_n9729, new_n9733);
nand_5 g09357(n5319, n3342, new_n9734);
and_5  g09358(n9457, n9111, new_n9735);
and_5  g09359(n9763, n4817, new_n9736);
xnor_4 g09360(new_n9736, new_n9735, new_n9737);
xnor_4 g09361(new_n9737, new_n9734, new_n9738);
xnor_4 g09362(new_n9738, new_n9733, new_n9739);
xnor_4 g09363(new_n9739, new_n9726, new_n9740);
xnor_4 g09364(new_n9740, new_n9722, new_n9741);
xnor_4 g09365(new_n9741, new_n9721, new_n9742);
xnor_4 g09366(new_n9742, new_n9718, new_n9743);
nor_5  g09367(new_n9547, new_n9522, new_n9744);
nor_5  g09368(new_n9548, new_n9521, new_n9745);
nor_5  g09369(new_n9745, new_n9744, new_n9746);
nor_5  g09370(new_n9571_1, new_n9570, new_n9747);
nor_5  g09371(new_n9573, new_n9568, new_n9748);
nor_5  g09372(new_n9748, new_n9747, new_n9749);
nor_5  g09373(new_n9507, new_n9506, new_n9750);
nor_5  g09374(new_n9509, new_n9504, new_n9751);
nor_5  g09375(new_n9751, new_n9750, new_n9752);
nor_5  g09376(new_n9588, new_n9583_1, new_n9753);
nor_5  g09377(new_n9598, new_n9589, new_n9754);
nor_5  g09378(new_n9754, new_n9753, new_n9755);
and_5  g09379(new_n9552, new_n9551, new_n9756_1);
nor_5  g09380(new_n9558, new_n9553, new_n9757);
nor_5  g09381(new_n9757, new_n9756_1, new_n9758);
and_5  g09382(n7891, n5798, new_n9759);
xnor_4 g09383(new_n9759, new_n9758, new_n9760);
and_5  g09384(n12391, n2347, new_n9761);
and_5  g09385(n7265, n2087, new_n9762);
xnor_4 g09386(new_n9762, new_n9761, new_n9763_1);
xnor_4 g09387(new_n9763_1, new_n9760, new_n9764);
xnor_4 g09388(new_n9764, new_n9755, new_n9765);
and_5  g09389(n2498, n1199, new_n9766);
and_5  g09390(n6578, n2558, new_n9767_1);
xnor_4 g09391(new_n9767_1, new_n9766, new_n9768);
xnor_4 g09392(new_n9768, new_n9765, new_n9769);
xnor_4 g09393(new_n9769, new_n9752, new_n9770);
xnor_4 g09394(new_n9770, new_n9749, new_n9771);
xnor_4 g09395(new_n9771, new_n9746, new_n9772);
xnor_4 g09396(new_n9772, new_n9743, new_n9773);
and_5  g09397(new_n9605, new_n9580, new_n9774);
nor_5  g09398(new_n9609, new_n9606, new_n9775);
nor_5  g09399(new_n9775, new_n9774, new_n9776);
nor_5  g09400(new_n9595, new_n9594, new_n9777);
nor_5  g09401(new_n9596, new_n9593, new_n9778);
nor_5  g09402(new_n9778, new_n9777, new_n9779);
nor_5  g09403(new_n9566, new_n9561, new_n9780);
and_5  g09404(new_n9567, new_n9559, new_n9781);
nor_5  g09405(new_n9781, new_n9780, new_n9782);
xnor_4 g09406(new_n9782, new_n9779, new_n9783);
xnor_4 g09407(new_n9783, new_n9776, new_n9784);
xnor_4 g09408(new_n9784, new_n9773, new_n9785);
xnor_4 g09409(new_n9785, new_n9631, new_n9786);
nor_5  g09410(new_n9510, new_n9485, new_n9787);
nor_5  g09411(new_n9514, new_n9511, new_n9788);
nor_5  g09412(new_n9788, new_n9787, new_n9789);
nor_5  g09413(new_n9574, new_n9550, new_n9790);
nor_5  g09414(new_n9578_1, new_n9575, new_n9791);
nor_5  g09415(new_n9791, new_n9790, new_n9792);
xnor_4 g09416(new_n9792, new_n9789, new_n9793);
xnor_4 g09417(new_n9793, new_n9786, new_n9794);
xnor_4 g09418(new_n9794, new_n9628, new_n9795);
xnor_4 g09419(new_n9795, new_n9624, n6192);
xor_4  g09420(new_n769, new_n745, n6273);
xnor_4 g09421(new_n5982, new_n5981, n6445);
xnor_4 g09422(new_n7439, new_n7438, n6645);
xnor_4 g09423(new_n6307, new_n6306, n6689);
xor_4  g09424(new_n1128, new_n1058, n6742);
xor_4  g09425(new_n1677, new_n1643, n6809);
xnor_4 g09426(new_n5351, new_n5347, n6822);
xnor_4 g09427(new_n8843, new_n8842, n6860);
xnor_4 g09428(new_n7434, new_n7427, n7193);
xor_4  g09429(new_n5985, new_n5984, n7568);
xnor_4 g09430(new_n1135, new_n1134, n7676);
nor_5  g09431(new_n774, new_n477, new_n9808);
nor_5  g09432(new_n881, new_n775, new_n9809);
nor_5  g09433(new_n9809, new_n9808, new_n9810);
nor_5  g09434(new_n876, new_n806_1, new_n9811);
nor_5  g09435(new_n880, new_n877, new_n9812);
nor_5  g09436(new_n9812, new_n9811, new_n9813);
nor_5  g09437(new_n870, new_n838, new_n9814);
nor_5  g09438(new_n875, new_n871, new_n9815);
nor_5  g09439(new_n9815, new_n9814, new_n9816);
nand_5 g09440(n9241, n1209, new_n9817);
and_5  g09441(new_n864, new_n839, new_n9818);
nor_5  g09442(new_n869, new_n865, new_n9819);
nor_5  g09443(new_n9819, new_n9818, new_n9820_1);
nor_5  g09444(new_n861, new_n860, new_n9821);
nor_5  g09445(new_n863, new_n858, new_n9822);
nor_5  g09446(new_n9822, new_n9821, new_n9823);
nor_5  g09447(new_n443, new_n438, new_n9824);
nor_5  g09448(new_n453, new_n444, new_n9825);
nor_5  g09449(new_n9825, new_n9824, new_n9826);
and_5  g09450(new_n446, new_n445, new_n9827);
nor_5  g09451(new_n452, new_n447_1, new_n9828);
nor_5  g09452(new_n9828, new_n9827, new_n9829);
and_5  g09453(n12705, n2508, new_n9830);
and_5  g09454(new_n441, new_n440, new_n9831);
nor_5  g09455(new_n441, new_n440, new_n9832);
nor_5  g09456(new_n9832, new_n439, new_n9833);
nor_5  g09457(new_n9833, new_n9831, new_n9834);
xnor_4 g09458(new_n9834, new_n9830, new_n9835);
and_5  g09459(n3986, n1980, new_n9836);
and_5  g09460(n10848, n5857, new_n9837);
xnor_4 g09461(new_n9837, new_n9836, new_n9838);
and_5  g09462(n11257, n2509, new_n9839);
and_5  g09463(n4005, n1097, new_n9840);
xnor_4 g09464(new_n9840, new_n9839, new_n9841);
xor_4  g09465(new_n9841, new_n9838, new_n9842);
xnor_4 g09466(new_n9842, new_n9835, new_n9843);
xnor_4 g09467(new_n9843, new_n9829, new_n9844);
and_5  g09468(n8028, n45, new_n9845);
nor_5  g09469(new_n782, new_n781, new_n9846);
nor_5  g09470(new_n783_1, new_n780, new_n9847);
nor_5  g09471(new_n9847, new_n9846, new_n9848);
xnor_4 g09472(new_n9848, new_n9845, new_n9849);
and_5  g09473(new_n791, new_n790, new_n9850);
nor_5  g09474(new_n791, new_n790, new_n9851);
nor_5  g09475(new_n9851, new_n789, new_n9852);
nor_5  g09476(new_n9852, new_n9850, new_n9853);
xnor_4 g09477(new_n9853, new_n9849, new_n9854);
nand_5 g09478(n4312, n2585, new_n9855);
nor_5  g09479(new_n450, new_n449, new_n9856);
nor_5  g09480(new_n451, new_n448, new_n9857);
nor_5  g09481(new_n9857, new_n9856, new_n9858);
nand_5 g09482(n10644, n7354, new_n9859);
and_5  g09483(n12706, n5964, new_n9860);
and_5  g09484(n12720, n12025, new_n9861);
xnor_4 g09485(new_n9861, new_n9860, new_n9862);
xnor_4 g09486(new_n9862, new_n9859, new_n9863);
xnor_4 g09487(new_n9863, new_n9858, new_n9864);
xnor_4 g09488(new_n9864, new_n9855, new_n9865);
xnor_4 g09489(new_n9865, new_n9854, new_n9866);
xnor_4 g09490(new_n9866, new_n9844, new_n9867);
xnor_4 g09491(new_n9867, new_n9826, new_n9868);
and_5  g09492(n7436, n4141, new_n9869);
and_5  g09493(new_n787, new_n786, new_n9870);
nor_5  g09494(new_n793, new_n788, new_n9871);
nor_5  g09495(new_n9871, new_n9870, new_n9872);
xnor_4 g09496(new_n9872, new_n9869, new_n9873);
xnor_4 g09497(new_n9873, new_n9868, new_n9874);
xnor_4 g09498(new_n9874, new_n9823, new_n9875);
xnor_4 g09499(new_n9875, new_n9820_1, new_n9876);
xnor_4 g09500(new_n9876, new_n9817, new_n9877);
xnor_4 g09501(new_n9877, new_n9816, new_n9878);
and_5  g09502(n10547, n6038, new_n9879);
nor_5  g09503(new_n813, new_n812, new_n9880);
nor_5  g09504(new_n814, new_n811, new_n9881);
nor_5  g09505(new_n9881, new_n9880, new_n9882);
xnor_4 g09506(new_n9882, new_n9879, new_n9883);
nor_5  g09507(new_n822, new_n821, new_n9884);
nor_5  g09508(new_n823, new_n820, new_n9885);
nor_5  g09509(new_n9885, new_n9884, new_n9886);
and_5  g09510(n12044, n8476, new_n9887);
and_5  g09511(n11892, n5814, new_n9888);
and_5  g09512(n3616, n1512, new_n9889);
xnor_4 g09513(new_n9889, new_n9888, new_n9890);
xnor_4 g09514(new_n9890, new_n9887, new_n9891);
xnor_4 g09515(new_n9891, new_n9886, new_n9892);
xnor_4 g09516(new_n9892, new_n9883, new_n9893);
nand_5 g09517(n12299, n4928, new_n9894);
nor_5  g09518(new_n854, new_n853, new_n9895);
nor_5  g09519(new_n855, new_n852, new_n9896);
nor_5  g09520(new_n9896, new_n9895, new_n9897);
xnor_4 g09521(new_n9897, new_n9894, new_n9898);
and_5  g09522(n5069, n2530, new_n9899);
and_5  g09523(n10545, n2802, new_n9900);
xnor_4 g09524(new_n9900, new_n9899, new_n9901);
xnor_4 g09525(new_n9901, new_n9898, new_n9902);
xnor_4 g09526(new_n9902, new_n9893, new_n9903);
nor_5  g09527(new_n815, new_n810, new_n9904);
nor_5  g09528(new_n825, new_n816, new_n9905);
nor_5  g09529(new_n9905, new_n9904, new_n9906);
and_5  g09530(new_n850, new_n849, new_n9907);
nor_5  g09531(new_n856, new_n851, new_n9908);
or_5   g09532(new_n9908, new_n9907, new_n9909);
and_5  g09533(new_n818, new_n817, new_n9910);
nor_5  g09534(new_n824, new_n819, new_n9911);
nor_5  g09535(new_n9911, new_n9910, new_n9912);
and_5  g09536(n7690, n533, new_n9913);
xnor_4 g09537(new_n9913, new_n9912, new_n9914);
xnor_4 g09538(new_n9914, new_n9909, new_n9915);
xnor_4 g09539(new_n9915, new_n9906, new_n9916);
xnor_4 g09540(new_n9916, new_n9903, new_n9917);
and_5  g09541(n12704, n2393, new_n9918);
and_5  g09542(n7294, n5860, new_n9919);
xnor_4 g09543(new_n9919, new_n9918, new_n9920_1);
and_5  g09544(n12648, n6806, new_n9921);
and_5  g09545(n4499, n1564, new_n9922);
xnor_4 g09546(new_n9922, new_n9921, new_n9923);
xnor_4 g09547(new_n9923, new_n9920_1, new_n9924);
nor_5  g09548(new_n845, new_n844_1, new_n9925);
nor_5  g09549(new_n846, new_n843, new_n9926);
nor_5  g09550(new_n9926, new_n9925, new_n9927);
and_5  g09551(n5694, n5331, new_n9928);
and_5  g09552(n7388, n4903, new_n9929);
xnor_4 g09553(new_n9929, new_n9928, new_n9930);
xnor_4 g09554(new_n9930, new_n9927, new_n9931);
xnor_4 g09555(new_n9931, new_n9924, new_n9932);
and_5  g09556(n8276, n5105, new_n9933);
and_5  g09557(n5305, n615, new_n9934);
xor_4  g09558(new_n9934, new_n9933, new_n9935);
xnor_4 g09559(new_n9935, new_n9932, new_n9936);
xnor_4 g09560(new_n9936, new_n9917, new_n9937);
nor_5  g09561(new_n798, new_n797, new_n9938_1);
nor_5  g09562(new_n800, new_n795, new_n9939);
nor_5  g09563(new_n9939, new_n9938_1, new_n9940);
nor_5  g09564(new_n829, new_n828, new_n9941);
nor_5  g09565(new_n831, new_n826, new_n9942);
nor_5  g09566(new_n9942, new_n9941, new_n9943);
xnor_4 g09567(new_n9943, new_n9940, new_n9944);
xnor_4 g09568(new_n9944, new_n9937, new_n9945);
and_5  g09569(n8759, n783, new_n9946);
and_5  g09570(n10510, n7500, new_n9947);
xor_4  g09571(new_n9947, new_n9946, new_n9948);
nor_5  g09572(new_n457, new_n456, new_n9949);
nor_5  g09573(new_n459, new_n454, new_n9950);
nor_5  g09574(new_n9950, new_n9949, new_n9951);
nor_5  g09575(new_n847, new_n842, new_n9952);
nor_5  g09576(new_n857, new_n848, new_n9953);
or_5   g09577(new_n9953, new_n9952, new_n9954);
xnor_4 g09578(new_n9954, new_n9951, new_n9955);
xnor_4 g09579(new_n9955, new_n9948, new_n9956_1);
xnor_4 g09580(new_n9956_1, new_n9945, new_n9957);
nor_5  g09581(new_n832, new_n807, new_n9958);
nor_5  g09582(new_n837_1, new_n833, new_n9959);
nor_5  g09583(new_n9959, new_n9958, new_n9960);
and_5  g09584(n7965, n1906, new_n9961);
xnor_4 g09585(new_n9961, new_n9960, new_n9962);
xnor_4 g09586(new_n9962, new_n9957, new_n9963);
and_5  g09587(new_n460, new_n435, new_n9964);
nor_5  g09588(new_n476, new_n461, new_n9965);
nor_5  g09589(new_n9965, new_n9964, new_n9966);
nor_5  g09590(new_n801, new_n776, new_n9967);
nor_5  g09591(new_n805, new_n802, new_n9968);
nor_5  g09592(new_n9968, new_n9967, new_n9969);
nor_5  g09593(new_n784, new_n779, new_n9970);
nor_5  g09594(new_n794, new_n785, new_n9971);
nor_5  g09595(new_n9971, new_n9970, new_n9972);
nand_5 g09596(n8236, n6776, new_n9973);
xnor_4 g09597(new_n9973, new_n9972, new_n9974);
xnor_4 g09598(new_n9974, new_n9969, new_n9975);
xnor_4 g09599(new_n9975, new_n9966, new_n9976);
xnor_4 g09600(new_n9976, new_n9963, new_n9977);
xnor_4 g09601(new_n9977, new_n9878, new_n9978);
xnor_4 g09602(new_n9978, new_n9813, new_n9979);
xnor_4 g09603(new_n9979, new_n9810, n7966);
xnor_4 g09604(new_n9622, new_n9621, n7981);
nor_5  g09605(new_n9288, new_n9096, new_n9982);
nor_5  g09606(new_n9298, new_n9289, new_n9983);
nor_5  g09607(new_n9983, new_n9982, new_n9984);
and_5  g09608(new_n9219, new_n9152, new_n9985);
nor_5  g09609(new_n9287, new_n9220, new_n9986);
nor_5  g09610(new_n9986, new_n9985, new_n9987);
nor_5  g09611(new_n9282, new_n9251, new_n9988);
nor_5  g09612(new_n9286, new_n9283, new_n9989);
nor_5  g09613(new_n9989, new_n9988, new_n9990);
nor_5  g09614(new_n9277, new_n9252, new_n9991);
nor_5  g09615(new_n9281, new_n9278, new_n9992);
nor_5  g09616(new_n9992, new_n9991, new_n9993);
nor_5  g09617(new_n9084, new_n9083, new_n9994);
nor_5  g09618(new_n9086, new_n9081, new_n9995);
nor_5  g09619(new_n9995, new_n9994, new_n9996);
and_5  g09620(new_n9267, new_n9266, new_n9997);
nor_5  g09621(new_n9267, new_n9266, new_n9998);
nor_5  g09622(new_n9998, new_n9265, new_n9999);
nor_5  g09623(new_n9999, new_n9997, new_n10000);
and_5  g09624(n8717, n6986, new_n10001);
and_5  g09625(n11222, n10022, new_n10002);
and_5  g09626(n12391, n1353, new_n10003);
xnor_4 g09627(new_n10003, new_n10002, new_n10004);
xnor_4 g09628(new_n10004, new_n10001, new_n10005);
xnor_4 g09629(new_n10005, new_n10000, new_n10006);
xnor_4 g09630(new_n10006, new_n9996, new_n10007);
xnor_4 g09631(new_n10007, new_n9993, new_n10008);
xnor_4 g09632(new_n10008, new_n9990, new_n10009);
nor_5  g09633(new_n9274, new_n9273, new_n10010);
nor_5  g09634(new_n9276, new_n9271, new_n10011);
nor_5  g09635(new_n10011, new_n10010, new_n10012);
nor_5  g09636(new_n9260, new_n9255, new_n10013);
nor_5  g09637(new_n9270, new_n9261, new_n10014);
nor_5  g09638(new_n10014, new_n10013, new_n10015);
and_5  g09639(n12069, n4436, new_n10016);
and_5  g09640(n11999, n11153, new_n10017);
xnor_4 g09641(new_n10017, new_n10016, new_n10018);
and_5  g09642(n7159, n1199, new_n10019);
and_5  g09643(n11967, n7160, new_n10020);
xnor_4 g09644(new_n10020, new_n10019, new_n10021);
xor_4  g09645(new_n10021, new_n10018, new_n10022_1);
and_5  g09646(new_n9258, new_n9257, new_n10023);
nor_5  g09647(new_n9258, new_n9257, new_n10024);
nor_5  g09648(new_n10024, new_n9256, new_n10025);
nor_5  g09649(new_n10025, new_n10023, new_n10026);
and_5  g09650(n6254, n4828, new_n10027);
and_5  g09651(n11407, n2087, new_n10028);
xor_4  g09652(new_n10028, new_n10027, new_n10029);
xnor_4 g09653(new_n10029, new_n10026, new_n10030);
xnor_4 g09654(new_n10030, new_n10022_1, new_n10031);
xnor_4 g09655(new_n10031, new_n10015, new_n10032);
xnor_4 g09656(new_n10032, new_n10012, new_n10033);
nor_5  g09657(new_n9229, new_n9224, new_n10034);
nor_5  g09658(new_n9239, new_n9230, new_n10035);
nor_5  g09659(new_n10035, new_n10034, new_n10036);
and_5  g09660(n12489, n6578, new_n10037);
and_5  g09661(n12947, n996, new_n10038);
and_5  g09662(n9457, n5760, new_n10039);
xnor_4 g09663(new_n10039, new_n10038, new_n10040);
xnor_4 g09664(new_n10040, new_n10037, new_n10041);
xnor_4 g09665(new_n10041, new_n10036, new_n10042);
and_5  g09666(new_n9263, new_n9262, new_n10043);
nor_5  g09667(new_n9269, new_n9264, new_n10044);
nor_5  g09668(new_n10044, new_n10043, new_n10045);
and_5  g09669(n7891, n447, new_n10046);
xnor_4 g09670(new_n10046, new_n10045, new_n10047);
and_5  g09671(n12777, n2515, new_n10048);
nor_5  g09672(new_n9236, new_n9235, new_n10049);
nor_5  g09673(new_n9237, new_n9234, new_n10050);
nor_5  g09674(new_n10050, new_n10049, new_n10051);
nor_5  g09675(new_n9227, new_n9226, new_n10052);
nor_5  g09676(new_n9228, new_n9225, new_n10053);
nor_5  g09677(new_n10053, new_n10052, new_n10054);
xnor_4 g09678(new_n10054, new_n10051, new_n10055);
xnor_4 g09679(new_n10055, new_n10048, new_n10056);
xnor_4 g09680(new_n10056, new_n10047, new_n10057);
and_5  g09681(n6441, n5314, new_n10058);
and_5  g09682(n11791, n5767, new_n10059);
xnor_4 g09683(new_n10059, new_n10058, new_n10060);
and_5  g09684(new_n9232, new_n9231, new_n10061);
nor_5  g09685(new_n9238, new_n9233, new_n10062);
nor_5  g09686(new_n10062, new_n10061, new_n10063);
nand_5 g09687(n6687, n6604, new_n10064);
xnor_4 g09688(new_n10064, new_n10063, new_n10065);
xnor_4 g09689(new_n10065, new_n10060, new_n10066);
xnor_4 g09690(new_n10066, new_n10057, new_n10067);
xnor_4 g09691(new_n10067, new_n10042, new_n10068);
xnor_4 g09692(new_n10068, new_n10033, new_n10069);
nor_5  g09693(new_n9147, new_n9146, new_n10070);
nor_5  g09694(new_n9149, new_n9144, new_n10071);
nor_5  g09695(new_n10071, new_n10070, new_n10072);
nor_5  g09696(new_n9133, new_n9128, new_n10073);
nor_5  g09697(new_n9143, new_n9134, new_n10074);
nor_5  g09698(new_n10074, new_n10073, new_n10075);
and_5  g09699(n10678, n6429, new_n10076);
xnor_4 g09700(new_n10076, new_n10075, new_n10077);
and_5  g09701(new_n9136, new_n9135, new_n10078);
nor_5  g09702(new_n9142, new_n9137_1, new_n10079);
nor_5  g09703(new_n10079, new_n10078, new_n10080);
nand_5 g09704(n2433, n2226, new_n10081);
and_5  g09705(n8819, n1094, new_n10082);
and_5  g09706(n10928, n7730, new_n10083);
xnor_4 g09707(new_n10083, new_n10082, new_n10084);
xnor_4 g09708(new_n10084, new_n10081, new_n10085);
xnor_4 g09709(new_n10085, new_n10080, new_n10086);
xnor_4 g09710(new_n10086, new_n10077, new_n10087);
xnor_4 g09711(new_n10087, new_n10072, new_n10088);
xnor_4 g09712(new_n10088, new_n10069, new_n10089);
nor_5  g09713(new_n9243, new_n9242, new_n10090);
nor_5  g09714(new_n9245, new_n9240, new_n10091);
or_5   g09715(new_n10091, new_n10090, new_n10092);
nor_5  g09716(new_n9087, new_n9062, new_n10093);
nor_5  g09717(new_n9095, new_n9088, new_n10094);
nor_5  g09718(new_n10094, new_n10093, new_n10095);
xnor_4 g09719(new_n10095, new_n10092, new_n10096);
xnor_4 g09720(new_n10096, new_n10089, new_n10097);
nor_5  g09721(new_n9246, new_n9221, new_n10098);
nor_5  g09722(new_n9250, new_n9247, new_n10099);
nor_5  g09723(new_n10099, new_n10098, new_n10100);
nor_5  g09724(new_n9150, new_n9125, new_n10101);
nor_5  g09725(new_n9151, new_n9124, new_n10102);
nor_5  g09726(new_n10102, new_n10101, new_n10103);
nor_5  g09727(new_n9070, new_n9065, new_n10104);
nor_5  g09728(new_n9080_1, new_n9071, new_n10105);
nor_5  g09729(new_n10105, new_n10104, new_n10106);
and_5  g09730(new_n9068, new_n9067, new_n10107);
nor_5  g09731(new_n9068, new_n9067, new_n10108);
nor_5  g09732(new_n10108, new_n9066, new_n10109);
nor_5  g09733(new_n10109, new_n10107, new_n10110);
and_5  g09734(n12709, n7523, new_n10111);
and_5  g09735(n12000, n4189, new_n10112);
xor_4  g09736(new_n10112, new_n10111, new_n10113);
xnor_4 g09737(new_n10113, new_n10110, new_n10114);
and_5  g09738(n9725, n2564, new_n10115);
and_5  g09739(n9920, n4370, new_n10116);
xnor_4 g09740(new_n10116, new_n10115, new_n10117);
nand_5 g09741(n5212, n4516, new_n10118);
and_5  g09742(n6770, n5320, new_n10119);
and_5  g09743(n5319, n1478, new_n10120);
xnor_4 g09744(new_n10120, new_n10119, new_n10121);
xnor_4 g09745(new_n10121, new_n10118, new_n10122);
xnor_4 g09746(new_n10122, new_n10117, new_n10123);
nand_5 g09747(n11728, n7320, new_n10124);
nor_5  g09748(new_n9140, new_n9139, new_n10125);
nor_5  g09749(new_n9141, new_n9138, new_n10126);
nor_5  g09750(new_n10126, new_n10125, new_n10127);
xnor_4 g09751(new_n10127, new_n10124, new_n10128);
xnor_4 g09752(new_n10128, new_n10123, new_n10129);
xnor_4 g09753(new_n10129, new_n10114, new_n10130);
and_5  g09754(new_n9077, new_n9076, new_n10131);
nor_5  g09755(new_n9077, new_n9076, new_n10132);
nor_5  g09756(new_n10132, new_n9075, new_n10133);
nor_5  g09757(new_n10133, new_n10131, new_n10134);
nand_5 g09758(n10990, n4817, new_n10135);
and_5  g09759(n11877, n3627, new_n10136);
and_5  g09760(n8336, n1198, new_n10137);
xnor_4 g09761(new_n10137, new_n10136, new_n10138);
xnor_4 g09762(new_n10138, new_n10135, new_n10139);
xnor_4 g09763(new_n10139, new_n10134, new_n10140);
and_5  g09764(new_n9073, new_n9072, new_n10141);
nor_5  g09765(new_n9079, new_n9074, new_n10142);
nor_5  g09766(new_n10142, new_n10141, new_n10143);
nor_5  g09767(new_n9131, new_n9130, new_n10144);
nor_5  g09768(new_n9132, new_n9129, new_n10145);
nor_5  g09769(new_n10145, new_n10144, new_n10146);
xnor_4 g09770(new_n10146, new_n10143, new_n10147);
xnor_4 g09771(new_n10147, new_n10140, new_n10148);
xnor_4 g09772(new_n10148, new_n10130, new_n10149);
xor_4  g09773(new_n10149, new_n10106, new_n10150);
xnor_4 g09774(new_n10150, new_n10103, new_n10151);
xnor_4 g09775(new_n10151, new_n10100, new_n10152);
xnor_4 g09776(new_n10152, new_n10097, new_n10153);
xnor_4 g09777(new_n10153, new_n10009, new_n10154);
xnor_4 g09778(new_n10154, new_n9987, new_n10155);
xnor_4 g09779(new_n10155, new_n9984, n8100);
xnor_4 g09780(new_n7432, new_n7431, n8138);
xnor_4 g09781(new_n4667, new_n4666, n8202);
xor_4  g09782(new_n2894, new_n2886, n8303);
xnor_4 g09783(new_n2335, new_n2334, n8398);
xnor_4 g09784(new_n3333, new_n3332, n9137);
xnor_4 g09785(new_n5442, new_n5441, n9387);
xnor_4 g09786(new_n8855, new_n8854, n9571);
xor_4  g09787(new_n772, new_n771, n9578);
xor_4  g09788(new_n981, new_n980, n9706);
xnor_4 g09789(new_n3335, new_n3327, n9756);
and_5  g09790(new_n5183, new_n4926, new_n10167);
nor_5  g09791(new_n5183, new_n4926, new_n10168);
nor_5  g09792(new_n5199, new_n10168, new_n10169);
nor_5  g09793(new_n10169, new_n10167, new_n10170);
nand_5 g09794(n12826, n7891, new_n10171);
nor_5  g09795(new_n4986, new_n4985, new_n10172);
nor_5  g09796(new_n4988, new_n4983, new_n10173);
nor_5  g09797(new_n10173, new_n10172, new_n10174_1);
xnor_4 g09798(new_n10174_1, new_n10171, new_n10175);
nor_5  g09799(new_n5164, new_n5000, new_n10176);
nor_5  g09800(new_n5182, new_n5165, new_n10177);
nor_5  g09801(new_n10177, new_n10176, new_n10178);
and_5  g09802(n8336, n2278, new_n10179);
nor_5  g09803(new_n4915, new_n4890, new_n10180);
nor_5  g09804(new_n4925, new_n4916, new_n10181);
nor_5  g09805(new_n10181, new_n10180, new_n10182);
xnor_4 g09806(new_n10182, new_n10179, new_n10183);
and_5  g09807(new_n5062, new_n5037, new_n10184);
nor_5  g09808(new_n5073, new_n5063, new_n10185);
nor_5  g09809(new_n10185, new_n10184, new_n10186);
and_5  g09810(new_n4901, new_n4900, new_n10187);
nor_5  g09811(new_n4907, new_n4902, new_n10188);
nor_5  g09812(new_n10188, new_n10187, new_n10189);
nor_5  g09813(new_n4972, new_n4967, new_n10190);
nor_5  g09814(new_n4982, new_n4973, new_n10191);
nor_5  g09815(new_n10191, new_n10190, new_n10192);
and_5  g09816(n11662, n6770, new_n10193);
and_5  g09817(n10451, n2226, new_n10194);
and_5  g09818(n5319, n3754, new_n10195);
xnor_4 g09819(new_n10195, new_n10194, new_n10196);
xnor_4 g09820(new_n10196, new_n10193, new_n10197);
nor_5  g09821(new_n4979, new_n4978, new_n10198);
nor_5  g09822(new_n4980, new_n4977, new_n10199);
nor_5  g09823(new_n10199, new_n10198, new_n10200);
xnor_4 g09824(new_n10200, new_n10197, new_n10201);
and_5  g09825(new_n4905, new_n4904, new_n10202);
nor_5  g09826(new_n4905, new_n4904, new_n10203);
nor_5  g09827(new_n10203, new_n4903_1, new_n10204);
nor_5  g09828(new_n10204, new_n10202, new_n10205);
and_5  g09829(n10278, n6986, new_n10206);
and_5  g09830(n10678, n3022, new_n10207);
xor_4  g09831(new_n10207, new_n10206, new_n10208);
xnor_4 g09832(new_n10208, new_n10205, new_n10209);
xnor_4 g09833(new_n10209, new_n10201, new_n10210);
and_5  g09834(new_n4975, new_n4974, new_n10211);
nor_5  g09835(new_n4981, new_n4976, new_n10212);
nor_5  g09836(new_n10212, new_n10211, new_n10213);
nor_5  g09837(new_n4970_1, new_n4969, new_n10214);
nor_5  g09838(new_n4971_1, new_n4968, new_n10215);
or_5   g09839(new_n10215, new_n10214, new_n10216);
xnor_4 g09840(new_n10216, new_n10213, new_n10217_1);
xnor_4 g09841(new_n10217_1, new_n10210, new_n10218);
xnor_4 g09842(new_n10218, new_n10192, new_n10219);
xnor_4 g09843(new_n10219, new_n10189, new_n10220);
nor_5  g09844(new_n4896, new_n4895, new_n10221);
nor_5  g09845(new_n4897, new_n4894, new_n10222);
nor_5  g09846(new_n10222, new_n10221, new_n10223_1);
nand_5 g09847(n8665, n2515, new_n10224);
and_5  g09848(n10898, n9457, new_n10225);
and_5  g09849(n12511, n11222, new_n10226);
xnor_4 g09850(new_n10226, new_n10225, new_n10227);
xnor_4 g09851(new_n10227, new_n10224, new_n10228);
xnor_4 g09852(new_n10228, new_n10223_1, new_n10229);
xnor_4 g09853(new_n10229, new_n10220, new_n10230);
nand_5 g09854(n12391, n4094, new_n10231);
nor_5  g09855(new_n4898, new_n4893, new_n10232);
nor_5  g09856(new_n4908, new_n4899, new_n10233);
nor_5  g09857(new_n10233, new_n10232, new_n10234);
and_5  g09858(n4516, n3932, new_n10235);
and_5  g09859(n7523, n6703, new_n10236);
xnor_4 g09860(new_n10236, new_n10235, new_n10237);
and_5  g09861(n11423, n10928, new_n10238);
and_5  g09862(n12591, n3627, new_n10239);
xnor_4 g09863(new_n10239, new_n10238, new_n10240);
xnor_4 g09864(new_n10240, new_n10237, new_n10241);
xnor_4 g09865(new_n10241, new_n10234, new_n10242);
and_5  g09866(n11876, n4817, new_n10243);
and_5  g09867(new_n5052, new_n5051, new_n10244);
nor_5  g09868(new_n5052, new_n5051, new_n10245);
nor_5  g09869(new_n10245, new_n5050, new_n10246);
nor_5  g09870(new_n10246, new_n10244, new_n10247);
and_5  g09871(n10327, n4189, new_n10248);
and_5  g09872(n9920, n7456, new_n10249);
xnor_4 g09873(new_n10249, new_n10248, new_n10250);
xnor_4 g09874(new_n10250, new_n10247, new_n10251);
xnor_4 g09875(new_n10251, new_n10243, new_n10252);
xnor_4 g09876(new_n10252, new_n10242, new_n10253);
xnor_4 g09877(new_n10253, new_n10231, new_n10254);
xnor_4 g09878(new_n10254, new_n10230, new_n10255);
xnor_4 g09879(new_n10255, new_n10186, new_n10256);
xnor_4 g09880(new_n10256, new_n10183, new_n10257);
nor_5  g09881(new_n4912, new_n4911, new_n10258);
nor_5  g09882(new_n4914, new_n4909, new_n10259);
nor_5  g09883(new_n10259, new_n10258, new_n10260);
nor_5  g09884(new_n5059, new_n5058, new_n10261);
nor_5  g09885(new_n5061, new_n5056, new_n10262);
nor_5  g09886(new_n10262, new_n10261, new_n10263);
xnor_4 g09887(new_n10263, new_n10260, new_n10264);
nor_5  g09888(new_n5113, new_n5112, new_n10265);
nor_5  g09889(new_n5134, new_n5115, new_n10266);
nor_5  g09890(new_n10266, new_n10265, new_n10267);
nand_5 g09891(n11023, n1094, new_n10268);
xnor_4 g09892(new_n10268, new_n10267, new_n10269);
nor_5  g09893(new_n5123, new_n5118, new_n10270);
nor_5  g09894(new_n5133, new_n5124, new_n10271);
nor_5  g09895(new_n10271, new_n10270, new_n10272);
and_5  g09896(new_n5048, new_n5047, new_n10273);
nor_5  g09897(new_n5054, new_n5049, new_n10274);
nor_5  g09898(new_n10274, new_n10273, new_n10275);
nor_5  g09899(new_n5121, new_n5120, new_n10276);
nor_5  g09900(new_n5122, new_n5119, new_n10277);
nor_5  g09901(new_n10277, new_n10276, new_n10278_1);
nor_5  g09902(new_n5130, new_n5129, new_n10279);
nor_5  g09903(new_n5131, new_n5128, new_n10280);
nor_5  g09904(new_n10280, new_n10279, new_n10281);
xnor_4 g09905(new_n10281, new_n10278_1, new_n10282);
and_5  g09906(n12069, n10685, new_n10283);
and_5  g09907(n6578, n5645, new_n10284);
xor_4  g09908(new_n10284, new_n10283, new_n10285);
nand_5 g09909(n5767, n2749, new_n10286);
and_5  g09910(n996, n159, new_n10287);
and_5  g09911(n5314, n1510, new_n10288);
xnor_4 g09912(new_n10288, new_n10287, new_n10289);
xnor_4 g09913(new_n10289, new_n10286, new_n10290);
xnor_4 g09914(new_n10290, new_n10285, new_n10291);
xnor_4 g09915(new_n10291, new_n10282, new_n10292);
and_5  g09916(new_n5126, new_n5125, new_n10293);
nor_5  g09917(new_n5132_1, new_n5127, new_n10294);
nor_5  g09918(new_n10294, new_n10293, new_n10295);
nand_5 g09919(n7160, n2551, new_n10296);
and_5  g09920(n9583, n2564, new_n10297);
and_5  g09921(n9640, n7320, new_n10298);
xnor_4 g09922(new_n10298, new_n10297, new_n10299);
xnor_4 g09923(new_n10299, new_n10296, new_n10300);
and_5  g09924(n1199, n1067, new_n10301);
and_5  g09925(n12247, n11153, new_n10302);
xnor_4 g09926(new_n10302, new_n10301, new_n10303);
xnor_4 g09927(new_n10303, new_n10300, new_n10304);
xnor_4 g09928(new_n10304, new_n10295, new_n10305);
xnor_4 g09929(new_n10305, new_n10292, new_n10306);
xnor_4 g09930(new_n10306, new_n10275, new_n10307);
nor_5  g09931(new_n5045, new_n5040, new_n10308);
nor_5  g09932(new_n5055, new_n5046, new_n10309);
nor_5  g09933(new_n10309, new_n10308, new_n10310);
nor_5  g09934(new_n5043, new_n5042, new_n10311);
nor_5  g09935(new_n5044, new_n5041, new_n10312);
nor_5  g09936(new_n10312, new_n10311, new_n10313);
and_5  g09937(n6687, n753, new_n10314);
and_5  g09938(n2087, n1798, new_n10315);
xnor_4 g09939(new_n10315, new_n10314, new_n10316);
xnor_4 g09940(new_n10316, new_n10313, new_n10317);
xnor_4 g09941(new_n10317, new_n10310, new_n10318);
xnor_4 g09942(new_n10318, new_n10307, new_n10319);
xnor_4 g09943(new_n10319, new_n10272, new_n10320);
xnor_4 g09944(new_n10320, new_n10269, new_n10321);
xnor_4 g09945(new_n10321, new_n10264, new_n10322);
nor_5  g09946(new_n5135, new_n5110, new_n10323);
nor_5  g09947(new_n5146, new_n5136, new_n10324);
nor_5  g09948(new_n10324, new_n10323, new_n10325);
nor_5  g09949(new_n4989, new_n4964, new_n10326);
nor_5  g09950(new_n4999, new_n4990, new_n10327_1);
nor_5  g09951(new_n10327_1, new_n10326, new_n10328);
xnor_4 g09952(new_n10328, new_n10325, new_n10329);
xnor_4 g09953(new_n10329, new_n10322, new_n10330);
xnor_4 g09954(new_n10330, new_n10257, new_n10331);
and_5  g09955(n11922, n4828, new_n10332);
nor_5  g09956(new_n5162, new_n5147, new_n10333);
nor_5  g09957(new_n5163, new_n5074, new_n10334);
nor_5  g09958(new_n10334, new_n10333, new_n10335);
xnor_4 g09959(new_n10335, new_n10332, new_n10336);
xnor_4 g09960(new_n10336, new_n10331, new_n10337);
xnor_4 g09961(new_n10337, new_n10178, new_n10338);
xnor_4 g09962(new_n10338, new_n10175, new_n10339);
xnor_4 g09963(new_n10339, new_n10170, n9767);
xnor_4 g09964(new_n1665, new_n1664, n9820);
xnor_4 g09965(new_n7447, new_n7446, n9938);
xor_4  g09966(new_n767, new_n766, n10476);
xnor_4 g09967(new_n764, new_n756, n10589);
xnor_4 g09968(new_n978, new_n977, n10695);
xnor_4 g09969(new_n2875, new_n2615, new_n10346);
xnor_4 g09970(new_n10346, new_n2909, n10789);
xor_4  g09971(new_n2330, new_n2322, n10851);
xnor_4 g09972(new_n3907, new_n3899, n10913);
xnor_4 g09973(new_n5552, new_n5446, n10949);
xnor_4 g09974(new_n8857, new_n8820, n11216);
xor_4  g09975(new_n3900, new_n3892, n11326);
nor_5  g09976(new_n4334, new_n4166, new_n10353);
nor_5  g09977(new_n4437, new_n4335, new_n10354);
nor_5  g09978(new_n10354, new_n10353, new_n10355);
nor_5  g09979(new_n4368, new_n4365, new_n10356);
nor_5  g09980(new_n4436_1, new_n4369, new_n10357);
nor_5  g09981(new_n10357, new_n10356, new_n10358);
nor_5  g09982(new_n4363, new_n4339, new_n10359);
nor_5  g09983(new_n4364, new_n4338, new_n10360);
nor_5  g09984(new_n10360, new_n10359, new_n10361);
nor_5  g09985(new_n4360, new_n4359, new_n10362);
nor_5  g09986(new_n4362, new_n4357, new_n10363);
nor_5  g09987(new_n10363, new_n10362, new_n10364);
and_5  g09988(n9763, n45, new_n10365);
and_5  g09989(n8759, n7823, new_n10366);
xor_4  g09990(new_n10366, new_n10365, new_n10367);
xnor_4 g09991(new_n10367, new_n10364, new_n10368);
nor_5  g09992(new_n4145, new_n4144, new_n10369);
nor_5  g09993(new_n4146, new_n4143, new_n10370);
nor_5  g09994(new_n10370, new_n10369, new_n10371);
and_5  g09995(n9241, n9189, new_n10372);
xnor_4 g09996(new_n10372, new_n10371, new_n10373);
and_5  g09997(n12705, n4634, new_n10374);
and_5  g09998(n12145, n7436, new_n10375);
xnor_4 g09999(new_n10375, new_n10374, new_n10376);
and_5  g10000(n9195, n4312, new_n10377);
and_5  g10001(n10217, n6776, new_n10378);
xnor_4 g10002(new_n10378, new_n10377, new_n10379);
xor_4  g10003(new_n10379, new_n10376, new_n10380);
xnor_4 g10004(new_n10380, new_n10373, new_n10381);
and_5  g10005(new_n4349, new_n4348, new_n10382);
nor_5  g10006(new_n4355, new_n4350, new_n10383);
nor_5  g10007(new_n10383, new_n10382, new_n10384);
nor_5  g10008(new_n4344, new_n4343, new_n10385);
nor_5  g10009(new_n4345, new_n4342, new_n10386);
or_5   g10010(new_n10386, new_n10385, new_n10387);
xnor_4 g10011(new_n10387, new_n10384, new_n10388);
xnor_4 g10012(new_n10388, new_n10381, new_n10389);
and_5  g10013(new_n4353, new_n4352, new_n10390);
nor_5  g10014(new_n4353, new_n4352, new_n10391_1);
nor_5  g10015(new_n10391_1, new_n4351, new_n10392);
nor_5  g10016(new_n10392, new_n10390, new_n10393);
xnor_4 g10017(new_n10393, new_n10389, new_n10394);
and_5  g10018(n3986, n3342, new_n10395);
and_5  g10019(n8276, n2522, new_n10396);
and_5  g10020(n12299, n12221, new_n10397);
xnor_4 g10021(new_n10397, new_n10396, new_n10398);
xnor_4 g10022(new_n10398, new_n10395, new_n10399);
xnor_4 g10023(new_n10399, new_n10394, new_n10400);
nor_5  g10024(new_n4346, new_n4341, new_n10401);
nor_5  g10025(new_n4356, new_n4347, new_n10402);
nor_5  g10026(new_n10402, new_n10401, new_n10403);
nor_5  g10027(new_n4423, new_n4422, new_n10404);
nor_5  g10028(new_n4425, new_n4420, new_n10405);
or_5   g10029(new_n10405, new_n10404, new_n10406);
xnor_4 g10030(new_n10406, new_n10403, new_n10407);
xnor_4 g10031(new_n10407, new_n10400, new_n10408);
xnor_4 g10032(new_n10408, new_n10368, new_n10409);
xnor_4 g10033(new_n10409, new_n10361, new_n10410);
nand_5 g10034(n12025, n10223, new_n10411);
and_5  g10035(new_n4141_1, new_n4140, new_n10412);
nor_5  g10036(new_n4147, new_n4142, new_n10413);
nor_5  g10037(new_n10413, new_n10412, new_n10414);
xnor_4 g10038(new_n10414, new_n10411, new_n10415);
xnor_4 g10039(new_n10415, new_n10410, new_n10416);
nor_5  g10040(new_n4409, new_n4404, new_n10417);
nor_5  g10041(new_n4419, new_n4410, new_n10418);
nor_5  g10042(new_n10418, new_n10417, new_n10419);
and_5  g10043(n7690, n5579, new_n10420);
and_5  g10044(n7388, n2507, new_n10421);
xnor_4 g10045(new_n10421, new_n10420, new_n10422);
and_5  g10046(n7270, n2393, new_n10423);
and_5  g10047(n5331, n1576, new_n10424);
xnor_4 g10048(new_n10424, new_n10423, new_n10425);
xnor_4 g10049(new_n10425, new_n10422, new_n10426);
and_5  g10050(n3616, n2498, new_n10427);
and_5  g10051(n12648, n6016, new_n10428);
xor_4  g10052(new_n10428, new_n10427, new_n10429);
xnor_4 g10053(new_n10429, new_n10426, new_n10430);
and_5  g10054(n5798, n2530, new_n10431);
and_5  g10055(n10644, n7946, new_n10432);
xor_4  g10056(new_n10432, new_n10431, new_n10433);
nor_5  g10057(new_n4407, new_n4406, new_n10434);
nor_5  g10058(new_n4408, new_n4405, new_n10435);
nor_5  g10059(new_n10435, new_n10434, new_n10436);
nor_5  g10060(new_n4136, new_n4135, new_n10437);
nor_5  g10061(new_n4137, new_n4134, new_n10438);
nor_5  g10062(new_n10438, new_n10437, new_n10439_1);
xnor_4 g10063(new_n10439_1, new_n10436, new_n10440);
xnor_4 g10064(new_n10440, new_n10433, new_n10441);
xnor_4 g10065(new_n10441, new_n10430, new_n10442);
xnor_4 g10066(new_n10442, new_n10419, new_n10443);
nor_5  g10067(new_n4392, new_n4391, new_n10444);
nor_5  g10068(new_n4394, new_n4389, new_n10445);
nor_5  g10069(new_n10445, new_n10444, new_n10446);
nor_5  g10070(new_n4416, new_n4415, new_n10447);
nor_5  g10071(new_n4417, new_n4414, new_n10448);
or_5   g10072(new_n10448, new_n10447, new_n10449);
and_5  g10073(new_n4412, new_n4411, new_n10450);
nor_5  g10074(new_n4418, new_n4413, new_n10451_1);
nor_5  g10075(new_n10451_1, new_n10450, new_n10452);
and_5  g10076(n7965, n6431, new_n10453);
and_5  g10077(n9111, n5857, new_n10454);
xnor_4 g10078(new_n10454, new_n10453, new_n10455);
and_5  g10079(n11892, n5153, new_n10456);
and_5  g10080(n5860, n806, new_n10457);
xnor_4 g10081(new_n10457, new_n10456, new_n10458);
and_5  g10082(n10545, n521, new_n10459);
and_5  g10083(n10547, n7265, new_n10460);
xnor_4 g10084(new_n10460, new_n10459, new_n10461);
xnor_4 g10085(new_n10461, new_n10458, new_n10462);
xnor_4 g10086(new_n10462, new_n10455, new_n10463);
xnor_4 g10087(new_n10463, new_n10452, new_n10464);
xnor_4 g10088(new_n10464, new_n10449, new_n10465);
xnor_4 g10089(new_n10465, new_n10446, new_n10466);
nor_5  g10090(new_n4138, new_n4133, new_n10467);
nor_5  g10091(new_n4148, new_n4139, new_n10468);
nor_5  g10092(new_n10468, new_n10467, new_n10469);
and_5  g10093(new_n4381, new_n4380, new_n10470);
nor_5  g10094(new_n4387, new_n4382, new_n10471);
or_5   g10095(new_n10471, new_n10470, new_n10472);
xnor_4 g10096(new_n10472, new_n10469, new_n10473);
xnor_4 g10097(new_n10473, new_n10466, new_n10474);
xnor_4 g10098(new_n10474, new_n10443, new_n10475);
nor_5  g10099(new_n4395, new_n4370_1, new_n10476_1);
nor_5  g10100(new_n4399, new_n4396, new_n10477);
nor_5  g10101(new_n10477, new_n10476_1, new_n10478);
nor_5  g10102(new_n4152, new_n4151, new_n10479);
nor_5  g10103(new_n4154, new_n4149, new_n10480);
nor_5  g10104(new_n10480, new_n10479, new_n10481);
nor_5  g10105(new_n4378_1, new_n4375, new_n10482);
nor_5  g10106(new_n4388, new_n4379, new_n10483);
nor_5  g10107(new_n10483, new_n10482, new_n10484);
nor_5  g10108(new_n4385, new_n4384, new_n10485);
nor_5  g10109(new_n4386, new_n4383, new_n10486);
nor_5  g10110(new_n10486, new_n10485, new_n10487);
and_5  g10111(n4499, n2558, new_n10488);
and_5  g10112(n5305, n2512, new_n10489);
xor_4  g10113(new_n10489, new_n10488, new_n10490);
xnor_4 g10114(new_n10490, new_n10487, new_n10491);
nor_5  g10115(new_n4374, new_n4371, new_n10492);
or_5   g10116(new_n10492, new_n4372, new_n10493);
nand_5 g10117(n8476, n2347, new_n10494);
nor_5  g10118(new_n10494, new_n10493, new_n10495);
or_5   g10119(new_n10494, new_n4265, new_n10496);
and_5  g10120(new_n10496, new_n10493, new_n10497);
nor_5  g10121(new_n10497, new_n10495, new_n10498);
and_5  g10122(n2253, n1097, new_n10499);
and_5  g10123(n5964, n3865, new_n10500);
xor_4  g10124(new_n10500, new_n10499, new_n10501);
xnor_4 g10125(new_n10501, new_n10498, new_n10502);
xnor_4 g10126(new_n10502, new_n10491, new_n10503);
xnor_4 g10127(new_n10503, new_n10484, new_n10504);
and_5  g10128(n10510, n2024, new_n10505);
and_5  g10129(n11257, n2879, new_n10506);
xnor_4 g10130(new_n10506, new_n10505, new_n10507);
xnor_4 g10131(new_n10507, new_n10504, new_n10508);
xnor_4 g10132(new_n10508, new_n10481, new_n10509);
xnor_4 g10133(new_n10509, new_n10478, new_n10510_1);
xnor_4 g10134(new_n10510_1, new_n10475, new_n10511);
xnor_4 g10135(new_n10511, new_n10416, new_n10512);
nor_5  g10136(new_n4431, new_n4400, new_n10513);
nor_5  g10137(new_n4435, new_n4432, new_n10514);
nor_5  g10138(new_n10514, new_n10513, new_n10515);
nor_5  g10139(new_n4155_1, new_n4131, new_n10516);
nor_5  g10140(new_n4165, new_n4156, new_n10517);
nor_5  g10141(new_n10517, new_n10516, new_n10518);
and_5  g10142(new_n4426, new_n4401, new_n10519);
nor_5  g10143(new_n4430, new_n4427, new_n10520);
nor_5  g10144(new_n10520, new_n10519, new_n10521);
xnor_4 g10145(new_n10521, new_n10518, new_n10522);
xnor_4 g10146(new_n10522, new_n10515, new_n10523);
xnor_4 g10147(new_n10523, new_n10512, new_n10524);
xnor_4 g10148(new_n10524, new_n10358, new_n10525);
xnor_4 g10149(new_n10525, new_n10355, n11707);
xnor_4 g10150(new_n4818, new_n4817_1, n11755);
xor_4  g10151(new_n2904, new_n2903, n11780);
xnor_4 g10152(new_n7765, new_n7764, n11919);
xor_4  g10153(new_n7767, new_n7754, n12005);
xnor_4 g10154(new_n8095, new_n8092, n12014);
xor_4  g10155(new_n6781, new_n6760, n12020);
xnor_4 g10156(new_n8850, new_n8825, n12076);
xnor_4 g10157(new_n9296, new_n9295, n12111);
xnor_4 g10158(new_n8097, new_n8088, n12444);
xnor_4 g10159(new_n4332, new_n4323, n12807);
endmodule


