// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Thu Jun 27 02:26:40 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095,
    new_n1096, new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269_1, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1318,
    new_n1319, new_n1320, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333_1, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355,
    new_n1356, new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471_1, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1,
    new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389,
    new_n2390, new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1,
    new_n2432, new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2462,
    new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1, new_n2510,
    new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339_1, new_n3340, new_n3342_1, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986_1, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992_1, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005_1,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086_1, new_n4087, new_n4088_1, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094_1, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155_1, new_n4156,
    new_n4157, new_n4158, new_n4159_1, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187_1, new_n4188, new_n4189_1, new_n4190_1, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203_1, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226_1, new_n4227, new_n4228,
    new_n4229, new_n4230_1, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300_1, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312_1, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326_1, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333_1, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370_1, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378_1, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397_1,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436_1, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499_1,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516_1, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553_1,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4624, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634_1, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686_1, new_n4687, new_n4688, new_n4689_1,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733_1, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757_1, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805_1, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817_1, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826_1, new_n4827,
    new_n4828_1, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212_1, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314_1, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1,
    new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481,
    new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487,
    new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493,
    new_n5494, new_n5495, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643, new_n5644,
    new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859, new_n5860_1,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934_1, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089_1,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254_1, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273_1, new_n6274, new_n6275,
    new_n6276, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294_1,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358_1, new_n6359_1, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429_1, new_n6430, new_n6431_1, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441_1, new_n6442, new_n6443, new_n6444,
    new_n6445_1, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6547, new_n6549,
    new_n6550, new_n6551, new_n6552, new_n6553, new_n6554, new_n6555,
    new_n6556, new_n6557, new_n6558, new_n6559, new_n6560, new_n6561,
    new_n6562, new_n6563, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578_1, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604_1, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611_1, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645_1,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687_1,
    new_n6688, new_n6689_1, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703_1, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742_1, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770_1, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776_1, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797_1, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806_1, new_n6807,
    new_n6808, new_n6809_1, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822_1, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860_1, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877_1, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986_1, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159_1, new_n7160_1, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193_1,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265_1,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270_1, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294_1, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320_1, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523_1,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7681,
    new_n7685, new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009,
    new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028_1, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100_1, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8202_1,
    new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208,
    new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214,
    new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220,
    new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303_1, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336_1, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8376, new_n8377, new_n8378, new_n8379,
    new_n8380, new_n8381, new_n8382, new_n8383, new_n8384_1, new_n8385,
    new_n8386, new_n8387, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398_1, new_n8399,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405,
    new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417,
    new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423,
    new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432, new_n8433_1, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8488, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595_1, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665_1, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717_1, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759_1, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819_1, new_n8820, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930,
    new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080_1,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111_1, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137_1, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189_1, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195_1, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241_1, new_n9242,
    new_n9243, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387_1, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400_1, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457_1, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571_1, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578_1, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583_1, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637_1, new_n9638, new_n9639, new_n9640_1, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706_1, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725_1,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756_1, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820_1, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920_1, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956_1, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022_1, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174_1, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217_1, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223_1, new_n10224, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278_1, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295, new_n10296, new_n10297,
    new_n10298, new_n10299, new_n10300, new_n10301, new_n10302, new_n10303,
    new_n10304, new_n10305, new_n10306, new_n10307, new_n10308, new_n10309,
    new_n10310, new_n10311, new_n10312, new_n10313, new_n10314, new_n10315,
    new_n10316, new_n10317, new_n10318, new_n10319, new_n10320, new_n10321,
    new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327_1, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391_1, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10409, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439_1, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451_1, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476_1,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510_1, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545_1, new_n10546,
    new_n10547_1, new_n10548, new_n10549, new_n10550, new_n10551,
    new_n10552, new_n10553, new_n10554, new_n10555, new_n10556, new_n10557,
    new_n10558, new_n10559, new_n10560, new_n10561, new_n10562, new_n10563,
    new_n10564, new_n10565, new_n10566, new_n10567, new_n10568, new_n10569,
    new_n10570, new_n10571, new_n10572, new_n10573, new_n10574, new_n10575,
    new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589_1, new_n10590, new_n10591, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616,
    new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622,
    new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628,
    new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644_1, new_n10645,
    new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651,
    new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678_1, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685_1,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695_1, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789_1, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848_1, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898_1, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913_1,
    new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943, new_n10944, new_n10945, new_n10946,
    new_n10947, new_n10948, new_n10949_1, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961, new_n10962, new_n10963,
    new_n10964, new_n10965_1, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990_1, new_n10991,
    new_n10992, new_n10993, new_n10994, new_n10995, new_n10996, new_n10997,
    new_n10998, new_n10999, new_n11000, new_n11001, new_n11002, new_n11003,
    new_n11004, new_n11005, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011, new_n11012, new_n11013, new_n11014, new_n11015,
    new_n11016, new_n11017, new_n11018, new_n11019, new_n11020, new_n11021,
    new_n11022, new_n11023_1, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11095, new_n11096, new_n11097, new_n11098, new_n11099,
    new_n11100, new_n11101, new_n11102, new_n11103, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120, new_n11121, new_n11122, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129,
    new_n11130, new_n11131, new_n11132, new_n11133, new_n11134, new_n11135,
    new_n11136, new_n11137, new_n11138, new_n11139, new_n11140, new_n11141,
    new_n11142, new_n11143, new_n11144, new_n11145, new_n11146, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153_1, new_n11154, new_n11155, new_n11156, new_n11157,
    new_n11158, new_n11159, new_n11160, new_n11161, new_n11162, new_n11163,
    new_n11164, new_n11165, new_n11166, new_n11167, new_n11168, new_n11169,
    new_n11170, new_n11171, new_n11172, new_n11173, new_n11174, new_n11175,
    new_n11176, new_n11177, new_n11178, new_n11179, new_n11180, new_n11181,
    new_n11182, new_n11183, new_n11184, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201, new_n11202, new_n11203, new_n11204, new_n11205,
    new_n11206, new_n11207, new_n11208, new_n11209, new_n11210, new_n11211,
    new_n11212, new_n11213, new_n11214, new_n11215, new_n11216_1,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221,
    new_n11222_1, new_n11223, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238,
    new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244,
    new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257_1, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311_1, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326_1, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407_1,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423_1, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478_1, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536_1, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612,
    new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662_1, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667, new_n11668, new_n11669, new_n11670, new_n11671,
    new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707_1, new_n11708, new_n11709, new_n11710, new_n11711,
    new_n11712, new_n11713, new_n11714, new_n11715, new_n11716, new_n11717,
    new_n11718, new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724, new_n11725, new_n11726, new_n11727, new_n11728_1,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755_1, new_n11756, new_n11757_1,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780_1,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791_1,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821_1, new_n11822, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843,
    new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855,
    new_n11856, new_n11857, new_n11858, new_n11859, new_n11860, new_n11861,
    new_n11862, new_n11863, new_n11864, new_n11865, new_n11866, new_n11867,
    new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873,
    new_n11874, new_n11875, new_n11876_1, new_n11877_1, new_n11878,
    new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884,
    new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891, new_n11892_1, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917_1, new_n11918,
    new_n11919_1, new_n11920, new_n11921, new_n11922_1, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11936, new_n11943, new_n11944, new_n11945, new_n11946,
    new_n11947, new_n11948, new_n11949, new_n11950, new_n11951, new_n11952,
    new_n11953, new_n11954, new_n11955, new_n11956, new_n11957, new_n11958,
    new_n11959, new_n11960, new_n11961, new_n11962, new_n11963, new_n11964,
    new_n11965, new_n11966, new_n11967_1, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980, new_n11981,
    new_n11982, new_n11983, new_n11984, new_n11985, new_n11986, new_n11987,
    new_n11988, new_n11989, new_n11990, new_n11991, new_n11992, new_n11993,
    new_n11994, new_n11995, new_n11996, new_n11997, new_n11998,
    new_n11999_1, new_n12000_1, new_n12001, new_n12002, new_n12003,
    new_n12004, new_n12005_1, new_n12006, new_n12007, new_n12008,
    new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014_1, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020_1, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025_1, new_n12026, new_n12027, new_n12028,
    new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044_1, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069_1, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076_1, new_n12077, new_n12078,
    new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108,
    new_n12109, new_n12110, new_n12111_1, new_n12112, new_n12113,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121, new_n12122, new_n12123, new_n12124, new_n12125,
    new_n12126, new_n12127, new_n12128, new_n12129, new_n12130, new_n12131,
    new_n12132, new_n12133, new_n12134, new_n12135, new_n12136, new_n12137,
    new_n12138, new_n12139, new_n12140, new_n12141, new_n12142, new_n12143,
    new_n12144, new_n12145_1, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221_1, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247_1, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299_1, new_n12300, new_n12301, new_n12302, new_n12303,
    new_n12304, new_n12305, new_n12306, new_n12307, new_n12308, new_n12309,
    new_n12310, new_n12311, new_n12312, new_n12313, new_n12314, new_n12315,
    new_n12316, new_n12317, new_n12318, new_n12319, new_n12320, new_n12321,
    new_n12322, new_n12323, new_n12324, new_n12325, new_n12326, new_n12327,
    new_n12328, new_n12329, new_n12330, new_n12331, new_n12332, new_n12333,
    new_n12334, new_n12335, new_n12336, new_n12337, new_n12338, new_n12339,
    new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12354, new_n12355, new_n12356, new_n12357,
    new_n12358, new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364, new_n12365, new_n12366, new_n12367, new_n12368, new_n12369,
    new_n12370, new_n12371, new_n12372, new_n12373, new_n12374, new_n12375,
    new_n12376, new_n12377, new_n12378, new_n12379, new_n12380, new_n12381,
    new_n12382, new_n12383, new_n12384, new_n12385, new_n12386, new_n12387,
    new_n12388, new_n12389, new_n12390, new_n12391_1, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404,
    new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444_1, new_n12445,
    new_n12446, new_n12447, new_n12448, new_n12449, new_n12450, new_n12451,
    new_n12452, new_n12453, new_n12454, new_n12455, new_n12456, new_n12457,
    new_n12458, new_n12459, new_n12460, new_n12461, new_n12462, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467, new_n12468, new_n12469,
    new_n12470, new_n12471, new_n12480, new_n12481, new_n12482, new_n12483,
    new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489_1, new_n12490, new_n12491, new_n12492, new_n12493,
    new_n12494, new_n12495, new_n12496, new_n12497, new_n12498, new_n12499,
    new_n12500, new_n12501, new_n12502, new_n12503, new_n12504, new_n12505,
    new_n12506, new_n12507, new_n12508, new_n12509, new_n12510,
    new_n12511_1, new_n12512, new_n12513, new_n12514, new_n12515,
    new_n12516, new_n12517, new_n12518, new_n12519, new_n12520, new_n12521,
    new_n12522, new_n12523, new_n12524, new_n12525, new_n12526, new_n12527,
    new_n12528, new_n12529, new_n12530, new_n12531, new_n12532, new_n12533,
    new_n12534, new_n12535, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545,
    new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591_1, new_n12592,
    new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598,
    new_n12599, new_n12600, new_n12601, new_n12602, new_n12603, new_n12604,
    new_n12605, new_n12606, new_n12607, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620, new_n12621, new_n12622,
    new_n12623, new_n12624, new_n12625, new_n12626, new_n12627, new_n12628,
    new_n12629, new_n12630, new_n12631, new_n12632, new_n12633, new_n12634,
    new_n12635, new_n12636, new_n12637, new_n12638, new_n12639, new_n12640,
    new_n12641, new_n12642, new_n12643, new_n12644, new_n12645, new_n12646,
    new_n12647, new_n12648_1, new_n12649, new_n12650, new_n12651,
    new_n12652, new_n12653, new_n12654, new_n12655, new_n12656, new_n12657,
    new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663,
    new_n12664, new_n12665, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670, new_n12671, new_n12672, new_n12673, new_n12674, new_n12675,
    new_n12676, new_n12677, new_n12678, new_n12679, new_n12680, new_n12681,
    new_n12682, new_n12683, new_n12684, new_n12685, new_n12686, new_n12687,
    new_n12688, new_n12689, new_n12690, new_n12691, new_n12692, new_n12693,
    new_n12694, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699,
    new_n12700, new_n12701, new_n12702, new_n12703, new_n12704_1,
    new_n12705_1, new_n12706_1, new_n12707, new_n12708, new_n12709_1,
    new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715,
    new_n12716, new_n12717, new_n12718, new_n12719, new_n12720_1,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753_1, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777_1, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807_1,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12839, new_n12840, new_n12845, new_n12850, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925_1,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947_1, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13039, new_n13040,
    new_n13041, new_n13042, new_n13043, new_n13044, new_n13045, new_n13046,
    new_n13047, new_n13048, new_n13049, new_n13050, new_n13051, new_n13052,
    new_n13053, new_n13054, new_n13055, new_n13056, new_n13057, new_n13058,
    new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064,
    new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13072, new_n13073, new_n13074, new_n13075, new_n13076,
    new_n13077, new_n13078, new_n13079, new_n13080, new_n13081, new_n13082,
    new_n13083, new_n13084, new_n13085, new_n13086, new_n13087, new_n13088,
    new_n13089, new_n13090, new_n13091, new_n13092, new_n13093, new_n13094,
    new_n13095, new_n13096, new_n13097, new_n13098, new_n13099, new_n13100,
    new_n13101, new_n13102, new_n13103, new_n13104, new_n13105, new_n13106,
    new_n13107, new_n13108, new_n13109, new_n13110, new_n13111, new_n13112,
    new_n13113, new_n13114, new_n13115, new_n13116, new_n13117, new_n13118,
    new_n13119, new_n13120, new_n13121, new_n13122, new_n13123, new_n13124,
    new_n13125, new_n13126, new_n13127, new_n13128, new_n13129, new_n13130,
    new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137, new_n13138, new_n13139, new_n13140, new_n13141, new_n13142,
    new_n13143, new_n13144, new_n13145, new_n13146, new_n13147, new_n13148,
    new_n13149, new_n13150, new_n13151, new_n13152, new_n13153, new_n13154,
    new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160,
    new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166,
    new_n13167, new_n13168, new_n13169, new_n13170, new_n13171, new_n13172,
    new_n13173, new_n13174, new_n13175, new_n13176, new_n13177, new_n13178,
    new_n13179, new_n13180, new_n13181, new_n13182, new_n13183, new_n13184,
    new_n13185, new_n13186, new_n13187, new_n13188, new_n13189, new_n13190,
    new_n13191, new_n13192, new_n13193, new_n13194, new_n13195, new_n13196,
    new_n13197, new_n13198, new_n13199, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13204, new_n13205, new_n13206, new_n13207, new_n13208,
    new_n13209, new_n13210, new_n13211, new_n13212, new_n13213, new_n13214,
    new_n13215, new_n13216, new_n13217, new_n13218, new_n13219, new_n13220,
    new_n13221, new_n13222, new_n13223, new_n13224, new_n13236, new_n13237,
    new_n13238, new_n13239, new_n13240, new_n13241, new_n13242, new_n13243,
    new_n13244, new_n13245, new_n13246, new_n13247, new_n13248, new_n13249,
    new_n13250, new_n13251, new_n13252, new_n13253, new_n13254, new_n13255,
    new_n13256, new_n13257, new_n13258, new_n13259, new_n13260, new_n13261,
    new_n13262, new_n13263, new_n13264, new_n13265, new_n13266, new_n13267,
    new_n13268, new_n13269, new_n13270, new_n13271, new_n13272, new_n13273,
    new_n13274, new_n13275, new_n13276, new_n13277, new_n13278, new_n13279,
    new_n13280, new_n13281, new_n13282, new_n13283, new_n13284, new_n13285,
    new_n13286, new_n13287, new_n13288, new_n13289, new_n13290, new_n13291,
    new_n13292, new_n13293, new_n13294, new_n13295, new_n13296, new_n13297,
    new_n13298, new_n13299, new_n13300, new_n13301, new_n13302, new_n13303,
    new_n13304, new_n13305, new_n13306, new_n13307, new_n13308, new_n13309,
    new_n13310, new_n13311, new_n13312, new_n13313, new_n13314, new_n13315,
    new_n13316, new_n13317, new_n13318, new_n13319, new_n13320, new_n13321,
    new_n13322, new_n13323, new_n13324, new_n13325, new_n13326, new_n13327,
    new_n13328, new_n13329, new_n13330, new_n13331, new_n13332, new_n13333,
    new_n13334, new_n13335, new_n13336, new_n13337, new_n13338, new_n13339,
    new_n13340, new_n13341, new_n13342, new_n13343, new_n13344, new_n13345,
    new_n13346, new_n13347, new_n13348, new_n13349, new_n13350, new_n13351,
    new_n13352, new_n13353, new_n13354, new_n13355, new_n13356, new_n13357,
    new_n13358, new_n13359, new_n13360, new_n13361, new_n13362, new_n13363,
    new_n13364, new_n13365, new_n13366, new_n13367, new_n13368, new_n13369,
    new_n13370, new_n13371, new_n13372, new_n13373, new_n13374, new_n13375,
    new_n13376, new_n13377, new_n13378, new_n13379, new_n13380, new_n13381,
    new_n13382, new_n13383, new_n13384, new_n13385, new_n13386, new_n13387,
    new_n13388, new_n13389, new_n13390, new_n13391, new_n13392, new_n13393,
    new_n13394, new_n13395, new_n13396, new_n13397, new_n13398, new_n13399,
    new_n13400, new_n13401, new_n13402, new_n13403, new_n13404, new_n13405,
    new_n13406, new_n13407, new_n13408, new_n13409, new_n13410, new_n13411,
    new_n13412, new_n13413, new_n13414, new_n13415, new_n13416, new_n13417,
    new_n13424, new_n13425, new_n13432, new_n13433, new_n13434, new_n13435,
    new_n13436, new_n13437, new_n13438, new_n13439, new_n13440, new_n13441,
    new_n13442, new_n13443, new_n13444, new_n13445, new_n13446, new_n13447,
    new_n13448, new_n13449, new_n13450, new_n13451, new_n13452, new_n13453,
    new_n13454, new_n13455, new_n13456, new_n13457, new_n13458, new_n13459,
    new_n13460, new_n13461, new_n13462, new_n13463, new_n13464, new_n13465,
    new_n13466, new_n13467, new_n13468, new_n13469, new_n13470, new_n13471,
    new_n13472, new_n13473, new_n13474, new_n13475, new_n13476, new_n13477,
    new_n13478, new_n13479, new_n13480, new_n13481, new_n13482, new_n13483,
    new_n13484, new_n13485, new_n13486, new_n13487, new_n13488, new_n13489,
    new_n13490, new_n13491, new_n13492, new_n13493, new_n13494, new_n13495,
    new_n13496, new_n13497, new_n13498, new_n13499, new_n13500, new_n13501,
    new_n13502, new_n13503, new_n13504, new_n13505, new_n13506, new_n13507,
    new_n13508, new_n13509, new_n13510, new_n13511, new_n13512, new_n13513,
    new_n13514, new_n13515, new_n13516, new_n13517, new_n13518, new_n13519,
    new_n13520, new_n13521, new_n13522, new_n13523, new_n13524, new_n13525,
    new_n13526, new_n13527, new_n13528, new_n13529, new_n13530, new_n13531,
    new_n13532, new_n13533, new_n13534, new_n13535, new_n13536, new_n13537,
    new_n13538, new_n13539, new_n13540, new_n13541, new_n13542, new_n13543,
    new_n13544, new_n13545, new_n13546, new_n13547, new_n13548, new_n13549,
    new_n13550, new_n13551, new_n13552, new_n13553, new_n13554, new_n13555,
    new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561,
    new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13625;
not_1  g00000(n6038, new_n377);
not_1  g00001(n6687, new_n378);
nor_1  g00002(new_n378, new_n377, new_n379);
not_1  g00003(new_n379, new_n380);
not_1  g00004(n7354, new_n381_1);
not_1  g00005(n8336, new_n382);
nor_1  g00006(new_n382, new_n381_1, new_n383);
not_1  g00007(n8028, new_n384);
not_1  g00008(n11222, new_n385);
nor_1  g00009(new_n385, new_n384, new_n386);
not_1  g00010(new_n386, new_n387);
nand_1 g00011(n12069, n1564, new_n388);
nor_1  g00012(new_n388, new_n387, new_n389);
not_1  g00013(new_n389, new_n390);
nand_1 g00014(new_n388, new_n387, new_n391);
nand_1 g00015(new_n391, new_n390, new_n392);
xnor_1 g00016(new_n392, new_n383, new_n393);
xnor_1 g00017(new_n393, new_n380, n112);
not_1  g00018(n4312, new_n395);
not_1  g00019(n12720, new_n396);
nor_1  g00020(new_n396, new_n395, new_n397_1);
not_1  g00021(new_n397_1, new_n398);
nand_1 g00022(n12025, n6038, new_n399);
nand_1 g00023(n12705, n2509, new_n400);
nand_1 g00024(new_n400, new_n399, new_n401);
nor_1  g00025(new_n400, new_n399, new_n402);
not_1  g00026(new_n402, new_n403);
nand_1 g00027(new_n403, new_n401, new_n404);
nor_1  g00028(new_n404, new_n398, new_n405_1);
not_1  g00029(new_n405_1, new_n406);
nand_1 g00030(new_n404, new_n398, new_n407);
nand_1 g00031(new_n407, new_n406, new_n408);
nand_1 g00032(n12705, n6038, new_n409);
nand_1 g00033(n12720, n1097, new_n410);
nand_1 g00034(new_n410, new_n409, new_n411);
not_1  g00035(new_n411, new_n412);
not_1  g00036(n2509, new_n413);
nor_1  g00037(new_n395, new_n413, new_n414);
xnor_1 g00038(new_n410, new_n409, new_n415);
nor_1  g00039(new_n415, new_n414, new_n416);
nor_1  g00040(new_n416, new_n412, new_n417);
xnor_1 g00041(new_n417, new_n408, new_n418);
not_1  g00042(n1097, new_n419);
not_1  g00043(n2508, new_n420);
nor_1  g00044(new_n420, new_n419, new_n421);
not_1  g00045(new_n421, new_n422);
not_1  g00046(n2585, new_n423);
not_1  g00047(n5964, new_n424);
nor_1  g00048(new_n424, new_n423, new_n425);
not_1  g00049(new_n425, new_n426);
nand_1 g00050(new_n426, new_n422, new_n427);
nor_1  g00051(new_n426, new_n422, new_n428);
not_1  g00052(new_n428, new_n429);
nand_1 g00053(new_n429, new_n427, new_n430);
xnor_1 g00054(new_n430, new_n418, new_n431);
nor_1  g00055(new_n424, new_n420, new_n432);
not_1  g00056(new_n432, new_n433);
not_1  g00057(new_n414, new_n434);
xnor_1 g00058(new_n415, new_n434, new_n435);
nand_1 g00059(new_n435, new_n433, new_n436);
not_1  g00060(new_n436, new_n437);
xnor_1 g00061(new_n435, new_n433, new_n438);
nor_1  g00062(new_n377, new_n395, new_n439);
not_1  g00063(new_n439, new_n440);
nor_1  g00064(new_n396, new_n424, new_n441);
not_1  g00065(new_n441, new_n442);
nand_1 g00066(new_n442, new_n440, new_n443);
not_1  g00067(new_n443, new_n444);
nor_1  g00068(new_n442, new_n440, new_n445);
nor_1  g00069(new_n413, new_n419, new_n446);
nor_1  g00070(new_n446, new_n445, new_n447_1);
nor_1  g00071(new_n447_1, new_n444, new_n448);
nor_1  g00072(new_n448, new_n438, new_n449);
nor_1  g00073(new_n449, new_n437, new_n450);
nand_1 g00074(new_n450, new_n431, new_n451);
not_1  g00075(new_n451, new_n452);
nor_1  g00076(new_n450, new_n431, new_n453);
nor_1  g00077(new_n453, new_n452, new_n454);
not_1  g00078(new_n454, new_n455);
not_1  g00079(n5305, new_n456);
nor_1  g00080(new_n456, new_n423, new_n457);
xnor_1 g00081(new_n448, new_n438, new_n458);
nor_1  g00082(new_n458, new_n457, new_n459);
not_1  g00083(new_n459, new_n460);
nand_1 g00084(new_n458, new_n457, new_n461);
nand_1 g00085(new_n461, new_n460, new_n462);
not_1  g00086(new_n462, new_n463);
nor_1  g00087(new_n456, new_n420, new_n464);
not_1  g00088(new_n464, new_n465);
nor_1  g00089(new_n377, new_n419, new_n466);
not_1  g00090(new_n466, new_n467);
nor_1  g00091(new_n396, new_n456, new_n468);
not_1  g00092(new_n468, new_n469);
nor_1  g00093(new_n469, new_n467, new_n470);
nand_1 g00094(new_n469, new_n467, new_n471);
not_1  g00095(new_n471, new_n472);
nor_1  g00096(new_n424, new_n413, new_n473);
not_1  g00097(new_n473, new_n474);
nor_1  g00098(new_n474, new_n472, new_n475);
nor_1  g00099(new_n475, new_n470, new_n476);
nor_1  g00100(new_n476, new_n465, new_n477);
xnor_1 g00101(new_n476, new_n464, new_n478);
not_1  g00102(new_n445, new_n479);
nand_1 g00103(new_n479, new_n443, new_n480);
xnor_1 g00104(new_n480, new_n446, new_n481);
nand_1 g00105(new_n481, new_n478, new_n482);
not_1  g00106(new_n482, new_n483);
nor_1  g00107(new_n483, new_n477, new_n484);
nand_1 g00108(new_n484, new_n463, new_n485);
nand_1 g00109(new_n485, new_n460, new_n486);
nor_1  g00110(new_n486, new_n455, new_n487);
not_1  g00111(new_n487, new_n488);
not_1  g00112(new_n408, new_n489);
nand_1 g00113(new_n417, new_n489, new_n490);
nand_1 g00114(new_n490, new_n406, new_n491);
not_1  g00115(n4005, new_n492);
nor_1  g00116(new_n424, new_n492, new_n493);
nor_1  g00117(new_n423, new_n419, new_n494);
not_1  g00118(new_n494, new_n495);
not_1  g00119(n12706, new_n496);
nor_1  g00120(new_n496, new_n456, new_n497);
not_1  g00121(new_n497, new_n498);
nand_1 g00122(new_n498, new_n495, new_n499);
nand_1 g00123(new_n497, new_n494, new_n500);
nand_1 g00124(new_n500, new_n499, new_n501);
xnor_1 g00125(new_n501, new_n493, new_n502);
nand_1 g00126(new_n502, new_n491, new_n503_1);
not_1  g00127(new_n491, new_n504);
not_1  g00128(new_n502, new_n505);
nand_1 g00129(new_n505, new_n504, new_n506);
nand_1 g00130(new_n506, new_n503_1, new_n507);
not_1  g00131(new_n507, new_n508);
nand_1 g00132(n4312, n2508, new_n509);
xnor_1 g00133(new_n509, new_n402, new_n510);
not_1  g00134(n12025, new_n511);
nor_1  g00135(new_n511, new_n413, new_n512);
nand_1 g00136(n12720, n12705, new_n513);
nand_1 g00137(n11257, n6038, new_n514);
xnor_1 g00138(new_n514, new_n513, new_n515);
xor_1  g00139(new_n515, new_n512, new_n516);
xnor_1 g00140(new_n516, new_n510, new_n517);
not_1  g00141(new_n517, new_n518);
nand_1 g00142(new_n518, new_n508, new_n519);
nand_1 g00143(new_n517, new_n507, new_n520);
nand_1 g00144(new_n520, new_n519, new_n521_1);
not_1  g00145(new_n521_1, new_n522);
not_1  g00146(new_n430, new_n523);
nand_1 g00147(new_n523, new_n418, new_n524);
nand_1 g00148(new_n452, new_n428, new_n525);
nand_1 g00149(new_n451, new_n429, new_n526);
nand_1 g00150(new_n526, new_n525, new_n527);
nand_1 g00151(new_n527, new_n524, new_n528);
xnor_1 g00152(new_n528, new_n522, new_n529);
xnor_1 g00153(new_n529, new_n488, new_n530);
nor_1  g00154(new_n456, new_n492, new_n531);
nand_1 g00155(new_n486, new_n455, new_n532);
nand_1 g00156(new_n532, new_n488, new_n533_1);
not_1  g00157(new_n533_1, new_n534);
nand_1 g00158(new_n534, new_n531, new_n535);
not_1  g00159(new_n531, new_n536);
nand_1 g00160(new_n533_1, new_n536, new_n537);
nor_1  g00161(new_n481, new_n478, new_n538);
nor_1  g00162(new_n538, new_n483, new_n539);
nor_1  g00163(new_n472, new_n470, new_n540);
nor_1  g00164(new_n377, new_n424, new_n541);
nor_1  g00165(new_n456, new_n413, new_n542);
nand_1 g00166(new_n542, new_n541, new_n543);
nor_1  g00167(new_n543, new_n540, new_n544);
nand_1 g00168(new_n544, new_n539, new_n545);
xnor_1 g00169(new_n484, new_n462, new_n546);
nor_1  g00170(new_n546, new_n545, new_n547);
nand_1 g00171(new_n547, new_n537, new_n548);
nand_1 g00172(new_n548, new_n535, new_n549);
xnor_1 g00173(new_n549, new_n530, new_n550);
not_1  g00174(n5105, new_n551);
not_1  g00175(n8759, new_n552);
nor_1  g00176(new_n552, new_n551, new_n553);
not_1  g00177(n12299, new_n554);
nor_1  g00178(new_n554, new_n381_1, new_n555);
not_1  g00179(new_n555, new_n556);
not_1  g00180(n1209, new_n557);
nor_1  g00181(new_n552, new_n557, new_n558);
not_1  g00182(new_n558, new_n559);
nand_1 g00183(new_n559, new_n556, new_n560);
not_1  g00184(new_n560, new_n561);
nor_1  g00185(new_n559, new_n556, new_n562);
not_1  g00186(n6776, new_n563);
not_1  g00187(n7500, new_n564);
nor_1  g00188(new_n564, new_n563, new_n565);
nor_1  g00189(new_n565, new_n562, new_n566);
nor_1  g00190(new_n566, new_n561, new_n567);
xnor_1 g00191(new_n567, new_n553, new_n568);
nor_1  g00192(new_n554, new_n564, new_n569);
nand_1 g00193(n7436, n7354, new_n570);
nand_1 g00194(n6776, n1209, new_n571);
xnor_1 g00195(new_n571, new_n570, new_n572);
xnor_1 g00196(new_n572, new_n569, new_n573);
not_1  g00197(new_n573, new_n574);
nor_1  g00198(new_n574, new_n568, new_n575);
not_1  g00199(new_n575, new_n576);
nand_1 g00200(new_n574, new_n568, new_n577);
nand_1 g00201(new_n577, new_n576, new_n578);
not_1  g00202(new_n578, new_n579);
not_1  g00203(new_n565, new_n580);
nor_1  g00204(new_n552, new_n381_1, new_n581);
nor_1  g00205(new_n581, new_n580, new_n582);
nor_1  g00206(new_n582, new_n560, new_n583);
nor_1  g00207(new_n583, new_n562, new_n584);
nor_1  g00208(new_n584, new_n580, new_n585);
nand_1 g00209(new_n585, new_n579, new_n586);
not_1  g00210(new_n586, new_n587);
not_1  g00211(n4141, new_n588);
nor_1  g00212(new_n552, new_n588, new_n589);
nor_1  g00213(new_n563, new_n551, new_n590);
nand_1 g00214(new_n571, new_n570, new_n591);
not_1  g00215(new_n591, new_n592);
nor_1  g00216(new_n572, new_n569, new_n593);
nor_1  g00217(new_n593, new_n592, new_n594);
nand_1 g00218(new_n594, new_n590, new_n595);
not_1  g00219(new_n595, new_n596);
nor_1  g00220(new_n594, new_n590, new_n597);
nor_1  g00221(new_n597, new_n596, new_n598);
not_1  g00222(n7436, new_n599);
nor_1  g00223(new_n564, new_n599, new_n600);
nand_1 g00224(n12299, n1209, new_n601);
nand_1 g00225(n8276, n7354, new_n602);
xnor_1 g00226(new_n602, new_n601, new_n603);
xnor_1 g00227(new_n603, new_n600, new_n604);
nand_1 g00228(new_n604, new_n598, new_n605);
not_1  g00229(new_n605, new_n606);
nor_1  g00230(new_n604, new_n598, new_n607);
nor_1  g00231(new_n607, new_n606, new_n608);
nand_1 g00232(new_n608, new_n589, new_n609);
not_1  g00233(new_n609, new_n610);
nor_1  g00234(new_n608, new_n589, new_n611);
nor_1  g00235(new_n611, new_n610, new_n612);
nand_1 g00236(new_n567, new_n553, new_n613);
nand_1 g00237(new_n576, new_n613, new_n614);
nand_1 g00238(new_n614, new_n612, new_n615_1);
not_1  g00239(new_n615_1, new_n616);
nor_1  g00240(new_n614, new_n612, new_n617);
nor_1  g00241(new_n617, new_n616, new_n618);
nand_1 g00242(new_n618, new_n587, new_n619);
not_1  g00243(new_n619, new_n620);
not_1  g00244(n4928, new_n621);
nor_1  g00245(new_n552, new_n621, new_n622);
not_1  g00246(new_n622, new_n623);
nor_1  g00247(new_n599, new_n557, new_n624);
not_1  g00248(new_n624, new_n625);
nand_1 g00249(n8276, n7500, new_n626);
nand_1 g00250(n9241, n7354, new_n627);
xnor_1 g00251(new_n627, new_n626, new_n628);
xnor_1 g00252(new_n628, new_n625, new_n629);
not_1  g00253(new_n629, new_n630);
nand_1 g00254(new_n602, new_n601, new_n631);
not_1  g00255(new_n631, new_n632);
nor_1  g00256(new_n603, new_n600, new_n633);
nor_1  g00257(new_n633, new_n632, new_n634);
nand_1 g00258(new_n634, new_n630, new_n635);
not_1  g00259(new_n635, new_n636);
nor_1  g00260(new_n634, new_n630, new_n637);
nor_1  g00261(new_n637, new_n636, new_n638);
nor_1  g00262(new_n563, new_n588, new_n639);
not_1  g00263(new_n639, new_n640);
nor_1  g00264(new_n554, new_n551, new_n641);
not_1  g00265(new_n641, new_n642);
nand_1 g00266(new_n642, new_n640, new_n643);
nor_1  g00267(new_n642, new_n640, new_n644);
not_1  g00268(new_n644, new_n645);
nand_1 g00269(new_n645, new_n643, new_n646);
xnor_1 g00270(new_n646, new_n638, new_n647);
nand_1 g00271(new_n605, new_n595, new_n648);
nand_1 g00272(new_n648, new_n647, new_n649);
not_1  g00273(new_n649, new_n650);
nor_1  g00274(new_n648, new_n647, new_n651);
nor_1  g00275(new_n651, new_n650, new_n652);
nand_1 g00276(new_n615_1, new_n609, new_n653);
nand_1 g00277(new_n653, new_n652, new_n654);
not_1  g00278(new_n654, new_n655);
nor_1  g00279(new_n653, new_n652, new_n656);
nor_1  g00280(new_n656, new_n655, new_n657);
xnor_1 g00281(new_n657, new_n623, new_n658_1);
xnor_1 g00282(new_n658_1, new_n620, new_n659);
nor_1  g00283(new_n618, new_n587, new_n660);
nor_1  g00284(new_n660, new_n620, new_n661);
not_1  g00285(new_n661, new_n662);
nor_1  g00286(new_n585, new_n579, new_n663);
nor_1  g00287(new_n663, new_n587, new_n664);
not_1  g00288(new_n664, new_n665);
not_1  g00289(new_n581, new_n666);
not_1  g00290(n1564, new_n667);
not_1  g00291(n5331, new_n668);
nor_1  g00292(new_n668, new_n667, new_n669);
nand_1 g00293(n8028, n7965, new_n670);
not_1  g00294(new_n670, new_n671_1);
nand_1 g00295(new_n671_1, new_n669, new_n672);
not_1  g00296(new_n669, new_n673);
nand_1 g00297(new_n670, new_n673, new_n674);
nand_1 g00298(new_n674, new_n672, new_n675);
nor_1  g00299(new_n675, new_n666, new_n676);
not_1  g00300(new_n676, new_n677);
nand_1 g00301(n7354, n6776, new_n678);
nand_1 g00302(n8759, n7500, new_n679);
xnor_1 g00303(new_n679, new_n678, new_n680);
nand_1 g00304(new_n680, new_n677, new_n681);
nand_1 g00305(n5331, n1512, new_n682);
nand_1 g00306(n8476, n1564, new_n683);
xnor_1 g00307(new_n683, new_n682, new_n684);
xnor_1 g00308(new_n684, new_n672, new_n685);
nand_1 g00309(n8028, n7388, new_n686);
nand_1 g00310(n10848, n7965, new_n687);
xnor_1 g00311(new_n687, new_n686, new_n688);
xnor_1 g00312(new_n688, new_n685, new_n689);
xnor_1 g00313(new_n680, new_n676, new_n690);
nand_1 g00314(new_n690, new_n689, new_n691);
nand_1 g00315(new_n691, new_n681, new_n692);
nand_1 g00316(new_n582, new_n560, new_n693);
nand_1 g00317(new_n693, new_n584, new_n694);
nand_1 g00318(new_n694, new_n692, new_n695);
not_1  g00319(n7388, new_n696);
not_1  g00320(n10848, new_n697);
nor_1  g00321(new_n697, new_n696, new_n698);
nand_1 g00322(new_n698, new_n670, new_n699);
not_1  g00323(new_n699, new_n700);
nand_1 g00324(n11892, n8028, new_n701);
nand_1 g00325(n7965, n1980, new_n702);
nand_1 g00326(new_n702, new_n701, new_n703);
not_1  g00327(new_n703, new_n704);
nand_1 g00328(n11892, n1980, new_n705);
nor_1  g00329(new_n705, new_n670, new_n706);
nor_1  g00330(new_n706, new_n704, new_n707);
nor_1  g00331(new_n707, new_n700, new_n708);
nor_1  g00332(new_n704, new_n699, new_n709);
nor_1  g00333(new_n709, new_n708, new_n710);
not_1  g00334(n1512, new_n711);
not_1  g00335(n8476, new_n712);
nor_1  g00336(new_n712, new_n711, new_n713);
nand_1 g00337(new_n713, new_n673, new_n714);
nand_1 g00338(n2530, n1564, new_n715);
nand_1 g00339(n5331, n533, new_n716);
nand_1 g00340(new_n716, new_n715, new_n717);
not_1  g00341(new_n717, new_n718);
nand_1 g00342(new_n718, new_n714, new_n719);
nor_1  g00343(new_n716, new_n715, new_n720);
not_1  g00344(new_n720, new_n721);
nand_1 g00345(new_n721, new_n719, new_n722);
nor_1  g00346(new_n718, new_n714, new_n723);
nor_1  g00347(new_n723, new_n722, new_n724);
xnor_1 g00348(new_n724, new_n710, new_n725);
nor_1  g00349(new_n684, new_n672, new_n726);
nor_1  g00350(new_n688, new_n685, new_n727);
nor_1  g00351(new_n727, new_n726, new_n728);
xnor_1 g00352(new_n728, new_n725, new_n729);
not_1  g00353(new_n694, new_n730);
xnor_1 g00354(new_n730, new_n692, new_n731);
nand_1 g00355(new_n731, new_n729, new_n732);
nand_1 g00356(new_n732, new_n695, new_n733);
nand_1 g00357(new_n733, new_n665, new_n734);
not_1  g00358(n2802, new_n735);
nor_1  g00359(new_n668, new_n735, new_n736);
nor_1  g00360(new_n720, new_n713, new_n737);
nor_1  g00361(new_n737, new_n718, new_n738);
xnor_1 g00362(new_n738, new_n736, new_n739);
not_1  g00363(n2530, new_n740);
nor_1  g00364(new_n740, new_n711, new_n741);
not_1  g00365(new_n741, new_n742);
nand_1 g00366(n12648, n1564, new_n743);
nand_1 g00367(n8476, n533, new_n744);
xnor_1 g00368(new_n744, new_n743, new_n745);
xnor_1 g00369(new_n745, new_n742, new_n746);
xnor_1 g00370(new_n746, new_n739, new_n747);
nand_1 g00371(new_n722, new_n713, new_n748);
nand_1 g00372(new_n748, new_n747, new_n749);
nor_1  g00373(new_n748, new_n747, new_n750);
not_1  g00374(new_n750, new_n751);
nand_1 g00375(new_n751, new_n749, new_n752);
not_1  g00376(n7294, new_n753_1);
not_1  g00377(n7965, new_n754);
nor_1  g00378(new_n754, new_n753_1, new_n755);
nor_1  g00379(new_n706, new_n698, new_n756);
nor_1  g00380(new_n756, new_n704, new_n757);
nand_1 g00381(new_n757, new_n755, new_n758);
not_1  g00382(new_n758, new_n759);
nor_1  g00383(new_n757, new_n755, new_n760);
nor_1  g00384(new_n760, new_n759, new_n761);
not_1  g00385(n11892, new_n762);
nor_1  g00386(new_n762, new_n697, new_n763);
not_1  g00387(n1980, new_n764);
nor_1  g00388(new_n696, new_n764, new_n765);
not_1  g00389(new_n765, new_n766);
not_1  g00390(n2393, new_n767);
nor_1  g00391(new_n384, new_n767, new_n768);
not_1  g00392(new_n768, new_n769);
nand_1 g00393(new_n769, new_n766, new_n770);
nor_1  g00394(new_n769, new_n766, new_n771);
not_1  g00395(new_n771, new_n772);
nand_1 g00396(new_n772, new_n770, new_n773);
xnor_1 g00397(new_n773, new_n763, new_n774);
xnor_1 g00398(new_n774, new_n761, new_n775);
nand_1 g00399(new_n708, new_n698, new_n776);
xnor_1 g00400(new_n776, new_n775, new_n777);
xnor_1 g00401(new_n777, new_n752, new_n778);
and_1  g00402(new_n724, new_n710, new_n779);
nor_1  g00403(new_n728, new_n725, new_n780);
nor_1  g00404(new_n780, new_n779, new_n781);
xnor_1 g00405(new_n781, new_n778, new_n782);
xnor_1 g00406(new_n733, new_n664, new_n783_1);
nand_1 g00407(new_n783_1, new_n782, new_n784);
nand_1 g00408(new_n784, new_n734, new_n785);
nand_1 g00409(new_n785, new_n662, new_n786);
nor_1  g00410(new_n776, new_n775, new_n787);
nand_1 g00411(new_n774, new_n761, new_n788);
nand_1 g00412(new_n788, new_n758, new_n789);
not_1  g00413(n12704, new_n790);
nor_1  g00414(new_n790, new_n754, new_n791);
not_1  g00415(new_n791, new_n792);
nor_1  g00416(new_n696, new_n753_1, new_n793);
not_1  g00417(new_n770, new_n794);
nor_1  g00418(new_n771, new_n763, new_n795);
nor_1  g00419(new_n795, new_n794, new_n796);
nand_1 g00420(new_n796, new_n793, new_n797);
not_1  g00421(new_n797, new_n798);
nor_1  g00422(new_n796, new_n793, new_n799);
nor_1  g00423(new_n799, new_n798, new_n800);
nor_1  g00424(new_n697, new_n767, new_n801);
not_1  g00425(n5860, new_n802);
nor_1  g00426(new_n384, new_n802, new_n803);
not_1  g00427(new_n803, new_n804);
nand_1 g00428(new_n804, new_n705, new_n805);
not_1  g00429(new_n705, new_n806_1);
nand_1 g00430(new_n803, new_n806_1, new_n807);
nand_1 g00431(new_n807, new_n805, new_n808);
xnor_1 g00432(new_n808, new_n801, new_n809);
nand_1 g00433(new_n809, new_n800, new_n810);
not_1  g00434(new_n810, new_n811);
nor_1  g00435(new_n809, new_n800, new_n812);
nor_1  g00436(new_n812, new_n811, new_n813);
not_1  g00437(new_n813, new_n814);
nand_1 g00438(new_n814, new_n792, new_n815);
nand_1 g00439(new_n813, new_n791, new_n816);
nand_1 g00440(new_n816, new_n815, new_n817);
xnor_1 g00441(new_n817, new_n789, new_n818);
xnor_1 g00442(new_n818, new_n787, new_n819);
not_1  g00443(n6806, new_n820);
nor_1  g00444(new_n820, new_n668, new_n821);
nor_1  g00445(new_n712, new_n735, new_n822);
not_1  g00446(new_n822, new_n823);
nand_1 g00447(new_n744, new_n743, new_n824);
not_1  g00448(new_n824, new_n825);
nor_1  g00449(new_n745, new_n741, new_n826);
nor_1  g00450(new_n826, new_n825, new_n827);
xnor_1 g00451(new_n827, new_n823, new_n828);
not_1  g00452(n12648, new_n829);
nor_1  g00453(new_n829, new_n711, new_n830);
not_1  g00454(new_n830, new_n831);
nand_1 g00455(n2530, n533, new_n832);
nand_1 g00456(n10545, n1564, new_n833);
xnor_1 g00457(new_n833, new_n832, new_n834);
xnor_1 g00458(new_n834, new_n831, new_n835);
xnor_1 g00459(new_n835, new_n828, new_n836);
nand_1 g00460(new_n836, new_n821, new_n837_1);
not_1  g00461(new_n837_1, new_n838);
nor_1  g00462(new_n836, new_n821, new_n839);
nor_1  g00463(new_n839, new_n838, new_n840);
nand_1 g00464(new_n738, new_n736, new_n841);
not_1  g00465(new_n841, new_n842);
nor_1  g00466(new_n746, new_n739, new_n843);
nor_1  g00467(new_n843, new_n842, new_n844_1);
xnor_1 g00468(new_n844_1, new_n840, new_n845);
nand_1 g00469(new_n845, new_n750, new_n846);
not_1  g00470(new_n846, new_n847);
nor_1  g00471(new_n845, new_n750, new_n848);
nor_1  g00472(new_n848, new_n847, new_n849);
nand_1 g00473(new_n777, new_n752, new_n850);
not_1  g00474(new_n778, new_n851);
nand_1 g00475(new_n781, new_n851, new_n852);
nand_1 g00476(new_n852, new_n850, new_n853);
xnor_1 g00477(new_n853, new_n849, new_n854);
nor_1  g00478(new_n854, new_n819, new_n855);
nand_1 g00479(new_n854, new_n819, new_n856);
not_1  g00480(new_n856, new_n857);
nor_1  g00481(new_n857, new_n855, new_n858);
xnor_1 g00482(new_n785, new_n661, new_n859);
nand_1 g00483(new_n859, new_n858, new_n860);
nand_1 g00484(new_n860, new_n786, new_n861);
xnor_1 g00485(new_n861, new_n659, new_n862);
not_1  g00486(new_n849, new_n863);
nand_1 g00487(new_n853, new_n863, new_n864);
nand_1 g00488(new_n856, new_n864, new_n865);
not_1  g00489(new_n865, new_n866);
not_1  g00490(n5069, new_n867);
nor_1  g00491(new_n668, new_n867, new_n868);
not_1  g00492(n533, new_n869);
nor_1  g00493(new_n829, new_n869, new_n870);
not_1  g00494(new_n870, new_n871);
nand_1 g00495(n10545, n1512, new_n872);
nand_1 g00496(n7690, n1564, new_n873);
xnor_1 g00497(new_n873, new_n872, new_n874);
xnor_1 g00498(new_n874, new_n871, new_n875);
not_1  g00499(new_n875, new_n876);
nand_1 g00500(new_n833, new_n832, new_n877);
not_1  g00501(new_n877, new_n878);
nor_1  g00502(new_n834, new_n830, new_n879);
nor_1  g00503(new_n879, new_n878, new_n880);
nand_1 g00504(new_n880, new_n876, new_n881);
not_1  g00505(new_n881, new_n882);
nor_1  g00506(new_n880, new_n876, new_n883);
nor_1  g00507(new_n883, new_n882, new_n884);
nand_1 g00508(n8476, n6806, new_n885);
nand_1 g00509(n2802, n2530, new_n886);
nand_1 g00510(new_n886, new_n885, new_n887);
nor_1  g00511(new_n886, new_n885, new_n888);
not_1  g00512(new_n888, new_n889);
nand_1 g00513(new_n889, new_n887, new_n890);
xnor_1 g00514(new_n890, new_n884, new_n891);
nand_1 g00515(new_n827, new_n822, new_n892);
not_1  g00516(new_n835, new_n893);
nand_1 g00517(new_n893, new_n828, new_n894);
nand_1 g00518(new_n894, new_n892, new_n895);
nand_1 g00519(new_n895, new_n891, new_n896);
not_1  g00520(new_n896, new_n897);
nor_1  g00521(new_n895, new_n891, new_n898);
nor_1  g00522(new_n898, new_n897, new_n899);
not_1  g00523(new_n844_1, new_n900);
nand_1 g00524(new_n900, new_n840, new_n901);
nand_1 g00525(new_n901, new_n837_1, new_n902);
xnor_1 g00526(new_n902, new_n899, new_n903);
not_1  g00527(new_n903, new_n904);
nand_1 g00528(new_n904, new_n868, new_n905);
not_1  g00529(new_n868, new_n906);
nand_1 g00530(new_n903, new_n906, new_n907);
nand_1 g00531(new_n907, new_n905, new_n908);
xnor_1 g00532(new_n908, new_n846, new_n909);
not_1  g00533(new_n909, new_n910);
nand_1 g00534(new_n910, new_n866, new_n911_1);
nand_1 g00535(new_n909, new_n865, new_n912);
nand_1 g00536(new_n912, new_n911_1, new_n913);
nand_1 g00537(new_n818, new_n787, new_n914);
not_1  g00538(n5814, new_n915);
nor_1  g00539(new_n754, new_n915, new_n916);
nor_1  g00540(new_n767, new_n764, new_n917);
not_1  g00541(new_n917, new_n918);
nand_1 g00542(n8028, n3986, new_n919);
nand_1 g00543(n10848, n5860, new_n920);
nand_1 g00544(new_n920, new_n919, new_n921);
nor_1  g00545(new_n920, new_n919, new_n922);
not_1  g00546(new_n922, new_n923);
nand_1 g00547(new_n923, new_n921, new_n924);
nor_1  g00548(new_n924, new_n918, new_n925);
not_1  g00549(new_n925, new_n926);
nand_1 g00550(new_n924, new_n918, new_n927);
nand_1 g00551(new_n927, new_n926, new_n928);
not_1  g00552(new_n928, new_n929);
not_1  g00553(new_n805, new_n930);
not_1  g00554(new_n807, new_n931);
nor_1  g00555(new_n931, new_n801, new_n932);
nor_1  g00556(new_n932, new_n930, new_n933);
xnor_1 g00557(new_n933, new_n929, new_n934);
nor_1  g00558(new_n790, new_n696, new_n935);
not_1  g00559(new_n935, new_n936);
nor_1  g00560(new_n762, new_n753_1, new_n937);
not_1  g00561(new_n937, new_n938);
nand_1 g00562(new_n938, new_n936, new_n939);
nor_1  g00563(new_n938, new_n936, new_n940);
not_1  g00564(new_n940, new_n941);
nand_1 g00565(new_n941, new_n939, new_n942);
not_1  g00566(new_n942, new_n943);
xnor_1 g00567(new_n943, new_n934, new_n944);
nor_1  g00568(new_n811, new_n798, new_n945);
xnor_1 g00569(new_n945, new_n944, new_n946);
not_1  g00570(new_n789, new_n947);
nand_1 g00571(new_n816, new_n947, new_n948);
nand_1 g00572(new_n948, new_n815, new_n949);
xnor_1 g00573(new_n949, new_n946, new_n950);
xnor_1 g00574(new_n950, new_n916, new_n951);
xnor_1 g00575(new_n951, new_n914, new_n952);
xnor_1 g00576(new_n952, new_n913, new_n953);
xnor_1 g00577(new_n953, new_n862, new_n954);
not_1  g00578(new_n954, new_n955);
nand_1 g00579(new_n537, new_n535, new_n956);
xnor_1 g00580(new_n956, new_n547, new_n957);
nand_1 g00581(new_n957, new_n955, new_n958);
xor_1  g00582(new_n546, new_n545, new_n959);
not_1  g00583(new_n859, new_n960);
xnor_1 g00584(new_n960, new_n858, new_n961);
not_1  g00585(new_n961, new_n962);
nand_1 g00586(new_n962, new_n959, new_n963);
xnor_1 g00587(new_n961, new_n959, new_n964);
xor_1  g00588(new_n544, new_n539, new_n965);
xnor_1 g00589(new_n783_1, new_n782, new_n966);
nand_1 g00590(new_n966, new_n965, new_n967);
xnor_1 g00591(new_n731, new_n729, new_n968);
nor_1  g00592(new_n377, new_n456, new_n969);
nor_1  g00593(new_n969, new_n474, new_n970);
nor_1  g00594(new_n970, new_n540, new_n971);
not_1  g00595(new_n969, new_n972);
and_1  g00596(new_n972, new_n475, new_n973);
nor_1  g00597(new_n973, new_n971, new_n974);
nor_1  g00598(new_n974, new_n968, new_n975);
xnor_1 g00599(new_n974, new_n968, new_n976);
xnor_1 g00600(new_n675, new_n581, new_n977);
nand_1 g00601(new_n977, new_n969, new_n978);
not_1  g00602(new_n541, new_n979);
xnor_1 g00603(new_n542, new_n979, new_n980);
not_1  g00604(new_n980, new_n981);
nand_1 g00605(new_n981, new_n978, new_n982);
not_1  g00606(new_n982, new_n983);
xor_1  g00607(new_n690, new_n689, new_n984);
not_1  g00608(new_n984, new_n985);
nor_1  g00609(new_n981, new_n978, new_n986);
nor_1  g00610(new_n986, new_n983, new_n987);
not_1  g00611(new_n987, new_n988);
nor_1  g00612(new_n988, new_n985, new_n989);
nor_1  g00613(new_n989, new_n983, new_n990);
nor_1  g00614(new_n990, new_n976, new_n991);
nor_1  g00615(new_n991, new_n975, new_n992_1);
xnor_1 g00616(new_n966, new_n965, new_n993);
not_1  g00617(new_n993, new_n994);
nand_1 g00618(new_n994, new_n992_1, new_n995);
nand_1 g00619(new_n995, new_n967, new_n996_1);
nand_1 g00620(new_n996_1, new_n964, new_n997);
nand_1 g00621(new_n997, new_n963, new_n998);
xnor_1 g00622(new_n957, new_n954, new_n999);
nand_1 g00623(new_n999, new_n998, new_n1000);
nand_1 g00624(new_n1000, new_n958, new_n1001);
xnor_1 g00625(new_n1001, new_n550, new_n1002);
not_1  g00626(new_n1002, new_n1003);
nor_1  g00627(new_n628, new_n625, new_n1004);
nor_1  g00628(new_n636, new_n1004, new_n1005);
nor_1  g00629(new_n563, new_n621, new_n1006);
nand_1 g00630(n12299, n4141, new_n1007);
nand_1 g00631(n8759, n8236, new_n1008);
xnor_1 g00632(new_n1008, new_n1007, new_n1009);
xor_1  g00633(new_n1009, new_n1006, new_n1010);
xnor_1 g00634(new_n1010, new_n1005, new_n1011);
nor_1  g00635(new_n627, new_n626, new_n1012);
nor_1  g00636(new_n599, new_n551, new_n1013);
xor_1  g00637(new_n1013, new_n1012, new_n1014);
nand_1 g00638(n9241, n7500, new_n1015);
nand_1 g00639(n8276, n1209, new_n1016);
nand_1 g00640(n10510, n7354, new_n1017);
xnor_1 g00641(new_n1017, new_n1016, new_n1018);
xnor_1 g00642(new_n1018, new_n1015, new_n1019);
xnor_1 g00643(new_n1019, new_n1014, new_n1020_1);
not_1  g00644(new_n1020_1, new_n1021);
xnor_1 g00645(new_n1021, new_n1011, new_n1022);
not_1  g00646(new_n646, new_n1023);
nand_1 g00647(new_n1023, new_n638, new_n1024);
nand_1 g00648(new_n650, new_n644, new_n1025);
nand_1 g00649(new_n649, new_n645, new_n1026);
nand_1 g00650(new_n1026, new_n1025, new_n1027);
nand_1 g00651(new_n1027, new_n1024, new_n1028);
xnor_1 g00652(new_n1028, new_n1022, new_n1029);
xnor_1 g00653(new_n1029, new_n654, new_n1030);
nand_1 g00654(new_n657, new_n622, new_n1031);
nand_1 g00655(new_n658_1, new_n620, new_n1032);
nand_1 g00656(new_n1032, new_n1031, new_n1033);
xnor_1 g00657(new_n1033, new_n1030, new_n1034);
nand_1 g00658(new_n902, new_n899, new_n1035);
nor_1  g00659(new_n874, new_n871, new_n1036);
nor_1  g00660(new_n882, new_n1036, new_n1037);
not_1  g00661(new_n1037, new_n1038);
nor_1  g00662(new_n712, new_n867, new_n1039);
nand_1 g00663(n6806, n2530, new_n1040);
nand_1 g00664(n12044, n5331, new_n1041);
xnor_1 g00665(new_n1041, new_n1040, new_n1042);
xor_1  g00666(new_n1042, new_n1039, new_n1043);
xnor_1 g00667(new_n1043, new_n1038, new_n1044);
nor_1  g00668(new_n873, new_n872, new_n1045);
nor_1  g00669(new_n829, new_n735, new_n1046);
xnor_1 g00670(new_n1046, new_n1045, new_n1047);
not_1  g00671(n7690, new_n1048);
nor_1  g00672(new_n1048, new_n711, new_n1049);
nand_1 g00673(n10545, n533, new_n1050);
nand_1 g00674(n3616, n1564, new_n1051);
xnor_1 g00675(new_n1051, new_n1050, new_n1052);
xnor_1 g00676(new_n1052, new_n1049, new_n1053);
not_1  g00677(new_n1053, new_n1054);
nand_1 g00678(new_n1054, new_n1047, new_n1055);
not_1  g00679(new_n1047, new_n1056);
nand_1 g00680(new_n1053, new_n1056, new_n1057);
nand_1 g00681(new_n1057, new_n1055, new_n1058);
not_1  g00682(new_n1058, new_n1059);
xnor_1 g00683(new_n1059, new_n1044, new_n1060);
not_1  g00684(new_n890, new_n1061);
nand_1 g00685(new_n1061, new_n884, new_n1062);
nand_1 g00686(new_n897, new_n888, new_n1063);
nand_1 g00687(new_n896, new_n889, new_n1064);
nand_1 g00688(new_n1064, new_n1063, new_n1065);
nand_1 g00689(new_n1065, new_n1062, new_n1066);
xnor_1 g00690(new_n1066, new_n1060, new_n1067_1);
xnor_1 g00691(new_n1067_1, new_n1035, new_n1068);
nand_1 g00692(new_n907, new_n847, new_n1069);
nand_1 g00693(new_n1069, new_n905, new_n1070);
xnor_1 g00694(new_n1070, new_n1068, new_n1071);
not_1  g00695(new_n946, new_n1072);
nor_1  g00696(new_n949, new_n1072, new_n1073);
nand_1 g00697(new_n933, new_n929, new_n1074);
nand_1 g00698(new_n1074, new_n926, new_n1075);
nor_1  g00699(new_n696, new_n915, new_n1076);
nand_1 g00700(n12704, n11892, new_n1077);
nand_1 g00701(n7965, n4903, new_n1078);
xnor_1 g00702(new_n1078, new_n1077, new_n1079);
xor_1  g00703(new_n1079, new_n1076, new_n1080);
xnor_1 g00704(new_n1080, new_n1075, new_n1081);
nand_1 g00705(n7294, n2393, new_n1082);
xnor_1 g00706(new_n1082, new_n922, new_n1083);
not_1  g00707(n3986, new_n1084);
nor_1  g00708(new_n697, new_n1084, new_n1085);
nand_1 g00709(n5860, n1980, new_n1086);
nand_1 g00710(n8028, n5857, new_n1087);
xnor_1 g00711(new_n1087, new_n1086, new_n1088);
xor_1  g00712(new_n1088, new_n1085, new_n1089);
xnor_1 g00713(new_n1089, new_n1083, new_n1090);
xnor_1 g00714(new_n1090, new_n1081, new_n1091);
nor_1  g00715(new_n942, new_n934, new_n1092);
not_1  g00716(new_n945, new_n1093);
nand_1 g00717(new_n1093, new_n944, new_n1094_1);
xnor_1 g00718(new_n1094_1, new_n940, new_n1095);
nor_1  g00719(new_n1095, new_n1092, new_n1096);
not_1  g00720(new_n1096, new_n1097_1);
xnor_1 g00721(new_n1097_1, new_n1091, new_n1098);
xnor_1 g00722(new_n1098, new_n1073, new_n1099);
nor_1  g00723(new_n950, new_n916, new_n1100);
not_1  g00724(new_n914, new_n1101);
not_1  g00725(new_n916, new_n1102);
not_1  g00726(new_n950, new_n1103);
nor_1  g00727(new_n1103, new_n1102, new_n1104);
nor_1  g00728(new_n1104, new_n1101, new_n1105);
nor_1  g00729(new_n1105, new_n1100, new_n1106);
xnor_1 g00730(new_n1106, new_n1099, new_n1107);
xnor_1 g00731(new_n1107, new_n1071, new_n1108);
not_1  g00732(new_n952, new_n1109);
nand_1 g00733(new_n1109, new_n912, new_n1110);
nand_1 g00734(new_n1110, new_n911_1, new_n1111);
xnor_1 g00735(new_n1111, new_n1108, new_n1112);
xnor_1 g00736(new_n1112, new_n1034, new_n1113);
not_1  g00737(new_n1113, new_n1114);
nand_1 g00738(new_n861, new_n659, new_n1115);
not_1  g00739(new_n862, new_n1116);
nand_1 g00740(new_n953, new_n1116, new_n1117);
nand_1 g00741(new_n1117, new_n1115, new_n1118);
xnor_1 g00742(new_n1118, new_n1114, new_n1119);
xnor_1 g00743(new_n1119, new_n1003, n226);
not_1  g00744(n4634, new_n1121);
nor_1  g00745(new_n456, new_n1121, new_n1122);
nand_1 g00746(n10223, n5305, new_n1123);
nand_1 g00747(n7265, n1097, new_n1124);
nand_1 g00748(new_n1124, new_n1123, new_n1125);
not_1  g00749(new_n1125, new_n1126);
nand_1 g00750(n7265, n5305, new_n1127);
nand_1 g00751(n10223, n1097, new_n1128);
nor_1  g00752(new_n1128, new_n1127, new_n1129);
not_1  g00753(n2879, new_n1130);
nor_1  g00754(new_n424, new_n1130, new_n1131);
nor_1  g00755(new_n1131, new_n1129, new_n1132);
nor_1  g00756(new_n1132, new_n1126, new_n1133);
nand_1 g00757(new_n1133, new_n1122, new_n1134);
not_1  g00758(new_n1134, new_n1135);
nor_1  g00759(new_n1133, new_n1122, new_n1136_1);
nor_1  g00760(new_n1136_1, new_n1135, new_n1137);
nor_1  g00761(new_n1130, new_n419, new_n1138_1);
not_1  g00762(n10223, new_n1139);
nor_1  g00763(new_n1139, new_n424, new_n1140);
not_1  g00764(new_n1140, new_n1141);
not_1  g00765(n7265, new_n1142);
nor_1  g00766(new_n1142, new_n395, new_n1143);
not_1  g00767(new_n1143, new_n1144);
nand_1 g00768(new_n1144, new_n1141, new_n1145);
nor_1  g00769(new_n1144, new_n1141, new_n1146);
not_1  g00770(new_n1146, new_n1147);
nand_1 g00771(new_n1147, new_n1145, new_n1148);
xnor_1 g00772(new_n1148, new_n1138_1, new_n1149);
nand_1 g00773(new_n1149, new_n1137, new_n1150);
not_1  g00774(new_n1150, new_n1151);
nor_1  g00775(new_n1149, new_n1137, new_n1152);
nor_1  g00776(new_n1152, new_n1151, new_n1153);
not_1  g00777(new_n1131, new_n1154);
not_1  g00778(new_n1127, new_n1155);
nor_1  g00779(new_n1154, new_n1155, new_n1156);
nor_1  g00780(new_n1129, new_n1126, new_n1157);
nor_1  g00781(new_n1157, new_n1156, new_n1158);
not_1  g00782(new_n1158, new_n1159);
nor_1  g00783(new_n1159, new_n1154, new_n1160);
xor_1  g00784(new_n1160, new_n1153, new_n1161);
nand_1 g00785(new_n1156, new_n1125, new_n1162);
nand_1 g00786(new_n1162, new_n1159, new_n1163);
nand_1 g00787(n8759, n7946, new_n1164);
nand_1 g00788(n5331, n2558, new_n1165);
nand_1 g00789(n9763, n7965, new_n1166);
nor_1  g00790(new_n1166, new_n1165, new_n1167);
not_1  g00791(new_n1167, new_n1168);
nand_1 g00792(new_n1166, new_n1165, new_n1169);
nand_1 g00793(new_n1169, new_n1168, new_n1170);
nor_1  g00794(new_n1170, new_n1164, new_n1171);
nand_1 g00795(n7946, n6776, new_n1172);
nand_1 g00796(n8759, n2024, new_n1173);
xnor_1 g00797(new_n1173, new_n1172, new_n1174);
not_1  g00798(new_n1174, new_n1175);
nand_1 g00799(new_n1175, new_n1171, new_n1176);
nand_1 g00800(n9111, n7965, new_n1177);
nand_1 g00801(n9763, n7388, new_n1178);
xnor_1 g00802(new_n1178, new_n1177, new_n1179);
xnor_1 g00803(new_n1179, new_n1167, new_n1180);
nand_1 g00804(n5331, n2498, new_n1181);
nand_1 g00805(n8476, n2558, new_n1182);
nand_1 g00806(new_n1182, new_n1181, new_n1183);
nor_1  g00807(new_n1182, new_n1181, new_n1184);
not_1  g00808(new_n1184, new_n1185);
nand_1 g00809(new_n1185, new_n1183, new_n1186);
xnor_1 g00810(new_n1186, new_n1180, new_n1187);
xnor_1 g00811(new_n1174, new_n1171, new_n1188);
nand_1 g00812(new_n1188, new_n1187, new_n1189);
nand_1 g00813(new_n1189, new_n1176, new_n1190);
not_1  g00814(new_n1164, new_n1191);
not_1  g00815(n2024, new_n1192);
nor_1  g00816(new_n563, new_n1192, new_n1193);
not_1  g00817(new_n1193, new_n1194);
nor_1  g00818(new_n1194, new_n1191, new_n1195);
not_1  g00819(n7946, new_n1196);
nor_1  g00820(new_n554, new_n1196, new_n1197);
not_1  g00821(new_n1197, new_n1198_1);
not_1  g00822(n9189, new_n1199_1);
nor_1  g00823(new_n1199_1, new_n552, new_n1200);
not_1  g00824(new_n1200, new_n1201);
nand_1 g00825(new_n1201, new_n1198_1, new_n1202);
not_1  g00826(new_n1202, new_n1203);
nor_1  g00827(new_n1201, new_n1198_1, new_n1204);
nor_1  g00828(new_n1204, new_n1203, new_n1205);
nor_1  g00829(new_n1205, new_n1195, new_n1206);
not_1  g00830(new_n1206, new_n1207);
nand_1 g00831(new_n1202, new_n1195, new_n1208);
nand_1 g00832(new_n1208, new_n1207, new_n1209_1);
xnor_1 g00833(new_n1209_1, new_n1190, new_n1210);
nand_1 g00834(new_n1179, new_n1168, new_n1211);
nand_1 g00835(new_n1186, new_n1180, new_n1212);
nand_1 g00836(new_n1212, new_n1211, new_n1213);
not_1  g00837(new_n1166, new_n1214);
not_1  g00838(n9111, new_n1215);
nor_1  g00839(new_n1215, new_n696, new_n1216);
not_1  g00840(new_n1216, new_n1217);
nor_1  g00841(new_n1217, new_n1214, new_n1218);
not_1  g00842(n3342, new_n1219);
nor_1  g00843(new_n762, new_n1219, new_n1220);
nand_1 g00844(new_n1220, new_n1214, new_n1221);
not_1  g00845(new_n1221, new_n1222);
nand_1 g00846(n11892, n9763, new_n1223);
nand_1 g00847(n7965, n3342, new_n1224);
nand_1 g00848(new_n1224, new_n1223, new_n1225);
not_1  g00849(new_n1225, new_n1226);
nor_1  g00850(new_n1226, new_n1222, new_n1227);
nor_1  g00851(new_n1227, new_n1218, new_n1228);
nand_1 g00852(new_n1225, new_n1218, new_n1229);
not_1  g00853(new_n1229, new_n1230);
nor_1  g00854(new_n1230, new_n1228, new_n1231);
xnor_1 g00855(new_n1231, new_n1213, new_n1232);
not_1  g00856(new_n1232, new_n1233);
not_1  g00857(new_n1165, new_n1234);
not_1  g00858(n2498, new_n1235);
nor_1  g00859(new_n712, new_n1235, new_n1236);
not_1  g00860(new_n1236, new_n1237);
nor_1  g00861(new_n1237, new_n1234, new_n1238);
nand_1 g00862(n2558, n2530, new_n1239);
nand_1 g00863(n5579, n5331, new_n1240);
nand_1 g00864(new_n1240, new_n1239, new_n1241);
not_1  g00865(new_n1241, new_n1242);
and_1  g00866(new_n1242, new_n1238, new_n1243);
not_1  g00867(n5579, new_n1244);
nor_1  g00868(new_n1244, new_n740, new_n1245);
not_1  g00869(new_n1245, new_n1246);
nor_1  g00870(new_n1246, new_n1165, new_n1247);
nor_1  g00871(new_n1247, new_n1242, new_n1248);
not_1  g00872(new_n1248, new_n1249);
nor_1  g00873(new_n1249, new_n1238, new_n1250);
nor_1  g00874(new_n1250, new_n1243, new_n1251);
xnor_1 g00875(new_n1251, new_n1233, new_n1252);
nand_1 g00876(new_n1252, new_n1210, new_n1253);
not_1  g00877(new_n1253, new_n1254);
nor_1  g00878(new_n1252, new_n1210, new_n1255);
nor_1  g00879(new_n1255, new_n1254, new_n1256);
nor_1  g00880(new_n1256, new_n1163, new_n1257);
not_1  g00881(new_n1257, new_n1258);
xnor_1 g00882(new_n1170, new_n1191, new_n1259);
nand_1 g00883(new_n1259, new_n1155, new_n1260);
nand_1 g00884(n7265, n5964, new_n1261);
nor_1  g00885(new_n456, new_n1130, new_n1262);
xnor_1 g00886(new_n1262, new_n1261, new_n1263);
not_1  g00887(new_n1263, new_n1264);
nand_1 g00888(new_n1264, new_n1260, new_n1265);
not_1  g00889(new_n1265, new_n1266);
xor_1  g00890(new_n1188, new_n1187, new_n1267);
nor_1  g00891(new_n1264, new_n1260, new_n1268);
nor_1  g00892(new_n1268, new_n1266, new_n1269_1);
not_1  g00893(new_n1269_1, new_n1270);
nor_1  g00894(new_n1270, new_n1267, new_n1271);
nor_1  g00895(new_n1271, new_n1266, new_n1272);
not_1  g00896(new_n1163, new_n1273);
xnor_1 g00897(new_n1256, new_n1273, new_n1274);
nand_1 g00898(new_n1274, new_n1272, new_n1275);
nand_1 g00899(new_n1275, new_n1258, new_n1276);
xnor_1 g00900(new_n1276, new_n1161, new_n1277);
not_1  g00901(n2522, new_n1278);
nor_1  g00902(new_n552, new_n1278, new_n1279);
nor_1  g00903(new_n1204, new_n1193, new_n1280);
nor_1  g00904(new_n1280, new_n1203, new_n1281);
nand_1 g00905(new_n1281, new_n1279, new_n1282);
not_1  g00906(new_n1282, new_n1283);
nor_1  g00907(new_n1281, new_n1279, new_n1284);
nor_1  g00908(new_n1284, new_n1283, new_n1285);
nor_1  g00909(new_n554, new_n1192, new_n1286);
not_1  g00910(new_n1286, new_n1287);
nand_1 g00911(n7946, n7436, new_n1288);
nand_1 g00912(n9189, n6776, new_n1289);
nand_1 g00913(new_n1289, new_n1288, new_n1290);
not_1  g00914(new_n1290, new_n1291);
nor_1  g00915(new_n1289, new_n1288, new_n1292);
nor_1  g00916(new_n1292, new_n1291, new_n1293);
xnor_1 g00917(new_n1293, new_n1287, new_n1294);
nand_1 g00918(new_n1294, new_n1285, new_n1295);
not_1  g00919(new_n1295, new_n1296);
nor_1  g00920(new_n1294, new_n1285, new_n1297);
nor_1  g00921(new_n1297, new_n1296, new_n1298);
nor_1  g00922(new_n1207, new_n1194, new_n1299);
nor_1  g00923(new_n1299, new_n1298, new_n1300);
not_1  g00924(new_n1298, new_n1301);
not_1  g00925(new_n1299, new_n1302);
nor_1  g00926(new_n1302, new_n1301, new_n1303);
nor_1  g00927(new_n1303, new_n1300, new_n1304);
not_1  g00928(new_n1209_1, new_n1305);
nor_1  g00929(new_n1305, new_n1190, new_n1306);
not_1  g00930(new_n1306, new_n1307);
nand_1 g00931(new_n1253, new_n1307, new_n1308);
xnor_1 g00932(new_n1308, new_n1304, new_n1309);
not_1  g00933(n521, new_n1310);
nor_1  g00934(new_n668, new_n1310, new_n1311);
nor_1  g00935(new_n1247, new_n1236, new_n1312);
nor_1  g00936(new_n1312, new_n1242, new_n1313);
xnor_1 g00937(new_n1313, new_n1311, new_n1314);
nor_1  g00938(new_n740, new_n1235, new_n1315);
not_1  g00939(new_n1315, new_n1316);
nand_1 g00940(n12648, n2558, new_n1317);
nand_1 g00941(n8476, n5579, new_n1318);
xnor_1 g00942(new_n1318, new_n1317, new_n1319);
xnor_1 g00943(new_n1319, new_n1316, new_n1320);
not_1  g00944(new_n1320, new_n1321);
xnor_1 g00945(new_n1321, new_n1314, new_n1322);
nor_1  g00946(new_n1248, new_n1185, new_n1323);
xnor_1 g00947(new_n1323, new_n1322, new_n1324);
not_1  g00948(n806, new_n1325);
nor_1  g00949(new_n754, new_n1325, new_n1326);
nand_1 g00950(new_n1225, new_n1216, new_n1327);
nand_1 g00951(new_n1327, new_n1221, new_n1328);
xnor_1 g00952(new_n1328, new_n1326, new_n1329);
nor_1  g00953(new_n762, new_n1215, new_n1330);
not_1  g00954(new_n1330, new_n1331);
nand_1 g00955(n9763, n2393, new_n1332);
nand_1 g00956(n7388, n3342, new_n1333_1);
xnor_1 g00957(new_n1333_1, new_n1332, new_n1334);
xnor_1 g00958(new_n1334, new_n1331, new_n1335);
xnor_1 g00959(new_n1335, new_n1329, new_n1336);
nand_1 g00960(new_n1228, new_n1216, new_n1337);
not_1  g00961(new_n1337, new_n1338);
xnor_1 g00962(new_n1338, new_n1336, new_n1339);
xnor_1 g00963(new_n1339, new_n1324, new_n1340);
not_1  g00964(new_n1231, new_n1341);
nand_1 g00965(new_n1341, new_n1213, new_n1342);
nand_1 g00966(new_n1251, new_n1232, new_n1343);
nand_1 g00967(new_n1343, new_n1342, new_n1344);
xnor_1 g00968(new_n1344, new_n1340, new_n1345);
xnor_1 g00969(new_n1345, new_n1309, new_n1346);
xor_1  g00970(new_n1346, new_n1277, n381);
not_1  g00971(n7862, new_n1348);
nor_1  g00972(new_n1348, new_n377, new_n1349);
not_1  g00973(n6877, new_n1350);
nor_1  g00974(new_n381_1, new_n1350, new_n1351);
not_1  g00975(new_n1351, new_n1352);
nand_1 g00976(n4805, n1564, new_n1353_1);
nand_1 g00977(n8028, n7236, new_n1354);
not_1  g00978(new_n1354, new_n1355);
xnor_1 g00979(new_n1355, new_n1353_1, new_n1356);
not_1  g00980(new_n1356, new_n1357_1);
nor_1  g00981(new_n1357_1, new_n1352, new_n1358);
nor_1  g00982(new_n1356, new_n1351, new_n1359);
nor_1  g00983(new_n1359, new_n1358, new_n1360);
nand_1 g00984(new_n1360, new_n1349, new_n1361);
not_1  g00985(new_n1361, new_n1362);
nor_1  g00986(new_n1360, new_n1349, new_n1363);
nor_1  g00987(new_n1363, new_n1362, n397);
not_1  g00988(n4370, new_n1365);
nor_1  g00989(new_n378, new_n1365, new_n1366);
not_1  g00990(n4189, new_n1367);
not_1  g00991(n11407, new_n1368);
nor_1  g00992(new_n1368, new_n1367, new_n1369);
not_1  g00993(new_n1369, new_n1370);
not_1  g00994(n11877, new_n1371);
nor_1  g00995(new_n1371, new_n378, new_n1372);
not_1  g00996(new_n1372, new_n1373);
nand_1 g00997(new_n1373, new_n1370, new_n1374);
not_1  g00998(new_n1374, new_n1375);
nor_1  g00999(new_n1373, new_n1370, new_n1376);
not_1  g01000(n2564, new_n1377);
not_1  g01001(n5212, new_n1378);
nor_1  g01002(new_n1378, new_n1377, new_n1379);
nor_1  g01003(new_n1379, new_n1376, new_n1380);
nor_1  g01004(new_n1380, new_n1375, new_n1381);
nand_1 g01005(new_n1381, new_n1366, new_n1382);
not_1  g01006(new_n1382, new_n1383);
nor_1  g01007(new_n1381, new_n1366, new_n1384);
nor_1  g01008(new_n1384, new_n1383, new_n1385);
nor_1  g01009(new_n1378, new_n1367, new_n1386);
nand_1 g01010(n11407, n6770, new_n1387);
nand_1 g01011(n11877, n2564, new_n1388);
xnor_1 g01012(new_n1388, new_n1387, new_n1389);
xnor_1 g01013(new_n1389, new_n1386, new_n1390);
nand_1 g01014(new_n1390, new_n1385, new_n1391);
not_1  g01015(new_n1391, new_n1392);
nor_1  g01016(new_n1390, new_n1385, new_n1393);
nor_1  g01017(new_n1393, new_n1392, new_n1394);
not_1  g01018(new_n1379, new_n1395);
nor_1  g01019(new_n1368, new_n378, new_n1396);
nor_1  g01020(new_n1396, new_n1395, new_n1397);
nor_1  g01021(new_n1397, new_n1374, new_n1398);
nor_1  g01022(new_n1398, new_n1376, new_n1399);
nor_1  g01023(new_n1399, new_n1395, new_n1400);
xor_1  g01024(new_n1400, new_n1394, new_n1401);
not_1  g01025(n12709, new_n1402);
nor_1  g01026(new_n1402, new_n382, new_n1403);
not_1  g01027(new_n1403, new_n1404);
nand_1 g01028(n11222, n10990, new_n1405);
nand_1 g01029(n12489, n12069, new_n1406);
nor_1  g01030(new_n1406, new_n1405, new_n1407);
not_1  g01031(new_n1407, new_n1408);
nand_1 g01032(new_n1406, new_n1405, new_n1409);
nand_1 g01033(new_n1409, new_n1408, new_n1410);
nor_1  g01034(new_n1410, new_n1404, new_n1411);
nand_1 g01035(n11728, n8336, new_n1412);
nand_1 g01036(n12709, n10928, new_n1413);
xnor_1 g01037(new_n1413, new_n1412, new_n1414);
not_1  g01038(new_n1414, new_n1415);
nor_1  g01039(new_n1415, new_n1411, new_n1416);
not_1  g01040(new_n1416, new_n1417);
nand_1 g01041(n11222, n5760, new_n1418);
nand_1 g01042(n11153, n10990, new_n1419);
xnor_1 g01043(new_n1419, new_n1418, new_n1420);
xnor_1 g01044(new_n1420, new_n1408, new_n1421);
nand_1 g01045(n12069, n7159, new_n1422);
nand_1 g01046(n12489, n12391, new_n1423);
xnor_1 g01047(new_n1423, new_n1422, new_n1424);
nand_1 g01048(new_n1424, new_n1421, new_n1425);
nor_1  g01049(new_n1424, new_n1421, new_n1426);
not_1  g01050(new_n1426, new_n1427);
nand_1 g01051(new_n1427, new_n1425, new_n1428);
nand_1 g01052(new_n1415, new_n1411, new_n1429);
nand_1 g01053(new_n1429, new_n1417, new_n1430);
not_1  g01054(new_n1430, new_n1431);
nand_1 g01055(new_n1431, new_n1428, new_n1432);
nand_1 g01056(new_n1432, new_n1417, new_n1433);
not_1  g01057(n10928, new_n1434);
not_1  g01058(n11728, new_n1435);
nor_1  g01059(new_n1435, new_n1434, new_n1436);
not_1  g01060(new_n1436, new_n1437);
nor_1  g01061(new_n1437, new_n1403, new_n1438);
nand_1 g01062(n6986, n6429, new_n1439);
nor_1  g01063(new_n1439, new_n1404, new_n1440);
nand_1 g01064(n12709, n6986, new_n1441);
nand_1 g01065(n8336, n6429, new_n1442);
nand_1 g01066(new_n1442, new_n1441, new_n1443);
not_1  g01067(new_n1443, new_n1444);
nor_1  g01068(new_n1444, new_n1440, new_n1445);
nor_1  g01069(new_n1445, new_n1438, new_n1446);
not_1  g01070(new_n1446, new_n1447);
nand_1 g01071(new_n1443, new_n1438, new_n1448);
nand_1 g01072(new_n1448, new_n1447, new_n1449);
xnor_1 g01073(new_n1449, new_n1433, new_n1450);
not_1  g01074(n7159, new_n1451);
not_1  g01075(n12391, new_n1452);
nor_1  g01076(new_n1452, new_n1451, new_n1453);
nand_1 g01077(new_n1453, new_n1406, new_n1454);
nand_1 g01078(n12489, n7891, new_n1455);
nand_1 g01079(n12777, n12069, new_n1456);
nand_1 g01080(new_n1456, new_n1455, new_n1457);
not_1  g01081(new_n1457, new_n1458);
nand_1 g01082(new_n1458, new_n1454, new_n1459);
not_1  g01083(new_n1459, new_n1460);
nor_1  g01084(new_n1456, new_n1455, new_n1461);
nor_1  g01085(new_n1461, new_n1460, new_n1462);
not_1  g01086(new_n1462, new_n1463);
nor_1  g01087(new_n1458, new_n1454, new_n1464);
nor_1  g01088(new_n1464, new_n1463, new_n1465);
not_1  g01089(n5760, new_n1466);
not_1  g01090(n11153, new_n1467);
nor_1  g01091(new_n1467, new_n1466, new_n1468);
nand_1 g01092(new_n1468, new_n1405, new_n1469);
not_1  g01093(new_n1469, new_n1470);
nand_1 g01094(n10990, n5314, new_n1471_1);
nand_1 g01095(n11222, n1478, new_n1472);
nand_1 g01096(new_n1472, new_n1471_1, new_n1473);
not_1  g01097(new_n1473, new_n1474);
nor_1  g01098(new_n1472, new_n1471_1, new_n1475);
nor_1  g01099(new_n1475, new_n1474, new_n1476);
nor_1  g01100(new_n1476, new_n1470, new_n1477);
nor_1  g01101(new_n1474, new_n1469, new_n1478_1);
nor_1  g01102(new_n1478_1, new_n1477, new_n1479);
xnor_1 g01103(new_n1479, new_n1465, new_n1480);
nor_1  g01104(new_n1420, new_n1408, new_n1481);
nor_1  g01105(new_n1426, new_n1481, new_n1482);
xnor_1 g01106(new_n1482, new_n1480, new_n1483);
not_1  g01107(new_n1483, new_n1484);
xnor_1 g01108(new_n1484, new_n1450, new_n1485);
nand_1 g01109(new_n1397, new_n1374, new_n1486);
nand_1 g01110(new_n1486, new_n1399, new_n1487);
not_1  g01111(new_n1487, new_n1488);
nor_1  g01112(new_n1488, new_n1485, new_n1489);
not_1  g01113(new_n1489, new_n1490);
xnor_1 g01114(new_n1487, new_n1485, new_n1491);
xnor_1 g01115(new_n1410, new_n1403, new_n1492);
nand_1 g01116(new_n1492, new_n1396, new_n1493);
nand_1 g01117(n11407, n2564, new_n1494);
nor_1  g01118(new_n378, new_n1378, new_n1495);
xnor_1 g01119(new_n1495, new_n1494, new_n1496);
not_1  g01120(new_n1496, new_n1497);
nand_1 g01121(new_n1497, new_n1493, new_n1498);
xnor_1 g01122(new_n1430, new_n1428, new_n1499);
xnor_1 g01123(new_n1496, new_n1493, new_n1500);
nand_1 g01124(new_n1500, new_n1499, new_n1501);
nand_1 g01125(new_n1501, new_n1498, new_n1502);
nand_1 g01126(new_n1502, new_n1491, new_n1503);
nand_1 g01127(new_n1503, new_n1490, new_n1504);
xnor_1 g01128(new_n1504, new_n1401, new_n1505);
not_1  g01129(n8819, new_n1506);
nor_1  g01130(new_n1506, new_n382, new_n1507);
not_1  g01131(n6986, new_n1508);
nor_1  g01132(new_n1435, new_n1508, new_n1509);
nand_1 g01133(n10928, n6429, new_n1510_1);
nand_1 g01134(n12709, n2226, new_n1511);
nand_1 g01135(new_n1511, new_n1510_1, new_n1512_1);
nor_1  g01136(new_n1511, new_n1510_1, new_n1513);
not_1  g01137(new_n1513, new_n1514);
nand_1 g01138(new_n1514, new_n1512_1, new_n1515);
xnor_1 g01139(new_n1515, new_n1509, new_n1516);
nand_1 g01140(new_n1516, new_n1507, new_n1517);
not_1  g01141(new_n1517, new_n1518);
nor_1  g01142(new_n1516, new_n1507, new_n1519);
nor_1  g01143(new_n1519, new_n1518, new_n1520);
nor_1  g01144(new_n1444, new_n1437, new_n1521);
nor_1  g01145(new_n1521, new_n1440, new_n1522);
not_1  g01146(new_n1522, new_n1523_1);
xnor_1 g01147(new_n1523_1, new_n1520, new_n1524);
not_1  g01148(new_n1524, new_n1525);
nor_1  g01149(new_n1447, new_n1437, new_n1526);
nor_1  g01150(new_n1526, new_n1525, new_n1527);
nand_1 g01151(new_n1526, new_n1525, new_n1528);
not_1  g01152(new_n1528, new_n1529);
nor_1  g01153(new_n1529, new_n1527, new_n1530);
not_1  g01154(new_n1530, new_n1531);
not_1  g01155(n6254, new_n1532);
not_1  g01156(n12069, new_n1533);
nor_1  g01157(new_n1533, new_n1532, new_n1534);
nor_1  g01158(new_n1461, new_n1453, new_n1535);
nor_1  g01159(new_n1535, new_n1458, new_n1536);
xnor_1 g01160(new_n1536, new_n1534, new_n1537);
not_1  g01161(n7160, new_n1538);
not_1  g01162(n12489, new_n1539);
nor_1  g01163(new_n1539, new_n1538, new_n1540);
not_1  g01164(new_n1540, new_n1541);
nand_1 g01165(n12777, n12391, new_n1542);
nand_1 g01166(n7891, n7159, new_n1543);
xnor_1 g01167(new_n1543, new_n1542, new_n1544);
xnor_1 g01168(new_n1544, new_n1541, new_n1545);
not_1  g01169(new_n1545, new_n1546);
xnor_1 g01170(new_n1546, new_n1537, new_n1547);
not_1  g01171(new_n1453, new_n1548);
nor_1  g01172(new_n1462, new_n1548, new_n1549);
nor_1  g01173(new_n1549, new_n1547, new_n1550);
nand_1 g01174(new_n1549, new_n1547, new_n1551);
not_1  g01175(new_n1551, new_n1552);
nor_1  g01176(new_n1552, new_n1550, new_n1553);
nand_1 g01177(n11791, n11222, new_n1554);
not_1  g01178(new_n1554, new_n1555);
nor_1  g01179(new_n1475, new_n1468, new_n1556);
nor_1  g01180(new_n1556, new_n1474, new_n1557);
nand_1 g01181(new_n1557, new_n1555, new_n1558);
not_1  g01182(new_n1558, new_n1559);
nor_1  g01183(new_n1557, new_n1555, new_n1560);
nor_1  g01184(new_n1560, new_n1559, new_n1561);
not_1  g01185(n5314, new_n1562);
nor_1  g01186(new_n1466, new_n1562, new_n1563);
not_1  g01187(new_n1563, new_n1564_1);
nand_1 g01188(n10990, n996, new_n1565);
nand_1 g01189(n11153, n1478, new_n1566);
xnor_1 g01190(new_n1566, new_n1565, new_n1567);
xnor_1 g01191(new_n1567, new_n1564_1, new_n1568);
xnor_1 g01192(new_n1568, new_n1561, new_n1569);
nand_1 g01193(new_n1477, new_n1468, new_n1570);
xnor_1 g01194(new_n1570, new_n1569, new_n1571);
not_1  g01195(new_n1571, new_n1572);
xnor_1 g01196(new_n1572, new_n1553, new_n1573);
nand_1 g01197(new_n1479, new_n1465, new_n1574);
not_1  g01198(new_n1574, new_n1575);
nor_1  g01199(new_n1482, new_n1480, new_n1576_1);
nor_1  g01200(new_n1576_1, new_n1575, new_n1577);
xnor_1 g01201(new_n1577, new_n1573, new_n1578);
xnor_1 g01202(new_n1578, new_n1531, new_n1579);
nand_1 g01203(new_n1449, new_n1433, new_n1580);
not_1  g01204(new_n1580, new_n1581);
nor_1  g01205(new_n1484, new_n1450, new_n1582);
nor_1  g01206(new_n1582, new_n1581, new_n1583);
nand_1 g01207(new_n1583, new_n1579, new_n1584);
not_1  g01208(new_n1584, new_n1585);
nor_1  g01209(new_n1583, new_n1579, new_n1586);
nor_1  g01210(new_n1586, new_n1585, new_n1587);
xor_1  g01211(new_n1587, new_n1505, n658);
nor_1  g01212(new_n1348, new_n423, new_n1589);
not_1  g01213(n1333, new_n1590);
nor_1  g01214(new_n420, new_n1590, new_n1591);
not_1  g01215(n11757, new_n1592);
nor_1  g01216(new_n1592, new_n377, new_n1593);
not_1  g01217(new_n1593, new_n1594);
nor_1  g01218(new_n396, new_n1590, new_n1595);
not_1  g01219(new_n1595, new_n1596);
nand_1 g01220(new_n1596, new_n1594, new_n1597);
not_1  g01221(new_n1597, new_n1598);
nor_1  g01222(new_n1596, new_n1594, new_n1599);
not_1  g01223(n3172, new_n1600);
nor_1  g01224(new_n1600, new_n413, new_n1601);
nor_1  g01225(new_n1601, new_n1599, new_n1602);
nor_1  g01226(new_n1602, new_n1598, new_n1603);
xnor_1 g01227(new_n1603, new_n1591, new_n1604);
nor_1  g01228(new_n1592, new_n413, new_n1605);
nand_1 g01229(n6038, n5240, new_n1606);
nand_1 g01230(n12720, n3172, new_n1607);
nand_1 g01231(new_n1607, new_n1606, new_n1608);
not_1  g01232(new_n1608, new_n1609);
nor_1  g01233(new_n1607, new_n1606, new_n1610);
nor_1  g01234(new_n1610, new_n1609, new_n1611);
xnor_1 g01235(new_n1611, new_n1605, new_n1612);
not_1  g01236(new_n1612, new_n1613);
xnor_1 g01237(new_n1613, new_n1604, new_n1614);
nor_1  g01238(new_n1614, new_n1589, new_n1615);
not_1  g01239(new_n1615, new_n1616);
not_1  g01240(new_n1589, new_n1617);
xnor_1 g01241(new_n1614, new_n1617, new_n1618);
nor_1  g01242(new_n1348, new_n420, new_n1619);
not_1  g01243(new_n1619, new_n1620);
nor_1  g01244(new_n413, new_n1590, new_n1621);
not_1  g01245(new_n1621, new_n1622);
nor_1  g01246(new_n377, new_n1600, new_n1623);
not_1  g01247(new_n1623, new_n1624);
nor_1  g01248(new_n396, new_n1348, new_n1625);
not_1  g01249(new_n1625, new_n1626);
nand_1 g01250(new_n1626, new_n1624, new_n1627);
not_1  g01251(new_n1627, new_n1628);
nor_1  g01252(new_n1628, new_n1622, new_n1629);
nor_1  g01253(new_n1626, new_n1624, new_n1630);
nor_1  g01254(new_n1630, new_n1629, new_n1631);
nor_1  g01255(new_n1631, new_n1620, new_n1632);
xnor_1 g01256(new_n1631, new_n1620, new_n1633);
not_1  g01257(new_n1599, new_n1634);
nand_1 g01258(new_n1634, new_n1597, new_n1635);
xnor_1 g01259(new_n1635, new_n1601, new_n1636);
not_1  g01260(new_n1636, new_n1637);
nor_1  g01261(new_n1637, new_n1633, new_n1638);
nor_1  g01262(new_n1638, new_n1632, new_n1639);
nand_1 g01263(new_n1639, new_n1618, new_n1640);
nand_1 g01264(new_n1640, new_n1616, new_n1641);
not_1  g01265(new_n1641, new_n1642);
nor_1  g01266(new_n396, new_n1592, new_n1643);
not_1  g01267(new_n1643, new_n1644);
nand_1 g01268(n5240, n2509, new_n1645);
nand_1 g01269(n11821, n6038, new_n1646);
xnor_1 g01270(new_n1646, new_n1645, new_n1647);
xnor_1 g01271(new_n1647, new_n1644, new_n1648);
not_1  g01272(new_n1648, new_n1649);
not_1  g01273(new_n1611, new_n1650);
nor_1  g01274(new_n1650, new_n1605, new_n1651);
nor_1  g01275(new_n1651, new_n1609, new_n1652);
nand_1 g01276(new_n1652, new_n1649, new_n1653);
not_1  g01277(new_n1653, new_n1654);
nor_1  g01278(new_n1652, new_n1649, new_n1655);
nor_1  g01279(new_n1655, new_n1654, new_n1656);
nand_1 g01280(new_n1603, new_n1591, new_n1657);
nor_1  g01281(new_n1612, new_n1604, new_n1658_1);
not_1  g01282(new_n1658_1, new_n1659);
nand_1 g01283(new_n1659, new_n1657, new_n1660);
not_1  g01284(new_n1660, new_n1661);
nor_1  g01285(new_n423, new_n1590, new_n1662);
not_1  g01286(new_n1662, new_n1663);
nor_1  g01287(new_n1600, new_n420, new_n1664);
not_1  g01288(new_n1664, new_n1665);
nor_1  g01289(new_n1665, new_n1663, new_n1666);
not_1  g01290(new_n1666, new_n1667);
nand_1 g01291(new_n1665, new_n1663, new_n1668);
nand_1 g01292(new_n1668, new_n1667, new_n1669);
nand_1 g01293(new_n1669, new_n1661, new_n1670);
nor_1  g01294(new_n1669, new_n1661, new_n1671);
not_1  g01295(new_n1671, new_n1672);
nand_1 g01296(new_n1672, new_n1670, new_n1673);
xnor_1 g01297(new_n1673, new_n1656, new_n1674);
nand_1 g01298(new_n1674, new_n1642, new_n1675);
nand_1 g01299(new_n1670, new_n1656, new_n1676);
xnor_1 g01300(new_n1676, new_n1666, new_n1677);
nor_1  g01301(new_n1677, new_n1671, new_n1678);
nor_1  g01302(new_n1646, new_n1645, new_n1679);
nor_1  g01303(new_n1592, new_n420, new_n1680);
xor_1  g01304(new_n1680, new_n1679, new_n1681);
not_1  g01305(n11821, new_n1682);
nor_1  g01306(new_n1682, new_n413, new_n1683);
nand_1 g01307(n12720, n5240, new_n1684);
nand_1 g01308(n9080, n6038, new_n1685);
xnor_1 g01309(new_n1685, new_n1684, new_n1686);
xnor_1 g01310(new_n1686, new_n1683, new_n1687);
xnor_1 g01311(new_n1687, new_n1681, new_n1688);
nor_1  g01312(new_n1647, new_n1644, new_n1689);
nor_1  g01313(new_n1654, new_n1689, new_n1690);
not_1  g01314(new_n1690, new_n1691);
nor_1  g01315(new_n492, new_n1590, new_n1692);
nor_1  g01316(new_n1600, new_n423, new_n1693);
not_1  g01317(new_n1693, new_n1694);
nor_1  g01318(new_n496, new_n1348, new_n1695);
not_1  g01319(new_n1695, new_n1696);
nand_1 g01320(new_n1696, new_n1694, new_n1697);
nand_1 g01321(new_n1695, new_n1693, new_n1698);
nand_1 g01322(new_n1698, new_n1697, new_n1699);
xor_1  g01323(new_n1699, new_n1692, new_n1700);
xnor_1 g01324(new_n1700, new_n1691, new_n1701);
xnor_1 g01325(new_n1701, new_n1688, new_n1702);
xnor_1 g01326(new_n1702, new_n1678, new_n1703);
xnor_1 g01327(new_n1703, new_n1675, new_n1704);
nor_1  g01328(new_n1348, new_n492, new_n1705);
not_1  g01329(new_n1675, new_n1706);
nor_1  g01330(new_n1674, new_n1642, new_n1707);
nor_1  g01331(new_n1707, new_n1706, new_n1708);
nand_1 g01332(new_n1708, new_n1705, new_n1709);
xnor_1 g01333(new_n1636, new_n1633, new_n1710);
nor_1  g01334(new_n1630, new_n1628, new_n1711);
nor_1  g01335(new_n377, new_n1590, new_n1712);
nor_1  g01336(new_n1348, new_n413, new_n1713);
nand_1 g01337(new_n1713, new_n1712, new_n1714);
nor_1  g01338(new_n1714, new_n1711, new_n1715);
nand_1 g01339(new_n1715, new_n1710, new_n1716);
xnor_1 g01340(new_n1639, new_n1618, new_n1717);
not_1  g01341(new_n1717, new_n1718);
nor_1  g01342(new_n1718, new_n1716, new_n1719);
not_1  g01343(new_n1705, new_n1720);
xnor_1 g01344(new_n1708, new_n1720, new_n1721);
nand_1 g01345(new_n1721, new_n1719, new_n1722);
nand_1 g01346(new_n1722, new_n1709, new_n1723);
xnor_1 g01347(new_n1723, new_n1704, new_n1724);
not_1  g01348(new_n1724, new_n1725);
nand_1 g01349(n6877, n5105, new_n1726);
not_1  g01350(new_n1726, new_n1727);
nor_1  g01351(new_n1350, new_n557, new_n1728);
not_1  g01352(n2464, new_n1729);
nor_1  g01353(new_n381_1, new_n1729, new_n1730);
nand_1 g01354(new_n1730, new_n1728, new_n1731);
not_1  g01355(new_n1728, new_n1732);
not_1  g01356(new_n1730, new_n1733);
nand_1 g01357(new_n1733, new_n1732, new_n1734);
not_1  g01358(n9400, new_n1735);
nor_1  g01359(new_n1735, new_n564, new_n1736);
nand_1 g01360(new_n1736, new_n1734, new_n1737);
nand_1 g01361(new_n1737, new_n1731, new_n1738);
nand_1 g01362(new_n1738, new_n1727, new_n1739);
not_1  g01363(new_n1739, new_n1740);
nor_1  g01364(new_n1738, new_n1727, new_n1741);
nor_1  g01365(new_n1741, new_n1740, new_n1742);
not_1  g01366(new_n1742, new_n1743);
nor_1  g01367(new_n564, new_n1729, new_n1744);
nor_1  g01368(new_n1735, new_n557, new_n1745);
not_1  g01369(new_n1745, new_n1746);
not_1  g01370(n11311, new_n1747);
nor_1  g01371(new_n1747, new_n381_1, new_n1748);
not_1  g01372(new_n1748, new_n1749);
nand_1 g01373(new_n1749, new_n1746, new_n1750);
nor_1  g01374(new_n1749, new_n1746, new_n1751);
not_1  g01375(new_n1751, new_n1752);
nand_1 g01376(new_n1752, new_n1750, new_n1753);
xnor_1 g01377(new_n1753, new_n1744, new_n1754);
not_1  g01378(new_n1754, new_n1755);
nor_1  g01379(new_n1755, new_n1743, new_n1756);
nor_1  g01380(new_n1754, new_n1742, new_n1757);
nor_1  g01381(new_n1757, new_n1756, new_n1758);
nand_1 g01382(new_n1734, new_n1731, new_n1759);
not_1  g01383(new_n1759, new_n1760);
nor_1  g01384(new_n1735, new_n381_1, new_n1761);
nor_1  g01385(new_n564, new_n1350, new_n1762);
nand_1 g01386(new_n1762, new_n1761, new_n1763);
nor_1  g01387(new_n1763, new_n1760, new_n1764);
nand_1 g01388(new_n1764, new_n1758, new_n1765);
nor_1  g01389(new_n1747, new_n564, new_n1766);
nand_1 g01390(n2464, n1209, new_n1767);
nand_1 g01391(n7354, n4187, new_n1768);
xnor_1 g01392(new_n1768, new_n1767, new_n1769);
nor_1  g01393(new_n1769, new_n1766, new_n1770);
not_1  g01394(new_n1770, new_n1771);
nand_1 g01395(new_n1769, new_n1766, new_n1772);
nand_1 g01396(new_n1772, new_n1771, new_n1773);
not_1  g01397(new_n1773, new_n1774);
nand_1 g01398(n9400, n5105, new_n1775);
not_1  g01399(new_n1775, new_n1776);
not_1  g01400(new_n1750, new_n1777);
nor_1  g01401(new_n1751, new_n1744, new_n1778);
nor_1  g01402(new_n1778, new_n1777, new_n1779);
nand_1 g01403(new_n1779, new_n1776, new_n1780);
not_1  g01404(new_n1780, new_n1781);
nor_1  g01405(new_n1779, new_n1776, new_n1782);
nor_1  g01406(new_n1782, new_n1781, new_n1783);
not_1  g01407(new_n1783, new_n1784);
nor_1  g01408(new_n1784, new_n1774, new_n1785);
not_1  g01409(new_n1785, new_n1786);
nand_1 g01410(new_n1784, new_n1774, new_n1787);
nand_1 g01411(new_n1787, new_n1786, new_n1788);
nor_1  g01412(new_n1350, new_n588, new_n1789);
nor_1  g01413(new_n1756, new_n1740, new_n1790);
xnor_1 g01414(new_n1790, new_n1789, new_n1791);
nand_1 g01415(new_n1791, new_n1788, new_n1792);
not_1  g01416(new_n1792, new_n1793);
nor_1  g01417(new_n1791, new_n1788, new_n1794);
nor_1  g01418(new_n1794, new_n1793, new_n1795);
nor_1  g01419(new_n1795, new_n1765, new_n1796);
nor_1  g01420(new_n1350, new_n621, new_n1797);
not_1  g01421(new_n1797, new_n1798_1);
not_1  g01422(new_n1789, new_n1799);
nand_1 g01423(new_n1790, new_n1799, new_n1800);
nand_1 g01424(new_n1792, new_n1800, new_n1801);
not_1  g01425(new_n1801, new_n1802);
nor_1  g01426(new_n1747, new_n557, new_n1803);
nand_1 g01427(n7500, n4187, new_n1804);
nand_1 g01428(n7354, n4203, new_n1805);
xnor_1 g01429(new_n1805, new_n1804, new_n1806);
xnor_1 g01430(new_n1806, new_n1803, new_n1807);
nand_1 g01431(new_n1768, new_n1767, new_n1808);
and_1  g01432(new_n1771, new_n1808, new_n1809);
xnor_1 g01433(new_n1809, new_n1807, new_n1810);
not_1  g01434(new_n1810, new_n1811);
nor_1  g01435(new_n1785, new_n1781, new_n1812);
nor_1  g01436(new_n1735, new_n588, new_n1813);
not_1  g01437(new_n1813, new_n1814);
nor_1  g01438(new_n551, new_n1729, new_n1815);
not_1  g01439(new_n1815, new_n1816);
nor_1  g01440(new_n1816, new_n1814, new_n1817);
not_1  g01441(new_n1817, new_n1818);
nand_1 g01442(new_n1816, new_n1814, new_n1819);
nand_1 g01443(new_n1819, new_n1818, new_n1820);
nand_1 g01444(new_n1820, new_n1812, new_n1821);
not_1  g01445(new_n1812, new_n1822);
not_1  g01446(new_n1820, new_n1823);
nand_1 g01447(new_n1823, new_n1822, new_n1824);
nand_1 g01448(new_n1824, new_n1821, new_n1825);
xnor_1 g01449(new_n1825, new_n1811, new_n1826);
nand_1 g01450(new_n1826, new_n1802, new_n1827);
not_1  g01451(new_n1827, new_n1828);
nor_1  g01452(new_n1826, new_n1802, new_n1829);
nor_1  g01453(new_n1829, new_n1828, new_n1830);
xnor_1 g01454(new_n1830, new_n1798_1, new_n1831);
xnor_1 g01455(new_n1831, new_n1796, new_n1832);
not_1  g01456(n7236, new_n1833);
nor_1  g01457(new_n753_1, new_n1833, new_n1834);
not_1  g01458(n3992, new_n1835_1);
nor_1  g01459(new_n697, new_n1835_1, new_n1836);
not_1  g01460(n8384, new_n1837);
nor_1  g01461(new_n1837, new_n384, new_n1838);
not_1  g01462(new_n1838, new_n1839);
nor_1  g01463(new_n1833, new_n764, new_n1840);
not_1  g01464(new_n1840, new_n1841);
nand_1 g01465(new_n1841, new_n1839, new_n1842);
nand_1 g01466(new_n1842, new_n1836, new_n1843);
nand_1 g01467(new_n1840, new_n1838, new_n1844);
nand_1 g01468(new_n1844, new_n1843, new_n1845);
xnor_1 g01469(new_n1845, new_n1834, new_n1846);
not_1  g01470(new_n1846, new_n1847_1);
nand_1 g01471(n8028, n6358, new_n1848);
nand_1 g01472(n10848, n8384, new_n1849);
nand_1 g01473(n3992, n1980, new_n1850);
xnor_1 g01474(new_n1850, new_n1849, new_n1851);
xnor_1 g01475(new_n1851, new_n1848, new_n1852);
not_1  g01476(new_n1852, new_n1853);
nand_1 g01477(new_n1853, new_n1847_1, new_n1854);
nand_1 g01478(new_n1852, new_n1846, new_n1855);
nand_1 g01479(new_n1855, new_n1854, new_n1856);
not_1  g01480(new_n1856, new_n1857);
and_1  g01481(new_n1844, new_n1842, new_n1858);
nand_1 g01482(n10848, n7236, new_n1859);
not_1  g01483(new_n1859, new_n1860);
nand_1 g01484(n8028, n3992, new_n1861);
not_1  g01485(new_n1861, new_n1862);
nand_1 g01486(new_n1862, new_n1860, new_n1863);
nor_1  g01487(new_n1863, new_n1858, new_n1864);
nand_1 g01488(new_n1864, new_n1857, new_n1865);
not_1  g01489(n6358, new_n1866);
nor_1  g01490(new_n697, new_n1866, new_n1867);
nand_1 g01491(n8384, n1980, new_n1868);
nand_1 g01492(n8028, n5198, new_n1869);
xnor_1 g01493(new_n1869, new_n1868, new_n1870);
xnor_1 g01494(new_n1870, new_n1867, new_n1871);
nor_1  g01495(new_n753_1, new_n1835_1, new_n1872);
not_1  g01496(new_n1872, new_n1873);
nand_1 g01497(new_n1850, new_n1849, new_n1874);
not_1  g01498(new_n1874, new_n1875);
not_1  g01499(new_n1848, new_n1876);
nor_1  g01500(new_n1851, new_n1876, new_n1877);
nor_1  g01501(new_n1877, new_n1875, new_n1878);
xnor_1 g01502(new_n1878, new_n1873, new_n1879);
xnor_1 g01503(new_n1879, new_n1871, new_n1880);
not_1  g01504(new_n1880, new_n1881);
nor_1  g01505(new_n790, new_n1833, new_n1882);
nand_1 g01506(new_n1845, new_n1834, new_n1883);
nand_1 g01507(new_n1854, new_n1883, new_n1884);
xnor_1 g01508(new_n1884, new_n1882, new_n1885);
nor_1  g01509(new_n1885, new_n1881, new_n1886);
not_1  g01510(new_n1886, new_n1887);
nand_1 g01511(new_n1885, new_n1881, new_n1888);
nand_1 g01512(new_n1888, new_n1887, new_n1889);
not_1  g01513(new_n1889, new_n1890);
nor_1  g01514(new_n1890, new_n1865, new_n1891);
nor_1  g01515(new_n1833, new_n915, new_n1892);
not_1  g01516(new_n1892, new_n1893);
nand_1 g01517(new_n1878, new_n1872, new_n1894);
nand_1 g01518(new_n1879, new_n1871, new_n1895);
nand_1 g01519(new_n1895, new_n1894, new_n1896);
nor_1  g01520(new_n1837, new_n753_1, new_n1897);
not_1  g01521(new_n1897, new_n1898);
nor_1  g01522(new_n790, new_n1835_1, new_n1899);
not_1  g01523(new_n1899, new_n1900);
nor_1  g01524(new_n1900, new_n1898, new_n1901);
not_1  g01525(new_n1901, new_n1902);
nand_1 g01526(new_n1900, new_n1898, new_n1903);
nand_1 g01527(new_n1903, new_n1902, new_n1904);
xnor_1 g01528(new_n1904, new_n1896, new_n1905);
nand_1 g01529(n6358, n1980, new_n1906_1);
nand_1 g01530(new_n1869, new_n1868, new_n1907);
not_1  g01531(new_n1907, new_n1908);
nor_1  g01532(new_n1870, new_n1867, new_n1909);
nor_1  g01533(new_n1909, new_n1908, new_n1910);
xnor_1 g01534(new_n1910, new_n1906_1, new_n1911);
nand_1 g01535(n10848, n5198, new_n1912);
nand_1 g01536(n8028, n1471, new_n1913);
xnor_1 g01537(new_n1913, new_n1912, new_n1914);
xnor_1 g01538(new_n1914, new_n1911, new_n1915);
xnor_1 g01539(new_n1915, new_n1905, new_n1916);
nor_1  g01540(new_n1884, new_n1882, new_n1917);
nor_1  g01541(new_n1886, new_n1917, new_n1918);
xnor_1 g01542(new_n1918, new_n1916, new_n1919);
xnor_1 g01543(new_n1919, new_n1893, new_n1920);
xnor_1 g01544(new_n1920, new_n1891, new_n1921);
nand_1 g01545(n4805, n2802, new_n1922);
not_1  g01546(n5283, new_n1923);
nor_1  g01547(new_n1923, new_n667, new_n1924);
not_1  g01548(n4805, new_n1925);
nor_1  g01549(new_n1925, new_n869, new_n1926);
nand_1 g01550(new_n1926, new_n1924, new_n1927);
not_1  g01551(new_n1924, new_n1928);
not_1  g01552(new_n1926, new_n1929);
nand_1 g01553(new_n1929, new_n1928, new_n1930);
not_1  g01554(n11478, new_n1931);
nor_1  g01555(new_n1931, new_n711, new_n1932);
nand_1 g01556(new_n1932, new_n1930, new_n1933);
nand_1 g01557(new_n1933, new_n1927, new_n1934);
xnor_1 g01558(new_n1934, new_n1922, new_n1935);
nand_1 g01559(n1564, n137, new_n1936);
nand_1 g01560(n5283, n1512, new_n1937);
nand_1 g01561(n11478, n533, new_n1938);
xnor_1 g01562(new_n1938, new_n1937, new_n1939);
xnor_1 g01563(new_n1939, new_n1936, new_n1940);
xnor_1 g01564(new_n1940, new_n1935, new_n1941);
xnor_1 g01565(new_n1926, new_n1928, new_n1942);
nand_1 g01566(n4805, n1512, new_n1943);
not_1  g01567(new_n1943, new_n1944);
nand_1 g01568(n11478, n1564, new_n1945);
not_1  g01569(new_n1945, new_n1946);
nand_1 g01570(new_n1946, new_n1944, new_n1947);
nor_1  g01571(new_n1947, new_n1942, new_n1948);
nand_1 g01572(new_n1948, new_n1941, new_n1949);
nor_1  g01573(new_n820, new_n1925, new_n1950);
not_1  g01574(new_n1950, new_n1951);
nor_1  g01575(new_n1931, new_n735, new_n1952);
nand_1 g01576(new_n1938, new_n1937, new_n1953);
not_1  g01577(new_n1953, new_n1954);
not_1  g01578(new_n1936, new_n1955);
nor_1  g01579(new_n1939, new_n1955, new_n1956);
nor_1  g01580(new_n1956, new_n1954, new_n1957);
xnor_1 g01581(new_n1957, new_n1952, new_n1958);
not_1  g01582(n137, new_n1959);
nor_1  g01583(new_n711, new_n1959, new_n1960);
nand_1 g01584(n5283, n533, new_n1961);
nand_1 g01585(n6294, n1564, new_n1962);
xnor_1 g01586(new_n1962, new_n1961, new_n1963);
nor_1  g01587(new_n1963, new_n1960, new_n1964);
not_1  g01588(new_n1964, new_n1965);
nand_1 g01589(new_n1963, new_n1960, new_n1966);
nand_1 g01590(new_n1966, new_n1965, new_n1967);
xnor_1 g01591(new_n1967, new_n1958, new_n1968);
xnor_1 g01592(new_n1968, new_n1951, new_n1969);
not_1  g01593(new_n1922, new_n1970);
nand_1 g01594(new_n1934, new_n1970, new_n1971);
not_1  g01595(new_n1971, new_n1972);
not_1  g01596(new_n1935, new_n1973);
nor_1  g01597(new_n1940, new_n1973, new_n1974);
nor_1  g01598(new_n1974, new_n1972, new_n1975);
nand_1 g01599(new_n1975, new_n1969, new_n1976);
not_1  g01600(new_n1976, new_n1977);
nor_1  g01601(new_n1975, new_n1969, new_n1978);
nor_1  g01602(new_n1978, new_n1977, new_n1979);
nor_1  g01603(new_n1979, new_n1949, new_n1980_1);
nor_1  g01604(new_n867, new_n1925, new_n1981);
nor_1  g01605(new_n869, new_n1959, new_n1982);
not_1  g01606(new_n1982, new_n1983);
nand_1 g01607(n6294, n1512, new_n1984);
nand_1 g01608(n6797, n1564, new_n1985);
xnor_1 g01609(new_n1985, new_n1984, new_n1986);
xnor_1 g01610(new_n1986, new_n1983, new_n1987);
not_1  g01611(new_n1987, new_n1988);
nand_1 g01612(new_n1962, new_n1961, new_n1989);
nand_1 g01613(new_n1965, new_n1989, new_n1990);
xnor_1 g01614(new_n1990, new_n1988, new_n1991);
nand_1 g01615(n11478, n6806, new_n1992);
nand_1 g01616(n5283, n2802, new_n1993);
nor_1  g01617(new_n1993, new_n1992, new_n1994);
not_1  g01618(new_n1994, new_n1995);
nand_1 g01619(new_n1993, new_n1992, new_n1996);
nand_1 g01620(new_n1996, new_n1995, new_n1997);
xnor_1 g01621(new_n1997, new_n1991, new_n1998);
nand_1 g01622(new_n1957, new_n1952, new_n1999);
not_1  g01623(new_n1967, new_n2000);
nor_1  g01624(new_n2000, new_n1958, new_n2001);
not_1  g01625(new_n2001, new_n2002);
nand_1 g01626(new_n2002, new_n1999, new_n2003);
nand_1 g01627(new_n2003, new_n1998, new_n2004);
not_1  g01628(new_n2004, new_n2005);
nor_1  g01629(new_n2003, new_n1998, new_n2006);
nor_1  g01630(new_n2006, new_n2005, new_n2007);
nor_1  g01631(new_n1968, new_n1950, new_n2008);
not_1  g01632(new_n2008, new_n2009);
nand_1 g01633(new_n1976, new_n2009, new_n2010);
xnor_1 g01634(new_n2010, new_n2007, new_n2011);
xnor_1 g01635(new_n2011, new_n1981, new_n2012);
xnor_1 g01636(new_n2012, new_n1980_1, new_n2013);
xnor_1 g01637(new_n2013, new_n1921, new_n2014);
not_1  g01638(new_n2014, new_n2015);
xnor_1 g01639(new_n1889, new_n1865, new_n2016);
not_1  g01640(new_n2016, new_n2017);
xnor_1 g01641(new_n1948, new_n1941, new_n2018);
xnor_1 g01642(new_n1864, new_n1856, new_n2019);
not_1  g01643(new_n2019, new_n2020);
nand_1 g01644(new_n2020, new_n2018, new_n2021);
nor_1  g01645(new_n1354, new_n1353_1, new_n2022);
not_1  g01646(new_n2022, new_n2023);
nand_1 g01647(new_n1945, new_n1943, new_n2024_1);
nand_1 g01648(new_n2024_1, new_n1947, new_n2025);
nand_1 g01649(new_n2025, new_n2023, new_n2026);
xnor_1 g01650(new_n2025, new_n2022, new_n2027);
nand_1 g01651(new_n1861, new_n1859, new_n2028);
nand_1 g01652(new_n2028, new_n1863, new_n2029);
nand_1 g01653(new_n2029, new_n2027, new_n2030);
nand_1 g01654(new_n2030, new_n2026, new_n2031);
and_1  g01655(new_n1932, new_n1353_1, new_n2032);
nor_1  g01656(new_n2032, new_n1942, new_n2033);
not_1  g01657(new_n1353_1, new_n2034);
nor_1  g01658(new_n1933, new_n2034, new_n2035);
nor_1  g01659(new_n2035, new_n2033, new_n2036);
not_1  g01660(new_n2036, new_n2037);
nand_1 g01661(new_n2037, new_n2031, new_n2038);
xnor_1 g01662(new_n2036, new_n2031, new_n2039);
nand_1 g01663(new_n1836, new_n1354, new_n2040);
not_1  g01664(new_n2040, new_n2041);
nor_1  g01665(new_n2041, new_n1858, new_n2042);
nor_1  g01666(new_n1843, new_n1355, new_n2043);
nor_1  g01667(new_n2043, new_n2042, new_n2044);
not_1  g01668(new_n2044, new_n2045);
nand_1 g01669(new_n2045, new_n2039, new_n2046);
nand_1 g01670(new_n2046, new_n2038, new_n2047);
xnor_1 g01671(new_n2019, new_n2018, new_n2048);
nand_1 g01672(new_n2048, new_n2047, new_n2049);
nand_1 g01673(new_n2049, new_n2021, new_n2050);
nand_1 g01674(new_n2050, new_n2017, new_n2051);
xnor_1 g01675(new_n1979, new_n1949, new_n2052);
xnor_1 g01676(new_n2050, new_n2016, new_n2053);
nand_1 g01677(new_n2053, new_n2052, new_n2054);
nand_1 g01678(new_n2054, new_n2051, new_n2055);
xnor_1 g01679(new_n2055, new_n2015, new_n2056);
nand_1 g01680(new_n2056, new_n1832, new_n2057);
not_1  g01681(new_n1832, new_n2058);
xnor_1 g01682(new_n2056, new_n2058, new_n2059);
xnor_1 g01683(new_n1795, new_n1765, new_n2060);
not_1  g01684(new_n2052, new_n2061);
xnor_1 g01685(new_n2053, new_n2061, new_n2062);
nor_1  g01686(new_n2062, new_n2060, new_n2063);
not_1  g01687(new_n2063, new_n2064);
not_1  g01688(new_n2060, new_n2065);
xnor_1 g01689(new_n2062, new_n2065, new_n2066);
xor_1  g01690(new_n1764, new_n1758, new_n2067);
not_1  g01691(new_n2067, new_n2068);
xnor_1 g01692(new_n2048, new_n2047, new_n2069);
not_1  g01693(new_n2069, new_n2070);
nor_1  g01694(new_n2070, new_n2068, new_n2071);
not_1  g01695(new_n2071, new_n2072);
nor_1  g01696(new_n2069, new_n2067, new_n2073);
nor_1  g01697(new_n2073, new_n2071, new_n2074);
xnor_1 g01698(new_n2044, new_n2039, new_n2075);
not_1  g01699(new_n2075, new_n2076);
nand_1 g01700(new_n1736, new_n1352, new_n2077);
nor_1  g01701(new_n2077, new_n1734, new_n2078);
not_1  g01702(new_n2078, new_n2079);
nand_1 g01703(new_n2077, new_n1760, new_n2080);
nand_1 g01704(new_n2080, new_n2079, new_n2081);
and_1  g01705(new_n2081, new_n2076, new_n2082);
xnor_1 g01706(new_n2081, new_n2076, new_n2083);
xnor_1 g01707(new_n2029, new_n2027, new_n2084);
not_1  g01708(new_n2084, new_n2085);
xnor_1 g01709(new_n1762, new_n1761, new_n2086);
nor_1  g01710(new_n2086, new_n2085, new_n2087_1);
xnor_1 g01711(new_n2086, new_n2084, new_n2088);
nand_1 g01712(new_n2088, new_n1358, new_n2089);
not_1  g01713(new_n2089, new_n2090);
nor_1  g01714(new_n2090, new_n2087_1, new_n2091);
nor_1  g01715(new_n2091, new_n2083, new_n2092);
nor_1  g01716(new_n2092, new_n2082, new_n2093);
not_1  g01717(new_n2093, new_n2094);
nand_1 g01718(new_n2094, new_n2074, new_n2095);
nand_1 g01719(new_n2095, new_n2072, new_n2096_1);
nand_1 g01720(new_n2096_1, new_n2066, new_n2097);
nand_1 g01721(new_n2097, new_n2064, new_n2098);
not_1  g01722(new_n2098, new_n2099);
nand_1 g01723(new_n2099, new_n2059, new_n2100);
nand_1 g01724(new_n2100, new_n2057, new_n2101);
not_1  g01725(new_n1803, new_n2102);
nor_1  g01726(new_n1806, new_n2102, new_n2103);
not_1  g01727(new_n2103, new_n2104);
nand_1 g01728(new_n1809, new_n1807, new_n2105);
nand_1 g01729(new_n2105, new_n2104, new_n2106);
nand_1 g01730(n9400, n4928, new_n2107);
nand_1 g01731(n4141, n2464, new_n2108);
nand_1 g01732(n8236, n6877, new_n2109);
nor_1  g01733(new_n2109, new_n2108, new_n2110);
nand_1 g01734(new_n2109, new_n2108, new_n2111);
not_1  g01735(new_n2111, new_n2112);
nor_1  g01736(new_n2112, new_n2110, new_n2113);
xor_1  g01737(new_n2113, new_n2107, new_n2114);
xnor_1 g01738(new_n2114, new_n2106, new_n2115);
nor_1  g01739(new_n1805, new_n1804, new_n2116);
nor_1  g01740(new_n1747, new_n551, new_n2117);
xor_1  g01741(new_n2117, new_n2116, new_n2118);
not_1  g01742(n4203, new_n2119);
nor_1  g01743(new_n564, new_n2119, new_n2120);
nand_1 g01744(n4187, n1209, new_n2121);
nand_1 g01745(n12753, n7354, new_n2122);
xnor_1 g01746(new_n2122, new_n2121, new_n2123);
xor_1  g01747(new_n2123, new_n2120, new_n2124);
xnor_1 g01748(new_n2124, new_n2118, new_n2125);
xnor_1 g01749(new_n2125, new_n2115, new_n2126);
nand_1 g01750(new_n1821, new_n1811, new_n2127);
not_1  g01751(new_n2127, new_n2128);
nand_1 g01752(new_n2128, new_n1817, new_n2129);
nand_1 g01753(new_n2127, new_n1818, new_n2130);
nand_1 g01754(new_n2130, new_n2129, new_n2131_1);
nand_1 g01755(new_n2131_1, new_n1824, new_n2132);
xnor_1 g01756(new_n2132, new_n2126, new_n2133);
xnor_1 g01757(new_n2133, new_n1827, new_n2134);
nand_1 g01758(new_n1830, new_n1797, new_n2135);
nand_1 g01759(new_n1831, new_n1796, new_n2136);
nand_1 g01760(new_n2136, new_n2135, new_n2137);
xnor_1 g01761(new_n2137, new_n2134, new_n2138);
not_1  g01762(new_n1918, new_n2139);
nor_1  g01763(new_n2139, new_n1916, new_n2140);
not_1  g01764(new_n1910, new_n2141);
nand_1 g01765(new_n2141, new_n1906_1, new_n2142);
nand_1 g01766(new_n1914, new_n1911, new_n2143);
nand_1 g01767(new_n2143, new_n2142, new_n2144);
nor_1  g01768(new_n915, new_n1835_1, new_n2145);
nand_1 g01769(n12704, n8384, new_n2146);
nand_1 g01770(n7236, n4903, new_n2147);
xnor_1 g01771(new_n2147, new_n2146, new_n2148);
xnor_1 g01772(new_n2148, new_n2145, new_n2149);
xnor_1 g01773(new_n2149, new_n2144, new_n2150);
nor_1  g01774(new_n1913, new_n1912, new_n2151);
nor_1  g01775(new_n753_1, new_n1866, new_n2152);
xor_1  g01776(new_n2152, new_n2151, new_n2153);
not_1  g01777(n1471, new_n2154);
nor_1  g01778(new_n697, new_n2154, new_n2155);
nand_1 g01779(n5198, n1980, new_n2156);
nand_1 g01780(n8028, n7646, new_n2157);
xnor_1 g01781(new_n2157, new_n2156, new_n2158);
xnor_1 g01782(new_n2158, new_n2155, new_n2159);
not_1  g01783(new_n2159, new_n2160);
xnor_1 g01784(new_n2160, new_n2153, new_n2161);
xnor_1 g01785(new_n2161, new_n2150, new_n2162);
not_1  g01786(new_n1904, new_n2163);
nand_1 g01787(new_n2163, new_n1896, new_n2164);
nand_1 g01788(new_n1915, new_n1905, new_n2165);
not_1  g01789(new_n2165, new_n2166);
nand_1 g01790(new_n2166, new_n1901, new_n2167);
nand_1 g01791(new_n2165, new_n1902, new_n2168);
nand_1 g01792(new_n2168, new_n2167, new_n2169);
nand_1 g01793(new_n2169, new_n2164, new_n2170);
xnor_1 g01794(new_n2170, new_n2162, new_n2171);
xnor_1 g01795(new_n2171, new_n2140, new_n2172);
nand_1 g01796(new_n1919, new_n1892, new_n2173);
nand_1 g01797(new_n1920, new_n1891, new_n2174);
nand_1 g01798(new_n2174, new_n2173, new_n2175);
xnor_1 g01799(new_n2175, new_n2172, new_n2176);
not_1  g01800(new_n2176, new_n2177);
nand_1 g01801(new_n2011, new_n1981, new_n2178);
not_1  g01802(new_n2012, new_n2179);
nand_1 g01803(new_n2179, new_n1980_1, new_n2180);
nand_1 g01804(new_n2180, new_n2178, new_n2181);
not_1  g01805(new_n2007, new_n2182);
nor_1  g01806(new_n2010, new_n2182, new_n2183);
nor_1  g01807(new_n1986, new_n1983, new_n2184);
nor_1  g01808(new_n1990, new_n1987, new_n2185);
nor_1  g01809(new_n2185, new_n2184, new_n2186);
nor_1  g01810(new_n1931, new_n867, new_n2187);
nor_1  g01811(new_n820, new_n1923, new_n2188);
not_1  g01812(new_n2188, new_n2189);
not_1  g01813(n12044, new_n2190);
nor_1  g01814(new_n2190, new_n1925, new_n2191);
not_1  g01815(new_n2191, new_n2192);
nand_1 g01816(new_n2192, new_n2189, new_n2193);
nand_1 g01817(new_n2191, new_n2188, new_n2194);
nand_1 g01818(new_n2194, new_n2193, new_n2195);
xnor_1 g01819(new_n2195, new_n2187, new_n2196);
not_1  g01820(new_n2196, new_n2197);
nand_1 g01821(new_n2197, new_n2186, new_n2198);
not_1  g01822(new_n2186, new_n2199);
nand_1 g01823(new_n2196, new_n2199, new_n2200);
nand_1 g01824(new_n2200, new_n2198, new_n2201);
nor_1  g01825(new_n1985, new_n1984, new_n2202);
nor_1  g01826(new_n735, new_n1959, new_n2203);
xnor_1 g01827(new_n2203, new_n2202, new_n2204);
not_1  g01828(n6797, new_n2205);
nor_1  g01829(new_n2205, new_n711, new_n2206);
nand_1 g01830(n6294, n533, new_n2207);
nand_1 g01831(n3146, n1564, new_n2208);
xnor_1 g01832(new_n2208, new_n2207, new_n2209);
xor_1  g01833(new_n2209, new_n2206, new_n2210);
nand_1 g01834(new_n2210, new_n2204, new_n2211);
not_1  g01835(new_n2204, new_n2212);
not_1  g01836(new_n2210, new_n2213);
nand_1 g01837(new_n2213, new_n2212, new_n2214);
nand_1 g01838(new_n2214, new_n2211, new_n2215);
xnor_1 g01839(new_n2215, new_n2201, new_n2216);
not_1  g01840(new_n1997, new_n2217);
nand_1 g01841(new_n2217, new_n1991, new_n2218);
nand_1 g01842(new_n2005, new_n1994, new_n2219);
nand_1 g01843(new_n2004, new_n1995, new_n2220);
nand_1 g01844(new_n2220, new_n2219, new_n2221);
nand_1 g01845(new_n2221, new_n2218, new_n2222);
xnor_1 g01846(new_n2222, new_n2216, new_n2223);
xnor_1 g01847(new_n2223, new_n2183, new_n2224);
xnor_1 g01848(new_n2224, new_n2181, new_n2225);
not_1  g01849(new_n2225, new_n2226_1);
nand_1 g01850(new_n2226_1, new_n2177, new_n2227);
nand_1 g01851(new_n2225, new_n2176, new_n2228);
nand_1 g01852(new_n2228, new_n2227, new_n2229);
not_1  g01853(new_n2013, new_n2230);
nand_1 g01854(new_n2230, new_n1921, new_n2231);
nand_1 g01855(new_n2055, new_n2014, new_n2232);
nand_1 g01856(new_n2232, new_n2231, new_n2233);
xnor_1 g01857(new_n2233, new_n2229, new_n2234);
xnor_1 g01858(new_n2234, new_n2138, new_n2235);
xnor_1 g01859(new_n2235, new_n2101, new_n2236);
not_1  g01860(new_n2236, new_n2237);
nand_1 g01861(new_n2237, new_n1725, new_n2238);
xnor_1 g01862(new_n2236, new_n1725, new_n2239);
xor_1  g01863(new_n1721, new_n1719, new_n2240);
xnor_1 g01864(new_n2098, new_n2059, new_n2241);
not_1  g01865(new_n2241, new_n2242);
nand_1 g01866(new_n2242, new_n2240, new_n2243);
xnor_1 g01867(new_n1717, new_n1716, new_n2244);
not_1  g01868(new_n2097, new_n2245);
nor_1  g01869(new_n2096_1, new_n2066, new_n2246);
nor_1  g01870(new_n2246, new_n2245, new_n2247);
nor_1  g01871(new_n2247, new_n2244, new_n2248);
xnor_1 g01872(new_n2247, new_n2244, new_n2249);
xor_1  g01873(new_n1715, new_n1710, new_n2250);
xnor_1 g01874(new_n2093, new_n2074, new_n2251);
nor_1  g01875(new_n2251, new_n2250, new_n2252);
xor_1  g01876(new_n2091, new_n2083, new_n2253_1);
nor_1  g01877(new_n1622, new_n1349, new_n2254);
nor_1  g01878(new_n2254, new_n1711, new_n2255);
not_1  g01879(new_n1629, new_n2256);
nor_1  g01880(new_n2256, new_n1349, new_n2257);
nor_1  g01881(new_n2257, new_n2255, new_n2258);
nor_1  g01882(new_n2258, new_n2253_1, new_n2259);
xnor_1 g01883(new_n2258, new_n2253_1, new_n2260);
not_1  g01884(new_n1712, new_n2261);
xnor_1 g01885(new_n1713, new_n2261, new_n2262);
nor_1  g01886(new_n2262, new_n1362, new_n2263);
nor_1  g01887(new_n2088, new_n1358, new_n2264);
nor_1  g01888(new_n2264, new_n2090, new_n2265);
xnor_1 g01889(new_n2262, new_n1362, new_n2266);
nor_1  g01890(new_n2266, new_n2265, new_n2267);
nor_1  g01891(new_n2267, new_n2263, new_n2268);
nor_1  g01892(new_n2268, new_n2260, new_n2269);
nor_1  g01893(new_n2269, new_n2259, new_n2270);
xnor_1 g01894(new_n2251, new_n2250, new_n2271);
nor_1  g01895(new_n2271, new_n2270, new_n2272);
nor_1  g01896(new_n2272, new_n2252, new_n2273);
nor_1  g01897(new_n2273, new_n2249, new_n2274);
nor_1  g01898(new_n2274, new_n2248, new_n2275);
xnor_1 g01899(new_n2241, new_n2240, new_n2276);
nand_1 g01900(new_n2276, new_n2275, new_n2277);
nand_1 g01901(new_n2277, new_n2243, new_n2278_1);
nand_1 g01902(new_n2278_1, new_n2239, new_n2279);
nand_1 g01903(new_n2279, new_n2238, new_n2280);
nand_1 g01904(new_n2234, new_n2138, new_n2281);
not_1  g01905(new_n2235, new_n2282);
nand_1 g01906(new_n2282, new_n2101, new_n2283);
nand_1 g01907(new_n2283, new_n2281, new_n2284);
not_1  g01908(new_n2229, new_n2285);
nand_1 g01909(new_n2233, new_n2285, new_n2286);
nand_1 g01910(new_n2286, new_n2227, new_n2287);
nand_1 g01911(new_n1703, new_n1706, new_n2288);
nand_1 g01912(new_n1723, new_n1704, new_n2289);
nand_1 g01913(new_n2289, new_n2288, new_n2290);
nand_1 g01914(new_n2171, new_n2140, new_n2291);
not_1  g01915(new_n2172, new_n2292);
nand_1 g01916(new_n2175, new_n2292, new_n2293);
nand_1 g01917(new_n2293, new_n2291, new_n2294);
xnor_1 g01918(new_n2294, new_n2290, new_n2295);
not_1  g01919(new_n2162, new_n2296);
nand_1 g01920(new_n2170, new_n2296, new_n2297);
nand_1 g01921(new_n2297, new_n2167, new_n2298);
nand_1 g01922(new_n2203, new_n2202, new_n2299);
nand_1 g01923(new_n2214, new_n2299, new_n2300);
nand_1 g01924(n7862, n615, new_n2301_1);
nand_1 g01925(n4903, n3992, new_n2302);
nand_1 g01926(n6806, n137, new_n2303);
xnor_1 g01927(new_n2303, new_n2302, new_n2304);
xor_1  g01928(new_n2304, new_n2301_1, new_n2305);
xnor_1 g01929(new_n2305, new_n2300, new_n2306);
nand_1 g01930(n6797, n533, new_n2307);
nand_1 g01931(n8384, n5814, new_n2308);
xnor_1 g01932(new_n2308, new_n2307, new_n2309);
nand_1 g01933(n12044, n11478, new_n2310);
nand_1 g01934(n7294, n5198, new_n2311);
xnor_1 g01935(new_n2311, new_n2310, new_n2312);
xnor_1 g01936(new_n2312, new_n2309, new_n2313);
nand_1 g01937(new_n2193, new_n2187, new_n2314);
nand_1 g01938(new_n2314, new_n2194, new_n2315);
xnor_1 g01939(new_n2315, new_n2313, new_n2316_1);
nand_1 g01940(n10174, n7354, new_n2317);
nand_1 g01941(n4928, n2464, new_n2318);
nand_1 g01942(n11311, n4141, new_n2319);
xnor_1 g01943(new_n2319, new_n2318, new_n2320);
nand_1 g01944(n4005, n3172, new_n2321);
nand_1 g01945(n7236, n1906, new_n2322);
xnor_1 g01946(new_n2322, new_n2321, new_n2323);
xnor_1 g01947(new_n2323, new_n2320, new_n2324);
xor_1  g01948(new_n2324, new_n2317, new_n2325);
xnor_1 g01949(new_n2325, new_n2316_1, new_n2326);
xnor_1 g01950(new_n2326, new_n2306, new_n2327);
xnor_1 g01951(new_n2327, new_n2298, new_n2328);
not_1  g01952(new_n2149, new_n2329);
nand_1 g01953(new_n2329, new_n2144, new_n2330);
not_1  g01954(new_n2161, new_n2331);
nand_1 g01955(new_n2331, new_n2150, new_n2332);
nand_1 g01956(new_n2332, new_n2330, new_n2333);
not_1  g01957(n9080, new_n2334);
nor_1  g01958(new_n2334, new_n413, new_n2335);
nand_1 g01959(new_n1685, new_n1684, new_n2336);
not_1  g01960(new_n2336, new_n2337);
nor_1  g01961(new_n1686, new_n1683, new_n2338);
nor_1  g01962(new_n2338, new_n2337, new_n2339);
nand_1 g01963(n5240, n2508, new_n2340);
nand_1 g01964(n11757, n2585, new_n2341);
nand_1 g01965(n12706, n1333, new_n2342);
xnor_1 g01966(new_n2342, new_n2341, new_n2343);
xnor_1 g01967(new_n2343, new_n2340, new_n2344);
xnor_1 g01968(new_n2344, new_n2339, new_n2345);
xnor_1 g01969(new_n2345, new_n2335, new_n2346);
xnor_1 g01970(new_n2346, new_n2333, new_n2347_1);
xnor_1 g01971(new_n2347_1, new_n2328, new_n2348);
not_1  g01972(new_n2126, new_n2349);
nand_1 g01973(new_n2132, new_n2349, new_n2350);
nand_1 g01974(new_n2350, new_n2129, new_n2351);
nor_1  g01975(new_n1676, new_n1667, new_n2352);
not_1  g01976(new_n1702, new_n2353);
nor_1  g01977(new_n2353, new_n1678, new_n2354);
nor_1  g01978(new_n2354, new_n2352, new_n2355);
xnor_1 g01979(new_n2355, new_n2351, new_n2356);
not_1  g01980(new_n2106, new_n2357);
nand_1 g01981(new_n2114, new_n2357, new_n2358);
not_1  g01982(new_n2125, new_n2359);
nand_1 g01983(new_n2359, new_n2115, new_n2360);
nand_1 g01984(new_n2360, new_n2358, new_n2361);
nand_1 g01985(n12704, n6358, new_n2362);
not_1  g01986(n3146, new_n2363);
nor_1  g01987(new_n2363, new_n711, new_n2364);
xnor_1 g01988(new_n2364, new_n2362, new_n2365);
nand_1 g01989(n5105, n4187, new_n2366);
nand_1 g01990(n6294, n2802, new_n2367);
xnor_1 g01991(new_n2367, new_n2366, new_n2368);
nand_1 g01992(n9400, n8236, new_n2369);
nand_1 g01993(n1980, n1471, new_n2370);
xnor_1 g01994(new_n2370, new_n2369, new_n2371);
xnor_1 g01995(new_n2371, new_n2368, new_n2372);
xnor_1 g01996(new_n2372, new_n2365, new_n2373);
nand_1 g01997(n12720, n11821, new_n2374);
nand_1 g01998(n4938, n1564, new_n2375);
nand_1 g01999(n5694, n4805, new_n2376);
xnor_1 g02000(new_n2376, new_n2375, new_n2377);
xnor_1 g02001(new_n2377, new_n2374, new_n2378);
xnor_1 g02002(new_n2378, new_n2373, new_n2379);
nand_1 g02003(new_n2147, new_n2146, new_n2380);
not_1  g02004(new_n2380, new_n2381);
nor_1  g02005(new_n2148, new_n2145, new_n2382);
nor_1  g02006(new_n2382, new_n2381, new_n2383_1);
nand_1 g02007(new_n1680, new_n1679, new_n2384);
nand_1 g02008(new_n1687, new_n1681, new_n2385);
nand_1 g02009(new_n2385, new_n2384, new_n2386);
xnor_1 g02010(new_n2386, new_n2383_1, new_n2387);
xnor_1 g02011(new_n2387, new_n2379, new_n2388);
xnor_1 g02012(new_n2388, new_n2361, new_n2389);
not_1  g02013(new_n2216, new_n2390);
nand_1 g02014(new_n2222, new_n2390, new_n2391);
nand_1 g02015(new_n2391, new_n2219, new_n2392);
not_1  g02016(new_n2201, new_n2393_1);
nand_1 g02017(new_n2215, new_n2393_1, new_n2394);
nand_1 g02018(new_n2394, new_n2198, new_n2395);
nand_1 g02019(new_n2152, new_n2151, new_n2396);
nand_1 g02020(new_n2159, new_n2153, new_n2397);
nand_1 g02021(new_n2397, new_n2396, new_n2398);
nor_1  g02022(new_n2119, new_n557, new_n2399);
nand_1 g02023(n6826, n6038, new_n2400);
nand_1 g02024(n5283, n5069, new_n2401);
xnor_1 g02025(new_n2401, new_n2400, new_n2402);
xnor_1 g02026(new_n2402, new_n2399, new_n2403);
xnor_1 g02027(new_n2403, new_n2398, new_n2404);
nand_1 g02028(new_n2208, new_n2207, new_n2405);
not_1  g02029(new_n2405, new_n2406);
nor_1  g02030(new_n2209, new_n2206, new_n2407);
nor_1  g02031(new_n2407, new_n2406, new_n2408);
nand_1 g02032(new_n2157, new_n2156, new_n2409);
not_1  g02033(new_n2409, new_n2410);
nor_1  g02034(new_n2158, new_n2155, new_n2411);
nor_1  g02035(new_n2411, new_n2410, new_n2412);
nor_1  g02036(new_n2112, new_n2107, new_n2413);
nor_1  g02037(new_n2413, new_n2110, new_n2414);
xnor_1 g02038(new_n2414, new_n2412, new_n2415);
xnor_1 g02039(new_n2415, new_n2408, new_n2416);
xnor_1 g02040(new_n2416, new_n2404, new_n2417);
xnor_1 g02041(new_n2417, new_n2395, new_n2418);
xnor_1 g02042(new_n2418, new_n2392, new_n2419);
xnor_1 g02043(new_n2419, new_n2389, new_n2420);
xnor_1 g02044(new_n2420, new_n2356, new_n2421);
xnor_1 g02045(new_n2421, new_n2348, new_n2422);
xnor_1 g02046(new_n2422, new_n2295, new_n2423);
xnor_1 g02047(new_n2423, new_n2287, new_n2424);
nand_1 g02048(new_n2117, new_n2116, new_n2425_1);
not_1  g02049(new_n2124, new_n2426);
nand_1 g02050(new_n2426, new_n2118, new_n2427);
nand_1 g02051(new_n2427, new_n2425_1, new_n2428);
nand_1 g02052(n6877, n783, new_n2429);
nand_1 g02053(n8028, n4722, new_n2430);
xnor_1 g02054(new_n2430, new_n2429, new_n2431_1);
xnor_1 g02055(new_n2431_1, new_n2428, new_n2432);
nand_1 g02056(new_n2133, new_n1828, new_n2433_1);
nand_1 g02057(new_n2137, new_n2134, new_n2434_1);
nand_1 g02058(new_n2434_1, new_n2433_1, new_n2435);
nand_1 g02059(n10848, n7646, new_n2436);
xnor_1 g02060(new_n2436, new_n2435, new_n2437);
xnor_1 g02061(new_n2437, new_n2432, new_n2438);
nand_1 g02062(new_n2223, new_n2183, new_n2439);
not_1  g02063(new_n2224, new_n2440);
nand_1 g02064(new_n2440, new_n2181, new_n2441);
nand_1 g02065(new_n2441, new_n2439, new_n2442);
nand_1 g02066(new_n1700, new_n1690, new_n2443);
nand_1 g02067(new_n1701, new_n1688, new_n2444);
nand_1 g02068(new_n2444, new_n2443, new_n2445);
nand_1 g02069(new_n2122, new_n2121, new_n2446);
not_1  g02070(new_n2446, new_n2447);
nor_1  g02071(new_n2123, new_n2120, new_n2448);
nor_1  g02072(new_n2448, new_n2447, new_n2449);
not_1  g02073(n12753, new_n2450);
nor_1  g02074(new_n2450, new_n564, new_n2451);
nand_1 g02075(new_n1697, new_n1692, new_n2452);
nand_1 g02076(new_n2452, new_n1698, new_n2453);
xnor_1 g02077(new_n2453, new_n2451, new_n2454);
xnor_1 g02078(new_n2454, new_n2449, new_n2455);
xnor_1 g02079(new_n2455, new_n2445, new_n2456);
xnor_1 g02080(new_n2456, new_n2442, new_n2457);
xnor_1 g02081(new_n2457, new_n2438, new_n2458);
xnor_1 g02082(new_n2458, new_n2424, new_n2459);
xnor_1 g02083(new_n2459, new_n2284, new_n2460);
xnor_1 g02084(new_n2460, new_n2280, n671);
not_1  g02085(n11917, new_n2462);
nor_1  g02086(new_n2462, new_n395, new_n2463);
nand_1 g02087(n12705, n4921, new_n2464_1);
nand_1 g02088(n12025, n9956, new_n2465);
nand_1 g02089(new_n2465, new_n2464_1, new_n2466);
nor_1  g02090(new_n2465, new_n2464_1, new_n2467);
not_1  g02091(new_n2467, new_n2468);
nand_1 g02092(new_n2468, new_n2466, new_n2469);
xnor_1 g02093(new_n2469, new_n2463, new_n2470);
nand_1 g02094(n12705, n9956, new_n2471);
nand_1 g02095(n11917, n1097, new_n2472);
nand_1 g02096(new_n2472, new_n2471, new_n2473);
not_1  g02097(new_n2473, new_n2474);
nor_1  g02098(new_n2472, new_n2471, new_n2475);
not_1  g02099(n4921, new_n2476);
nor_1  g02100(new_n2476, new_n395, new_n2477);
nor_1  g02101(new_n2477, new_n2475, new_n2478);
nor_1  g02102(new_n2478, new_n2474, new_n2479);
xnor_1 g02103(new_n2479, new_n2470, new_n2480);
not_1  g02104(n2577, new_n2481);
nor_1  g02105(new_n424, new_n2481, new_n2482);
not_1  g02106(new_n2482, new_n2483);
not_1  g02107(n3842, new_n2484);
nor_1  g02108(new_n2484, new_n419, new_n2485);
not_1  g02109(new_n2485, new_n2486);
nor_1  g02110(new_n2486, new_n2483, new_n2487);
not_1  g02111(new_n2487, new_n2488);
nand_1 g02112(new_n2486, new_n2483, new_n2489);
nand_1 g02113(new_n2489, new_n2488, new_n2490);
xor_1  g02114(new_n2490, new_n2480, new_n2491);
nor_1  g02115(new_n424, new_n2484, new_n2492);
not_1  g02116(n9956, new_n2493);
nor_1  g02117(new_n2493, new_n395, new_n2494);
not_1  g02118(new_n2494, new_n2495);
nor_1  g02119(new_n2462, new_n424, new_n2496);
not_1  g02120(new_n2496, new_n2497);
nand_1 g02121(new_n2497, new_n2495, new_n2498_1);
not_1  g02122(new_n2498_1, new_n2499);
nor_1  g02123(new_n2497, new_n2495, new_n2500);
nor_1  g02124(new_n2476, new_n419, new_n2501);
nor_1  g02125(new_n2501, new_n2500, new_n2502);
nor_1  g02126(new_n2502, new_n2499, new_n2503);
nand_1 g02127(new_n2503, new_n2492, new_n2504);
not_1  g02128(new_n2504, new_n2505);
nor_1  g02129(new_n2503, new_n2492, new_n2506);
nor_1  g02130(new_n2506, new_n2505, new_n2507_1);
not_1  g02131(new_n2507_1, new_n2508_1);
not_1  g02132(new_n2475, new_n2509_1);
nand_1 g02133(new_n2509_1, new_n2473, new_n2510);
xnor_1 g02134(new_n2510, new_n2477, new_n2511);
not_1  g02135(new_n2511, new_n2512_1);
nor_1  g02136(new_n2512_1, new_n2508_1, new_n2513);
nor_1  g02137(new_n2513, new_n2505, new_n2514);
xnor_1 g02138(new_n2514, new_n2491, new_n2515_1);
nor_1  g02139(new_n456, new_n2481, new_n2516);
nor_1  g02140(new_n2511, new_n2507_1, new_n2517);
nor_1  g02141(new_n2517, new_n2513, new_n2518);
nor_1  g02142(new_n2518, new_n2516, new_n2519);
not_1  g02143(new_n2519, new_n2520);
not_1  g02144(new_n2516, new_n2521);
xnor_1 g02145(new_n2518, new_n2521, new_n2522_1);
nor_1  g02146(new_n456, new_n2484, new_n2523);
not_1  g02147(new_n2523, new_n2524);
nor_1  g02148(new_n2493, new_n419, new_n2525);
not_1  g02149(new_n2525, new_n2526);
nor_1  g02150(new_n2462, new_n456, new_n2527);
not_1  g02151(new_n2527, new_n2528);
nor_1  g02152(new_n2528, new_n2526, new_n2529);
nand_1 g02153(new_n2528, new_n2526, new_n2530_1);
not_1  g02154(new_n2530_1, new_n2531);
nor_1  g02155(new_n424, new_n2476, new_n2532);
not_1  g02156(new_n2532, new_n2533);
nor_1  g02157(new_n2533, new_n2531, new_n2534);
nor_1  g02158(new_n2534, new_n2529, new_n2535);
nor_1  g02159(new_n2535, new_n2524, new_n2536);
xnor_1 g02160(new_n2535, new_n2524, new_n2537);
nor_1  g02161(new_n2500, new_n2499, new_n2538);
xnor_1 g02162(new_n2538, new_n2501, new_n2539);
nor_1  g02163(new_n2539, new_n2537, new_n2540);
nor_1  g02164(new_n2540, new_n2536, new_n2541);
nand_1 g02165(new_n2541, new_n2522_1, new_n2542);
nand_1 g02166(new_n2542, new_n2520, new_n2543);
not_1  g02167(new_n2543, new_n2544);
nand_1 g02168(new_n2544, new_n2515_1, new_n2545);
not_1  g02169(new_n2463, new_n2546);
nand_1 g02170(new_n2469, new_n2546, new_n2547);
not_1  g02171(new_n2479, new_n2548);
nand_1 g02172(new_n2548, new_n2470, new_n2549);
nand_1 g02173(new_n2549, new_n2547, new_n2550);
not_1  g02174(n9637, new_n2551_1);
nor_1  g02175(new_n2551_1, new_n424, new_n2552);
nand_1 g02176(n2577, n1097, new_n2553);
nand_1 g02177(n5305, n1835, new_n2554);
xnor_1 g02178(new_n2554, new_n2553, new_n2555);
xnor_1 g02179(new_n2555, new_n2552, new_n2556);
xnor_1 g02180(new_n2556, new_n2550, new_n2557);
nor_1  g02181(new_n395, new_n2484, new_n2558_1);
not_1  g02182(new_n2558_1, new_n2559);
nand_1 g02183(new_n2559, new_n2468, new_n2560);
nand_1 g02184(new_n2558_1, new_n2467, new_n2561);
and_1  g02185(new_n2561, new_n2560, new_n2562);
not_1  g02186(new_n2562, new_n2563);
nor_1  g02187(new_n511, new_n2476, new_n2564_1);
nand_1 g02188(n12705, n11917, new_n2565);
nand_1 g02189(n11257, n9956, new_n2566);
xnor_1 g02190(new_n2566, new_n2565, new_n2567);
and_1  g02191(new_n2567, new_n2564_1, new_n2568);
nor_1  g02192(new_n2567, new_n2564_1, new_n2569);
nor_1  g02193(new_n2569, new_n2568, new_n2570);
xnor_1 g02194(new_n2570, new_n2563, new_n2571);
xor_1  g02195(new_n2571, new_n2557, new_n2572);
not_1  g02196(new_n2572, new_n2573);
nor_1  g02197(new_n2490, new_n2480, new_n2574);
not_1  g02198(new_n2514, new_n2575);
nand_1 g02199(new_n2575, new_n2491, new_n2576);
xnor_1 g02200(new_n2576, new_n2487, new_n2577_1);
nor_1  g02201(new_n2577_1, new_n2574, new_n2578);
xnor_1 g02202(new_n2578, new_n2573, new_n2579);
xnor_1 g02203(new_n2579, new_n2545, new_n2580);
nor_1  g02204(new_n2551_1, new_n456, new_n2581_1);
not_1  g02205(new_n2545, new_n2582);
nor_1  g02206(new_n2544, new_n2515_1, new_n2583);
nor_1  g02207(new_n2583, new_n2582, new_n2584);
nand_1 g02208(new_n2584, new_n2581_1, new_n2585_1);
xnor_1 g02209(new_n2539, new_n2537, new_n2586);
not_1  g02210(new_n2586, new_n2587);
nor_1  g02211(new_n2531, new_n2529, new_n2588);
nor_1  g02212(new_n2493, new_n424, new_n2589);
nor_1  g02213(new_n456, new_n2476, new_n2590);
nand_1 g02214(new_n2590, new_n2589, new_n2591);
nor_1  g02215(new_n2591, new_n2588, new_n2592);
nand_1 g02216(new_n2592, new_n2587, new_n2593);
not_1  g02217(new_n2522_1, new_n2594);
xnor_1 g02218(new_n2541, new_n2594, new_n2595);
nor_1  g02219(new_n2595, new_n2593, new_n2596);
not_1  g02220(new_n2581_1, new_n2597);
xnor_1 g02221(new_n2584, new_n2597, new_n2598);
nand_1 g02222(new_n2598, new_n2596, new_n2599);
nand_1 g02223(new_n2599, new_n2585_1, new_n2600);
xnor_1 g02224(new_n2600, new_n2580, new_n2601);
not_1  g02225(new_n2601, new_n2602);
not_1  g02226(n8065, new_n2603);
nor_1  g02227(new_n552, new_n2603, new_n2604);
nand_1 g02228(n7436, n6126, new_n2605);
nand_1 g02229(n9241, n3719, new_n2606);
nand_1 g02230(n8276, n3602, new_n2607);
xnor_1 g02231(new_n2607, new_n2606, new_n2608);
nor_1  g02232(new_n2608, new_n2605, new_n2609);
not_1  g02233(new_n2609, new_n2610);
nand_1 g02234(new_n2608, new_n2605, new_n2611);
nand_1 g02235(new_n2611, new_n2610, new_n2612);
nand_1 g02236(n8276, n3719, new_n2613);
nand_1 g02237(n12299, n6126, new_n2614);
nand_1 g02238(new_n2614, new_n2613, new_n2615);
not_1  g02239(new_n2615, new_n2616);
nor_1  g02240(new_n2614, new_n2613, new_n2617);
not_1  g02241(n3602, new_n2618);
nor_1  g02242(new_n599, new_n2618, new_n2619);
nor_1  g02243(new_n2619, new_n2617, new_n2620);
nor_1  g02244(new_n2620, new_n2616, new_n2621);
xnor_1 g02245(new_n2621, new_n2612, new_n2622);
not_1  g02246(n10439, new_n2623);
nor_1  g02247(new_n2623, new_n563, new_n2624_1);
not_1  g02248(new_n2624_1, new_n2625);
not_1  g02249(n8595, new_n2626);
nor_1  g02250(new_n554, new_n2626, new_n2627);
not_1  g02251(new_n2627, new_n2628);
nand_1 g02252(new_n2628, new_n2625, new_n2629);
nor_1  g02253(new_n2628, new_n2625, new_n2630);
not_1  g02254(new_n2630, new_n2631);
nand_1 g02255(new_n2631, new_n2629, new_n2632);
xnor_1 g02256(new_n2632, new_n2622, new_n2633);
nand_1 g02257(n8595, n6776, new_n2634);
not_1  g02258(new_n2634, new_n2635);
nand_1 g02259(n7436, n3719, new_n2636);
nand_1 g02260(n6776, n6126, new_n2637);
nand_1 g02261(new_n2637, new_n2636, new_n2638);
not_1  g02262(new_n2638, new_n2639);
nor_1  g02263(new_n2637, new_n2636, new_n2640);
nor_1  g02264(new_n554, new_n2618, new_n2641);
nor_1  g02265(new_n2641, new_n2640, new_n2642);
nor_1  g02266(new_n2642, new_n2639, new_n2643);
nand_1 g02267(new_n2643, new_n2635, new_n2644);
not_1  g02268(new_n2644, new_n2645);
xnor_1 g02269(new_n2643, new_n2635, new_n2646);
not_1  g02270(new_n2619, new_n2647);
xnor_1 g02271(new_n2614, new_n2613, new_n2648);
xnor_1 g02272(new_n2648, new_n2647, new_n2649);
nor_1  g02273(new_n2649, new_n2646, new_n2650);
nor_1  g02274(new_n2650, new_n2645, new_n2651);
not_1  g02275(new_n2651, new_n2652);
nand_1 g02276(new_n2652, new_n2633, new_n2653);
not_1  g02277(new_n2653, new_n2654);
nor_1  g02278(new_n2652, new_n2633, new_n2655);
nor_1  g02279(new_n2655, new_n2654, new_n2656);
nor_1  g02280(new_n2623, new_n552, new_n2657);
not_1  g02281(new_n2657, new_n2658);
xnor_1 g02282(new_n2649, new_n2646, new_n2659);
nand_1 g02283(new_n2659, new_n2658, new_n2660);
xnor_1 g02284(new_n2659, new_n2657, new_n2661);
nor_1  g02285(new_n552, new_n2626, new_n2662);
nand_1 g02286(n12299, n3719, new_n2663);
not_1  g02287(new_n2663, new_n2664);
nand_1 g02288(n8759, n6126, new_n2665);
not_1  g02289(new_n2665, new_n2666);
nand_1 g02290(new_n2666, new_n2664, new_n2667);
nand_1 g02291(new_n2665, new_n2663, new_n2668);
nor_1  g02292(new_n563, new_n2618, new_n2669);
nand_1 g02293(new_n2669, new_n2668, new_n2670);
nand_1 g02294(new_n2670, new_n2667, new_n2671);
nand_1 g02295(new_n2671, new_n2662, new_n2672);
not_1  g02296(new_n2672, new_n2673);
xnor_1 g02297(new_n2671, new_n2662, new_n2674);
xnor_1 g02298(new_n2637, new_n2636, new_n2675);
xnor_1 g02299(new_n2675, new_n2641, new_n2676);
not_1  g02300(new_n2676, new_n2677);
nor_1  g02301(new_n2677, new_n2674, new_n2678);
nor_1  g02302(new_n2678, new_n2673, new_n2679_1);
nand_1 g02303(new_n2679_1, new_n2661, new_n2680);
nand_1 g02304(new_n2680, new_n2660, new_n2681);
not_1  g02305(new_n2681, new_n2682);
nand_1 g02306(new_n2682, new_n2656, new_n2683);
not_1  g02307(new_n2683, new_n2684);
nor_1  g02308(new_n2682, new_n2656, new_n2685);
nor_1  g02309(new_n2685, new_n2684, new_n2686);
nand_1 g02310(new_n2686, new_n2604, new_n2687);
xnor_1 g02311(new_n2676, new_n2674, new_n2688);
nand_1 g02312(new_n2668, new_n2667, new_n2689);
not_1  g02313(new_n2689, new_n2690);
not_1  g02314(n3719, new_n2691);
nor_1  g02315(new_n563, new_n2691, new_n2692);
nor_1  g02316(new_n552, new_n2618, new_n2693);
nand_1 g02317(new_n2693, new_n2692, new_n2694);
nor_1  g02318(new_n2694, new_n2690, new_n2695);
nand_1 g02319(new_n2695, new_n2688, new_n2696);
not_1  g02320(new_n2680, new_n2697);
nor_1  g02321(new_n2679_1, new_n2661, new_n2698);
nor_1  g02322(new_n2698, new_n2697, new_n2699);
nor_1  g02323(new_n2699, new_n2696, new_n2700);
not_1  g02324(new_n2604, new_n2701);
xnor_1 g02325(new_n2686, new_n2701, new_n2702);
nand_1 g02326(new_n2702, new_n2700, new_n2703);
nand_1 g02327(new_n2703, new_n2687, new_n2704);
not_1  g02328(new_n2612, new_n2705);
nand_1 g02329(new_n2621, new_n2705, new_n2706);
nand_1 g02330(new_n2706, new_n2610, new_n2707);
not_1  g02331(new_n2707, new_n2708_1);
nor_1  g02332(new_n2603, new_n563, new_n2709);
nand_1 g02333(n12299, n10439, new_n2710);
nand_1 g02334(n10391, n8759, new_n2711);
xnor_1 g02335(new_n2711, new_n2710, new_n2712);
xnor_1 g02336(new_n2712, new_n2709, new_n2713);
not_1  g02337(new_n2713, new_n2714);
nand_1 g02338(new_n2714, new_n2708_1, new_n2715);
nand_1 g02339(new_n2713, new_n2707, new_n2716);
nand_1 g02340(new_n2716, new_n2715, new_n2717);
not_1  g02341(new_n2717, new_n2718);
nor_1  g02342(new_n2607, new_n2606, new_n2719);
nor_1  g02343(new_n2626, new_n599, new_n2720);
xnor_1 g02344(new_n2720, new_n2719, new_n2721);
not_1  g02345(new_n2721, new_n2722);
not_1  g02346(n9241, new_n2723);
nor_1  g02347(new_n2723, new_n2618, new_n2724);
not_1  g02348(n6126, new_n2725);
not_1  g02349(n8276, new_n2726);
nor_1  g02350(new_n2726, new_n2725, new_n2727);
not_1  g02351(new_n2727, new_n2728);
not_1  g02352(n10510, new_n2729);
nor_1  g02353(new_n2729, new_n2691, new_n2730);
not_1  g02354(new_n2730, new_n2731);
nand_1 g02355(new_n2731, new_n2728, new_n2732);
nand_1 g02356(new_n2730, new_n2727, new_n2733);
nand_1 g02357(new_n2733, new_n2732, new_n2734);
xor_1  g02358(new_n2734, new_n2724, new_n2735);
xnor_1 g02359(new_n2735, new_n2722, new_n2736);
xnor_1 g02360(new_n2736, new_n2718, new_n2737);
not_1  g02361(new_n2632, new_n2738);
nand_1 g02362(new_n2738, new_n2622, new_n2739);
nand_1 g02363(new_n2654, new_n2630, new_n2740);
nand_1 g02364(new_n2653, new_n2631, new_n2741);
nand_1 g02365(new_n2741, new_n2740, new_n2742);
nand_1 g02366(new_n2742, new_n2739, new_n2743);
xnor_1 g02367(new_n2743, new_n2737, new_n2744);
xnor_1 g02368(new_n2744, new_n2683, new_n2745);
xnor_1 g02369(new_n2745, new_n2704, new_n2746);
not_1  g02370(new_n2746, new_n2747);
not_1  g02371(n4826, new_n2748);
nor_1  g02372(new_n829, new_n2748, new_n2749_1);
nand_1 g02373(n10545, n7733, new_n2750);
nand_1 g02374(n12925, n7690, new_n2751);
nor_1  g02375(new_n2751, new_n2750, new_n2752);
not_1  g02376(new_n2752, new_n2753);
nand_1 g02377(new_n2751, new_n2750, new_n2754);
nand_1 g02378(new_n2754, new_n2753, new_n2755);
xnor_1 g02379(new_n2755, new_n2749_1, new_n2756);
nand_1 g02380(n12925, n10545, new_n2757);
nand_1 g02381(n4826, n2530, new_n2758);
nand_1 g02382(new_n2758, new_n2757, new_n2759);
not_1  g02383(new_n2759, new_n2760);
not_1  g02384(n7733, new_n2761);
nor_1  g02385(new_n829, new_n2761, new_n2762);
xnor_1 g02386(new_n2758, new_n2757, new_n2763);
nor_1  g02387(new_n2763, new_n2762, new_n2764);
nor_1  g02388(new_n2764, new_n2760, new_n2765);
xnor_1 g02389(new_n2765, new_n2756, new_n2766);
not_1  g02390(n4970, new_n2767);
nor_1  g02391(new_n712, new_n2767, new_n2768);
not_1  g02392(new_n2768, new_n2769);
not_1  g02393(n7610, new_n2770);
nor_1  g02394(new_n2770, new_n740, new_n2771);
not_1  g02395(new_n2771, new_n2772);
nand_1 g02396(new_n2772, new_n2769, new_n2773);
nor_1  g02397(new_n2772, new_n2769, new_n2774);
not_1  g02398(new_n2774, new_n2775);
nand_1 g02399(new_n2775, new_n2773, new_n2776);
not_1  g02400(new_n2776, new_n2777);
xnor_1 g02401(new_n2777, new_n2766, new_n2778);
nor_1  g02402(new_n712, new_n2770, new_n2779);
nand_1 g02403(n12925, n12648, new_n2780);
nand_1 g02404(n8476, n4826, new_n2781);
nand_1 g02405(new_n2781, new_n2780, new_n2782);
not_1  g02406(new_n2782, new_n2783);
nor_1  g02407(new_n2761, new_n740, new_n2784);
xnor_1 g02408(new_n2781, new_n2780, new_n2785);
nor_1  g02409(new_n2785, new_n2784, new_n2786);
nor_1  g02410(new_n2786, new_n2783, new_n2787);
nand_1 g02411(new_n2787, new_n2779, new_n2788);
not_1  g02412(new_n2788, new_n2789);
xnor_1 g02413(new_n2787, new_n2779, new_n2790);
not_1  g02414(new_n2762, new_n2791);
xnor_1 g02415(new_n2763, new_n2791, new_n2792);
nor_1  g02416(new_n2792, new_n2790, new_n2793);
nor_1  g02417(new_n2793, new_n2789, new_n2794);
not_1  g02418(new_n2794, new_n2795);
nand_1 g02419(new_n2795, new_n2778, new_n2796);
not_1  g02420(new_n2796, new_n2797);
nor_1  g02421(new_n2795, new_n2778, new_n2798);
nor_1  g02422(new_n2798, new_n2797, new_n2799);
not_1  g02423(new_n2799, new_n2800);
nor_1  g02424(new_n668, new_n2767, new_n2801);
nand_1 g02425(n7610, n5331, new_n2802_1);
not_1  g02426(new_n2802_1, new_n2803);
nand_1 g02427(n12925, n2530, new_n2804);
nand_1 g02428(n5331, n4826, new_n2805);
nand_1 g02429(new_n2805, new_n2804, new_n2806);
not_1  g02430(new_n2806, new_n2807);
nor_1  g02431(new_n2805, new_n2804, new_n2808);
nor_1  g02432(new_n712, new_n2761, new_n2809);
nor_1  g02433(new_n2809, new_n2808, new_n2810);
nor_1  g02434(new_n2810, new_n2807, new_n2811);
nand_1 g02435(new_n2811, new_n2803, new_n2812);
xnor_1 g02436(new_n2811, new_n2802_1, new_n2813);
xnor_1 g02437(new_n2785, new_n2784, new_n2814);
nand_1 g02438(new_n2814, new_n2813, new_n2815);
nand_1 g02439(new_n2815, new_n2812, new_n2816);
nor_1  g02440(new_n2816, new_n2801, new_n2817);
not_1  g02441(new_n2817, new_n2818_1);
not_1  g02442(new_n2792, new_n2819);
xnor_1 g02443(new_n2819, new_n2790, new_n2820);
not_1  g02444(new_n2820, new_n2821);
not_1  g02445(new_n2801, new_n2822);
xnor_1 g02446(new_n2816, new_n2822, new_n2823);
nand_1 g02447(new_n2823, new_n2821, new_n2824);
nand_1 g02448(new_n2824, new_n2818_1, new_n2825);
nor_1  g02449(new_n2825, new_n2800, new_n2826);
not_1  g02450(new_n2826, new_n2827);
not_1  g02451(new_n2766, new_n2828);
nand_1 g02452(new_n2777, new_n2828, new_n2829);
nand_1 g02453(new_n2797, new_n2774, new_n2830);
nand_1 g02454(new_n2796, new_n2775, new_n2831);
nand_1 g02455(new_n2831, new_n2830, new_n2832);
nand_1 g02456(new_n2832, new_n2829, new_n2833);
nand_1 g02457(n12648, n7610, new_n2834);
xnor_1 g02458(new_n2834, new_n2752, new_n2835);
nor_1  g02459(new_n2761, new_n1048, new_n2836);
nand_1 g02460(n10545, n4826, new_n2837);
nand_1 g02461(n12925, n3616, new_n2838);
xnor_1 g02462(new_n2838, new_n2837, new_n2839);
xor_1  g02463(new_n2839, new_n2836, new_n2840);
xnor_1 g02464(new_n2840, new_n2835, new_n2841);
not_1  g02465(new_n2755, new_n2842);
nand_1 g02466(new_n2842, new_n2749_1, new_n2843);
nand_1 g02467(new_n2765, new_n2756, new_n2844);
nand_1 g02468(new_n2844, new_n2843, new_n2845);
not_1  g02469(n503, new_n2846);
nor_1  g02470(new_n712, new_n2846, new_n2847);
nand_1 g02471(n4970, n2530, new_n2848);
nand_1 g02472(n10965, n5331, new_n2849);
xnor_1 g02473(new_n2849, new_n2848, new_n2850);
xor_1  g02474(new_n2850, new_n2847, new_n2851);
xnor_1 g02475(new_n2851, new_n2845, new_n2852);
xnor_1 g02476(new_n2852, new_n2841, new_n2853);
xnor_1 g02477(new_n2853, new_n2833, new_n2854);
xnor_1 g02478(new_n2854, new_n2827, new_n2855);
nor_1  g02479(new_n668, new_n2846, new_n2856);
xnor_1 g02480(new_n2825, new_n2799, new_n2857);
nand_1 g02481(new_n2857, new_n2856, new_n2858);
not_1  g02482(new_n2815, new_n2859);
nor_1  g02483(new_n2814, new_n2813, new_n2860);
nor_1  g02484(new_n2860, new_n2859, new_n2861);
not_1  g02485(new_n2808, new_n2862);
nand_1 g02486(n12925, n5331, new_n2863);
nand_1 g02487(new_n2863, new_n2809, new_n2864);
nand_1 g02488(new_n2864, new_n2807, new_n2865);
nand_1 g02489(new_n2865, new_n2862, new_n2866);
nand_1 g02490(new_n2866, new_n2809, new_n2867);
not_1  g02491(new_n2867, new_n2868);
nand_1 g02492(new_n2868, new_n2861, new_n2869);
xnor_1 g02493(new_n2823, new_n2820, new_n2870);
nor_1  g02494(new_n2870, new_n2869, new_n2871);
not_1  g02495(new_n2856, new_n2872);
xnor_1 g02496(new_n2857, new_n2872, new_n2873);
nand_1 g02497(new_n2873, new_n2871, new_n2874);
nand_1 g02498(new_n2874, new_n2858, new_n2875);
xnor_1 g02499(new_n2875, new_n2855, new_n2876);
nand_1 g02500(n4086, n2393, new_n2877);
nand_1 g02501(n5860, n405, new_n2878);
nand_1 g02502(n8433, n3986, new_n2879_1);
xnor_1 g02503(new_n2879_1, new_n2878, new_n2880);
nor_1  g02504(new_n2880, new_n2877, new_n2881);
not_1  g02505(new_n2881, new_n2882);
nand_1 g02506(new_n2880, new_n2877, new_n2883);
nand_1 g02507(new_n2883, new_n2882, new_n2884);
nand_1 g02508(n8433, n5860, new_n2885);
nand_1 g02509(n11892, n4086, new_n2886);
nand_1 g02510(new_n2886, new_n2885, new_n2887);
not_1  g02511(new_n2887, new_n2888);
not_1  g02512(n405, new_n2889);
nor_1  g02513(new_n767, new_n2889, new_n2890);
xnor_1 g02514(new_n2886, new_n2885, new_n2891);
nor_1  g02515(new_n2891, new_n2890, new_n2892);
nor_1  g02516(new_n2892, new_n2888, new_n2893);
xnor_1 g02517(new_n2893, new_n2884, new_n2894);
not_1  g02518(n6611, new_n2895);
nor_1  g02519(new_n696, new_n2895, new_n2896);
not_1  g02520(new_n2896, new_n2897);
not_1  g02521(n217, new_n2898);
nor_1  g02522(new_n762, new_n2898, new_n2899);
not_1  g02523(new_n2899, new_n2900);
nor_1  g02524(new_n2900, new_n2897, new_n2901);
not_1  g02525(new_n2901, new_n2902_1);
nand_1 g02526(new_n2900, new_n2897, new_n2903);
nand_1 g02527(new_n2903, new_n2902_1, new_n2904);
xnor_1 g02528(new_n2904, new_n2894, new_n2905);
nor_1  g02529(new_n696, new_n2898, new_n2906);
nand_1 g02530(n8433, n2393, new_n2907);
nand_1 g02531(n7388, n4086, new_n2908);
nand_1 g02532(new_n2908, new_n2907, new_n2909);
not_1  g02533(new_n2909, new_n2910);
nor_1  g02534(new_n762, new_n2889, new_n2911);
xnor_1 g02535(new_n2908, new_n2907, new_n2912);
nor_1  g02536(new_n2912, new_n2911, new_n2913);
nor_1  g02537(new_n2913, new_n2910, new_n2914);
nand_1 g02538(new_n2914, new_n2906, new_n2915);
not_1  g02539(new_n2906, new_n2916);
xnor_1 g02540(new_n2914, new_n2916, new_n2917);
xnor_1 g02541(new_n2891, new_n2890, new_n2918);
nand_1 g02542(new_n2918, new_n2917, new_n2919);
nand_1 g02543(new_n2919, new_n2915, new_n2920);
xnor_1 g02544(new_n2920, new_n2905, new_n2921);
not_1  g02545(new_n2921, new_n2922);
nor_1  g02546(new_n754, new_n2895, new_n2923);
not_1  g02547(new_n2919, new_n2924);
nor_1  g02548(new_n2918, new_n2917, new_n2925);
nor_1  g02549(new_n2925, new_n2924, new_n2926);
nand_1 g02550(new_n2926, new_n2923, new_n2927);
not_1  g02551(new_n2927, new_n2928);
nor_1  g02552(new_n2926, new_n2923, new_n2929);
nor_1  g02553(new_n2929, new_n2928, new_n2930);
nor_1  g02554(new_n754, new_n2898, new_n2931);
not_1  g02555(new_n2931, new_n2932);
nand_1 g02556(n11892, n8433, new_n2933);
nand_1 g02557(n7965, n4086, new_n2934);
nor_1  g02558(new_n2934, new_n2933, new_n2935);
nand_1 g02559(new_n2934, new_n2933, new_n2936);
not_1  g02560(new_n2936, new_n2937);
nor_1  g02561(new_n696, new_n2889, new_n2938);
not_1  g02562(new_n2938, new_n2939);
nor_1  g02563(new_n2939, new_n2937, new_n2940);
nor_1  g02564(new_n2940, new_n2935, new_n2941);
nor_1  g02565(new_n2941, new_n2932, new_n2942);
xnor_1 g02566(new_n2941, new_n2932, new_n2943);
xnor_1 g02567(new_n2912, new_n2911, new_n2944);
not_1  g02568(new_n2944, new_n2945);
nor_1  g02569(new_n2945, new_n2943, new_n2946);
nor_1  g02570(new_n2946, new_n2942, new_n2947);
not_1  g02571(new_n2947, new_n2948);
nand_1 g02572(new_n2948, new_n2930, new_n2949);
nand_1 g02573(new_n2949, new_n2927, new_n2950);
nand_1 g02574(new_n2950, new_n2922, new_n2951);
not_1  g02575(new_n2904, new_n2952);
nand_1 g02576(new_n2952, new_n2894, new_n2953);
nand_1 g02577(new_n2920, new_n2905, new_n2954);
xnor_1 g02578(new_n2954, new_n2902_1, new_n2955);
nand_1 g02579(new_n2955, new_n2953, new_n2956);
nor_1  g02580(new_n2879_1, new_n2878, new_n2957);
nor_1  g02581(new_n767, new_n2898, new_n2958);
xor_1  g02582(new_n2958, new_n2957, new_n2959);
nor_1  g02583(new_n1084, new_n2889, new_n2960);
nand_1 g02584(n5860, n4086, new_n2961);
nand_1 g02585(n8433, n5857, new_n2962);
xnor_1 g02586(new_n2962, new_n2961, new_n2963);
xor_1  g02587(new_n2963, new_n2960, new_n2964);
xnor_1 g02588(new_n2964, new_n2959, new_n2965);
not_1  g02589(new_n2884, new_n2966);
nand_1 g02590(new_n2893, new_n2966, new_n2967);
nand_1 g02591(new_n2967, new_n2882, new_n2968);
not_1  g02592(n11296, new_n2969);
nor_1  g02593(new_n2969, new_n754, new_n2970);
nand_1 g02594(n11892, n6611, new_n2971);
nand_1 g02595(n7388, n6359, new_n2972);
xnor_1 g02596(new_n2972, new_n2971, new_n2973);
xor_1  g02597(new_n2973, new_n2970, new_n2974);
xnor_1 g02598(new_n2974, new_n2968, new_n2975);
xnor_1 g02599(new_n2975, new_n2965, new_n2976);
xnor_1 g02600(new_n2976, new_n2956, new_n2977);
xnor_1 g02601(new_n2977, new_n2951, new_n2978);
not_1  g02602(new_n2978, new_n2979);
not_1  g02603(n6359, new_n2980);
nor_1  g02604(new_n754, new_n2980, new_n2981);
xnor_1 g02605(new_n2950, new_n2921, new_n2982);
nand_1 g02606(new_n2982, new_n2981, new_n2983);
xnor_1 g02607(new_n2944, new_n2943, new_n2984);
nor_1  g02608(new_n2937, new_n2935, new_n2985);
not_1  g02609(new_n2985, new_n2986);
nand_1 g02610(n8433, n7388, new_n2987);
nand_1 g02611(n7965, n405, new_n2988);
nor_1  g02612(new_n2988, new_n2987, new_n2989);
and_1  g02613(new_n2989, new_n2986, new_n2990);
nand_1 g02614(new_n2990, new_n2984, new_n2991);
xnor_1 g02615(new_n2948, new_n2930, new_n2992);
nor_1  g02616(new_n2992, new_n2991, new_n2993);
not_1  g02617(new_n2981, new_n2994);
xnor_1 g02618(new_n2982, new_n2994, new_n2995);
nand_1 g02619(new_n2995, new_n2993, new_n2996);
nand_1 g02620(new_n2996, new_n2983, new_n2997);
xnor_1 g02621(new_n2997, new_n2979, new_n2998);
xnor_1 g02622(new_n2998, new_n2876, new_n2999);
not_1  g02623(new_n2871, new_n3000);
xnor_1 g02624(new_n2873, new_n3000, new_n3001);
not_1  g02625(new_n3001, new_n3002);
xnor_1 g02626(new_n2995, new_n2993, new_n3003);
nand_1 g02627(new_n3003, new_n3002, new_n3004);
xnor_1 g02628(new_n2992, new_n2991, new_n3005);
xnor_1 g02629(new_n2868, new_n2861, new_n3006);
not_1  g02630(new_n2984, new_n3007);
xnor_1 g02631(new_n2990, new_n3007, new_n3008);
not_1  g02632(new_n3008, new_n3009);
nand_1 g02633(new_n3009, new_n3006, new_n3010);
nand_1 g02634(n8433, n7965, new_n3011);
nor_1  g02635(new_n3011, new_n2863, new_n3012);
not_1  g02636(new_n3012, new_n3013);
xnor_1 g02637(new_n2988, new_n2987, new_n3014);
nand_1 g02638(new_n3014, new_n3013, new_n3015);
xnor_1 g02639(new_n3014, new_n3012, new_n3016);
nand_1 g02640(n12925, n8476, new_n3017);
nand_1 g02641(n7733, n5331, new_n3018);
xnor_1 g02642(new_n3018, new_n3017, new_n3019);
nand_1 g02643(new_n3019, new_n3016, new_n3020);
nand_1 g02644(new_n3020, new_n3015, new_n3021);
nor_1  g02645(new_n2864, new_n2807, new_n3022_1);
nor_1  g02646(new_n3022_1, new_n2866, new_n3023);
not_1  g02647(new_n3023, new_n3024);
nand_1 g02648(new_n3024, new_n3021, new_n3025);
xnor_1 g02649(new_n3023, new_n3021, new_n3026);
nand_1 g02650(new_n3011, new_n2938, new_n3027);
not_1  g02651(new_n3027, new_n3028);
nor_1  g02652(new_n3028, new_n2985, new_n3029);
nor_1  g02653(new_n3027, new_n2937, new_n3030);
nor_1  g02654(new_n3030, new_n3029, new_n3031);
not_1  g02655(new_n3031, new_n3032);
nand_1 g02656(new_n3032, new_n3026, new_n3033);
nand_1 g02657(new_n3033, new_n3025, new_n3034);
xnor_1 g02658(new_n3008, new_n3006, new_n3035);
nand_1 g02659(new_n3035, new_n3034, new_n3036);
nand_1 g02660(new_n3036, new_n3010, new_n3037);
nand_1 g02661(new_n3037, new_n3005, new_n3038);
nand_1 g02662(new_n2870, new_n2869, new_n3039);
nand_1 g02663(new_n3039, new_n3000, new_n3040);
not_1  g02664(new_n3005, new_n3041);
xnor_1 g02665(new_n3037, new_n3041, new_n3042);
nand_1 g02666(new_n3042, new_n3040, new_n3043);
nand_1 g02667(new_n3043, new_n3038, new_n3044);
xnor_1 g02668(new_n3003, new_n3001, new_n3045);
nand_1 g02669(new_n3045, new_n3044, new_n3046);
nand_1 g02670(new_n3046, new_n3004, new_n3047);
xnor_1 g02671(new_n3047, new_n2999, new_n3048);
xnor_1 g02672(new_n3048, new_n2747, new_n3049);
xnor_1 g02673(new_n2702, new_n2700, new_n3050);
xnor_1 g02674(new_n3003, new_n3002, new_n3051);
xnor_1 g02675(new_n3051, new_n3044, new_n3052);
nand_1 g02676(new_n3052, new_n3050, new_n3053);
not_1  g02677(new_n3053, new_n3054);
xnor_1 g02678(new_n3052, new_n3050, new_n3055);
xnor_1 g02679(new_n2699, new_n2696, new_n3056);
not_1  g02680(new_n3056, new_n3057);
xnor_1 g02681(new_n3042, new_n3040, new_n3058);
nand_1 g02682(new_n3058, new_n3057, new_n3059);
xnor_1 g02683(new_n3058, new_n3056, new_n3060);
xor_1  g02684(new_n2695, new_n2688, new_n3061);
not_1  g02685(new_n3061, new_n3062);
xnor_1 g02686(new_n3035, new_n3034, new_n3063);
not_1  g02687(new_n3063, new_n3064);
nor_1  g02688(new_n3064, new_n3062, new_n3065);
not_1  g02689(new_n3065, new_n3066);
nor_1  g02690(new_n3063, new_n3061, new_n3067);
nor_1  g02691(new_n3067, new_n3065, new_n3068);
xnor_1 g02692(new_n3031, new_n3026, new_n3069);
not_1  g02693(new_n3069, new_n3070);
nor_1  g02694(new_n552, new_n2691, new_n3071_1);
not_1  g02695(new_n3071_1, new_n3072);
nand_1 g02696(new_n3072, new_n2669, new_n3073);
not_1  g02697(new_n3073, new_n3074);
nor_1  g02698(new_n3074, new_n2690, new_n3075);
nand_1 g02699(new_n3074, new_n2668, new_n3076);
not_1  g02700(new_n3076, new_n3077);
nor_1  g02701(new_n3077, new_n3075, new_n3078);
and_1  g02702(new_n3078, new_n3070, new_n3079);
not_1  g02703(new_n3079, new_n3080);
nor_1  g02704(new_n3078, new_n3070, new_n3081);
nor_1  g02705(new_n3081, new_n3079, new_n3082);
xnor_1 g02706(new_n3019, new_n3016, new_n3083);
not_1  g02707(new_n3083, new_n3084);
xnor_1 g02708(new_n2693, new_n2692, new_n3085);
nor_1  g02709(new_n3085, new_n3084, new_n3086);
not_1  g02710(new_n3086, new_n3087);
nand_1 g02711(new_n3011, new_n2863, new_n3088);
and_1  g02712(new_n3088, new_n3013, new_n3089);
not_1  g02713(new_n3089, new_n3090);
nor_1  g02714(new_n3090, new_n3072, new_n3091);
xnor_1 g02715(new_n3085, new_n3083, new_n3092);
nand_1 g02716(new_n3092, new_n3091, new_n3093);
and_1  g02717(new_n3093, new_n3087, new_n3094);
not_1  g02718(new_n3094, new_n3095);
nand_1 g02719(new_n3095, new_n3082, new_n3096);
nand_1 g02720(new_n3096, new_n3080, new_n3097);
nand_1 g02721(new_n3097, new_n3068, new_n3098);
nand_1 g02722(new_n3098, new_n3066, new_n3099);
nand_1 g02723(new_n3099, new_n3060, new_n3100);
nand_1 g02724(new_n3100, new_n3059, new_n3101);
nor_1  g02725(new_n3101, new_n3055, new_n3102);
nor_1  g02726(new_n3102, new_n3054, new_n3103);
xnor_1 g02727(new_n3103, new_n3049, new_n3104);
nand_1 g02728(new_n3104, new_n2602, new_n3105);
xnor_1 g02729(new_n3104, new_n2601, new_n3106);
xnor_1 g02730(new_n2598, new_n2596, new_n3107);
not_1  g02731(new_n3107, new_n3108);
xnor_1 g02732(new_n3101, new_n3055, new_n3109);
nand_1 g02733(new_n3109, new_n3108, new_n3110);
xor_1  g02734(new_n2595, new_n2593, new_n3111);
not_1  g02735(new_n3099, new_n3112);
xnor_1 g02736(new_n3112, new_n3060, new_n3113);
nor_1  g02737(new_n3113, new_n3111, new_n3114);
xnor_1 g02738(new_n3113, new_n3111, new_n3115);
xnor_1 g02739(new_n2592, new_n2586, new_n3116);
not_1  g02740(new_n3098, new_n3117);
nor_1  g02741(new_n3097, new_n3068, new_n3118);
nor_1  g02742(new_n3118, new_n3117, new_n3119);
nor_1  g02743(new_n3119, new_n3116, new_n3120);
xnor_1 g02744(new_n3094, new_n3082, new_n3121);
nor_1  g02745(new_n2493, new_n456, new_n3122);
nor_1  g02746(new_n3122, new_n2533, new_n3123);
nor_1  g02747(new_n3123, new_n2588, new_n3124_1);
and_1  g02748(new_n3123, new_n2530_1, new_n3125);
nor_1  g02749(new_n3125, new_n3124_1, new_n3126);
nor_1  g02750(new_n3126, new_n3121, new_n3127);
xnor_1 g02751(new_n3126, new_n3121, new_n3128);
nor_1  g02752(new_n3089, new_n3071_1, new_n3129);
nor_1  g02753(new_n3129, new_n3091, new_n3130);
nand_1 g02754(new_n3130, new_n3122, new_n3131);
not_1  g02755(new_n2589, new_n3132);
xnor_1 g02756(new_n2590, new_n3132, new_n3133);
not_1  g02757(new_n3133, new_n3134);
nand_1 g02758(new_n3134, new_n3131, new_n3135);
not_1  g02759(new_n3135, new_n3136);
xor_1  g02760(new_n3092, new_n3091, new_n3137);
nor_1  g02761(new_n3134, new_n3131, new_n3138);
nor_1  g02762(new_n3138, new_n3136, new_n3139);
not_1  g02763(new_n3139, new_n3140);
nor_1  g02764(new_n3140, new_n3137, new_n3141);
nor_1  g02765(new_n3141, new_n3136, new_n3142);
nor_1  g02766(new_n3142, new_n3128, new_n3143);
nor_1  g02767(new_n3143, new_n3127, new_n3144);
xnor_1 g02768(new_n3119, new_n3116, new_n3145);
nor_1  g02769(new_n3145, new_n3144, new_n3146_1);
nor_1  g02770(new_n3146_1, new_n3120, new_n3147);
nor_1  g02771(new_n3147, new_n3115, new_n3148);
nor_1  g02772(new_n3148, new_n3114, new_n3149);
xnor_1 g02773(new_n3109, new_n3107, new_n3150);
nand_1 g02774(new_n3150, new_n3149, new_n3151);
nand_1 g02775(new_n3151, new_n3110, new_n3152);
nand_1 g02776(new_n3152, new_n3106, new_n3153);
nand_1 g02777(new_n3153, new_n3105, new_n3154);
nand_1 g02778(new_n3048, new_n2747, new_n3155);
xnor_1 g02779(new_n3048, new_n2746, new_n3156);
nand_1 g02780(new_n3103, new_n3156, new_n3157);
nand_1 g02781(new_n3157, new_n3155, new_n3158);
nor_1  g02782(new_n2834, new_n2753, new_n3159);
not_1  g02783(new_n2835, new_n3160);
nor_1  g02784(new_n2840, new_n3160, new_n3161);
nor_1  g02785(new_n3161, new_n3159, new_n3162);
nand_1 g02786(new_n2838, new_n2837, new_n3163);
not_1  g02787(new_n3163, new_n3164);
nor_1  g02788(new_n2839, new_n2836, new_n3165);
nor_1  g02789(new_n3165, new_n3164, new_n3166);
nand_1 g02790(n12648, n4970, new_n3167);
nand_1 g02791(n11296, n7388, new_n3168);
nand_1 g02792(n9241, n6126, new_n3169);
xnor_1 g02793(new_n3169, new_n3168, new_n3170);
xnor_1 g02794(new_n3170, new_n3167, new_n3171);
xnor_1 g02795(new_n3171, new_n3166, new_n3172_1);
xnor_1 g02796(new_n3172_1, new_n3162, new_n3173);
nand_1 g02797(new_n2962, new_n2961, new_n3174);
not_1  g02798(new_n3174, new_n3175);
nor_1  g02799(new_n2963, new_n2960, new_n3176);
nor_1  g02800(new_n3176, new_n3175, new_n3177);
nand_1 g02801(new_n2972, new_n2971, new_n3178);
not_1  g02802(new_n3178, new_n3179);
nor_1  g02803(new_n2973, new_n2970, new_n3180);
nor_1  g02804(new_n3180, new_n3179, new_n3181);
xnor_1 g02805(new_n3181, new_n3177, new_n3182);
nor_1  g02806(new_n762, new_n2980, new_n3183);
nand_1 g02807(n7546, n5331, new_n3184);
xnor_1 g02808(new_n3184, new_n3183, new_n3185);
xnor_1 g02809(new_n3185, new_n3182, new_n3186);
nand_1 g02810(new_n2720, new_n2719, new_n3187);
not_1  g02811(new_n2735, new_n3188);
nand_1 g02812(new_n3188, new_n2722, new_n3189);
nand_1 g02813(new_n3189, new_n3187, new_n3190);
nand_1 g02814(n8595, n8276, new_n3191);
nand_1 g02815(n6611, n2393, new_n3192);
xnor_1 g02816(new_n3192, new_n3191, new_n3193);
nand_1 g02817(n12925, n4499, new_n3194);
nand_1 g02818(n11536, n5305, new_n3195);
xnor_1 g02819(new_n3195, new_n3194, new_n3196);
xnor_1 g02820(new_n3196, new_n3193, new_n3197);
xnor_1 g02821(new_n3197, new_n3190, new_n3198);
xnor_1 g02822(new_n3198, new_n3186, new_n3199);
nand_1 g02823(new_n2958, new_n2957, new_n3200);
not_1  g02824(new_n2964, new_n3201);
nand_1 g02825(new_n3201, new_n2959, new_n3202);
nand_1 g02826(new_n3202, new_n3200, new_n3203);
nand_1 g02827(new_n2849, new_n2848, new_n3204);
not_1  g02828(new_n3204, new_n3205);
nor_1  g02829(new_n2850, new_n2847, new_n3206);
nor_1  g02830(new_n3206, new_n3205, new_n3207);
nand_1 g02831(n4086, n3986, new_n3208);
nand_1 g02832(n7733, n3616, new_n3209);
xnor_1 g02833(new_n3209, new_n3208, new_n3210);
xnor_1 g02834(new_n3210, new_n3207, new_n3211);
xnor_1 g02835(new_n3211, new_n3203, new_n3212);
xnor_1 g02836(new_n3212, new_n3199, new_n3213);
xnor_1 g02837(new_n3213, new_n3173, new_n3214_1);
not_1  g02838(new_n2951, new_n3215);
nand_1 g02839(new_n2977, new_n3215, new_n3216);
nand_1 g02840(new_n2997, new_n2978, new_n3217);
nand_1 g02841(new_n3217, new_n3216, new_n3218);
nor_1  g02842(new_n802, new_n2898, new_n3219);
xnor_1 g02843(new_n3219, new_n3218, new_n3220);
nand_1 g02844(new_n2744, new_n2684, new_n3221);
nand_1 g02845(new_n2745, new_n2704, new_n3222);
nand_1 g02846(new_n3222, new_n3221, new_n3223);
not_1  g02847(new_n2851, new_n3224);
nand_1 g02848(new_n3224, new_n2845, new_n3225);
nand_1 g02849(new_n2852, new_n2841, new_n3226);
nand_1 g02850(new_n3226, new_n3225, new_n3227);
nand_1 g02851(n12299, n8065, new_n3228);
nor_1  g02852(new_n2729, new_n2618, new_n3229);
xnor_1 g02853(new_n3229, new_n3228, new_n3230_1);
nand_1 g02854(n10644, n3719, new_n3231);
nand_1 g02855(n7965, n1357, new_n3232);
xnor_1 g02856(new_n3232, new_n3231, new_n3233);
nand_1 g02857(n10439, n7436, new_n3234);
nand_1 g02858(n8759, n4190, new_n3235);
xnor_1 g02859(new_n3235, new_n3234, new_n3236);
xnor_1 g02860(new_n3236, new_n3233, new_n3237);
xnor_1 g02861(new_n3237, new_n3230_1, new_n3238);
nand_1 g02862(new_n2554, new_n2553, new_n3239);
not_1  g02863(new_n3239, new_n3240);
nor_1  g02864(new_n2555, new_n2552, new_n3241);
nor_1  g02865(new_n3241, new_n3240, new_n3242);
nand_1 g02866(n9637, n1097, new_n3243);
xnor_1 g02867(new_n3243, new_n3242, new_n3244);
xnor_1 g02868(new_n3244, new_n3238, new_n3245);
xnor_1 g02869(new_n3245, new_n3227, new_n3246);
xnor_1 g02870(new_n2735, new_n2721, new_n3247);
nand_1 g02871(new_n3247, new_n2718, new_n3248);
nand_1 g02872(new_n3248, new_n2715, new_n3249);
not_1  g02873(new_n2556, new_n3250);
nand_1 g02874(new_n3250, new_n2550, new_n3251);
nand_1 g02875(new_n2571, new_n2557, new_n3252);
nand_1 g02876(new_n3252, new_n3251, new_n3253);
xnor_1 g02877(new_n3253, new_n3249, new_n3254);
xnor_1 g02878(new_n3254, new_n3246, new_n3255);
nand_1 g02879(new_n2736, new_n2717, new_n3256);
nand_1 g02880(new_n3256, new_n3248, new_n3257);
nand_1 g02881(new_n2743, new_n3257, new_n3258);
nand_1 g02882(new_n3258, new_n2740, new_n3259);
nand_1 g02883(new_n2711, new_n2710, new_n3260);
not_1  g02884(new_n3260, new_n3261);
nor_1  g02885(new_n2712, new_n2709, new_n3262);
nor_1  g02886(new_n3262, new_n3261, new_n3263);
nand_1 g02887(n4312, n2577, new_n3264);
xnor_1 g02888(new_n3264, new_n3263, new_n3265);
nand_1 g02889(new_n2732, new_n2724, new_n3266);
nand_1 g02890(new_n3266, new_n2733, new_n3267);
nand_1 g02891(n11257, n4921, new_n3268);
nand_1 g02892(n12705, n3842, new_n3269);
xnor_1 g02893(new_n3269, new_n3268, new_n3270);
xnor_1 g02894(new_n3270, new_n3267, new_n3271);
xnor_1 g02895(new_n3271, new_n3265, new_n3272_1);
nand_1 g02896(n8433, n45, new_n3273);
nor_1  g02897(new_n511, new_n2462, new_n3274);
xnor_1 g02898(new_n3274, new_n3273, new_n3275);
nand_1 g02899(new_n2566, new_n2565, new_n3276);
not_1  g02900(new_n3276, new_n3277);
nor_1  g02901(new_n2569, new_n3277, new_n3278);
nand_1 g02902(n5964, n1835, new_n3279);
not_1  g02903(n5857, new_n3280);
nor_1  g02904(new_n3280, new_n2889, new_n3281);
xnor_1 g02905(new_n3281, new_n3279, new_n3282);
xnor_1 g02906(new_n3282, new_n3278, new_n3283);
xnor_1 g02907(new_n3283, new_n3275, new_n3284);
nand_1 g02908(new_n2570, new_n2562, new_n3285);
nand_1 g02909(new_n3285, new_n2560, new_n3286);
not_1  g02910(n10391, new_n3287_1);
nor_1  g02911(new_n3287_1, new_n563, new_n3288);
xnor_1 g02912(new_n3288, new_n3286, new_n3289);
xnor_1 g02913(new_n3289, new_n3284, new_n3290);
xnor_1 g02914(new_n3290, new_n3272_1, new_n3291);
xnor_1 g02915(new_n3291, new_n3259, new_n3292);
xnor_1 g02916(new_n3292, new_n3255, new_n3293);
xnor_1 g02917(new_n3293, new_n3223, new_n3294);
xnor_1 g02918(new_n3294, new_n3220, new_n3295);
xnor_1 g02919(new_n3295, new_n3214_1, new_n3296);
not_1  g02920(new_n2998, new_n3297);
nand_1 g02921(new_n3297, new_n2876, new_n3298);
nand_1 g02922(new_n3047, new_n2999, new_n3299);
nand_1 g02923(new_n3299, new_n3298, new_n3300);
or_1   g02924(new_n2954, new_n2902_1, new_n3301);
not_1  g02925(new_n2976, new_n3302);
nand_1 g02926(new_n3302, new_n2956, new_n3303);
nand_1 g02927(new_n3303, new_n3301, new_n3304);
nor_1  g02928(new_n2576, new_n2488, new_n3305);
nor_1  g02929(new_n2578, new_n2572, new_n3306);
nor_1  g02930(new_n3306, new_n3305, new_n3307);
xnor_1 g02931(new_n3307, new_n3304, new_n3308);
xnor_1 g02932(new_n3308, new_n3300, new_n3309);
xnor_1 g02933(new_n3309, new_n3296, new_n3310);
xnor_1 g02934(new_n3310, new_n3158, new_n3311);
nand_1 g02935(new_n2854, new_n2826, new_n3312);
nand_1 g02936(new_n2875, new_n2855, new_n3313);
nand_1 g02937(new_n3313, new_n3312, new_n3314);
nand_1 g02938(new_n2579, new_n2582, new_n3315);
nand_1 g02939(new_n2600, new_n2580, new_n3316);
nand_1 g02940(new_n3316, new_n3315, new_n3317);
xnor_1 g02941(new_n3317, new_n3314, new_n3318);
not_1  g02942(new_n2853, new_n3319);
nand_1 g02943(new_n3319, new_n2833, new_n3320);
nand_1 g02944(new_n3320, new_n2830, new_n3321);
not_1  g02945(new_n2968, new_n3322);
nand_1 g02946(new_n2974, new_n3322, new_n3323);
not_1  g02947(new_n2965, new_n3324);
nand_1 g02948(new_n2975, new_n3324, new_n3325);
nand_1 g02949(new_n3325, new_n3323, new_n3326);
not_1  g02950(n10547, new_n3327);
nor_1  g02951(new_n3327, new_n2493, new_n3328);
nand_1 g02952(n10965, n8476, new_n3329);
nand_1 g02953(n7690, n4826, new_n3330);
xnor_1 g02954(new_n3330, new_n3329, new_n3331);
nand_1 g02955(n10545, n7610, new_n3332);
nand_1 g02956(n2530, n503, new_n3333);
xnor_1 g02957(new_n3333, new_n3332, new_n3334);
xnor_1 g02958(new_n3334, new_n3331, new_n3335);
xnor_1 g02959(new_n3335, new_n3328, new_n3336);
xnor_1 g02960(new_n3336, new_n3326, new_n3337);
xnor_1 g02961(new_n3337, new_n3321, new_n3338);
xnor_1 g02962(new_n3338, new_n3318, new_n3339_1);
xnor_1 g02963(new_n3339_1, new_n3311, new_n3340);
xnor_1 g02964(new_n3340, new_n3154, n837);
nor_1  g02965(new_n2462, new_n1592, new_n3342_1);
nand_1 g02966(n9956, n5240, new_n3343);
nor_1  g02967(new_n1592, new_n2476, new_n3344);
nand_1 g02968(n11917, n3172, new_n3345);
xnor_1 g02969(new_n3345, new_n3343, new_n3346);
nor_1  g02970(new_n3346, new_n3344, new_n3347);
nor_1  g02971(new_n3347, new_n3343, new_n3348);
nor_1  g02972(new_n3348, new_n3342_1, new_n3349);
not_1  g02973(new_n3342_1, new_n3350);
nor_1  g02974(new_n2476, new_n1600, new_n3351);
nor_1  g02975(new_n3351, new_n3348, new_n3352);
nor_1  g02976(new_n3352, new_n3350, new_n3353);
nor_1  g02977(new_n3353, new_n3349, new_n3354);
nand_1 g02978(n5240, n4921, new_n3355);
nand_1 g02979(n11821, n9956, new_n3356);
xnor_1 g02980(new_n3356, new_n3355, new_n3357);
not_1  g02981(new_n3357, new_n3358);
nor_1  g02982(new_n3358, new_n3354, new_n3359);
nand_1 g02983(new_n3358, new_n3354, new_n3360);
not_1  g02984(new_n3360, new_n3361);
nor_1  g02985(new_n3361, new_n3359, new_n3362);
nor_1  g02986(new_n2481, new_n1590, new_n3363);
not_1  g02987(new_n3363, new_n3364);
nor_1  g02988(new_n2484, new_n1600, new_n3365);
not_1  g02989(new_n3365, new_n3366);
nand_1 g02990(new_n3366, new_n3364, new_n3367);
nor_1  g02991(new_n3366, new_n3364, new_n3368);
not_1  g02992(new_n3368, new_n3369);
nand_1 g02993(new_n3369, new_n3367, new_n3370);
xnor_1 g02994(new_n3370, new_n3362, new_n3371);
nor_1  g02995(new_n2484, new_n1590, new_n3372);
nand_1 g02996(n11757, n9956, new_n3373);
nand_1 g02997(n11917, n1333, new_n3374);
nand_1 g02998(new_n3374, new_n3373, new_n3375);
not_1  g02999(new_n3375, new_n3376);
nor_1  g03000(new_n3374, new_n3373, new_n3377);
nor_1  g03001(new_n3377, new_n3351, new_n3378);
nor_1  g03002(new_n3378, new_n3376, new_n3379);
nand_1 g03003(new_n3379, new_n3372, new_n3380);
xnor_1 g03004(new_n3346, new_n3344, new_n3381);
not_1  g03005(new_n3380, new_n3382);
nor_1  g03006(new_n3379, new_n3372, new_n3383);
nor_1  g03007(new_n3383, new_n3382, new_n3384);
nand_1 g03008(new_n3384, new_n3381, new_n3385);
nand_1 g03009(new_n3385, new_n3380, new_n3386);
nand_1 g03010(new_n3386, new_n3371, new_n3387);
not_1  g03011(new_n3387, new_n3388);
nor_1  g03012(new_n3386, new_n3371, new_n3389);
nor_1  g03013(new_n3389, new_n3388, new_n3390);
nor_1  g03014(new_n1348, new_n2481, new_n3391);
not_1  g03015(new_n3391, new_n3392);
xnor_1 g03016(new_n3384, new_n3381, new_n3393);
nor_1  g03017(new_n3393, new_n3392, new_n3394);
nor_1  g03018(new_n1348, new_n2484, new_n3395);
nor_1  g03019(new_n2493, new_n1600, new_n3396);
not_1  g03020(new_n3396, new_n3397);
nor_1  g03021(new_n2462, new_n1348, new_n3398);
not_1  g03022(new_n3398, new_n3399);
nor_1  g03023(new_n3399, new_n3397, new_n3400);
not_1  g03024(new_n3400, new_n3401);
nand_1 g03025(new_n3399, new_n3397, new_n3402);
not_1  g03026(new_n3402, new_n3403);
nor_1  g03027(new_n2476, new_n1590, new_n3404);
not_1  g03028(new_n3404, new_n3405);
nor_1  g03029(new_n3405, new_n3403, new_n3406);
not_1  g03030(new_n3406, new_n3407);
nand_1 g03031(new_n3407, new_n3401, new_n3408);
nand_1 g03032(new_n3408, new_n3395, new_n3409);
not_1  g03033(new_n3409, new_n3410);
xnor_1 g03034(new_n3408, new_n3395, new_n3411);
not_1  g03035(new_n3377, new_n3412);
nand_1 g03036(new_n3412, new_n3375, new_n3413);
xnor_1 g03037(new_n3413, new_n3351, new_n3414);
not_1  g03038(new_n3414, new_n3415);
nor_1  g03039(new_n3415, new_n3411, new_n3416);
nor_1  g03040(new_n3416, new_n3410, new_n3417);
xnor_1 g03041(new_n3393, new_n3392, new_n3418);
nor_1  g03042(new_n3418, new_n3417, new_n3419);
nor_1  g03043(new_n3419, new_n3394, new_n3420);
not_1  g03044(new_n3420, new_n3421);
nand_1 g03045(new_n3421, new_n3390, new_n3422);
nor_1  g03046(new_n3361, new_n3353, new_n3423);
nand_1 g03047(n9637, n1333, new_n3424);
nand_1 g03048(n3172, n2577, new_n3425);
nand_1 g03049(n7862, n1835, new_n3426);
nand_1 g03050(new_n3426, new_n3425, new_n3427);
not_1  g03051(new_n3427, new_n3428);
nor_1  g03052(new_n3426, new_n3425, new_n3429);
nor_1  g03053(new_n3429, new_n3428, new_n3430);
xor_1  g03054(new_n3430, new_n3424, new_n3431);
xnor_1 g03055(new_n3431, new_n3423, new_n3432);
not_1  g03056(new_n3432, new_n3433);
nor_1  g03057(new_n3356, new_n3355, new_n3434);
nor_1  g03058(new_n1592, new_n2484, new_n3435);
xor_1  g03059(new_n3435, new_n3434, new_n3436);
nor_1  g03060(new_n1682, new_n2476, new_n3437);
nand_1 g03061(n9956, n9080, new_n3438);
nand_1 g03062(n11917, n5240, new_n3439);
xnor_1 g03063(new_n3439, new_n3438, new_n3440);
xnor_1 g03064(new_n3440, new_n3437, new_n3441);
xnor_1 g03065(new_n3441, new_n3436, new_n3442);
nand_1 g03066(new_n3442, new_n3433, new_n3443);
not_1  g03067(new_n3442, new_n3444);
nand_1 g03068(new_n3444, new_n3432, new_n3445);
nand_1 g03069(new_n3445, new_n3443, new_n3446);
not_1  g03070(new_n3446, new_n3447);
not_1  g03071(new_n3370, new_n3448);
nand_1 g03072(new_n3448, new_n3362, new_n3449);
nand_1 g03073(new_n3388, new_n3368, new_n3450);
nand_1 g03074(new_n3387, new_n3369, new_n3451);
nand_1 g03075(new_n3451, new_n3450, new_n3452);
nand_1 g03076(new_n3452, new_n3449, new_n3453);
xnor_1 g03077(new_n3453, new_n3447, new_n3454);
xnor_1 g03078(new_n3454, new_n3422, new_n3455);
nor_1  g03079(new_n2551_1, new_n1348, new_n3456_1);
not_1  g03080(new_n3422, new_n3457);
nor_1  g03081(new_n3421, new_n3390, new_n3458);
nor_1  g03082(new_n3458, new_n3457, new_n3459);
nand_1 g03083(new_n3459, new_n3456_1, new_n3460);
xnor_1 g03084(new_n3414, new_n3411, new_n3461);
nor_1  g03085(new_n3403, new_n3400, new_n3462);
nor_1  g03086(new_n2493, new_n1590, new_n3463);
nor_1  g03087(new_n1348, new_n2476, new_n3464);
nand_1 g03088(new_n3464, new_n3463, new_n3465);
nor_1  g03089(new_n3465, new_n3462, new_n3466);
nand_1 g03090(new_n3466, new_n3461, new_n3467);
xnor_1 g03091(new_n3418, new_n3417, new_n3468);
nor_1  g03092(new_n3468, new_n3467, new_n3469);
not_1  g03093(new_n3456_1, new_n3470);
xnor_1 g03094(new_n3459, new_n3470, new_n3471);
nand_1 g03095(new_n3471, new_n3469, new_n3472);
nand_1 g03096(new_n3472, new_n3460, new_n3473);
xnor_1 g03097(new_n3473, new_n3455, new_n3474);
not_1  g03098(new_n3474, new_n3475);
xnor_1 g03099(new_n3471, new_n3469, new_n3476);
not_1  g03100(new_n3476, new_n3477);
nor_1  g03101(new_n2626, new_n1350, new_n3478);
nand_1 g03102(n6877, n6126, new_n3479);
nand_1 g03103(n3719, n2464, new_n3480);
nand_1 g03104(new_n3480, new_n3479, new_n3481);
not_1  g03105(new_n3481, new_n3482);
nand_1 g03106(n6877, n3719, new_n3483);
nand_1 g03107(n6126, n2464, new_n3484);
nor_1  g03108(new_n3484, new_n3483, new_n3485);
nor_1  g03109(new_n1735, new_n2618, new_n3486);
nor_1  g03110(new_n3486, new_n3485, new_n3487);
nor_1  g03111(new_n3487, new_n3482, new_n3488);
nand_1 g03112(new_n3488, new_n3478, new_n3489);
not_1  g03113(new_n3489, new_n3490);
nor_1  g03114(new_n3488, new_n3478, new_n3491);
nor_1  g03115(new_n3491, new_n3490, new_n3492);
nor_1  g03116(new_n2618, new_n1729, new_n3493);
nand_1 g03117(n9400, n6126, new_n3494);
nand_1 g03118(n11311, n3719, new_n3495);
nand_1 g03119(new_n3495, new_n3494, new_n3496);
nor_1  g03120(new_n3495, new_n3494, new_n3497);
not_1  g03121(new_n3497, new_n3498);
nand_1 g03122(new_n3498, new_n3496, new_n3499);
xnor_1 g03123(new_n3499, new_n3493, new_n3500);
nand_1 g03124(new_n3500, new_n3492, new_n3501);
not_1  g03125(new_n3501, new_n3502);
nor_1  g03126(new_n3500, new_n3492, new_n3503);
nor_1  g03127(new_n3503, new_n3502, new_n3504);
not_1  g03128(new_n3486, new_n3505);
not_1  g03129(new_n3483, new_n3506);
nor_1  g03130(new_n3505, new_n3506, new_n3507);
nor_1  g03131(new_n3485, new_n3482, new_n3508);
nor_1  g03132(new_n3508, new_n3507, new_n3509);
not_1  g03133(new_n3509, new_n3510);
nor_1  g03134(new_n3510, new_n3505, new_n3511);
nand_1 g03135(new_n3511, new_n3504, new_n3512);
not_1  g03136(new_n3512, new_n3513);
nor_1  g03137(new_n2623, new_n1350, new_n3514);
nand_1 g03138(n9400, n8595, new_n3515);
not_1  g03139(new_n3515, new_n3516);
not_1  g03140(new_n3496, new_n3517);
nor_1  g03141(new_n3497, new_n3493, new_n3518);
nor_1  g03142(new_n3518, new_n3517, new_n3519);
xnor_1 g03143(new_n3519, new_n3516, new_n3520);
nand_1 g03144(n11311, n3602, new_n3521);
nand_1 g03145(n4187, n3719, new_n3522);
xnor_1 g03146(new_n3522, new_n3484, new_n3523);
xnor_1 g03147(new_n3523, new_n3521, new_n3524);
not_1  g03148(new_n3524, new_n3525);
xnor_1 g03149(new_n3525, new_n3520, new_n3526);
nand_1 g03150(new_n3526, new_n3514, new_n3527);
not_1  g03151(new_n3527, new_n3528);
nor_1  g03152(new_n3526, new_n3514, new_n3529);
nor_1  g03153(new_n3529, new_n3528, new_n3530);
nand_1 g03154(new_n3501, new_n3489, new_n3531);
nor_1  g03155(new_n3531, new_n3530, new_n3532);
nand_1 g03156(new_n3531, new_n3530, new_n3533);
not_1  g03157(new_n3533, new_n3534);
nor_1  g03158(new_n3534, new_n3532, new_n3535);
nand_1 g03159(new_n3535, new_n3513, new_n3536);
nor_1  g03160(new_n2603, new_n1350, new_n3537);
not_1  g03161(new_n3537, new_n3538);
nor_1  g03162(new_n1747, new_n2725, new_n3539);
nand_1 g03163(n4203, n3719, new_n3540);
nand_1 g03164(n4187, n3602, new_n3541);
xnor_1 g03165(new_n3541, new_n3540, new_n3542);
xnor_1 g03166(new_n3542, new_n3539, new_n3543);
nand_1 g03167(new_n3522, new_n3484, new_n3544);
not_1  g03168(new_n3544, new_n3545);
not_1  g03169(new_n3521, new_n3546);
nor_1  g03170(new_n3523, new_n3546, new_n3547);
nor_1  g03171(new_n3547, new_n3545, new_n3548);
nand_1 g03172(new_n3548, new_n3543, new_n3549);
not_1  g03173(new_n3549, new_n3550);
nor_1  g03174(new_n3548, new_n3543, new_n3551);
nor_1  g03175(new_n3551, new_n3550, new_n3552);
nor_1  g03176(new_n2623, new_n1735, new_n3553);
not_1  g03177(new_n3553, new_n3554);
nor_1  g03178(new_n2626, new_n1729, new_n3555);
not_1  g03179(new_n3555, new_n3556);
nand_1 g03180(new_n3556, new_n3554, new_n3557);
nor_1  g03181(new_n3556, new_n3554, new_n3558);
not_1  g03182(new_n3558, new_n3559);
nand_1 g03183(new_n3559, new_n3557, new_n3560);
xnor_1 g03184(new_n3560, new_n3552, new_n3561);
nand_1 g03185(new_n3519, new_n3516, new_n3562);
not_1  g03186(new_n3562, new_n3563);
nor_1  g03187(new_n3524, new_n3520, new_n3564);
nor_1  g03188(new_n3564, new_n3563, new_n3565);
not_1  g03189(new_n3565, new_n3566);
xnor_1 g03190(new_n3566, new_n3561, new_n3567);
not_1  g03191(new_n3567, new_n3568);
nand_1 g03192(new_n3533, new_n3527, new_n3569);
nand_1 g03193(new_n3569, new_n3568, new_n3570);
not_1  g03194(new_n3570, new_n3571);
nor_1  g03195(new_n3569, new_n3568, new_n3572);
nor_1  g03196(new_n3572, new_n3571, new_n3573);
xnor_1 g03197(new_n3573, new_n3538, new_n3574);
nor_1  g03198(new_n3574, new_n3536, new_n3575);
nand_1 g03199(new_n3574, new_n3536, new_n3576);
not_1  g03200(new_n3576, new_n3577);
nor_1  g03201(new_n3577, new_n3575, new_n3578);
not_1  g03202(new_n3578, new_n3579);
xnor_1 g03203(new_n3535, new_n3512, new_n3580);
not_1  g03204(new_n3580, new_n3581);
nor_1  g03205(new_n3511, new_n3504, new_n3582);
nor_1  g03206(new_n3582, new_n3513, new_n3583);
nand_1 g03207(new_n3507, new_n3481, new_n3584);
nand_1 g03208(new_n3584, new_n3510, new_n3585);
not_1  g03209(new_n3585, new_n3586);
nand_1 g03210(n8433, n7236, new_n3587);
nand_1 g03211(n12925, n4805, new_n3588);
nor_1  g03212(new_n3588, new_n3587, new_n3589);
not_1  g03213(new_n3589, new_n3590);
nand_1 g03214(n7733, n4805, new_n3591);
nand_1 g03215(n12925, n11478, new_n3592);
nand_1 g03216(new_n3592, new_n3591, new_n3593);
nor_1  g03217(new_n3592, new_n3591, new_n3594);
not_1  g03218(new_n3594, new_n3595);
nand_1 g03219(new_n3595, new_n3593, new_n3596);
nand_1 g03220(new_n3596, new_n3590, new_n3597);
xnor_1 g03221(new_n3596, new_n3589, new_n3598);
nand_1 g03222(n7236, n405, new_n3599);
nand_1 g03223(n8433, n3992, new_n3600);
xnor_1 g03224(new_n3600, new_n3599, new_n3601);
nand_1 g03225(new_n3601, new_n3598, new_n3602_1);
nand_1 g03226(new_n3602_1, new_n3597, new_n3603);
nor_1  g03227(new_n1835_1, new_n2889, new_n3604);
nand_1 g03228(new_n3604, new_n3587, new_n3605);
nand_1 g03229(n8433, n8384, new_n3606);
nand_1 g03230(n7236, n4086, new_n3607);
nand_1 g03231(new_n3607, new_n3606, new_n3608);
not_1  g03232(new_n3608, new_n3609);
nand_1 g03233(new_n3609, new_n3605, new_n3610);
nor_1  g03234(new_n3607, new_n3606, new_n3611);
not_1  g03235(new_n3611, new_n3612);
nand_1 g03236(new_n3612, new_n3610, new_n3613);
nor_1  g03237(new_n3609, new_n3605, new_n3614);
nor_1  g03238(new_n3614, new_n3613, new_n3615);
xnor_1 g03239(new_n3615, new_n3603, new_n3616_1);
nor_1  g03240(new_n1931, new_n2761, new_n3617);
nand_1 g03241(new_n3617, new_n3588, new_n3618);
nand_1 g03242(n12925, n5283, new_n3619);
nand_1 g03243(n4826, n4805, new_n3620);
nand_1 g03244(new_n3620, new_n3619, new_n3621);
nor_1  g03245(new_n3621, new_n3618, new_n3622);
not_1  g03246(new_n3622, new_n3623);
not_1  g03247(new_n3621, new_n3624);
nor_1  g03248(new_n3620, new_n3619, new_n3625);
nor_1  g03249(new_n3625, new_n3624, new_n3626);
nand_1 g03250(new_n3626, new_n3618, new_n3627_1);
nand_1 g03251(new_n3627_1, new_n3623, new_n3628);
not_1  g03252(new_n3628, new_n3629);
xnor_1 g03253(new_n3629, new_n3616_1, new_n3630);
nand_1 g03254(new_n3630, new_n3586, new_n3631);
not_1  g03255(new_n3631, new_n3632);
nor_1  g03256(new_n3630, new_n3586, new_n3633);
nor_1  g03257(new_n3633, new_n3632, new_n3634);
xnor_1 g03258(new_n3601, new_n3598, new_n3635);
not_1  g03259(new_n3635, new_n3636);
nand_1 g03260(n9400, n3719, new_n3637);
nand_1 g03261(n6877, n3602, new_n3638);
xnor_1 g03262(new_n3638, new_n3637, new_n3639);
nor_1  g03263(new_n3639, new_n3636, new_n3640);
not_1  g03264(new_n3640, new_n3641);
nand_1 g03265(new_n3588, new_n3587, new_n3642);
nand_1 g03266(new_n3642, new_n3590, new_n3643);
nor_1  g03267(new_n3643, new_n3483, new_n3644);
xnor_1 g03268(new_n3639, new_n3635, new_n3645);
nand_1 g03269(new_n3645, new_n3644, new_n3646);
nand_1 g03270(new_n3646, new_n3641, new_n3647);
nand_1 g03271(new_n3647, new_n3634, new_n3648);
nand_1 g03272(new_n3648, new_n3631, new_n3649);
nor_1  g03273(new_n3649, new_n3583, new_n3650);
nor_1  g03274(new_n2770, new_n1925, new_n3651);
not_1  g03275(new_n3625, new_n3652);
nand_1 g03276(new_n3621, new_n3617, new_n3653);
nand_1 g03277(new_n3653, new_n3652, new_n3654_1);
nand_1 g03278(new_n3654_1, new_n3651, new_n3655);
not_1  g03279(new_n3655, new_n3656);
nor_1  g03280(new_n3654_1, new_n3651, new_n3657);
nor_1  g03281(new_n3657, new_n3656, new_n3658);
not_1  g03282(new_n3658, new_n3659);
nor_1  g03283(new_n2761, new_n1923, new_n3660);
nand_1 g03284(n12925, n137, new_n3661_1);
nand_1 g03285(n11478, n4826, new_n3662);
xnor_1 g03286(new_n3662, new_n3661_1, new_n3663);
nand_1 g03287(new_n3663, new_n3660, new_n3664);
nor_1  g03288(new_n3663, new_n3660, new_n3665);
not_1  g03289(new_n3665, new_n3666);
nand_1 g03290(new_n3666, new_n3664, new_n3667);
not_1  g03291(new_n3667, new_n3668);
nor_1  g03292(new_n3668, new_n3659, new_n3669);
nor_1  g03293(new_n3667, new_n3658, new_n3670);
nor_1  g03294(new_n3670, new_n3669, new_n3671);
nor_1  g03295(new_n3626, new_n3595, new_n3672);
xnor_1 g03296(new_n3672, new_n3671, new_n3673);
nor_1  g03297(new_n1833, new_n2898, new_n3674);
nor_1  g03298(new_n3611, new_n3604, new_n3675);
nor_1  g03299(new_n3675, new_n3609, new_n3676);
xnor_1 g03300(new_n3676, new_n3674, new_n3677_1);
nor_1  g03301(new_n1837, new_n2889, new_n3678);
nand_1 g03302(n8433, n6358, new_n3679);
nand_1 g03303(n4086, n3992, new_n3680);
xnor_1 g03304(new_n3680, new_n3679, new_n3681);
xnor_1 g03305(new_n3681, new_n3678, new_n3682);
not_1  g03306(new_n3682, new_n3683);
nor_1  g03307(new_n3683, new_n3677_1, new_n3684);
not_1  g03308(new_n3684, new_n3685);
nand_1 g03309(new_n3683, new_n3677_1, new_n3686);
nand_1 g03310(new_n3686, new_n3685, new_n3687);
nand_1 g03311(new_n3613, new_n3604, new_n3688);
not_1  g03312(new_n3688, new_n3689);
xnor_1 g03313(new_n3689, new_n3687, new_n3690);
xnor_1 g03314(new_n3690, new_n3673, new_n3691);
not_1  g03315(new_n3615, new_n3692);
nand_1 g03316(new_n3692, new_n3603, new_n3693);
nand_1 g03317(new_n3629, new_n3616_1, new_n3694);
nand_1 g03318(new_n3694, new_n3693, new_n3695);
xnor_1 g03319(new_n3695, new_n3691, new_n3696);
not_1  g03320(new_n3650, new_n3697);
nand_1 g03321(new_n3649, new_n3583, new_n3698);
nand_1 g03322(new_n3698, new_n3697, new_n3699);
nor_1  g03323(new_n3699, new_n3696, new_n3700);
nor_1  g03324(new_n3700, new_n3650, new_n3701);
not_1  g03325(new_n3701, new_n3702);
nand_1 g03326(new_n3702, new_n3581, new_n3703);
nand_1 g03327(new_n3701, new_n3580, new_n3704);
nor_1  g03328(new_n3688, new_n3687, new_n3705);
nor_1  g03329(new_n1833, new_n2895, new_n3706);
nor_1  g03330(new_n1835_1, new_n2898, new_n3707);
not_1  g03331(new_n3707, new_n3708);
nand_1 g03332(new_n3680, new_n3679, new_n3709);
not_1  g03333(new_n3709, new_n3710);
nor_1  g03334(new_n3681, new_n3678, new_n3711);
nor_1  g03335(new_n3711, new_n3710, new_n3712);
xnor_1 g03336(new_n3712, new_n3708, new_n3713);
nor_1  g03337(new_n1866, new_n2889, new_n3714);
nand_1 g03338(n8384, n4086, new_n3715);
nand_1 g03339(n8433, n5198, new_n3716);
xnor_1 g03340(new_n3716, new_n3715, new_n3717);
xnor_1 g03341(new_n3717, new_n3714, new_n3718);
xnor_1 g03342(new_n3718, new_n3713, new_n3719_1);
xnor_1 g03343(new_n3719_1, new_n3706, new_n3720);
nand_1 g03344(new_n3676, new_n3674, new_n3721);
nand_1 g03345(new_n3685, new_n3721, new_n3722);
nand_1 g03346(new_n3722, new_n3720, new_n3723);
not_1  g03347(new_n3723, new_n3724);
nor_1  g03348(new_n3722, new_n3720, new_n3725);
nor_1  g03349(new_n3725, new_n3724, new_n3726);
nand_1 g03350(new_n3726, new_n3705, new_n3727);
not_1  g03351(new_n3727, new_n3728);
nor_1  g03352(new_n3726, new_n3705, new_n3729);
nor_1  g03353(new_n3729, new_n3728, new_n3730);
nand_1 g03354(new_n3672, new_n3671, new_n3731);
not_1  g03355(new_n3731, new_n3732);
nor_1  g03356(new_n2767, new_n1925, new_n3733);
nor_1  g03357(new_n1931, new_n2770, new_n3734);
nand_1 g03358(new_n3662, new_n3661_1, new_n3735);
not_1  g03359(new_n3735, new_n3736);
nor_1  g03360(new_n3665, new_n3736, new_n3737);
nand_1 g03361(new_n3737, new_n3734, new_n3738);
not_1  g03362(new_n3738, new_n3739);
nor_1  g03363(new_n3737, new_n3734, new_n3740);
nor_1  g03364(new_n3740, new_n3739, new_n3741);
nor_1  g03365(new_n2761, new_n1959, new_n3742);
nand_1 g03366(n5283, n4826, new_n3743);
nand_1 g03367(n12925, n6294, new_n3744);
xnor_1 g03368(new_n3744, new_n3743, new_n3745);
xnor_1 g03369(new_n3745, new_n3742, new_n3746);
nand_1 g03370(new_n3746, new_n3741, new_n3747);
not_1  g03371(new_n3747, new_n3748);
nor_1  g03372(new_n3746, new_n3741, new_n3749);
nor_1  g03373(new_n3749, new_n3748, new_n3750);
nand_1 g03374(new_n3750, new_n3733, new_n3751);
not_1  g03375(new_n3751, new_n3752);
nor_1  g03376(new_n3750, new_n3733, new_n3753);
nor_1  g03377(new_n3753, new_n3752, new_n3754_1);
nor_1  g03378(new_n3669, new_n3656, new_n3755);
xnor_1 g03379(new_n3755, new_n3754_1, new_n3756);
nand_1 g03380(new_n3756, new_n3732, new_n3757);
not_1  g03381(new_n3757, new_n3758);
nor_1  g03382(new_n3756, new_n3732, new_n3759);
nor_1  g03383(new_n3759, new_n3758, new_n3760);
not_1  g03384(new_n3690, new_n3761);
nand_1 g03385(new_n3761, new_n3673, new_n3762);
nand_1 g03386(new_n3695, new_n3691, new_n3763);
nand_1 g03387(new_n3763, new_n3762, new_n3764);
xnor_1 g03388(new_n3764, new_n3760, new_n3765);
xnor_1 g03389(new_n3765, new_n3730, new_n3766);
nand_1 g03390(new_n3766, new_n3704, new_n3767);
nand_1 g03391(new_n3767, new_n3703, new_n3768);
xnor_1 g03392(new_n3768, new_n3579, new_n3769);
not_1  g03393(new_n3769, new_n3770);
nand_1 g03394(n7236, n6359, new_n3771);
not_1  g03395(n4086, new_n3772);
nor_1  g03396(new_n1866, new_n3772, new_n3773);
nand_1 g03397(new_n3716, new_n3715, new_n3774);
not_1  g03398(new_n3774, new_n3775);
nor_1  g03399(new_n3717, new_n3714, new_n3776);
nor_1  g03400(new_n3776, new_n3775, new_n3777);
nand_1 g03401(new_n3777, new_n3773, new_n3778);
not_1  g03402(new_n3778, new_n3779);
nor_1  g03403(new_n3777, new_n3773, new_n3780);
nor_1  g03404(new_n3780, new_n3779, new_n3781);
nand_1 g03405(n5198, n405, new_n3782);
nand_1 g03406(n8433, n1471, new_n3783);
xnor_1 g03407(new_n3783, new_n3782, new_n3784);
xnor_1 g03408(new_n3784, new_n3781, new_n3785);
nor_1  g03409(new_n1837, new_n2898, new_n3786);
not_1  g03410(new_n3786, new_n3787);
nor_1  g03411(new_n2895, new_n1835_1, new_n3788);
not_1  g03412(new_n3788, new_n3789);
nand_1 g03413(new_n3789, new_n3787, new_n3790);
nor_1  g03414(new_n3789, new_n3787, new_n3791);
not_1  g03415(new_n3791, new_n3792);
nand_1 g03416(new_n3792, new_n3790, new_n3793);
xnor_1 g03417(new_n3793, new_n3785, new_n3794);
nand_1 g03418(new_n3712, new_n3707, new_n3795);
nand_1 g03419(new_n3718, new_n3713, new_n3796);
nand_1 g03420(new_n3796, new_n3795, new_n3797);
xnor_1 g03421(new_n3797, new_n3794, new_n3798);
not_1  g03422(new_n3798, new_n3799);
not_1  g03423(new_n3706, new_n3800);
nor_1  g03424(new_n3719_1, new_n3800, new_n3801);
not_1  g03425(new_n3801, new_n3802);
nand_1 g03426(new_n3723, new_n3802, new_n3803);
nand_1 g03427(new_n3803, new_n3799, new_n3804);
not_1  g03428(new_n3804, new_n3805);
nor_1  g03429(new_n3803, new_n3799, new_n3806);
nor_1  g03430(new_n3806, new_n3805, new_n3807);
xnor_1 g03431(new_n3807, new_n3771, new_n3808);
xnor_1 g03432(new_n3808, new_n3728, new_n3809);
nor_1  g03433(new_n1925, new_n2846, new_n3810);
nand_1 g03434(n4826, n137, new_n3811);
nand_1 g03435(n7733, n6294, new_n3812);
nand_1 g03436(n12925, n6797, new_n3813);
xnor_1 g03437(new_n3813, new_n3812, new_n3814);
nor_1  g03438(new_n3814, new_n3811, new_n3815);
not_1  g03439(new_n3815, new_n3816);
nand_1 g03440(new_n3814, new_n3811, new_n3817);
nand_1 g03441(new_n3817, new_n3816, new_n3818);
nand_1 g03442(new_n3744, new_n3743, new_n3819);
not_1  g03443(new_n3819, new_n3820);
nor_1  g03444(new_n3745, new_n3742, new_n3821);
nor_1  g03445(new_n3821, new_n3820, new_n3822);
xnor_1 g03446(new_n3822, new_n3818, new_n3823);
nor_1  g03447(new_n1931, new_n2767, new_n3824);
not_1  g03448(new_n3824, new_n3825);
nor_1  g03449(new_n2770, new_n1923, new_n3826);
not_1  g03450(new_n3826, new_n3827);
nand_1 g03451(new_n3827, new_n3825, new_n3828);
nor_1  g03452(new_n3827, new_n3825, new_n3829);
not_1  g03453(new_n3829, new_n3830);
nand_1 g03454(new_n3830, new_n3828, new_n3831);
xnor_1 g03455(new_n3831, new_n3823, new_n3832);
nand_1 g03456(new_n3747, new_n3738, new_n3833);
nand_1 g03457(new_n3833, new_n3832, new_n3834);
not_1  g03458(new_n3834, new_n3835);
nor_1  g03459(new_n3833, new_n3832, new_n3836);
nor_1  g03460(new_n3836, new_n3835, new_n3837);
not_1  g03461(new_n3755, new_n3838);
nand_1 g03462(new_n3838, new_n3754_1, new_n3839);
nand_1 g03463(new_n3839, new_n3751, new_n3840);
xnor_1 g03464(new_n3840, new_n3837, new_n3841);
xnor_1 g03465(new_n3841, new_n3810, new_n3842_1);
xnor_1 g03466(new_n3842_1, new_n3758, new_n3843);
xnor_1 g03467(new_n3843, new_n3809, new_n3844);
not_1  g03468(new_n3760, new_n3845);
nand_1 g03469(new_n3764, new_n3845, new_n3846);
not_1  g03470(new_n3730, new_n3847);
nand_1 g03471(new_n3765, new_n3847, new_n3848);
nand_1 g03472(new_n3848, new_n3846, new_n3849_1);
xnor_1 g03473(new_n3849_1, new_n3844, new_n3850);
nor_1  g03474(new_n3850, new_n3770, new_n3851);
not_1  g03475(new_n3850, new_n3852);
nor_1  g03476(new_n3852, new_n3769, new_n3853);
nor_1  g03477(new_n3853, new_n3851, new_n3854);
nor_1  g03478(new_n3854, new_n3477, new_n3855);
not_1  g03479(new_n3855, new_n3856);
nand_1 g03480(new_n3854, new_n3477, new_n3857);
xor_1  g03481(new_n3468, new_n3467, new_n3858);
not_1  g03482(new_n3858, new_n3859);
nand_1 g03483(new_n3704, new_n3703, new_n3860);
xnor_1 g03484(new_n3860, new_n3766, new_n3861);
nor_1  g03485(new_n3861, new_n3859, new_n3862);
xor_1  g03486(new_n3466, new_n3461, new_n3863);
not_1  g03487(new_n3863, new_n3864);
not_1  g03488(new_n3699, new_n3865_1);
xnor_1 g03489(new_n3865_1, new_n3696, new_n3866);
nor_1  g03490(new_n3866, new_n3864, new_n3867);
xnor_1 g03491(new_n3647, new_n3634, new_n3868);
not_1  g03492(new_n3868, new_n3869);
nor_1  g03493(new_n2493, new_n1348, new_n3870);
nor_1  g03494(new_n3870, new_n3405, new_n3871);
nor_1  g03495(new_n3871, new_n3462, new_n3872);
nand_1 g03496(new_n3871, new_n3402, new_n3873);
not_1  g03497(new_n3873, new_n3874);
nor_1  g03498(new_n3874, new_n3872, new_n3875);
nor_1  g03499(new_n3875, new_n3869, new_n3876);
not_1  g03500(new_n3876, new_n3877);
nand_1 g03501(new_n3875, new_n3869, new_n3878);
nand_1 g03502(new_n3878, new_n3877, new_n3879);
not_1  g03503(new_n3879, new_n3880);
xnor_1 g03504(new_n3643, new_n3506, new_n3881);
nand_1 g03505(new_n3881, new_n3870, new_n3882);
not_1  g03506(new_n3463, new_n3883);
xnor_1 g03507(new_n3464, new_n3883, new_n3884);
not_1  g03508(new_n3884, new_n3885);
nand_1 g03509(new_n3885, new_n3882, new_n3886);
xor_1  g03510(new_n3645, new_n3644, new_n3887);
not_1  g03511(new_n3887, new_n3888);
xnor_1 g03512(new_n3884, new_n3882, new_n3889);
nand_1 g03513(new_n3889, new_n3888, new_n3890);
nand_1 g03514(new_n3890, new_n3886, new_n3891);
nand_1 g03515(new_n3891, new_n3880, new_n3892);
nand_1 g03516(new_n3892, new_n3877, new_n3893);
xnor_1 g03517(new_n3866, new_n3864, new_n3894);
nor_1  g03518(new_n3894, new_n3893, new_n3895);
nor_1  g03519(new_n3895, new_n3867, new_n3896);
not_1  g03520(new_n3862, new_n3897);
nand_1 g03521(new_n3861, new_n3859, new_n3898);
nand_1 g03522(new_n3898, new_n3897, new_n3899);
nor_1  g03523(new_n3899, new_n3896, new_n3900);
nor_1  g03524(new_n3900, new_n3862, new_n3901);
nand_1 g03525(new_n3901, new_n3857, new_n3902);
nand_1 g03526(new_n3902, new_n3856, new_n3903);
not_1  g03527(new_n3903, new_n3904);
nor_1  g03528(new_n3904, new_n3475, new_n3905);
nor_1  g03529(new_n3903, new_n3474, new_n3906);
nor_1  g03530(new_n3906, new_n3905, new_n3907);
nor_1  g03531(new_n1735, new_n2603, new_n3908);
nor_1  g03532(new_n2623, new_n1729, new_n3909);
not_1  g03533(new_n3909, new_n3910);
nor_1  g03534(new_n3287_1, new_n1350, new_n3911);
xnor_1 g03535(new_n3911, new_n3910, new_n3912);
not_1  g03536(new_n3912, new_n3913);
nand_1 g03537(new_n3913, new_n3908, new_n3914);
nor_1  g03538(new_n3913, new_n3908, new_n3915);
not_1  g03539(new_n3915, new_n3916);
nand_1 g03540(new_n3916, new_n3914, new_n3917);
not_1  g03541(new_n3539, new_n3918);
nor_1  g03542(new_n3542, new_n3918, new_n3919);
nor_1  g03543(new_n3550, new_n3919, new_n3920);
not_1  g03544(new_n3920, new_n3921);
nand_1 g03545(new_n3921, new_n3917, new_n3922);
not_1  g03546(new_n3917, new_n3923);
nand_1 g03547(new_n3920, new_n3923, new_n3924);
nand_1 g03548(new_n3924, new_n3922, new_n3925);
not_1  g03549(new_n3925, new_n3926);
nor_1  g03550(new_n3541, new_n3540, new_n3927);
nor_1  g03551(new_n1747, new_n2626, new_n3928);
xor_1  g03552(new_n3928, new_n3927, new_n3929);
nor_1  g03553(new_n2119, new_n2618, new_n3930);
nand_1 g03554(n6126, n4187, new_n3931);
nand_1 g03555(n12753, n3719, new_n3932_1);
xnor_1 g03556(new_n3932_1, new_n3931, new_n3933);
xor_1  g03557(new_n3933, new_n3930, new_n3934);
xnor_1 g03558(new_n3934, new_n3929, new_n3935);
xnor_1 g03559(new_n3935, new_n3926, new_n3936);
not_1  g03560(new_n3560, new_n3937);
nand_1 g03561(new_n3937, new_n3552, new_n3938);
nand_1 g03562(new_n3566, new_n3561, new_n3939);
not_1  g03563(new_n3939, new_n3940);
nand_1 g03564(new_n3940, new_n3558, new_n3941);
nand_1 g03565(new_n3939, new_n3559, new_n3942);
nand_1 g03566(new_n3942, new_n3941, new_n3943);
nand_1 g03567(new_n3943, new_n3938, new_n3944);
xnor_1 g03568(new_n3944, new_n3936, new_n3945);
xnor_1 g03569(new_n3945, new_n3570, new_n3946);
nor_1  g03570(new_n3573, new_n3537, new_n3947);
not_1  g03571(new_n3947, new_n3948);
nand_1 g03572(new_n3576, new_n3948, new_n3949);
xnor_1 g03573(new_n3949, new_n3946, new_n3950);
nand_1 g03574(new_n3840, new_n3837, new_n3951);
not_1  g03575(n10965, new_n3952);
nor_1  g03576(new_n3952, new_n1925, new_n3953);
nand_1 g03577(n5283, n4970, new_n3954);
nand_1 g03578(n11478, n503, new_n3955);
xnor_1 g03579(new_n3955, new_n3954, new_n3956);
xor_1  g03580(new_n3956, new_n3953, new_n3957);
not_1  g03581(new_n3818, new_n3958);
nand_1 g03582(new_n3822, new_n3958, new_n3959);
nand_1 g03583(new_n3959, new_n3816, new_n3960);
xnor_1 g03584(new_n3960, new_n3957, new_n3961);
nor_1  g03585(new_n3813, new_n3812, new_n3962);
nor_1  g03586(new_n2770, new_n1959, new_n3963);
xor_1  g03587(new_n3963, new_n3962, new_n3964);
nor_1  g03588(new_n2761, new_n2205, new_n3965);
not_1  g03589(n6294, new_n3966);
nor_1  g03590(new_n3966, new_n2748, new_n3967);
not_1  g03591(new_n3967, new_n3968);
not_1  g03592(n12925, new_n3969);
nor_1  g03593(new_n3969, new_n2363, new_n3970);
not_1  g03594(new_n3970, new_n3971);
nand_1 g03595(new_n3971, new_n3968, new_n3972);
nand_1 g03596(new_n3970, new_n3967, new_n3973);
nand_1 g03597(new_n3973, new_n3972, new_n3974);
xnor_1 g03598(new_n3974, new_n3965, new_n3975);
xnor_1 g03599(new_n3975, new_n3964, new_n3976);
not_1  g03600(new_n3976, new_n3977);
xnor_1 g03601(new_n3977, new_n3961, new_n3978);
not_1  g03602(new_n3831, new_n3979);
nand_1 g03603(new_n3979, new_n3823, new_n3980);
nand_1 g03604(new_n3835, new_n3829, new_n3981);
nand_1 g03605(new_n3834, new_n3830, new_n3982);
nand_1 g03606(new_n3982, new_n3981, new_n3983);
nand_1 g03607(new_n3983, new_n3980, new_n3984);
xnor_1 g03608(new_n3984, new_n3978, new_n3985);
xnor_1 g03609(new_n3985, new_n3951, new_n3986_1);
not_1  g03610(new_n3810, new_n3987);
nand_1 g03611(new_n3841, new_n3987, new_n3988);
nand_1 g03612(new_n3842_1, new_n3757, new_n3989);
nand_1 g03613(new_n3989, new_n3988, new_n3990);
not_1  g03614(new_n3990, new_n3991);
xnor_1 g03615(new_n3991, new_n3986_1, new_n3992_1);
nor_1  g03616(new_n2969, new_n1833, new_n3993);
nand_1 g03617(n8384, n6611, new_n3994);
nand_1 g03618(n6359, n3992, new_n3995);
xnor_1 g03619(new_n3995, new_n3994, new_n3996);
xor_1  g03620(new_n3996, new_n3993, new_n3997);
not_1  g03621(new_n3784, new_n3998);
nand_1 g03622(new_n3998, new_n3781, new_n3999);
nand_1 g03623(new_n3999, new_n3778, new_n4000);
xnor_1 g03624(new_n4000, new_n3997, new_n4001);
nor_1  g03625(new_n3783, new_n3782, new_n4002);
nor_1  g03626(new_n1866, new_n2898, new_n4003);
xor_1  g03627(new_n4003, new_n4002, new_n4004);
nor_1  g03628(new_n2154, new_n2889, new_n4005_1);
not_1  g03629(n5198, new_n4006);
nor_1  g03630(new_n4006, new_n3772, new_n4007);
not_1  g03631(new_n4007, new_n4008);
not_1  g03632(n7646, new_n4009);
not_1  g03633(n8433, new_n4010);
nor_1  g03634(new_n4010, new_n4009, new_n4011);
not_1  g03635(new_n4011, new_n4012);
nand_1 g03636(new_n4012, new_n4008, new_n4013);
nand_1 g03637(new_n4011, new_n4007, new_n4014);
nand_1 g03638(new_n4014, new_n4013, new_n4015);
xnor_1 g03639(new_n4015, new_n4005_1, new_n4016);
not_1  g03640(new_n4016, new_n4017);
xnor_1 g03641(new_n4017, new_n4004, new_n4018);
xnor_1 g03642(new_n4018, new_n4001, new_n4019);
not_1  g03643(new_n3785, new_n4020);
nor_1  g03644(new_n3793, new_n4020, new_n4021);
not_1  g03645(new_n4021, new_n4022);
nand_1 g03646(new_n3797, new_n3794, new_n4023);
xnor_1 g03647(new_n4023, new_n3792, new_n4024);
nand_1 g03648(new_n4024, new_n4022, new_n4025);
xnor_1 g03649(new_n4025, new_n4019, new_n4026);
xnor_1 g03650(new_n4026, new_n3804, new_n4027);
not_1  g03651(new_n3807, new_n4028);
nand_1 g03652(new_n4028, new_n3771, new_n4029);
nand_1 g03653(new_n3808, new_n3727, new_n4030);
nand_1 g03654(new_n4030, new_n4029, new_n4031);
xnor_1 g03655(new_n4031, new_n4027, new_n4032);
xnor_1 g03656(new_n4032, new_n3992_1, new_n4033);
nand_1 g03657(new_n3843, new_n3809, new_n4034);
not_1  g03658(new_n3844, new_n4035);
nand_1 g03659(new_n3849_1, new_n4035, new_n4036);
nand_1 g03660(new_n4036, new_n4034, new_n4037);
xnor_1 g03661(new_n4037, new_n4033, new_n4038);
xnor_1 g03662(new_n4038, new_n3950, new_n4039);
nor_1  g03663(new_n3768, new_n3578, new_n4040);
nor_1  g03664(new_n3851, new_n4040, new_n4041);
xnor_1 g03665(new_n4041, new_n4039, new_n4042);
xnor_1 g03666(new_n4042, new_n3907, n844);
not_1  g03667(n7456, new_n4044);
nor_1  g03668(new_n4044, new_n378, new_n4045);
nand_1 g03669(n12591, n6687, new_n4046);
nand_1 g03670(n4189, n1798, new_n4047);
nand_1 g03671(new_n4047, new_n4046, new_n4048);
not_1  g03672(new_n4048, new_n4049);
nand_1 g03673(n6687, n1798, new_n4050);
nand_1 g03674(n12591, n4189, new_n4051);
nor_1  g03675(new_n4051, new_n4050, new_n4052);
not_1  g03676(n3932, new_n4053);
nor_1  g03677(new_n4053, new_n1377, new_n4054);
nor_1  g03678(new_n4054, new_n4052, new_n4055);
nor_1  g03679(new_n4055, new_n4049, new_n4056);
nand_1 g03680(new_n4056, new_n4045, new_n4057);
not_1  g03681(new_n4057, new_n4058);
nor_1  g03682(new_n4056, new_n4045, new_n4059);
nor_1  g03683(new_n4059, new_n4058, new_n4060);
nor_1  g03684(new_n1367, new_n4053, new_n4061);
not_1  g03685(new_n4061, new_n4062);
nand_1 g03686(n12591, n2564, new_n4063);
nand_1 g03687(n6770, n1798, new_n4064);
nand_1 g03688(new_n4064, new_n4063, new_n4065);
not_1  g03689(new_n4065, new_n4066);
nor_1  g03690(new_n4064, new_n4063, new_n4067);
nor_1  g03691(new_n4067, new_n4066, new_n4068);
xnor_1 g03692(new_n4068, new_n4062, new_n4069);
nand_1 g03693(new_n4069, new_n4060, new_n4070);
not_1  g03694(new_n4070, new_n4071);
nor_1  g03695(new_n4069, new_n4060, new_n4072);
nor_1  g03696(new_n4072, new_n4071, new_n4073);
not_1  g03697(new_n4054, new_n4074);
not_1  g03698(new_n4050, new_n4075);
nor_1  g03699(new_n4074, new_n4075, new_n4076);
nor_1  g03700(new_n4052, new_n4049, new_n4077);
nor_1  g03701(new_n4077, new_n4076, new_n4078);
not_1  g03702(new_n4078, new_n4079);
nor_1  g03703(new_n4079, new_n4074, new_n4080);
xor_1  g03704(new_n4080, new_n4073, new_n4081);
not_1  g03705(new_n4081, new_n4082);
nand_1 g03706(new_n4076, new_n4048, new_n4083);
nand_1 g03707(new_n4083, new_n4079, new_n4084);
not_1  g03708(n6703, new_n4085);
nor_1  g03709(new_n382, new_n4085, new_n4086_1);
not_1  g03710(new_n4086_1, new_n4087);
not_1  g03711(n11876, new_n4088_1);
nor_1  g03712(new_n4088_1, new_n385, new_n4089);
not_1  g03713(new_n4089, new_n4090);
nand_1 g03714(n12069, n5645, new_n4091);
nor_1  g03715(new_n4091, new_n4090, new_n4092);
not_1  g03716(new_n4092, new_n4093);
nand_1 g03717(new_n4091, new_n4090, new_n4094_1);
nand_1 g03718(new_n4094_1, new_n4093, new_n4095);
nor_1  g03719(new_n4095, new_n4087, new_n4096);
nand_1 g03720(n9640, n8336, new_n4097);
nand_1 g03721(n10928, n6703, new_n4098);
xnor_1 g03722(new_n4098, new_n4097, new_n4099);
not_1  g03723(new_n4099, new_n4100);
nand_1 g03724(new_n4100, new_n4096, new_n4101);
nand_1 g03725(n12391, n5645, new_n4102);
nand_1 g03726(n12069, n1067, new_n4103);
nand_1 g03727(new_n4103, new_n4102, new_n4104);
nor_1  g03728(new_n4103, new_n4102, new_n4105);
not_1  g03729(new_n4105, new_n4106);
nand_1 g03730(new_n4106, new_n4104, new_n4107);
xnor_1 g03731(new_n4107, new_n4092, new_n4108);
nand_1 g03732(n11222, n10898, new_n4109);
nand_1 g03733(n11876, n11153, new_n4110);
xnor_1 g03734(new_n4110, new_n4109, new_n4111);
xnor_1 g03735(new_n4111, new_n4108, new_n4112);
xnor_1 g03736(new_n4099, new_n4096, new_n4113);
nand_1 g03737(new_n4113, new_n4112, new_n4114);
nand_1 g03738(new_n4114, new_n4101, new_n4115);
not_1  g03739(n9640, new_n4116);
nor_1  g03740(new_n1434, new_n4116, new_n4117);
not_1  g03741(new_n4117, new_n4118);
nor_1  g03742(new_n4118, new_n4086_1, new_n4119);
nand_1 g03743(n6986, n6703, new_n4120);
nand_1 g03744(n8336, n3022, new_n4121);
nand_1 g03745(new_n4121, new_n4120, new_n4122);
not_1  g03746(new_n4122, new_n4123);
nand_1 g03747(n6986, n3022, new_n4124);
nor_1  g03748(new_n4124, new_n4087, new_n4125);
nor_1  g03749(new_n4125, new_n4123, new_n4126);
nor_1  g03750(new_n4126, new_n4119, new_n4127);
not_1  g03751(new_n4127, new_n4128);
nand_1 g03752(new_n4122, new_n4119, new_n4129);
nand_1 g03753(new_n4129, new_n4128, new_n4130);
xnor_1 g03754(new_n4130, new_n4115, new_n4131);
not_1  g03755(n8665, new_n4132);
nor_1  g03756(new_n1533, new_n4132, new_n4133);
not_1  g03757(new_n4133, new_n4134);
nand_1 g03758(n12391, n1067, new_n4135);
nand_1 g03759(n7891, n5645, new_n4136);
xnor_1 g03760(new_n4136, new_n4135, new_n4137);
xnor_1 g03761(new_n4137, new_n4134, new_n4138);
xnor_1 g03762(new_n4138, new_n4106, new_n4139);
nand_1 g03763(new_n4107, new_n4093, new_n4140);
nand_1 g03764(new_n4111, new_n4108, new_n4141_1);
nand_1 g03765(new_n4141_1, new_n4140, new_n4142);
not_1  g03766(n10898, new_n4143);
nor_1  g03767(new_n1467, new_n4143, new_n4144);
nand_1 g03768(new_n4144, new_n4090, new_n4145);
nand_1 g03769(n11876, n5314, new_n4146);
nand_1 g03770(n11222, n3754, new_n4147);
nand_1 g03771(new_n4147, new_n4146, new_n4148);
not_1  g03772(new_n4148, new_n4149);
nand_1 g03773(new_n4149, new_n4145, new_n4150);
nand_1 g03774(n5314, n3754, new_n4151);
nor_1  g03775(new_n4151, new_n4090, new_n4152);
not_1  g03776(new_n4152, new_n4153);
nand_1 g03777(new_n4153, new_n4150, new_n4154);
nor_1  g03778(new_n4149, new_n4145, new_n4155_1);
nor_1  g03779(new_n4155_1, new_n4154, new_n4156);
xnor_1 g03780(new_n4156, new_n4142, new_n4157);
nor_1  g03781(new_n4157, new_n4139, new_n4158);
nand_1 g03782(new_n4157, new_n4139, new_n4159_1);
not_1  g03783(new_n4159_1, new_n4160);
nor_1  g03784(new_n4160, new_n4158, new_n4161);
nand_1 g03785(new_n4161, new_n4131, new_n4162);
not_1  g03786(new_n4162, new_n4163);
nor_1  g03787(new_n4161, new_n4131, new_n4164);
nor_1  g03788(new_n4164, new_n4163, new_n4165);
nor_1  g03789(new_n4165, new_n4084, new_n4166);
xnor_1 g03790(new_n4095, new_n4086_1, new_n4167);
nand_1 g03791(new_n4167, new_n4075, new_n4168);
nand_1 g03792(n2564, n1798, new_n4169);
nor_1  g03793(new_n378, new_n4053, new_n4170);
xnor_1 g03794(new_n4170, new_n4169, new_n4171);
not_1  g03795(new_n4171, new_n4172);
nand_1 g03796(new_n4172, new_n4168, new_n4173);
not_1  g03797(new_n4173, new_n4174);
xor_1  g03798(new_n4113, new_n4112, new_n4175);
nor_1  g03799(new_n4172, new_n4168, new_n4176);
nor_1  g03800(new_n4176, new_n4174, new_n4177);
not_1  g03801(new_n4177, new_n4178);
nor_1  g03802(new_n4178, new_n4175, new_n4179);
nor_1  g03803(new_n4179, new_n4174, new_n4180);
not_1  g03804(new_n4180, new_n4181);
xnor_1 g03805(new_n4165, new_n4084, new_n4182);
nor_1  g03806(new_n4182, new_n4181, new_n4183);
nor_1  g03807(new_n4183, new_n4166, new_n4184);
xnor_1 g03808(new_n4184, new_n4082, new_n4185);
nor_1  g03809(new_n4138, new_n4106, new_n4186);
not_1  g03810(n11922, new_n4187_1);
nor_1  g03811(new_n1533, new_n4187_1, new_n4188);
not_1  g03812(new_n4188, new_n4189_1);
nand_1 g03813(new_n4136, new_n4135, new_n4190_1);
not_1  g03814(new_n4190_1, new_n4191);
nor_1  g03815(new_n4137, new_n4133, new_n4192);
nor_1  g03816(new_n4192, new_n4191, new_n4193);
xnor_1 g03817(new_n4193, new_n4189_1, new_n4194);
not_1  g03818(n5645, new_n4195);
nor_1  g03819(new_n1538, new_n4195, new_n4196);
not_1  g03820(new_n4196, new_n4197);
nand_1 g03821(n7891, n1067, new_n4198);
nand_1 g03822(n12391, n8665, new_n4199);
xnor_1 g03823(new_n4199, new_n4198, new_n4200);
xnor_1 g03824(new_n4200, new_n4197, new_n4201);
xnor_1 g03825(new_n4201, new_n4194, new_n4202);
xnor_1 g03826(new_n4202, new_n4186, new_n4203_1);
not_1  g03827(n2749, new_n4204);
nor_1  g03828(new_n385, new_n4204, new_n4205);
nor_1  g03829(new_n4152, new_n4144, new_n4206);
nor_1  g03830(new_n4206, new_n4149, new_n4207);
nand_1 g03831(new_n4207, new_n4205, new_n4208);
not_1  g03832(new_n4208, new_n4209);
nor_1  g03833(new_n4207, new_n4205, new_n4210);
nor_1  g03834(new_n4210, new_n4209, new_n4211);
nor_1  g03835(new_n4143, new_n1562, new_n4212);
not_1  g03836(new_n4212, new_n4213);
nand_1 g03837(n11153, n3754, new_n4214);
nand_1 g03838(n11876, n996, new_n4215);
xnor_1 g03839(new_n4215, new_n4214, new_n4216);
xnor_1 g03840(new_n4216, new_n4213, new_n4217);
not_1  g03841(new_n4217, new_n4218);
xnor_1 g03842(new_n4218, new_n4211, new_n4219);
nand_1 g03843(new_n4154, new_n4144, new_n4220);
not_1  g03844(new_n4220, new_n4221);
xnor_1 g03845(new_n4221, new_n4219, new_n4222);
xnor_1 g03846(new_n4222, new_n4203_1, new_n4223);
not_1  g03847(new_n4156, new_n4224);
nand_1 g03848(new_n4224, new_n4142, new_n4225);
nand_1 g03849(new_n4159_1, new_n4225, new_n4226_1);
nand_1 g03850(new_n4226_1, new_n4223, new_n4227);
not_1  g03851(new_n4227, new_n4228);
nor_1  g03852(new_n4226_1, new_n4223, new_n4229);
nor_1  g03853(new_n4229, new_n4228, new_n4230_1);
not_1  g03854(new_n4230_1, new_n4231);
not_1  g03855(n11023, new_n4232);
nor_1  g03856(new_n4232, new_n382, new_n4233);
nor_1  g03857(new_n4125, new_n4117, new_n4234);
nor_1  g03858(new_n4234, new_n4123, new_n4235);
xnor_1 g03859(new_n4235, new_n4233, new_n4236);
nor_1  g03860(new_n4116, new_n1508, new_n4237);
nand_1 g03861(n10928, n3022, new_n4238);
nand_1 g03862(n6703, n2226, new_n4239);
nand_1 g03863(new_n4239, new_n4238, new_n4240);
nor_1  g03864(new_n4239, new_n4238, new_n4241);
not_1  g03865(new_n4241, new_n4242);
nand_1 g03866(new_n4242, new_n4240, new_n4243);
xnor_1 g03867(new_n4243, new_n4237, new_n4244);
xnor_1 g03868(new_n4244, new_n4236, new_n4245);
nor_1  g03869(new_n4128, new_n4118, new_n4246);
nor_1  g03870(new_n4246, new_n4245, new_n4247);
nand_1 g03871(new_n4246, new_n4245, new_n4248);
not_1  g03872(new_n4248, new_n4249);
nor_1  g03873(new_n4249, new_n4247, new_n4250);
not_1  g03874(new_n4250, new_n4251);
not_1  g03875(new_n4130, new_n4252);
nor_1  g03876(new_n4252, new_n4115, new_n4253);
nor_1  g03877(new_n4163, new_n4253, new_n4254);
not_1  g03878(new_n4254, new_n4255);
nor_1  g03879(new_n4255, new_n4251, new_n4256);
nor_1  g03880(new_n4254, new_n4250, new_n4257);
nor_1  g03881(new_n4257, new_n4256, new_n4258);
nor_1  g03882(new_n4258, new_n4231, new_n4259);
nand_1 g03883(new_n4258, new_n4231, new_n4260);
not_1  g03884(new_n4260, new_n4261);
nor_1  g03885(new_n4261, new_n4259, new_n4262);
xnor_1 g03886(new_n4262, new_n4185, n911);
nor_1  g03887(new_n378, new_n2484, new_n4264);
nand_1 g03888(n11917, n6687, new_n4265);
nand_1 g03889(n9956, n4189, new_n4266);
nand_1 g03890(new_n4266, new_n4265, new_n4267);
not_1  g03891(new_n4267, new_n4268);
nor_1  g03892(new_n2493, new_n378, new_n4269);
not_1  g03893(new_n4269, new_n4270);
nand_1 g03894(n11917, n4189, new_n4271);
nor_1  g03895(new_n4271, new_n4270, new_n4272);
nor_1  g03896(new_n2476, new_n1377, new_n4273);
nor_1  g03897(new_n4273, new_n4272, new_n4274);
nor_1  g03898(new_n4274, new_n4268, new_n4275);
nand_1 g03899(new_n4275, new_n4264, new_n4276);
not_1  g03900(new_n4276, new_n4277);
nor_1  g03901(new_n4275, new_n4264, new_n4278);
nor_1  g03902(new_n4278, new_n4277, new_n4279);
nor_1  g03903(new_n2476, new_n1367, new_n4280);
nor_1  g03904(new_n2462, new_n1377, new_n4281);
not_1  g03905(new_n4281, new_n4282);
not_1  g03906(n6770, new_n4283);
nor_1  g03907(new_n2493, new_n4283, new_n4284);
not_1  g03908(new_n4284, new_n4285);
nand_1 g03909(new_n4285, new_n4282, new_n4286);
nor_1  g03910(new_n4285, new_n4282, new_n4287);
not_1  g03911(new_n4287, new_n4288);
nand_1 g03912(new_n4288, new_n4286, new_n4289);
xnor_1 g03913(new_n4289, new_n4280, new_n4290);
nand_1 g03914(new_n4290, new_n4279, new_n4291);
not_1  g03915(new_n4291, new_n4292);
nor_1  g03916(new_n4290, new_n4279, new_n4293);
nor_1  g03917(new_n4293, new_n4292, new_n4294);
nor_1  g03918(new_n4272, new_n4268, new_n4295);
not_1  g03919(new_n4295, new_n4296);
nor_1  g03920(new_n2493, new_n1377, new_n4297);
nor_1  g03921(new_n378, new_n2476, new_n4298);
and_1  g03922(new_n4298, new_n4297, new_n4299);
nand_1 g03923(new_n4299, new_n4296, new_n4300_1);
not_1  g03924(new_n4300_1, new_n4301);
and_1  g03925(new_n4301, new_n4294, new_n4302);
nor_1  g03926(new_n378, new_n2481, new_n4303);
nand_1 g03927(new_n4291, new_n4276, new_n4304);
nand_1 g03928(new_n4304, new_n4303, new_n4305);
not_1  g03929(new_n4305, new_n4306);
nor_1  g03930(new_n4304, new_n4303, new_n4307);
nor_1  g03931(new_n4307, new_n4306, new_n4308);
nor_1  g03932(new_n2484, new_n1377, new_n4309);
not_1  g03933(new_n4286, new_n4310);
nor_1  g03934(new_n4287, new_n4280, new_n4311);
nor_1  g03935(new_n4311, new_n4310, new_n4312_1);
nand_1 g03936(new_n4312_1, new_n4309, new_n4313);
not_1  g03937(new_n4313, new_n4314);
nor_1  g03938(new_n4312_1, new_n4309, new_n4315);
nor_1  g03939(new_n4315, new_n4314, new_n4316);
nor_1  g03940(new_n4283, new_n2476, new_n4317);
nand_1 g03941(n9956, n9920, new_n4318);
xnor_1 g03942(new_n4318, new_n4271, new_n4319);
xnor_1 g03943(new_n4319, new_n4317, new_n4320);
nand_1 g03944(new_n4320, new_n4316, new_n4321);
not_1  g03945(new_n4321, new_n4322);
nor_1  g03946(new_n4320, new_n4316, new_n4323);
nor_1  g03947(new_n4323, new_n4322, new_n4324);
nand_1 g03948(new_n4324, new_n4308, new_n4325);
not_1  g03949(new_n4325, new_n4326_1);
nor_1  g03950(new_n4324, new_n4308, new_n4327);
nor_1  g03951(new_n4327, new_n4326_1, new_n4328);
nand_1 g03952(new_n4328, new_n4302, new_n4329);
not_1  g03953(new_n4329, new_n4330);
nor_1  g03954(new_n4328, new_n4302, new_n4331);
nor_1  g03955(new_n4331, new_n4330, new_n4332);
nor_1  g03956(new_n4301, new_n4294, new_n4333_1);
nor_1  g03957(new_n4333_1, new_n4302, new_n4334);
not_1  g03958(new_n4334, new_n4335);
nor_1  g03959(new_n2626, new_n382, new_n4336);
nand_1 g03960(n8336, n6126, new_n4337);
nand_1 g03961(n6986, n3719, new_n4338);
nand_1 g03962(new_n4338, new_n4337, new_n4339);
not_1  g03963(new_n4339, new_n4340);
nand_1 g03964(n8336, n3719, new_n4341);
nand_1 g03965(n6986, n6126, new_n4342);
nor_1  g03966(new_n4342, new_n4341, new_n4343);
nor_1  g03967(new_n1434, new_n2618, new_n4344);
nor_1  g03968(new_n4344, new_n4343, new_n4345);
nor_1  g03969(new_n4345, new_n4340, new_n4346);
nand_1 g03970(new_n4346, new_n4336, new_n4347);
not_1  g03971(new_n4347, new_n4348);
nor_1  g03972(new_n4346, new_n4336, new_n4349);
nor_1  g03973(new_n4349, new_n4348, new_n4350);
nor_1  g03974(new_n1508, new_n2618, new_n4351);
nand_1 g03975(n10928, n6126, new_n4352);
nand_1 g03976(n3719, n2226, new_n4353);
nand_1 g03977(new_n4353, new_n4352, new_n4354);
not_1  g03978(new_n4352, new_n4355);
not_1  g03979(new_n4353, new_n4356);
nand_1 g03980(new_n4356, new_n4355, new_n4357);
nand_1 g03981(new_n4357, new_n4354, new_n4358);
xnor_1 g03982(new_n4358, new_n4351, new_n4359);
nand_1 g03983(new_n4359, new_n4350, new_n4360);
not_1  g03984(new_n4360, new_n4361);
nor_1  g03985(new_n4359, new_n4350, new_n4362);
nor_1  g03986(new_n4362, new_n4361, new_n4363);
not_1  g03987(new_n4344, new_n4364);
and_1  g03988(new_n4344, new_n4341, new_n4365);
nor_1  g03989(new_n4343, new_n4340, new_n4366);
nor_1  g03990(new_n4366, new_n4365, new_n4367);
not_1  g03991(new_n4367, new_n4368);
nor_1  g03992(new_n4368, new_n4364, new_n4369);
nor_1  g03993(new_n4369, new_n4363, new_n4370_1);
nand_1 g03994(new_n4369, new_n4363, new_n4371);
not_1  g03995(new_n4371, new_n4372);
nor_1  g03996(new_n4372, new_n4370_1, new_n4373);
nor_1  g03997(new_n1533, new_n2770, new_n4374);
nand_1 g03998(n12069, n4826, new_n4375);
nand_1 g03999(n12925, n7891, new_n4376);
nand_1 g04000(new_n4376, new_n4375, new_n4377);
not_1  g04001(new_n4377, new_n4378_1);
nand_1 g04002(n12925, n12069, new_n4379);
nand_1 g04003(n7891, n4826, new_n4380);
nor_1  g04004(new_n4380, new_n4379, new_n4381);
nor_1  g04005(new_n1452, new_n2761, new_n4382);
nor_1  g04006(new_n4382, new_n4381, new_n4383);
nor_1  g04007(new_n4383, new_n4378_1, new_n4384);
xnor_1 g04008(new_n4384, new_n4374, new_n4385);
not_1  g04009(n7891, new_n4386);
nor_1  g04010(new_n4386, new_n2761, new_n4387);
nand_1 g04011(n12925, n7160, new_n4388);
nand_1 g04012(n12391, n4826, new_n4389);
xnor_1 g04013(new_n4389, new_n4388, new_n4390);
xnor_1 g04014(new_n4390, new_n4387, new_n4391);
not_1  g04015(new_n4391, new_n4392);
nor_1  g04016(new_n4392, new_n4385, new_n4393);
not_1  g04017(new_n4393, new_n4394);
nand_1 g04018(new_n4392, new_n4385, new_n4395);
nand_1 g04019(new_n4395, new_n4394, new_n4396);
nor_1  g04020(new_n4381, new_n4378_1, new_n4397_1);
not_1  g04021(new_n4397_1, new_n4398);
nand_1 g04022(n12925, n12391, new_n4399);
nand_1 g04023(n12069, n7733, new_n4400);
nor_1  g04024(new_n4400, new_n4399, new_n4401);
nand_1 g04025(new_n4401, new_n4398, new_n4402);
not_1  g04026(new_n4402, new_n4403);
xnor_1 g04027(new_n4403, new_n4396, new_n4404);
nor_1  g04028(new_n385, new_n2898, new_n4405);
nand_1 g04029(n8433, n5314, new_n4406);
nand_1 g04030(n11222, n4086, new_n4407);
nand_1 g04031(new_n4407, new_n4406, new_n4408);
not_1  g04032(new_n4408, new_n4409);
nor_1  g04033(new_n4407, new_n4406, new_n4410);
nor_1  g04034(new_n1467, new_n2889, new_n4411);
nor_1  g04035(new_n4411, new_n4410, new_n4412);
nor_1  g04036(new_n4412, new_n4409, new_n4413);
nand_1 g04037(new_n4413, new_n4405, new_n4414);
not_1  g04038(new_n4414, new_n4415);
nor_1  g04039(new_n4413, new_n4405, new_n4416);
nor_1  g04040(new_n4416, new_n4415, new_n4417);
nand_1 g04041(n5314, n405, new_n4418);
nand_1 g04042(n8433, n996, new_n4419);
nand_1 g04043(n11153, n4086, new_n4420);
nand_1 g04044(new_n4420, new_n4419, new_n4421);
not_1  g04045(new_n4421, new_n4422);
nor_1  g04046(new_n4420, new_n4419, new_n4423);
nor_1  g04047(new_n4423, new_n4422, new_n4424);
xnor_1 g04048(new_n4424, new_n4418, new_n4425);
xnor_1 g04049(new_n4425, new_n4417, new_n4426);
not_1  g04050(new_n4426, new_n4427);
not_1  g04051(new_n4411, new_n4428);
nor_1  g04052(new_n385, new_n4010, new_n4429);
nor_1  g04053(new_n4429, new_n4428, new_n4430);
nor_1  g04054(new_n4430, new_n4408, new_n4431);
nor_1  g04055(new_n4431, new_n4410, new_n4432);
nor_1  g04056(new_n4432, new_n4428, new_n4433);
nand_1 g04057(new_n4433, new_n4427, new_n4434);
not_1  g04058(new_n4434, new_n4435);
nor_1  g04059(new_n4433, new_n4427, new_n4436_1);
nor_1  g04060(new_n4436_1, new_n4435, new_n4437);
nand_1 g04061(new_n4437, new_n4404, new_n4438);
not_1  g04062(new_n4404, new_n4439);
not_1  g04063(new_n4437, new_n4440);
nand_1 g04064(new_n4440, new_n4439, new_n4441);
nand_1 g04065(new_n4441, new_n4438, new_n4442);
not_1  g04066(new_n4379, new_n4443);
nand_1 g04067(new_n4429, new_n4443, new_n4444);
nand_1 g04068(n11153, n8433, new_n4445);
nand_1 g04069(n11222, n405, new_n4446);
xnor_1 g04070(new_n4446, new_n4445, new_n4447);
nand_1 g04071(new_n4447, new_n4444, new_n4448);
xnor_1 g04072(new_n4447, new_n4444, new_n4449);
not_1  g04073(new_n4449, new_n4450);
xnor_1 g04074(new_n4400, new_n4399, new_n4451);
nand_1 g04075(new_n4451, new_n4450, new_n4452);
nand_1 g04076(new_n4452, new_n4448, new_n4453);
nand_1 g04077(new_n4430, new_n4408, new_n4454);
nand_1 g04078(new_n4454, new_n4432, new_n4455);
nand_1 g04079(new_n4455, new_n4453, new_n4456);
not_1  g04080(new_n4455, new_n4457);
xnor_1 g04081(new_n4457, new_n4453, new_n4458);
nand_1 g04082(new_n4382, new_n4379, new_n4459);
and_1  g04083(new_n4459, new_n4398, new_n4460);
nor_1  g04084(new_n4459, new_n4378_1, new_n4461);
nor_1  g04085(new_n4461, new_n4460, new_n4462);
not_1  g04086(new_n4462, new_n4463);
nand_1 g04087(new_n4463, new_n4458, new_n4464);
nand_1 g04088(new_n4464, new_n4456, new_n4465);
xnor_1 g04089(new_n4465, new_n4442, new_n4466);
xnor_1 g04090(new_n4466, new_n4373, new_n4467);
nand_1 g04091(new_n4365, new_n4339, new_n4468);
nand_1 g04092(new_n4468, new_n4368, new_n4469);
xnor_1 g04093(new_n4462, new_n4458, new_n4470);
nor_1  g04094(new_n4470, new_n4469, new_n4471);
xnor_1 g04095(new_n4470, new_n4469, new_n4472);
xnor_1 g04096(new_n4451, new_n4449, new_n4473);
nand_1 g04097(n10928, n3719, new_n4474);
nand_1 g04098(n8336, n3602, new_n4475);
xnor_1 g04099(new_n4475, new_n4474, new_n4476);
nor_1  g04100(new_n4476, new_n4473, new_n4477);
not_1  g04101(new_n4429, new_n4478);
nand_1 g04102(new_n4478, new_n4379, new_n4479);
nand_1 g04103(new_n4479, new_n4444, new_n4480);
nor_1  g04104(new_n4480, new_n4341, new_n4481);
not_1  g04105(new_n4481, new_n4482);
xnor_1 g04106(new_n4476, new_n4473, new_n4483);
nor_1  g04107(new_n4483, new_n4482, new_n4484);
nor_1  g04108(new_n4484, new_n4477, new_n4485);
nor_1  g04109(new_n4485, new_n4472, new_n4486);
nor_1  g04110(new_n4486, new_n4471, new_n4487);
xnor_1 g04111(new_n4487, new_n4467, new_n4488);
not_1  g04112(new_n4488, new_n4489);
nand_1 g04113(new_n4489, new_n4335, new_n4490);
xnor_1 g04114(new_n4485, new_n4472, new_n4491);
not_1  g04115(new_n4491, new_n4492);
nand_1 g04116(new_n4273, new_n4270, new_n4493);
and_1  g04117(new_n4493, new_n4296, new_n4494);
nor_1  g04118(new_n4493, new_n4268, new_n4495);
nor_1  g04119(new_n4495, new_n4494, new_n4496);
nor_1  g04120(new_n4496, new_n4492, new_n4497);
not_1  g04121(new_n4497, new_n4498);
xnor_1 g04122(new_n4496, new_n4491, new_n4499_1);
and_1  g04123(new_n4480, new_n4341, new_n4500);
nor_1  g04124(new_n4500, new_n4481, new_n4501);
nand_1 g04125(new_n4501, new_n4269, new_n4502);
xor_1  g04126(new_n4298, new_n4297, new_n4503);
not_1  g04127(new_n4503, new_n4504);
nand_1 g04128(new_n4504, new_n4502, new_n4505);
xnor_1 g04129(new_n4483, new_n4481, new_n4506);
not_1  g04130(new_n4506, new_n4507);
xnor_1 g04131(new_n4503, new_n4502, new_n4508);
nand_1 g04132(new_n4508, new_n4507, new_n4509);
nand_1 g04133(new_n4509, new_n4505, new_n4510);
nand_1 g04134(new_n4510, new_n4499_1, new_n4511);
nand_1 g04135(new_n4511, new_n4498, new_n4512);
xnor_1 g04136(new_n4488, new_n4335, new_n4513);
nand_1 g04137(new_n4513, new_n4512, new_n4514);
nand_1 g04138(new_n4514, new_n4490, new_n4515);
xnor_1 g04139(new_n4515, new_n4332, new_n4516_1);
nor_1  g04140(new_n2623, new_n382, new_n4517);
nand_1 g04141(new_n4360, new_n4347, new_n4518);
nand_1 g04142(new_n4518, new_n4517, new_n4519);
not_1  g04143(new_n4519, new_n4520);
nor_1  g04144(new_n4518, new_n4517, new_n4521);
nor_1  g04145(new_n4521, new_n4520, new_n4522);
nor_1  g04146(new_n1434, new_n2626, new_n4523);
not_1  g04147(new_n4354, new_n4524);
not_1  g04148(new_n4357, new_n4525);
nor_1  g04149(new_n4525, new_n4351, new_n4526);
nor_1  g04150(new_n4526, new_n4524, new_n4527);
xnor_1 g04151(new_n4527, new_n4523, new_n4528);
not_1  g04152(n2226, new_n4529);
nor_1  g04153(new_n2618, new_n4529, new_n4530);
nand_1 g04154(n3719, n1094, new_n4531);
xnor_1 g04155(new_n4531, new_n4342, new_n4532);
nand_1 g04156(new_n4532, new_n4530, new_n4533);
nor_1  g04157(new_n4532, new_n4530, new_n4534);
not_1  g04158(new_n4534, new_n4535);
nand_1 g04159(new_n4535, new_n4533, new_n4536);
xnor_1 g04160(new_n4536, new_n4528, new_n4537);
xor_1  g04161(new_n4537, new_n4522, new_n4538);
xnor_1 g04162(new_n4538, new_n4371, new_n4539);
nor_1  g04163(new_n385, new_n2895, new_n4540);
nor_1  g04164(new_n1467, new_n2898, new_n4541);
not_1  g04165(n996, new_n4542);
nor_1  g04166(new_n4542, new_n2889, new_n4543);
not_1  g04167(new_n4543, new_n4544);
nand_1 g04168(n5314, n4086, new_n4545);
nand_1 g04169(n8433, n5767, new_n4546);
nand_1 g04170(new_n4546, new_n4545, new_n4547);
not_1  g04171(new_n4547, new_n4548);
nor_1  g04172(new_n4546, new_n4545, new_n4549);
nor_1  g04173(new_n4549, new_n4548, new_n4550);
xnor_1 g04174(new_n4550, new_n4544, new_n4551);
xnor_1 g04175(new_n4551, new_n4541, new_n4552);
nor_1  g04176(new_n1562, new_n2889, new_n4553_1);
nor_1  g04177(new_n4423, new_n4553_1, new_n4554);
nor_1  g04178(new_n4554, new_n4422, new_n4555);
xnor_1 g04179(new_n4555, new_n4552, new_n4556);
nand_1 g04180(new_n4556, new_n4540, new_n4557);
not_1  g04181(new_n4557, new_n4558);
nor_1  g04182(new_n4556, new_n4540, new_n4559);
nor_1  g04183(new_n4559, new_n4558, new_n4560);
nand_1 g04184(new_n4425, new_n4417, new_n4561);
nand_1 g04185(new_n4561, new_n4414, new_n4562);
xnor_1 g04186(new_n4562, new_n4560, new_n4563);
nand_1 g04187(new_n4563, new_n4434, new_n4564);
nor_1  g04188(new_n4563, new_n4434, new_n4565);
not_1  g04189(new_n4565, new_n4566);
nand_1 g04190(new_n4566, new_n4564, new_n4567);
not_1  g04191(new_n4567, new_n4568);
nor_1  g04192(new_n4402, new_n4396, new_n4569);
nor_1  g04193(new_n1533, new_n2767, new_n4570);
nand_1 g04194(n12391, n7610, new_n4571);
nand_1 g04195(new_n4389, new_n4388, new_n4572);
not_1  g04196(new_n4572, new_n4573);
nor_1  g04197(new_n4390, new_n4387, new_n4574);
nor_1  g04198(new_n4574, new_n4573, new_n4575);
xnor_1 g04199(new_n4575, new_n4571, new_n4576);
not_1  g04200(new_n4576, new_n4577);
nor_1  g04201(new_n2761, new_n1538, new_n4578);
nand_1 g04202(n12925, n4828, new_n4579);
xnor_1 g04203(new_n4579, new_n4380, new_n4580);
xnor_1 g04204(new_n4580, new_n4578, new_n4581);
xnor_1 g04205(new_n4581, new_n4577, new_n4582);
nand_1 g04206(new_n4582, new_n4570, new_n4583);
not_1  g04207(new_n4583, new_n4584);
nor_1  g04208(new_n4582, new_n4570, new_n4585);
nor_1  g04209(new_n4585, new_n4584, new_n4586);
nand_1 g04210(new_n4384, new_n4374, new_n4587);
nand_1 g04211(new_n4394, new_n4587, new_n4588);
nand_1 g04212(new_n4588, new_n4586, new_n4589);
not_1  g04213(new_n4589, new_n4590);
nor_1  g04214(new_n4588, new_n4586, new_n4591);
nor_1  g04215(new_n4591, new_n4590, new_n4592);
nand_1 g04216(new_n4592, new_n4569, new_n4593);
not_1  g04217(new_n4593, new_n4594);
nor_1  g04218(new_n4592, new_n4569, new_n4595);
nor_1  g04219(new_n4595, new_n4594, new_n4596);
not_1  g04220(new_n4442, new_n4597);
nand_1 g04221(new_n4465, new_n4597, new_n4598);
nand_1 g04222(new_n4598, new_n4441, new_n4599);
xnor_1 g04223(new_n4599, new_n4596, new_n4600);
xnor_1 g04224(new_n4600, new_n4568, new_n4601);
xnor_1 g04225(new_n4601, new_n4539, new_n4602);
not_1  g04226(new_n4373, new_n4603);
nor_1  g04227(new_n4466, new_n4603, new_n4604);
not_1  g04228(new_n4467, new_n4605);
nor_1  g04229(new_n4487, new_n4605, new_n4606);
nor_1  g04230(new_n4606, new_n4604, new_n4607);
xnor_1 g04231(new_n4607, new_n4602, new_n4608);
xor_1  g04232(new_n4608, new_n4516_1, n992);
nor_1  g04233(new_n1142, new_n378, new_n4610);
not_1  g04234(new_n4610, new_n4611);
nand_1 g04235(n8336, n7946, new_n4612);
not_1  g04236(new_n4612, new_n4613);
nand_1 g04237(n11222, n9763, new_n4614);
not_1  g04238(n2558, new_n4615);
nor_1  g04239(new_n1533, new_n4615, new_n4616);
not_1  g04240(new_n4616, new_n4617);
nor_1  g04241(new_n4617, new_n4614, new_n4618);
not_1  g04242(new_n4618, new_n4619);
nand_1 g04243(new_n4617, new_n4614, new_n4620);
nand_1 g04244(new_n4620, new_n4619, new_n4621);
xnor_1 g04245(new_n4621, new_n4613, new_n4622);
xnor_1 g04246(new_n4622, new_n4611, n1020);
not_1  g04247(new_n2276, new_n4624);
xnor_1 g04248(new_n4624, new_n2275, n1136);
xnor_1 g04249(new_n4513, new_n4512, n1138);
not_1  g04250(n12591, new_n4627);
nor_1  g04251(new_n4627, new_n1592, new_n4628);
not_1  g04252(new_n4628, new_n4629);
nand_1 g04253(n5240, n3932, new_n4630);
nand_1 g04254(n11821, n1798, new_n4631);
xnor_1 g04255(new_n4631, new_n4630, new_n4632);
nor_1  g04256(new_n4632, new_n4629, new_n4633);
not_1  g04257(new_n4633, new_n4634_1);
nand_1 g04258(new_n4632, new_n4629, new_n4635);
nand_1 g04259(new_n4635, new_n4634_1, new_n4636);
nand_1 g04260(n5240, n1798, new_n4637);
nand_1 g04261(n12591, n3172, new_n4638);
nand_1 g04262(new_n4638, new_n4637, new_n4639);
not_1  g04263(new_n4639, new_n4640);
nor_1  g04264(new_n4638, new_n4637, new_n4641);
nor_1  g04265(new_n1592, new_n4053, new_n4642);
nor_1  g04266(new_n4642, new_n4641, new_n4643);
nor_1  g04267(new_n4643, new_n4640, new_n4644);
xnor_1 g04268(new_n4644, new_n4636, new_n4645);
not_1  g04269(new_n4645, new_n4646);
nor_1  g04270(new_n4044, new_n1590, new_n4647);
nand_1 g04271(n11757, n1798, new_n4648);
nand_1 g04272(n12591, n1333, new_n4649);
nand_1 g04273(new_n4649, new_n4648, new_n4650);
not_1  g04274(new_n4650, new_n4651);
nor_1  g04275(new_n4649, new_n4648, new_n4652);
nor_1  g04276(new_n4053, new_n1600, new_n4653);
nor_1  g04277(new_n4653, new_n4652, new_n4654);
nor_1  g04278(new_n4654, new_n4651, new_n4655);
nand_1 g04279(new_n4655, new_n4647, new_n4656);
not_1  g04280(new_n4656, new_n4657);
nor_1  g04281(new_n4655, new_n4647, new_n4658);
nor_1  g04282(new_n4658, new_n4657, new_n4659);
not_1  g04283(new_n4641, new_n4660);
nand_1 g04284(new_n4660, new_n4639, new_n4661);
xnor_1 g04285(new_n4661, new_n4642, new_n4662);
nand_1 g04286(new_n4662, new_n4659, new_n4663);
nand_1 g04287(new_n4663, new_n4656, new_n4664);
not_1  g04288(n11662, new_n4665);
nor_1  g04289(new_n4665, new_n1590, new_n4666);
not_1  g04290(new_n4666, new_n4667);
nor_1  g04291(new_n4044, new_n1600, new_n4668);
not_1  g04292(new_n4668, new_n4669);
nand_1 g04293(new_n4669, new_n4667, new_n4670);
nor_1  g04294(new_n4669, new_n4667, new_n4671);
not_1  g04295(new_n4671, new_n4672);
nand_1 g04296(new_n4672, new_n4670, new_n4673);
xnor_1 g04297(new_n4673, new_n4664, new_n4674);
xnor_1 g04298(new_n4674, new_n4646, new_n4675);
nor_1  g04299(new_n4665, new_n1348, new_n4676);
not_1  g04300(new_n4676, new_n4677);
xnor_1 g04301(new_n4662, new_n4659, new_n4678);
nand_1 g04302(new_n4678, new_n4677, new_n4679);
xnor_1 g04303(new_n4678, new_n4676, new_n4680);
nor_1  g04304(new_n1348, new_n4044, new_n4681);
not_1  g04305(n1798, new_n4682);
nor_1  g04306(new_n1600, new_n4682, new_n4683);
not_1  g04307(new_n4683, new_n4684);
nor_1  g04308(new_n4627, new_n1348, new_n4685);
not_1  g04309(new_n4685, new_n4686_1);
nor_1  g04310(new_n4686_1, new_n4684, new_n4687);
not_1  g04311(new_n4687, new_n4688);
nand_1 g04312(new_n4686_1, new_n4684, new_n4689_1);
nor_1  g04313(new_n4053, new_n1590, new_n4690);
nand_1 g04314(new_n4690, new_n4689_1, new_n4691);
nand_1 g04315(new_n4691, new_n4688, new_n4692);
nand_1 g04316(new_n4692, new_n4681, new_n4693);
not_1  g04317(new_n4693, new_n4694);
xnor_1 g04318(new_n4692, new_n4681, new_n4695);
not_1  g04319(new_n4652, new_n4696);
nand_1 g04320(new_n4696, new_n4650, new_n4697);
xnor_1 g04321(new_n4697, new_n4653, new_n4698);
not_1  g04322(new_n4698, new_n4699);
nor_1  g04323(new_n4699, new_n4695, new_n4700);
nor_1  g04324(new_n4700, new_n4694, new_n4701);
nand_1 g04325(new_n4701, new_n4680, new_n4702);
nand_1 g04326(new_n4702, new_n4679, new_n4703);
not_1  g04327(new_n4703, new_n4704);
nand_1 g04328(new_n4704, new_n4675, new_n4705);
not_1  g04329(new_n4636, new_n4706);
nand_1 g04330(new_n4644, new_n4706, new_n4707);
nand_1 g04331(new_n4707, new_n4634_1, new_n4708);
not_1  g04332(n10327, new_n4709);
nor_1  g04333(new_n4709, new_n1590, new_n4710);
nand_1 g04334(n11662, n3172, new_n4711);
nand_1 g04335(n9583, n7862, new_n4712);
xnor_1 g04336(new_n4712, new_n4711, new_n4713);
xor_1  g04337(new_n4713, new_n4710, new_n4714);
xnor_1 g04338(new_n4714, new_n4708, new_n4715);
nor_1  g04339(new_n4631, new_n4630, new_n4716);
nor_1  g04340(new_n1592, new_n4044, new_n4717);
xor_1  g04341(new_n4717, new_n4716, new_n4718);
nor_1  g04342(new_n1682, new_n4053, new_n4719);
not_1  g04343(n5240, new_n4720);
nor_1  g04344(new_n4627, new_n4720, new_n4721);
not_1  g04345(new_n4721, new_n4722_1);
nor_1  g04346(new_n2334, new_n4682, new_n4723);
not_1  g04347(new_n4723, new_n4724);
nand_1 g04348(new_n4724, new_n4722_1, new_n4725);
nand_1 g04349(new_n4723, new_n4721, new_n4726);
nand_1 g04350(new_n4726, new_n4725, new_n4727);
xnor_1 g04351(new_n4727, new_n4719, new_n4728);
not_1  g04352(new_n4728, new_n4729);
xnor_1 g04353(new_n4729, new_n4718, new_n4730);
xnor_1 g04354(new_n4730, new_n4715, new_n4731);
not_1  g04355(new_n4673, new_n4732);
nand_1 g04356(new_n4732, new_n4664, new_n4733_1);
nand_1 g04357(new_n4674, new_n4645, new_n4734);
xnor_1 g04358(new_n4734, new_n4672, new_n4735);
nand_1 g04359(new_n4735, new_n4733_1, new_n4736);
xnor_1 g04360(new_n4736, new_n4731, new_n4737);
xnor_1 g04361(new_n4737, new_n4705, new_n4738);
nor_1  g04362(new_n4709, new_n1348, new_n4739);
not_1  g04363(new_n4705, new_n4740);
nor_1  g04364(new_n4704, new_n4675, new_n4741);
nor_1  g04365(new_n4741, new_n4740, new_n4742);
nand_1 g04366(new_n4742, new_n4739, new_n4743);
xnor_1 g04367(new_n4698, new_n4695, new_n4744);
not_1  g04368(new_n4689_1, new_n4745);
nor_1  g04369(new_n4745, new_n4687, new_n4746);
nor_1  g04370(new_n4682, new_n1590, new_n4747);
nor_1  g04371(new_n1348, new_n4053, new_n4748);
nand_1 g04372(new_n4748, new_n4747, new_n4749);
nor_1  g04373(new_n4749, new_n4746, new_n4750);
nand_1 g04374(new_n4750, new_n4744, new_n4751);
not_1  g04375(new_n4702, new_n4752);
nor_1  g04376(new_n4701, new_n4680, new_n4753);
nor_1  g04377(new_n4753, new_n4752, new_n4754);
nor_1  g04378(new_n4754, new_n4751, new_n4755);
not_1  g04379(new_n4739, new_n4756);
xnor_1 g04380(new_n4742, new_n4756, new_n4757_1);
nand_1 g04381(new_n4757_1, new_n4755, new_n4758);
nand_1 g04382(new_n4758, new_n4743, new_n4759);
xor_1  g04383(new_n4759, new_n4738, new_n4760);
not_1  g04384(n3022, new_n4761);
nor_1  g04385(new_n1747, new_n4761, new_n4762);
not_1  g04386(new_n4762, new_n4763);
nand_1 g04387(n9640, n4187, new_n4764);
nand_1 g04388(n6703, n4203, new_n4765);
xnor_1 g04389(new_n4765, new_n4764, new_n4766);
xnor_1 g04390(new_n4766, new_n4763, new_n4767);
not_1  g04391(new_n4767, new_n4768);
not_1  g04392(n4187, new_n4769);
nor_1  g04393(new_n4085, new_n4769, new_n4770);
not_1  g04394(new_n4770, new_n4771);
nor_1  g04395(new_n4761, new_n1729, new_n4772);
not_1  g04396(new_n4772, new_n4773);
nand_1 g04397(new_n4773, new_n4771, new_n4774);
not_1  g04398(new_n4774, new_n4775);
nor_1  g04399(new_n4773, new_n4771, new_n4776);
nor_1  g04400(new_n1747, new_n4116, new_n4777);
nor_1  g04401(new_n4777, new_n4776, new_n4778);
nor_1  g04402(new_n4778, new_n4775, new_n4779);
nand_1 g04403(new_n4779, new_n4768, new_n4780);
not_1  g04404(new_n4780, new_n4781);
nor_1  g04405(new_n4779, new_n4768, new_n4782);
nor_1  g04406(new_n4782, new_n4781, new_n4783);
nand_1 g04407(n10451, n9400, new_n4784);
nand_1 g04408(n11023, n2464, new_n4785);
xor_1  g04409(new_n4785, new_n4784, new_n4786);
xnor_1 g04410(new_n4786, new_n4783, new_n4787);
nor_1  g04411(new_n4232, new_n1735, new_n4788);
nor_1  g04412(new_n1747, new_n4085, new_n4789);
not_1  g04413(new_n4789, new_n4790);
nor_1  g04414(new_n1735, new_n4761, new_n4791);
not_1  g04415(new_n4791, new_n4792);
nand_1 g04416(new_n4792, new_n4790, new_n4793);
not_1  g04417(new_n4793, new_n4794);
nor_1  g04418(new_n4792, new_n4790, new_n4795);
nor_1  g04419(new_n4116, new_n1729, new_n4796);
nor_1  g04420(new_n4796, new_n4795, new_n4797);
nor_1  g04421(new_n4797, new_n4794, new_n4798);
nand_1 g04422(new_n4798, new_n4788, new_n4799);
not_1  g04423(new_n4799, new_n4800);
nor_1  g04424(new_n4798, new_n4788, new_n4801);
nor_1  g04425(new_n4801, new_n4800, new_n4802);
not_1  g04426(new_n4802, new_n4803);
not_1  g04427(new_n4776, new_n4804);
nand_1 g04428(new_n4804, new_n4774, new_n4805_1);
xnor_1 g04429(new_n4805_1, new_n4777, new_n4806);
not_1  g04430(new_n4806, new_n4807);
nor_1  g04431(new_n4807, new_n4803, new_n4808);
nor_1  g04432(new_n4808, new_n4800, new_n4809);
nor_1  g04433(new_n4809, new_n4787, new_n4810);
not_1  g04434(new_n4810, new_n4811);
nand_1 g04435(new_n4809, new_n4787, new_n4812);
nand_1 g04436(new_n4812, new_n4811, new_n4813);
not_1  g04437(new_n4813, new_n4814);
not_1  g04438(n10451, new_n4815);
nor_1  g04439(new_n4815, new_n1350, new_n4816);
nor_1  g04440(new_n4806, new_n4802, new_n4817_1);
nor_1  g04441(new_n4817_1, new_n4808, new_n4818);
nand_1 g04442(new_n4818, new_n4816, new_n4819);
nor_1  g04443(new_n4232, new_n1350, new_n4820);
nor_1  g04444(new_n4085, new_n1729, new_n4821);
not_1  g04445(new_n4821, new_n4822);
nor_1  g04446(new_n1350, new_n4761, new_n4823);
not_1  g04447(new_n4823, new_n4824);
nand_1 g04448(new_n4824, new_n4822, new_n4825);
not_1  g04449(new_n4825, new_n4826_1);
nor_1  g04450(new_n4824, new_n4822, new_n4827);
nor_1  g04451(new_n4116, new_n1735, new_n4828_1);
nor_1  g04452(new_n4828_1, new_n4827, new_n4829);
nor_1  g04453(new_n4829, new_n4826_1, new_n4830);
nand_1 g04454(new_n4830, new_n4820, new_n4831);
not_1  g04455(new_n4831, new_n4832);
nor_1  g04456(new_n4830, new_n4820, new_n4833);
nor_1  g04457(new_n4833, new_n4832, new_n4834);
not_1  g04458(new_n4834, new_n4835);
not_1  g04459(new_n4795, new_n4836);
nand_1 g04460(new_n4836, new_n4793, new_n4837);
xnor_1 g04461(new_n4837, new_n4796, new_n4838);
not_1  g04462(new_n4838, new_n4839);
nor_1  g04463(new_n4839, new_n4835, new_n4840);
nor_1  g04464(new_n4840, new_n4832, new_n4841);
not_1  g04465(new_n4841, new_n4842);
not_1  g04466(new_n4819, new_n4843);
nor_1  g04467(new_n4818, new_n4816, new_n4844);
nor_1  g04468(new_n4844, new_n4843, new_n4845);
nand_1 g04469(new_n4845, new_n4842, new_n4846);
nand_1 g04470(new_n4846, new_n4819, new_n4847);
nand_1 g04471(new_n4847, new_n4814, new_n4848);
nor_1  g04472(new_n4766, new_n4763, new_n4849);
nor_1  g04473(new_n4781, new_n4849, new_n4850);
not_1  g04474(new_n4850, new_n4851);
not_1  g04475(n10278, new_n4852);
nor_1  g04476(new_n4852, new_n1735, new_n4853);
nor_1  g04477(new_n4815, new_n1729, new_n4854);
nand_1 g04478(n11423, n6877, new_n4855);
not_1  g04479(new_n4855, new_n4856);
nand_1 g04480(new_n4856, new_n4854, new_n4857);
not_1  g04481(new_n4854, new_n4858);
nand_1 g04482(new_n4855, new_n4858, new_n4859);
nand_1 g04483(new_n4859, new_n4857, new_n4860);
xor_1  g04484(new_n4860, new_n4853, new_n4861);
xnor_1 g04485(new_n4861, new_n4851, new_n4862);
not_1  g04486(new_n4862, new_n4863);
nor_1  g04487(new_n4765, new_n4764, new_n4864);
nor_1  g04488(new_n1747, new_n4232, new_n4865);
xor_1  g04489(new_n4865, new_n4864, new_n4866);
not_1  g04490(new_n4866, new_n4867);
nor_1  g04491(new_n4116, new_n2119, new_n4868);
nor_1  g04492(new_n4769, new_n4761, new_n4869);
not_1  g04493(new_n4869, new_n4870);
nor_1  g04494(new_n2450, new_n4085, new_n4871);
not_1  g04495(new_n4871, new_n4872);
nand_1 g04496(new_n4872, new_n4870, new_n4873);
nand_1 g04497(new_n4871, new_n4869, new_n4874);
nand_1 g04498(new_n4874, new_n4873, new_n4875);
xor_1  g04499(new_n4875, new_n4868, new_n4876);
xnor_1 g04500(new_n4876, new_n4867, new_n4877);
xnor_1 g04501(new_n4877, new_n4863, new_n4878);
nand_1 g04502(new_n4786, new_n4783, new_n4879);
nor_1  g04503(new_n4785, new_n4784, new_n4880);
xnor_1 g04504(new_n4810, new_n4880, new_n4881);
nand_1 g04505(new_n4881, new_n4879, new_n4882);
xnor_1 g04506(new_n4882, new_n4878, new_n4883);
xnor_1 g04507(new_n4883, new_n4848, new_n4884);
nor_1  g04508(new_n4852, new_n1350, new_n4885);
not_1  g04509(new_n4848, new_n4886);
nor_1  g04510(new_n4847, new_n4814, new_n4887);
nor_1  g04511(new_n4887, new_n4886, new_n4888);
nand_1 g04512(new_n4888, new_n4885, new_n4889);
nor_1  g04513(new_n4838, new_n4834, new_n4890);
nor_1  g04514(new_n4890, new_n4840, new_n4891);
not_1  g04515(new_n4891, new_n4892);
not_1  g04516(new_n4828_1, new_n4893);
nor_1  g04517(new_n1350, new_n4085, new_n4894);
nor_1  g04518(new_n4894, new_n4893, new_n4895);
nor_1  g04519(new_n4827, new_n4826_1, new_n4896);
nor_1  g04520(new_n4896, new_n4895, new_n4897);
nand_1 g04521(new_n4897, new_n4828_1, new_n4898);
nor_1  g04522(new_n4898, new_n4892, new_n4899);
xnor_1 g04523(new_n4845, new_n4841, new_n4900);
nand_1 g04524(new_n4900, new_n4899, new_n4901);
not_1  g04525(new_n4901, new_n4902);
not_1  g04526(new_n4885, new_n4903_1);
xnor_1 g04527(new_n4888, new_n4903_1, new_n4904);
nand_1 g04528(new_n4904, new_n4902, new_n4905);
nand_1 g04529(new_n4905, new_n4889, new_n4906);
xnor_1 g04530(new_n4906, new_n4884, new_n4907);
not_1  g04531(n12826, new_n4908);
nor_1  g04532(new_n4908, new_n1925, new_n4909);
nor_1  g04533(new_n4132, new_n1959, new_n4910);
nand_1 g04534(n6294, n1067, new_n4911);
nand_1 g04535(n6797, n5645, new_n4912);
xnor_1 g04536(new_n4912, new_n4911, new_n4913);
xnor_1 g04537(new_n4913, new_n4910, new_n4914);
nand_1 g04538(n6294, n5645, new_n4915);
nand_1 g04539(n8665, n5283, new_n4916);
nand_1 g04540(new_n4916, new_n4915, new_n4917);
not_1  g04541(new_n4917, new_n4918);
not_1  g04542(n1067, new_n4919);
nor_1  g04543(new_n4919, new_n1959, new_n4920);
xnor_1 g04544(new_n4916, new_n4915, new_n4921_1);
nor_1  g04545(new_n4921_1, new_n4920, new_n4922);
nor_1  g04546(new_n4922, new_n4918, new_n4923);
nand_1 g04547(new_n4923, new_n4914, new_n4924);
not_1  g04548(new_n4924, new_n4925);
nor_1  g04549(new_n4923, new_n4914, new_n4926);
nor_1  g04550(new_n4926, new_n4925, new_n4927);
nand_1 g04551(n11922, n11478, new_n4928_1);
not_1  g04552(new_n4928_1, new_n4929);
nand_1 g04553(n5283, n1067, new_n4930);
nand_1 g04554(n11478, n8665, new_n4931);
nand_1 g04555(new_n4931, new_n4930, new_n4932);
not_1  g04556(new_n4932, new_n4933);
nor_1  g04557(new_n4195, new_n1959, new_n4934);
xnor_1 g04558(new_n4931, new_n4930, new_n4935);
nor_1  g04559(new_n4935, new_n4934, new_n4936);
nor_1  g04560(new_n4936, new_n4933, new_n4937);
nand_1 g04561(new_n4937, new_n4929, new_n4938_1);
xnor_1 g04562(new_n4921_1, new_n4920, new_n4939);
xnor_1 g04563(new_n4937, new_n4928_1, new_n4940);
nand_1 g04564(new_n4940, new_n4939, new_n4941);
nand_1 g04565(new_n4941, new_n4938_1, new_n4942);
nand_1 g04566(n11478, n2551, new_n4943);
nand_1 g04567(n11922, n5283, new_n4944);
nand_1 g04568(new_n4944, new_n4943, new_n4945);
nor_1  g04569(new_n4944, new_n4943, new_n4946);
not_1  g04570(new_n4946, new_n4947);
nand_1 g04571(new_n4947, new_n4945, new_n4948);
xnor_1 g04572(new_n4948, new_n4942, new_n4949);
xnor_1 g04573(new_n4949, new_n4927, new_n4950);
not_1  g04574(n2551, new_n4951);
nor_1  g04575(new_n1925, new_n4951, new_n4952);
nand_1 g04576(n11922, n4805, new_n4953);
not_1  g04577(new_n4953, new_n4954);
nand_1 g04578(n5645, n5283, new_n4955);
not_1  g04579(new_n4955, new_n4956);
nand_1 g04580(n8665, n4805, new_n4957);
not_1  g04581(new_n4957, new_n4958);
nand_1 g04582(new_n4958, new_n4956, new_n4959);
nand_1 g04583(new_n4957, new_n4955, new_n4960);
nor_1  g04584(new_n1931, new_n4919, new_n4961);
nand_1 g04585(new_n4961, new_n4960, new_n4962);
nand_1 g04586(new_n4962, new_n4959, new_n4963);
nand_1 g04587(new_n4963, new_n4954, new_n4964);
xnor_1 g04588(new_n4963, new_n4953, new_n4965);
xnor_1 g04589(new_n4935, new_n4934, new_n4966);
nand_1 g04590(new_n4966, new_n4965, new_n4967);
nand_1 g04591(new_n4967, new_n4964, new_n4968);
nor_1  g04592(new_n4968, new_n4952, new_n4969);
not_1  g04593(new_n4939, new_n4970_1);
xnor_1 g04594(new_n4940, new_n4970_1, new_n4971_1);
not_1  g04595(new_n4969, new_n4972);
nand_1 g04596(new_n4968, new_n4952, new_n4973);
nand_1 g04597(new_n4973, new_n4972, new_n4974);
nor_1  g04598(new_n4974, new_n4971_1, new_n4975);
nor_1  g04599(new_n4975, new_n4969, new_n4976);
xnor_1 g04600(new_n4976, new_n4950, new_n4977);
nand_1 g04601(new_n4977, new_n4909, new_n4978);
not_1  g04602(new_n4967, new_n4979);
nor_1  g04603(new_n4966, new_n4965, new_n4980);
nor_1  g04604(new_n4980, new_n4979, new_n4981);
nand_1 g04605(new_n4960, new_n4959, new_n4982);
nand_1 g04606(n4805, n1067, new_n4983);
nand_1 g04607(n11478, n5645, new_n4984);
nor_1  g04608(new_n4984, new_n4983, new_n4985);
and_1  g04609(new_n4985, new_n4982, new_n4986);
nand_1 g04610(new_n4986, new_n4981, new_n4987);
not_1  g04611(new_n4974, new_n4988);
xnor_1 g04612(new_n4988, new_n4971_1, new_n4989);
nor_1  g04613(new_n4989, new_n4987, new_n4990);
not_1  g04614(new_n4909, new_n4991);
xnor_1 g04615(new_n4977, new_n4991, new_n4992);
nand_1 g04616(new_n4992, new_n4990, new_n4993);
nand_1 g04617(new_n4993, new_n4978, new_n4994);
not_1  g04618(new_n4976, new_n4995);
nor_1  g04619(new_n4995, new_n4950, new_n4996);
nor_1  g04620(new_n4908, new_n1931, new_n4997);
nor_1  g04621(new_n1923, new_n4951, new_n4998);
nand_1 g04622(n4805, n4094, new_n4999);
xnor_1 g04623(new_n4999, new_n4998, new_n5000);
xnor_1 g04624(new_n5000, new_n4997, new_n5001);
not_1  g04625(new_n4910, new_n5002);
nor_1  g04626(new_n4913, new_n5002, new_n5003);
not_1  g04627(new_n5003, new_n5004);
nand_1 g04628(new_n4924, new_n5004, new_n5005);
xnor_1 g04629(new_n5005, new_n5001, new_n5006);
nor_1  g04630(new_n4912, new_n4911, new_n5007);
nor_1  g04631(new_n4187_1, new_n1959, new_n5008);
xor_1  g04632(new_n5008, new_n5007, new_n5009);
nor_1  g04633(new_n2205, new_n4919, new_n5010);
nand_1 g04634(n8665, n6294, new_n5011);
nand_1 g04635(n5645, n3146, new_n5012);
xnor_1 g04636(new_n5012, new_n5011, new_n5013);
xnor_1 g04637(new_n5013, new_n5010, new_n5014);
not_1  g04638(new_n5014, new_n5015);
xnor_1 g04639(new_n5015, new_n5009, new_n5016);
xnor_1 g04640(new_n5016, new_n5006, new_n5017);
not_1  g04641(new_n4948, new_n5018);
nand_1 g04642(new_n5018, new_n4942, new_n5019);
nand_1 g04643(new_n4949, new_n4927, new_n5020);
xnor_1 g04644(new_n5020, new_n4947, new_n5021);
nand_1 g04645(new_n5021, new_n5019, new_n5022);
xnor_1 g04646(new_n5022, new_n5017, new_n5023);
xnor_1 g04647(new_n5023, new_n4996, new_n5024);
xnor_1 g04648(new_n5024, new_n4994, new_n5025);
nand_1 g04649(n3992, n2749, new_n5026);
not_1  g04650(new_n5026, new_n5027);
nand_1 g04651(n11876, n6358, new_n5028);
nand_1 g04652(n3992, n3754, new_n5029);
nand_1 g04653(new_n5029, new_n5028, new_n5030_1);
not_1  g04654(new_n5030_1, new_n5031);
nor_1  g04655(new_n4143, new_n1837, new_n5032);
xnor_1 g04656(new_n5029, new_n5028, new_n5033);
nor_1  g04657(new_n5033, new_n5032, new_n5034_1);
nor_1  g04658(new_n5034_1, new_n5031, new_n5035);
nand_1 g04659(new_n5035, new_n5027, new_n5036);
xnor_1 g04660(new_n5035, new_n5026, new_n5037);
nor_1  g04661(new_n4143, new_n1866, new_n5038);
nand_1 g04662(n11876, n5198, new_n5039);
nand_1 g04663(n8384, n3754, new_n5040);
xnor_1 g04664(new_n5040, new_n5039, new_n5041);
xnor_1 g04665(new_n5041, new_n5038, new_n5042);
nand_1 g04666(new_n5042, new_n5037, new_n5043);
nand_1 g04667(new_n5043, new_n5036, new_n5044);
nand_1 g04668(n8384, n2749, new_n5045);
nand_1 g04669(n3992, n159, new_n5046);
nand_1 g04670(new_n5046, new_n5045, new_n5047);
nor_1  g04671(new_n5046, new_n5045, new_n5048);
not_1  g04672(new_n5048, new_n5049);
nand_1 g04673(new_n5049, new_n5047, new_n5050);
xnor_1 g04674(new_n5050, new_n5044, new_n5051);
not_1  g04675(n3754, new_n5052);
nor_1  g04676(new_n1866, new_n5052, new_n5053);
not_1  g04677(new_n5053, new_n5054);
nand_1 g04678(n10898, n5198, new_n5055);
nand_1 g04679(n11876, n1471, new_n5056);
xnor_1 g04680(new_n5056, new_n5055, new_n5057);
xnor_1 g04681(new_n5057, new_n5054, new_n5058);
nand_1 g04682(new_n5040, new_n5039, new_n5059);
not_1  g04683(new_n5059, new_n5060);
nor_1  g04684(new_n5041, new_n5038, new_n5061);
nor_1  g04685(new_n5061, new_n5060, new_n5062);
xnor_1 g04686(new_n5062, new_n5058, new_n5063);
xnor_1 g04687(new_n5063, new_n5051, new_n5064);
not_1  g04688(n159, new_n5065);
nor_1  g04689(new_n1833, new_n5065, new_n5066);
nand_1 g04690(n7236, n2749, new_n5067);
not_1  g04691(new_n5067, new_n5068);
nand_1 g04692(n11876, n8384, new_n5069_1);
nand_1 g04693(n7236, n3754, new_n5070);
nand_1 g04694(new_n5070, new_n5069_1, new_n5071);
not_1  g04695(new_n5071, new_n5072);
nand_1 g04696(n11876, n7236, new_n5073);
nor_1  g04697(new_n5073, new_n5040, new_n5074);
nor_1  g04698(new_n4143, new_n1835_1, new_n5075);
nor_1  g04699(new_n5075, new_n5074, new_n5076);
nor_1  g04700(new_n5076, new_n5072, new_n5077);
nand_1 g04701(new_n5077, new_n5068, new_n5078);
xnor_1 g04702(new_n5077, new_n5067, new_n5079);
xnor_1 g04703(new_n5033, new_n5032, new_n5080);
nand_1 g04704(new_n5080, new_n5079, new_n5081);
nand_1 g04705(new_n5081, new_n5078, new_n5082);
nor_1  g04706(new_n5082, new_n5066, new_n5083);
not_1  g04707(new_n5037, new_n5084);
xnor_1 g04708(new_n5042, new_n5084, new_n5085);
not_1  g04709(new_n5083, new_n5086);
nand_1 g04710(new_n5082, new_n5066, new_n5087);
nand_1 g04711(new_n5087, new_n5086, new_n5088);
nor_1  g04712(new_n5088, new_n5085, new_n5089);
nor_1  g04713(new_n5089, new_n5083, new_n5090);
not_1  g04714(new_n5090, new_n5091);
nor_1  g04715(new_n5091, new_n5064, new_n5092);
nor_1  g04716(new_n5056, new_n5055, new_n5093);
nor_1  g04717(new_n1866, new_n4204, new_n5094_1);
xor_1  g04718(new_n5094_1, new_n5093, new_n5095);
nor_1  g04719(new_n4143, new_n2154, new_n5096);
nand_1 g04720(n5198, n3754, new_n5097);
nand_1 g04721(n11876, n7646, new_n5098);
xnor_1 g04722(new_n5098, new_n5097, new_n5099);
xnor_1 g04723(new_n5099, new_n5096, new_n5100);
not_1  g04724(new_n5100, new_n5101);
xnor_1 g04725(new_n5101, new_n5095, new_n5102);
nand_1 g04726(new_n5057, new_n5054, new_n5103);
not_1  g04727(new_n5103, new_n5104);
nor_1  g04728(new_n5062, new_n5058, new_n5105_1);
nor_1  g04729(new_n5105_1, new_n5104, new_n5106);
not_1  g04730(n1510, new_n5107);
nor_1  g04731(new_n1835_1, new_n5107, new_n5108);
nand_1 g04732(n8384, n159, new_n5109);
nand_1 g04733(n12247, n7236, new_n5110);
xnor_1 g04734(new_n5110, new_n5109, new_n5111);
nor_1  g04735(new_n5111, new_n5108, new_n5112);
and_1  g04736(new_n5111, new_n5108, new_n5113);
nor_1  g04737(new_n5113, new_n5112, new_n5114);
xnor_1 g04738(new_n5114, new_n5106, new_n5115);
xnor_1 g04739(new_n5115, new_n5102, new_n5116);
not_1  g04740(new_n5050, new_n5117);
nand_1 g04741(new_n5117, new_n5044, new_n5118);
nand_1 g04742(new_n5063, new_n5051, new_n5119);
xnor_1 g04743(new_n5119, new_n5049, new_n5120);
nand_1 g04744(new_n5120, new_n5118, new_n5121);
xnor_1 g04745(new_n5121, new_n5116, new_n5122);
xnor_1 g04746(new_n5122, new_n5092, new_n5123);
nor_1  g04747(new_n1833, new_n5107, new_n5124);
xnor_1 g04748(new_n5090, new_n5064, new_n5125);
nand_1 g04749(new_n5125, new_n5124, new_n5126);
xnor_1 g04750(new_n5080, new_n5079, new_n5127);
nor_1  g04751(new_n5074, new_n5072, new_n5128);
not_1  g04752(new_n5128, new_n5129);
nand_1 g04753(n11876, n3992, new_n5130);
nand_1 g04754(n10898, n7236, new_n5131);
nor_1  g04755(new_n5131, new_n5130, new_n5132_1);
nand_1 g04756(new_n5132_1, new_n5129, new_n5133);
nor_1  g04757(new_n5133, new_n5127, new_n5134);
not_1  g04758(new_n5134, new_n5135);
not_1  g04759(new_n5085, new_n5136);
xnor_1 g04760(new_n5088, new_n5136, new_n5137);
nor_1  g04761(new_n5137, new_n5135, new_n5138);
not_1  g04762(new_n5124, new_n5139);
xnor_1 g04763(new_n5125, new_n5139, new_n5140);
nand_1 g04764(new_n5140, new_n5138, new_n5141);
nand_1 g04765(new_n5141, new_n5126, new_n5142);
xnor_1 g04766(new_n5142, new_n5123, new_n5143);
xnor_1 g04767(new_n5143, new_n5025, new_n5144);
xnor_1 g04768(new_n4992, new_n4990, new_n5145);
not_1  g04769(new_n5138, new_n5146);
xnor_1 g04770(new_n5140, new_n5146, new_n5147);
not_1  g04771(new_n5147, new_n5148);
nand_1 g04772(new_n5148, new_n5145, new_n5149);
xnor_1 g04773(new_n5147, new_n5145, new_n5150);
nand_1 g04774(new_n5137, new_n5135, new_n5151);
nand_1 g04775(new_n5151, new_n5146, new_n5152);
not_1  g04776(new_n5152, new_n5153_1);
xnor_1 g04777(new_n4986, new_n4981, new_n5154);
not_1  g04778(new_n5133, new_n5155);
xnor_1 g04779(new_n5155, new_n5127, new_n5156);
not_1  g04780(new_n5156, new_n5157);
nand_1 g04781(new_n5157, new_n5154, new_n5158);
not_1  g04782(new_n5158, new_n5159);
xnor_1 g04783(new_n5131, new_n5130, new_n5160);
xnor_1 g04784(new_n4984, new_n4983, new_n5161);
nand_1 g04785(new_n5161, new_n5160, new_n5162);
not_1  g04786(new_n5162, new_n5163);
nand_1 g04787(n5645, n4805, new_n5164);
nor_1  g04788(new_n5164, new_n5073, new_n5165);
xnor_1 g04789(new_n5161, new_n5160, new_n5166);
nor_1  g04790(new_n5166, new_n5165, new_n5167);
nor_1  g04791(new_n5167, new_n5163, new_n5168);
nand_1 g04792(new_n5164, new_n4961, new_n5169);
nor_1  g04793(new_n5169, new_n4960, new_n5170);
not_1  g04794(new_n5170, new_n5171);
not_1  g04795(new_n5169, new_n5172);
nor_1  g04796(new_n5172, new_n4982, new_n5173);
not_1  g04797(new_n5173, new_n5174);
nand_1 g04798(new_n5174, new_n5171, new_n5175);
nor_1  g04799(new_n5175, new_n5168, new_n5176);
not_1  g04800(new_n5176, new_n5177);
nand_1 g04801(new_n5175, new_n5168, new_n5178);
nand_1 g04802(new_n5178, new_n5177, new_n5179);
not_1  g04803(new_n5179, new_n5180);
nand_1 g04804(new_n5075, new_n5073, new_n5181);
not_1  g04805(new_n5181, new_n5182);
nor_1  g04806(new_n5182, new_n5128, new_n5183);
nor_1  g04807(new_n5181, new_n5072, new_n5184);
nor_1  g04808(new_n5184, new_n5183, new_n5185);
not_1  g04809(new_n5185, new_n5186);
nand_1 g04810(new_n5186, new_n5180, new_n5187);
nand_1 g04811(new_n5187, new_n5177, new_n5188);
not_1  g04812(new_n5188, new_n5189);
xnor_1 g04813(new_n5157, new_n5154, new_n5190);
nor_1  g04814(new_n5190, new_n5189, new_n5191_1);
nor_1  g04815(new_n5191_1, new_n5159, new_n5192);
nor_1  g04816(new_n5192, new_n5153_1, new_n5193);
xnor_1 g04817(new_n4989, new_n4987, new_n5194);
not_1  g04818(new_n5194, new_n5195);
not_1  g04819(new_n5192, new_n5196);
nand_1 g04820(new_n5196, new_n5152, new_n5197);
nand_1 g04821(new_n5192, new_n5153_1, new_n5198_1);
nand_1 g04822(new_n5198_1, new_n5197, new_n5199);
nor_1  g04823(new_n5199, new_n5195, new_n5200);
nor_1  g04824(new_n5200, new_n5193, new_n5201);
not_1  g04825(new_n5201, new_n5202);
nand_1 g04826(new_n5202, new_n5150, new_n5203);
nand_1 g04827(new_n5203, new_n5149, new_n5204);
xnor_1 g04828(new_n5204, new_n5144, new_n5205);
xnor_1 g04829(new_n5205, new_n4907, new_n5206);
xnor_1 g04830(new_n4904, new_n4902, new_n5207);
xnor_1 g04831(new_n5201, new_n5150, new_n5208);
nand_1 g04832(new_n5208, new_n5207, new_n5209);
xnor_1 g04833(new_n4900, new_n4899, new_n5210);
xnor_1 g04834(new_n4898, new_n4891, new_n5211);
xnor_1 g04835(new_n5190, new_n5189, new_n5212_1);
nand_1 g04836(new_n5212_1, new_n5211, new_n5213);
not_1  g04837(new_n5213, new_n5214);
nor_1  g04838(new_n5212_1, new_n5211, new_n5215);
nor_1  g04839(new_n5215, new_n5214, new_n5216);
nand_1 g04840(new_n5185, new_n5179, new_n5217);
nand_1 g04841(new_n5217, new_n5187, new_n5218);
and_1  g04842(new_n4895, new_n4825, new_n5219);
nor_1  g04843(new_n5219, new_n4897, new_n5220);
nand_1 g04844(new_n5220, new_n5218, new_n5221);
not_1  g04845(new_n5221, new_n5222);
nor_1  g04846(new_n5220, new_n5218, new_n5223);
nor_1  g04847(new_n5223, new_n5222, new_n5224);
xnor_1 g04848(new_n5166, new_n5165, new_n5225);
nand_1 g04849(n9400, n6703, new_n5226);
nand_1 g04850(n9640, n6877, new_n5227);
xnor_1 g04851(new_n5227, new_n5226, new_n5228);
not_1  g04852(new_n5228, new_n5229);
nand_1 g04853(new_n5229, new_n5225, new_n5230);
not_1  g04854(new_n4894, new_n5231);
xnor_1 g04855(new_n5164, new_n5073, new_n5232);
nor_1  g04856(new_n5232, new_n5231, new_n5233);
xnor_1 g04857(new_n5228, new_n5225, new_n5234);
nand_1 g04858(new_n5234, new_n5233, new_n5235);
nand_1 g04859(new_n5235, new_n5230, new_n5236);
nand_1 g04860(new_n5236, new_n5224, new_n5237);
nand_1 g04861(new_n5237, new_n5221, new_n5238);
nand_1 g04862(new_n5238, new_n5216, new_n5239);
nand_1 g04863(new_n5239, new_n5213, new_n5240_1);
not_1  g04864(new_n5240_1, new_n5241);
nand_1 g04865(new_n5241, new_n5210, new_n5242);
xnor_1 g04866(new_n5199, new_n5194, new_n5243);
xnor_1 g04867(new_n5240_1, new_n5210, new_n5244);
nand_1 g04868(new_n5244, new_n5243, new_n5245);
nand_1 g04869(new_n5245, new_n5242, new_n5246);
xnor_1 g04870(new_n4904, new_n4901, new_n5247);
xnor_1 g04871(new_n5208, new_n5247, new_n5248);
nand_1 g04872(new_n5248, new_n5246, new_n5249);
nand_1 g04873(new_n5249, new_n5209, new_n5250);
xnor_1 g04874(new_n5250, new_n5206, new_n5251);
not_1  g04875(new_n5251, new_n5252);
nand_1 g04876(new_n5252, new_n4760, new_n5253);
xnor_1 g04877(new_n5251, new_n4760, new_n5254);
xor_1  g04878(new_n4757_1, new_n4755, new_n5255);
xnor_1 g04879(new_n5208, new_n5207, new_n5256);
xnor_1 g04880(new_n5256, new_n5246, new_n5257_1);
not_1  g04881(new_n5257_1, new_n5258);
nand_1 g04882(new_n5258, new_n5255, new_n5259);
xnor_1 g04883(new_n4754, new_n4751, new_n5260);
not_1  g04884(new_n5260, new_n5261);
xnor_1 g04885(new_n5244, new_n5243, new_n5262);
nor_1  g04886(new_n5262, new_n5261, new_n5263);
xnor_1 g04887(new_n5262, new_n5261, new_n5264);
xor_1  g04888(new_n4750, new_n4744, new_n5265);
not_1  g04889(new_n5239, new_n5266);
nor_1  g04890(new_n5238, new_n5216, new_n5267);
nor_1  g04891(new_n5267, new_n5266, new_n5268);
nor_1  g04892(new_n5268, new_n5265, new_n5269);
not_1  g04893(new_n5237, new_n5270);
nor_1  g04894(new_n5236, new_n5224, new_n5271);
nor_1  g04895(new_n5271, new_n5270, new_n5272);
nor_1  g04896(new_n1348, new_n4682, new_n5273);
not_1  g04897(new_n5273, new_n5274);
nand_1 g04898(new_n5274, new_n4690, new_n5275);
not_1  g04899(new_n5275, new_n5276);
nor_1  g04900(new_n5276, new_n4746, new_n5277);
nor_1  g04901(new_n5275, new_n4745, new_n5278);
nor_1  g04902(new_n5278, new_n5277, new_n5279);
nor_1  g04903(new_n5279, new_n5272, new_n5280);
xnor_1 g04904(new_n5279, new_n5272, new_n5281);
xnor_1 g04905(new_n5232, new_n4894, new_n5282);
nand_1 g04906(new_n5282, new_n5273, new_n5283_1);
not_1  g04907(new_n4747, new_n5284);
xnor_1 g04908(new_n4748, new_n5284, new_n5285);
not_1  g04909(new_n5285, new_n5286);
nand_1 g04910(new_n5286, new_n5283_1, new_n5287);
not_1  g04911(new_n5287, new_n5288);
xor_1  g04912(new_n5234, new_n5233, new_n5289);
nor_1  g04913(new_n5286, new_n5283_1, new_n5290);
nor_1  g04914(new_n5290, new_n5288, new_n5291);
not_1  g04915(new_n5291, new_n5292);
nor_1  g04916(new_n5292, new_n5289, new_n5293);
nor_1  g04917(new_n5293, new_n5288, new_n5294);
nor_1  g04918(new_n5294, new_n5281, new_n5295);
nor_1  g04919(new_n5295, new_n5280, new_n5296);
xnor_1 g04920(new_n5268, new_n5265, new_n5297);
nor_1  g04921(new_n5297, new_n5296, new_n5298);
nor_1  g04922(new_n5298, new_n5269, new_n5299);
nor_1  g04923(new_n5299, new_n5264, new_n5300);
nor_1  g04924(new_n5300, new_n5263, new_n5301);
xnor_1 g04925(new_n5257_1, new_n5255, new_n5302);
nand_1 g04926(new_n5302, new_n5301, new_n5303);
nand_1 g04927(new_n5303, new_n5259, new_n5304);
nand_1 g04928(new_n5304, new_n5254, new_n5305_1);
nand_1 g04929(new_n5305_1, new_n5253, new_n5306);
nand_1 g04930(new_n4883, new_n4886, new_n5307);
nand_1 g04931(new_n4906, new_n4884, new_n5308);
nand_1 g04932(new_n5308, new_n5307, new_n5309);
nand_1 g04933(n7862, n753, new_n5310);
not_1  g04934(new_n5005, new_n5311);
nand_1 g04935(new_n5311, new_n5001, new_n5312);
not_1  g04936(new_n5016, new_n5313);
nand_1 g04937(new_n5313, new_n5006, new_n5314_1);
nand_1 g04938(new_n5314_1, new_n5312, new_n5315);
xor_1  g04939(new_n5315, new_n5310, new_n5316);
nand_1 g04940(new_n5008, new_n5007, new_n5317);
nand_1 g04941(new_n5014, new_n5009, new_n5318);
nand_1 g04942(new_n5318, new_n5317, new_n5319_1);
nand_1 g04943(n3146, n1067, new_n5320_1);
nand_1 g04944(n2551, n137, new_n5321);
xnor_1 g04945(new_n5321, new_n5320_1, new_n5322);
nand_1 g04946(n12826, n5283, new_n5323);
nand_1 g04947(n8665, n6797, new_n5324);
xnor_1 g04948(new_n5324, new_n5323, new_n5325);
xnor_1 g04949(new_n5325, new_n5322, new_n5326);
xnor_1 g04950(new_n5326, new_n5319_1, new_n5327);
nand_1 g04951(new_n5094_1, new_n5093, new_n5328);
nand_1 g04952(new_n5100, new_n5095, new_n5329);
nand_1 g04953(new_n5329, new_n5328, new_n5330);
nand_1 g04954(new_n5110, new_n5109, new_n5331_1);
not_1  g04955(new_n5331_1, new_n5332);
nor_1  g04956(new_n5112, new_n5332, new_n5333);
nand_1 g04957(n8384, n1510, new_n5334);
nor_1  g04958(new_n4006, new_n4204, new_n5335);
xnor_1 g04959(new_n5335, new_n5334, new_n5336);
xnor_1 g04960(new_n5336, new_n5333, new_n5337);
xnor_1 g04961(new_n5337, new_n5330, new_n5338);
xnor_1 g04962(new_n5338, new_n5327, new_n5339);
xnor_1 g04963(new_n5339, new_n5316, new_n5340);
xnor_1 g04964(new_n5340, new_n5309, new_n5341);
nor_1  g04965(new_n4734, new_n4672, new_n5342);
not_1  g04966(new_n4736, new_n5343);
nor_1  g04967(new_n5343, new_n4731, new_n5344);
nor_1  g04968(new_n5344, new_n5342, new_n5345);
not_1  g04969(new_n5020, new_n5346);
nand_1 g04970(new_n5346, new_n4946, new_n5347);
not_1  g04971(new_n5017, new_n5348);
nand_1 g04972(new_n5022, new_n5348, new_n5349);
nand_1 g04973(new_n5349, new_n5347, new_n5350);
xnor_1 g04974(new_n5350, new_n5345, new_n5351);
nand_1 g04975(n12511, n7236, new_n5352);
nand_1 g04976(n6826, n1798, new_n5353);
xor_1  g04977(new_n5353, new_n5352, new_n5354);
nand_1 g04978(new_n5012, new_n5011, new_n5355);
not_1  g04979(new_n5355, new_n5356);
nor_1  g04980(new_n5013, new_n5010, new_n5357);
nor_1  g04981(new_n5357, new_n5356, new_n5358);
nand_1 g04982(new_n5098, new_n5097, new_n5359);
not_1  g04983(new_n5359, new_n5360);
nor_1  g04984(new_n5099, new_n5096, new_n5361);
nor_1  g04985(new_n5361, new_n5360, new_n5362);
xnor_1 g04986(new_n5362, new_n5358, new_n5363);
xnor_1 g04987(new_n5363, new_n5354, new_n5364);
nor_1  g04988(new_n1866, new_n5065, new_n5365);
not_1  g04989(new_n4998, new_n5366);
not_1  g04990(new_n5000, new_n5367);
nor_1  g04991(new_n5367, new_n4997, new_n5368);
nor_1  g04992(new_n5368, new_n5366, new_n5369);
and_1  g04993(n11478, n4094, new_n5370);
nand_1 g04994(new_n5370, new_n5369, new_n5371);
not_1  g04995(new_n5369, new_n5372);
nand_1 g04996(new_n5370, new_n4991, new_n5373);
nand_1 g04997(new_n5373, new_n5372, new_n5374);
nand_1 g04998(new_n5374, new_n5371, new_n5375);
xnor_1 g04999(new_n5375, new_n5365, new_n5376);
xnor_1 g05000(new_n5376, new_n5364, new_n5377);
xnor_1 g05001(new_n5377, new_n5351, new_n5378);
xnor_1 g05002(new_n5378, new_n5341, new_n5379);
or_1   g05003(new_n5119, new_n5049, new_n5380);
not_1  g05004(new_n5116, new_n5381);
nand_1 g05005(new_n5121, new_n5381, new_n5382);
nand_1 g05006(new_n5382, new_n5380, new_n5383);
nand_1 g05007(n5645, n4938, new_n5384);
nand_1 g05008(n10898, n7646, new_n5385);
xnor_1 g05009(new_n5385, new_n5384, new_n5386);
xnor_1 g05010(new_n5386, new_n5383, new_n5387);
xnor_1 g05011(new_n5387, new_n5379, new_n5388);
not_1  g05012(new_n5025, new_n5389);
not_1  g05013(new_n5143, new_n5390);
nand_1 g05014(new_n5390, new_n5389, new_n5391);
not_1  g05015(new_n5144, new_n5392);
nand_1 g05016(new_n5204, new_n5392, new_n5393);
nand_1 g05017(new_n5393, new_n5391, new_n5394);
nand_1 g05018(n11922, n6294, new_n5395);
nand_1 g05019(new_n5023, new_n4996, new_n5396);
not_1  g05020(new_n5024, new_n5397);
nand_1 g05021(new_n5397, new_n4994, new_n5398);
nand_1 g05022(new_n5398, new_n5396, new_n5399);
xnor_1 g05023(new_n5399, new_n5395, new_n5400);
nand_1 g05024(new_n4737, new_n4740, new_n5401);
nand_1 g05025(new_n4759, new_n4738, new_n5402);
nand_1 g05026(new_n5402, new_n5401, new_n5403);
nand_1 g05027(new_n4810, new_n4880, new_n5404);
not_1  g05028(new_n4878, new_n5405);
nand_1 g05029(new_n4882, new_n5405, new_n5406);
nand_1 g05030(new_n5406, new_n5404, new_n5407);
nand_1 g05031(new_n4861, new_n4850, new_n5408);
nand_1 g05032(new_n4877, new_n4862, new_n5409);
nand_1 g05033(new_n5409, new_n5408, new_n5410);
nand_1 g05034(new_n4873, new_n4868, new_n5411_1);
nand_1 g05035(new_n5411_1, new_n4874, new_n5412);
nand_1 g05036(n4203, n3022, new_n5413);
nor_1  g05037(new_n4232, new_n4769, new_n5414);
xnor_1 g05038(new_n5414, new_n5413, new_n5415);
xnor_1 g05039(new_n5415, new_n5412, new_n5416);
nand_1 g05040(n7456, n5240, new_n5417);
nand_1 g05041(n12753, n9640, new_n5418);
xnor_1 g05042(new_n5418, new_n5417, new_n5419);
nand_1 g05043(n9583, n1333, new_n5420);
nand_1 g05044(n12591, n11821, new_n5421);
xnor_1 g05045(new_n5421, new_n5420, new_n5422);
xnor_1 g05046(new_n5422, new_n5419, new_n5423);
xnor_1 g05047(new_n5423, new_n5416, new_n5424);
xnor_1 g05048(new_n5424, new_n5410, new_n5425);
not_1  g05049(new_n4708, new_n5426);
nand_1 g05050(new_n4714, new_n5426, new_n5427);
not_1  g05051(new_n4730, new_n5428);
nand_1 g05052(new_n5428, new_n4715, new_n5429);
nand_1 g05053(new_n5429, new_n5427, new_n5430);
nand_1 g05054(n9080, n3932, new_n5431);
nand_1 g05055(n10174, n6703, new_n5432);
nand_1 g05056(n6877, n2278, new_n5433);
xnor_1 g05057(new_n5433, new_n5432, new_n5434);
xnor_1 g05058(new_n5434, new_n5431, new_n5435_1);
xnor_1 g05059(new_n5435_1, new_n5430, new_n5436);
xnor_1 g05060(new_n5436, new_n5425, new_n5437);
xnor_1 g05061(new_n5437, new_n5407, new_n5438);
xnor_1 g05062(new_n5438, new_n5403, new_n5439);
xnor_1 g05063(new_n5439, new_n5400, new_n5440);
xnor_1 g05064(new_n5440, new_n5394, new_n5441);
xnor_1 g05065(new_n5441, new_n5388, new_n5442);
xnor_1 g05066(new_n5442, new_n5306, new_n5443);
not_1  g05067(new_n5106, new_n5444);
nand_1 g05068(new_n5114, new_n5444, new_n5445);
not_1  g05069(new_n5102, new_n5446);
nand_1 g05070(new_n5115, new_n5446, new_n5447);
nand_1 g05071(new_n5447, new_n5445, new_n5448);
nand_1 g05072(new_n4717, new_n4716, new_n5449);
nand_1 g05073(new_n4728, new_n4718, new_n5450);
nand_1 g05074(new_n5450, new_n5449, new_n5451);
nand_1 g05075(new_n4859, new_n4853, new_n5452);
nand_1 g05076(new_n5452, new_n4857, new_n5453);
xnor_1 g05077(new_n5453, new_n5451, new_n5454);
nand_1 g05078(new_n4712, new_n4711, new_n5455);
not_1  g05079(new_n5455, new_n5456);
nor_1  g05080(new_n4713, new_n4710, new_n5457);
nor_1  g05081(new_n5457, new_n5456, new_n5458);
nand_1 g05082(new_n4725, new_n4719, new_n5459);
nand_1 g05083(new_n5459, new_n4726, new_n5460);
nand_1 g05084(n10278, n2464, new_n5461);
nand_1 g05085(n11757, n11662, new_n5462);
xnor_1 g05086(new_n5462, new_n5461, new_n5463);
nand_1 g05087(n10327, n3172, new_n5464);
nand_1 g05088(n11423, n9400, new_n5465);
xnor_1 g05089(new_n5465, new_n5464, new_n5466);
xnor_1 g05090(new_n5466, new_n5463, new_n5467);
xnor_1 g05091(new_n5467, new_n5460, new_n5468);
xnor_1 g05092(new_n5468, new_n5458, new_n5469);
xnor_1 g05093(new_n5469, new_n5454, new_n5470);
xnor_1 g05094(new_n5470, new_n5448, new_n5471);
nand_1 g05095(n3754, n1471, new_n5472);
nand_1 g05096(n11311, n10451, new_n5473);
xnor_1 g05097(new_n5473, new_n5472, new_n5474);
nand_1 g05098(new_n4865, new_n4864, new_n5475);
or_1   g05099(new_n4876, new_n4867, new_n5476);
nand_1 g05100(new_n5476, new_n5475, new_n5477);
nand_1 g05101(n11876, n4722, new_n5478);
nand_1 g05102(n10685, n4805, new_n5479);
nand_1 g05103(n12247, n3992, new_n5480);
xnor_1 g05104(new_n5480, new_n5479, new_n5481);
xnor_1 g05105(new_n5481, new_n5478, new_n5482);
xnor_1 g05106(new_n5482, new_n5477, new_n5483);
xnor_1 g05107(new_n5483, new_n5474, new_n5484);
xnor_1 g05108(new_n5484, new_n5471, new_n5485);
nand_1 g05109(new_n5122, new_n5092, new_n5486);
not_1  g05110(new_n5123, new_n5487);
nand_1 g05111(new_n5142, new_n5487, new_n5488);
and_1  g05112(new_n5488, new_n5486, new_n5489);
nand_1 g05113(new_n5205, new_n4907, new_n5490);
not_1  g05114(new_n5206, new_n5491);
nand_1 g05115(new_n5250, new_n5491, new_n5492);
nand_1 g05116(new_n5492, new_n5490, new_n5493);
xnor_1 g05117(new_n5493, new_n5489, new_n5494);
xnor_1 g05118(new_n5494, new_n5485, new_n5495);
xnor_1 g05119(new_n5495, new_n5443, n1269);
nor_1  g05120(new_n1139, new_n395, new_n5497);
nand_1 g05121(n12705, n7265, new_n5498);
nor_1  g05122(new_n395, new_n1130, new_n5499);
xnor_1 g05123(new_n5498, new_n1128, new_n5500);
nor_1  g05124(new_n5500, new_n5499, new_n5501);
nor_1  g05125(new_n5501, new_n5498, new_n5502);
nor_1  g05126(new_n5502, new_n5497, new_n5503);
not_1  g05127(new_n5497, new_n5504);
nor_1  g05128(new_n5502, new_n1138_1, new_n5505);
nor_1  g05129(new_n5505, new_n5504, new_n5506);
nor_1  g05130(new_n5506, new_n5503, new_n5507);
nand_1 g05131(n12025, n7265, new_n5508);
nand_1 g05132(n12705, n2879, new_n5509);
xnor_1 g05133(new_n5509, new_n5508, new_n5510);
not_1  g05134(new_n5510, new_n5511);
nor_1  g05135(new_n5511, new_n5507, new_n5512);
nand_1 g05136(new_n5511, new_n5507, new_n5513);
not_1  g05137(new_n5513, new_n5514);
nor_1  g05138(new_n5514, new_n5512, new_n5515);
not_1  g05139(n9195, new_n5516);
nor_1  g05140(new_n5516, new_n424, new_n5517);
not_1  g05141(new_n5517, new_n5518);
nor_1  g05142(new_n1121, new_n419, new_n5519);
not_1  g05143(new_n5519, new_n5520);
nand_1 g05144(new_n5520, new_n5518, new_n5521);
nor_1  g05145(new_n5520, new_n5518, new_n5522);
not_1  g05146(new_n5522, new_n5523);
nand_1 g05147(new_n5523, new_n5521, new_n5524);
xnor_1 g05148(new_n5524, new_n5515, new_n5525);
nor_1  g05149(new_n424, new_n1121, new_n5526);
not_1  g05150(new_n1145, new_n5527);
nor_1  g05151(new_n1146, new_n1138_1, new_n5528);
nor_1  g05152(new_n5528, new_n5527, new_n5529);
nand_1 g05153(new_n5529, new_n5526, new_n5530);
xnor_1 g05154(new_n5500, new_n5499, new_n5531);
not_1  g05155(new_n5530, new_n5532);
nor_1  g05156(new_n5529, new_n5526, new_n5533);
nor_1  g05157(new_n5533, new_n5532, new_n5534);
nand_1 g05158(new_n5534, new_n5531, new_n5535);
nand_1 g05159(new_n5535, new_n5530, new_n5536);
xnor_1 g05160(new_n5536, new_n5525, new_n5537);
not_1  g05161(new_n5537, new_n5538);
nor_1  g05162(new_n5516, new_n456, new_n5539);
nand_1 g05163(new_n1150, new_n1134, new_n5540);
nor_1  g05164(new_n5540, new_n5539, new_n5541);
xnor_1 g05165(new_n5534, new_n5531, new_n5542);
not_1  g05166(new_n5542, new_n5543);
xnor_1 g05167(new_n5540, new_n5539, new_n5544);
nor_1  g05168(new_n5544, new_n5543, new_n5545);
nor_1  g05169(new_n5545, new_n5541, new_n5546);
nand_1 g05170(new_n5546, new_n5538, new_n5547);
nor_1  g05171(new_n5514, new_n5506, new_n5548);
not_1  g05172(new_n5548, new_n5549);
not_1  g05173(n2253, new_n5550);
nor_1  g05174(new_n424, new_n5550, new_n5551);
nand_1 g05175(n9195, n1097, new_n5552);
nand_1 g05176(n5305, n3865, new_n5553);
xnor_1 g05177(new_n5553, new_n5552, new_n5554);
xor_1  g05178(new_n5554, new_n5551, new_n5555);
xnor_1 g05179(new_n5555, new_n5549, new_n5556);
nor_1  g05180(new_n5509, new_n5508, new_n5557);
nor_1  g05181(new_n1121, new_n395, new_n5558);
xor_1  g05182(new_n5558, new_n5557, new_n5559);
nor_1  g05183(new_n511, new_n1130, new_n5560);
nand_1 g05184(n11257, n7265, new_n5561);
nand_1 g05185(n12705, n10223, new_n5562);
xnor_1 g05186(new_n5562, new_n5561, new_n5563);
xor_1  g05187(new_n5563, new_n5560, new_n5564);
xnor_1 g05188(new_n5564, new_n5559, new_n5565);
xnor_1 g05189(new_n5565, new_n5556, new_n5566);
not_1  g05190(new_n5524, new_n5567);
nand_1 g05191(new_n5567, new_n5515, new_n5568);
nand_1 g05192(new_n5536, new_n5525, new_n5569);
not_1  g05193(new_n5569, new_n5570);
nand_1 g05194(new_n5570, new_n5522, new_n5571);
nand_1 g05195(new_n5569, new_n5523, new_n5572);
nand_1 g05196(new_n5572, new_n5571, new_n5573);
nand_1 g05197(new_n5573, new_n5568, new_n5574);
xnor_1 g05198(new_n5574, new_n5566, new_n5575);
xnor_1 g05199(new_n5575, new_n5547, new_n5576);
nor_1  g05200(new_n456, new_n5550, new_n5577);
not_1  g05201(new_n5547, new_n5578);
nor_1  g05202(new_n5546, new_n5538, new_n5579_1);
nor_1  g05203(new_n5579_1, new_n5578, new_n5580);
nand_1 g05204(new_n5580, new_n5577, new_n5581);
nand_1 g05205(new_n1160, new_n1153, new_n5582);
xnor_1 g05206(new_n5544, new_n5542, new_n5583);
nor_1  g05207(new_n5583, new_n5582, new_n5584);
not_1  g05208(new_n5577, new_n5585);
xnor_1 g05209(new_n5580, new_n5585, new_n5586);
nand_1 g05210(new_n5586, new_n5584, new_n5587);
nand_1 g05211(new_n5587, new_n5581, new_n5588);
xnor_1 g05212(new_n5588, new_n5576, new_n5589);
not_1  g05213(new_n5589, new_n5590);
xnor_1 g05214(new_n5586, new_n5584, new_n5591);
not_1  g05215(n12145, new_n5592);
nor_1  g05216(new_n5592, new_n552, new_n5593);
nand_1 g05217(new_n1295, new_n1282, new_n5594);
nand_1 g05218(new_n5594, new_n5593, new_n5595);
not_1  g05219(new_n5595, new_n5596);
nor_1  g05220(new_n5594, new_n5593, new_n5597);
nor_1  g05221(new_n5597, new_n5596, new_n5598);
nor_1  g05222(new_n563, new_n1278, new_n5599);
not_1  g05223(new_n5599, new_n5600);
nor_1  g05224(new_n1292, new_n1286, new_n5601);
nor_1  g05225(new_n5601, new_n1291, new_n5602);
xnor_1 g05226(new_n5602, new_n5600, new_n5603);
nor_1  g05227(new_n599, new_n1192, new_n5604);
nand_1 g05228(n12299, n9189, new_n5605);
nand_1 g05229(n8276, n7946, new_n5606);
not_1  g05230(new_n5606, new_n5607);
xnor_1 g05231(new_n5607, new_n5605, new_n5608);
xnor_1 g05232(new_n5608, new_n5604, new_n5609);
xnor_1 g05233(new_n5609, new_n5603, new_n5610);
xnor_1 g05234(new_n5610, new_n5598, new_n5611);
not_1  g05235(new_n5611, new_n5612);
nand_1 g05236(new_n5612, new_n1303, new_n5613);
not_1  g05237(new_n5613, new_n5614);
not_1  g05238(n12221, new_n5615);
nor_1  g05239(new_n5615, new_n552, new_n5616);
not_1  g05240(new_n5616, new_n5617);
nand_1 g05241(new_n5602, new_n5599, new_n5618);
not_1  g05242(new_n5609, new_n5619);
nand_1 g05243(new_n5619, new_n5603, new_n5620);
nand_1 g05244(new_n5620, new_n5618, new_n5621);
nor_1  g05245(new_n5592, new_n563, new_n5622);
not_1  g05246(new_n5622, new_n5623);
nor_1  g05247(new_n554, new_n1278, new_n5624);
not_1  g05248(new_n5624, new_n5625);
nand_1 g05249(new_n5625, new_n5623, new_n5626);
nor_1  g05250(new_n5625, new_n5623, new_n5627);
not_1  g05251(new_n5627, new_n5628);
nand_1 g05252(new_n5628, new_n5626, new_n5629);
xnor_1 g05253(new_n5629, new_n5621, new_n5630);
nor_1  g05254(new_n1199_1, new_n599, new_n5631);
not_1  g05255(new_n5608, new_n5632);
nor_1  g05256(new_n5632, new_n5604, new_n5633);
nor_1  g05257(new_n5633, new_n5606, new_n5634);
nor_1  g05258(new_n5634, new_n5631, new_n5635);
not_1  g05259(new_n5631, new_n5636);
nor_1  g05260(new_n5634, new_n1286, new_n5637);
nor_1  g05261(new_n5637, new_n5636, new_n5638);
nor_1  g05262(new_n5638, new_n5635, new_n5639);
nand_1 g05263(n8276, n2024, new_n5640);
nand_1 g05264(n9241, n7946, new_n5641_1);
xor_1  g05265(new_n5641_1, new_n5640, new_n5642);
nor_1  g05266(new_n5642, new_n5639, new_n5643);
nand_1 g05267(new_n5642, new_n5639, new_n5644);
not_1  g05268(new_n5644, new_n5645_1);
nor_1  g05269(new_n5645_1, new_n5643, new_n5646);
xnor_1 g05270(new_n5646, new_n5630, new_n5647);
nand_1 g05271(new_n5610, new_n5598, new_n5648);
nand_1 g05272(new_n5648, new_n5595, new_n5649);
xnor_1 g05273(new_n5649, new_n5647, new_n5650);
xnor_1 g05274(new_n5650, new_n5617, new_n5651);
xnor_1 g05275(new_n5651, new_n5614, new_n5652);
not_1  g05276(new_n5652, new_n5653);
xnor_1 g05277(new_n5612, new_n1303, new_n5654);
not_1  g05278(new_n5654, new_n5655);
nand_1 g05279(new_n1323, new_n1322, new_n5656);
not_1  g05280(new_n5656, new_n5657);
not_1  g05281(n6016, new_n5658);
nor_1  g05282(new_n5658, new_n668, new_n5659);
not_1  g05283(new_n5659, new_n5660);
nor_1  g05284(new_n712, new_n1310, new_n5661);
nand_1 g05285(new_n1318, new_n1317, new_n5662);
not_1  g05286(new_n5662, new_n5663);
nor_1  g05287(new_n1319, new_n1315, new_n5664);
nor_1  g05288(new_n5664, new_n5663, new_n5665);
xnor_1 g05289(new_n5665, new_n5661, new_n5666);
nor_1  g05290(new_n829, new_n1235, new_n5667);
not_1  g05291(n10545, new_n5668);
nor_1  g05292(new_n5668, new_n4615, new_n5669);
not_1  g05293(new_n5669, new_n5670_1);
nand_1 g05294(new_n5670_1, new_n1246, new_n5671);
nand_1 g05295(new_n5669, new_n1245, new_n5672);
nand_1 g05296(new_n5672, new_n5671, new_n5673);
xnor_1 g05297(new_n5673, new_n5667, new_n5674);
xnor_1 g05298(new_n5674, new_n5666, new_n5675);
xnor_1 g05299(new_n5675, new_n5660, new_n5676);
nand_1 g05300(new_n1313, new_n1311, new_n5677);
not_1  g05301(new_n5677, new_n5678);
nor_1  g05302(new_n1320, new_n1314, new_n5679);
nor_1  g05303(new_n5679, new_n5678, new_n5680);
xnor_1 g05304(new_n5680, new_n5676, new_n5681);
xnor_1 g05305(new_n5681, new_n5657, new_n5682);
nor_1  g05306(new_n1337, new_n1336, new_n5683);
not_1  g05307(new_n5683, new_n5684);
not_1  g05308(n7270, new_n5685);
nor_1  g05309(new_n754, new_n5685, new_n5686);
not_1  g05310(new_n5686, new_n5687);
nor_1  g05311(new_n696, new_n1325, new_n5688);
nand_1 g05312(new_n1333_1, new_n1332, new_n5689);
not_1  g05313(new_n5689, new_n5690);
nor_1  g05314(new_n1334, new_n1330, new_n5691);
nor_1  g05315(new_n5691, new_n5690, new_n5692);
xnor_1 g05316(new_n5692, new_n5688, new_n5693_1);
nor_1  g05317(new_n1215, new_n767, new_n5694_1);
not_1  g05318(new_n1220, new_n5695);
not_1  g05319(n9763, new_n5696);
nor_1  g05320(new_n5696, new_n802, new_n5697);
not_1  g05321(new_n5697, new_n5698);
nand_1 g05322(new_n5698, new_n5695, new_n5699);
nand_1 g05323(new_n5697, new_n1220, new_n5700);
nand_1 g05324(new_n5700, new_n5699, new_n5701);
xnor_1 g05325(new_n5701, new_n5694_1, new_n5702);
xnor_1 g05326(new_n5702, new_n5693_1, new_n5703);
xnor_1 g05327(new_n5703, new_n5687, new_n5704);
nand_1 g05328(new_n1328, new_n1326, new_n5705);
not_1  g05329(new_n5705, new_n5706);
nor_1  g05330(new_n1335, new_n1329, new_n5707);
nor_1  g05331(new_n5707, new_n5706, new_n5708);
xnor_1 g05332(new_n5708, new_n5704, new_n5709);
xnor_1 g05333(new_n5709, new_n5684, new_n5710);
xnor_1 g05334(new_n5710, new_n5682, new_n5711);
not_1  g05335(new_n1339, new_n5712);
nand_1 g05336(new_n5712, new_n1324, new_n5713);
nand_1 g05337(new_n1344, new_n1340, new_n5714);
nand_1 g05338(new_n5714, new_n5713, new_n5715);
xnor_1 g05339(new_n5715, new_n5711, new_n5716);
nand_1 g05340(new_n5716, new_n5655, new_n5717);
not_1  g05341(new_n1308, new_n5718);
nand_1 g05342(new_n5718, new_n1304, new_n5719);
nand_1 g05343(new_n1345, new_n1309, new_n5720);
nand_1 g05344(new_n5720, new_n5719, new_n5721);
xnor_1 g05345(new_n5716, new_n5654, new_n5722);
nand_1 g05346(new_n5722, new_n5721, new_n5723);
nand_1 g05347(new_n5723, new_n5717, new_n5724);
xnor_1 g05348(new_n5724, new_n5653, new_n5725);
nand_1 g05349(new_n5681, new_n5657, new_n5726);
not_1  g05350(n5798, new_n5727);
nor_1  g05351(new_n5727, new_n668, new_n5728);
not_1  g05352(new_n5728, new_n5729);
nor_1  g05353(new_n829, new_n1244, new_n5730);
not_1  g05354(new_n5730, new_n5731);
nand_1 g05355(n10545, n2498, new_n5732);
nand_1 g05356(n7690, n2558, new_n5733);
nand_1 g05357(new_n5733, new_n5732, new_n5734);
nor_1  g05358(new_n5733, new_n5732, new_n5735);
not_1  g05359(new_n5735, new_n5736);
nand_1 g05360(new_n5736, new_n5734, new_n5737);
nor_1  g05361(new_n5737, new_n5731, new_n5738);
not_1  g05362(new_n5738, new_n5739);
nand_1 g05363(new_n5737, new_n5731, new_n5740);
nand_1 g05364(new_n5740, new_n5739, new_n5741);
not_1  g05365(new_n5671, new_n5742);
not_1  g05366(new_n5672, new_n5743);
nor_1  g05367(new_n5743, new_n5667, new_n5744);
nor_1  g05368(new_n5744, new_n5742, new_n5745);
xnor_1 g05369(new_n5745, new_n5741, new_n5746);
nor_1  g05370(new_n712, new_n5658, new_n5747);
not_1  g05371(new_n5747, new_n5748);
nor_1  g05372(new_n740, new_n1310, new_n5749);
not_1  g05373(new_n5749, new_n5750);
nand_1 g05374(new_n5750, new_n5748, new_n5751);
nor_1  g05375(new_n5750, new_n5748, new_n5752);
not_1  g05376(new_n5752, new_n5753);
nand_1 g05377(new_n5753, new_n5751, new_n5754);
xnor_1 g05378(new_n5754, new_n5746, new_n5755);
nand_1 g05379(new_n5665, new_n5661, new_n5756);
not_1  g05380(new_n5666, new_n5757);
nand_1 g05381(new_n5674, new_n5757, new_n5758);
nand_1 g05382(new_n5758, new_n5756, new_n5759);
xnor_1 g05383(new_n5759, new_n5755, new_n5760_1);
not_1  g05384(new_n5760_1, new_n5761);
nand_1 g05385(new_n5675, new_n5659, new_n5762);
not_1  g05386(new_n5680, new_n5763);
nand_1 g05387(new_n5763, new_n5676, new_n5764);
nand_1 g05388(new_n5764, new_n5762, new_n5765);
nand_1 g05389(new_n5765, new_n5761, new_n5766);
not_1  g05390(new_n5766, new_n5767_1);
nor_1  g05391(new_n5765, new_n5761, new_n5768);
nor_1  g05392(new_n5768, new_n5767_1, new_n5769);
xnor_1 g05393(new_n5769, new_n5729, new_n5770);
xnor_1 g05394(new_n5770, new_n5726, new_n5771);
nand_1 g05395(new_n5709, new_n5683, new_n5772);
not_1  g05396(new_n5772, new_n5773);
nand_1 g05397(n7965, n5153, new_n5774);
nand_1 g05398(n3342, n2393, new_n5775);
nand_1 g05399(n9763, n3986, new_n5776);
nand_1 g05400(n9111, n5860, new_n5777);
xnor_1 g05401(new_n5777, new_n5776, new_n5778);
nor_1  g05402(new_n5778, new_n5775, new_n5779);
not_1  g05403(new_n5779, new_n5780);
nand_1 g05404(new_n5778, new_n5775, new_n5781);
nand_1 g05405(new_n5781, new_n5780, new_n5782);
not_1  g05406(new_n5699, new_n5783);
not_1  g05407(new_n5700, new_n5784);
nor_1  g05408(new_n5784, new_n5694_1, new_n5785);
nor_1  g05409(new_n5785, new_n5783, new_n5786);
xnor_1 g05410(new_n5786, new_n5782, new_n5787);
nor_1  g05411(new_n696, new_n5685, new_n5788);
not_1  g05412(new_n5788, new_n5789);
nor_1  g05413(new_n762, new_n1325, new_n5790);
not_1  g05414(new_n5790, new_n5791);
nand_1 g05415(new_n5791, new_n5789, new_n5792);
nor_1  g05416(new_n5791, new_n5789, new_n5793);
not_1  g05417(new_n5793, new_n5794);
nand_1 g05418(new_n5794, new_n5792, new_n5795);
xnor_1 g05419(new_n5795, new_n5787, new_n5796);
nand_1 g05420(new_n5692, new_n5688, new_n5797);
not_1  g05421(new_n5693_1, new_n5798_1);
nand_1 g05422(new_n5702, new_n5798_1, new_n5799);
nand_1 g05423(new_n5799, new_n5797, new_n5800);
xnor_1 g05424(new_n5800, new_n5796, new_n5801);
not_1  g05425(new_n5801, new_n5802);
nand_1 g05426(new_n5703, new_n5686, new_n5803);
not_1  g05427(new_n5708, new_n5804);
nand_1 g05428(new_n5804, new_n5704, new_n5805);
nand_1 g05429(new_n5805, new_n5803, new_n5806);
nand_1 g05430(new_n5806, new_n5802, new_n5807);
not_1  g05431(new_n5807, new_n5808);
nor_1  g05432(new_n5806, new_n5802, new_n5809);
nor_1  g05433(new_n5809, new_n5808, new_n5810);
xnor_1 g05434(new_n5810, new_n5774, new_n5811);
xnor_1 g05435(new_n5811, new_n5773, new_n5812);
xnor_1 g05436(new_n5812, new_n5771, new_n5813);
not_1  g05437(new_n5710, new_n5814_1);
nand_1 g05438(new_n5814_1, new_n5682, new_n5815);
nand_1 g05439(new_n5715, new_n5711, new_n5816);
nand_1 g05440(new_n5816, new_n5815, new_n5817);
xnor_1 g05441(new_n5817, new_n5813, new_n5818);
xnor_1 g05442(new_n5818, new_n5725, new_n5819);
not_1  g05443(new_n5819, new_n5820);
nand_1 g05444(new_n5820, new_n5591, new_n5821);
xnor_1 g05445(new_n5819, new_n5591, new_n5822);
xnor_1 g05446(new_n5583, new_n5582, new_n5823);
not_1  g05447(new_n5722, new_n5824);
xnor_1 g05448(new_n5824, new_n5721, new_n5825);
not_1  g05449(new_n5825, new_n5826);
nand_1 g05450(new_n5826, new_n5823, new_n5827);
and_1  g05451(new_n1276, new_n1161, new_n5828);
nor_1  g05452(new_n1346, new_n1277, new_n5829);
nor_1  g05453(new_n5829, new_n5828, new_n5830);
xnor_1 g05454(new_n5825, new_n5823, new_n5831);
nand_1 g05455(new_n5831, new_n5830, new_n5832);
nand_1 g05456(new_n5832, new_n5827, new_n5833);
nand_1 g05457(new_n5833, new_n5822, new_n5834);
nand_1 g05458(new_n5834, new_n5821, new_n5835);
xnor_1 g05459(new_n5835, new_n5590, new_n5836);
nand_1 g05460(new_n5650, new_n5616, new_n5837);
nand_1 g05461(new_n5651, new_n5614, new_n5838);
nand_1 g05462(new_n5838, new_n5837, new_n5839);
not_1  g05463(new_n5649, new_n5840);
nor_1  g05464(new_n5840, new_n5647, new_n5841);
not_1  g05465(new_n5638, new_n5842);
nand_1 g05466(new_n5644, new_n5842, new_n5843);
nor_1  g05467(new_n5615, new_n563, new_n5844);
nand_1 g05468(n12299, n12145, new_n5845);
nand_1 g05469(n10217, n8759, new_n5846);
xnor_1 g05470(new_n5846, new_n5845, new_n5847);
xor_1  g05471(new_n5847, new_n5844, new_n5848);
xnor_1 g05472(new_n5848, new_n5843, new_n5849);
nor_1  g05473(new_n5641_1, new_n5640, new_n5850);
nor_1  g05474(new_n599, new_n1278, new_n5851);
xor_1  g05475(new_n5851, new_n5850, new_n5852);
nor_1  g05476(new_n2723, new_n1192, new_n5853);
not_1  g05477(new_n5853, new_n5854);
nand_1 g05478(n10510, n7946, new_n5855);
nand_1 g05479(n9189, n8276, new_n5856);
xnor_1 g05480(new_n5856, new_n5855, new_n5857_1);
xnor_1 g05481(new_n5857_1, new_n5854, new_n5858);
xnor_1 g05482(new_n5858, new_n5852, new_n5859);
xnor_1 g05483(new_n5859, new_n5849, new_n5860_1);
not_1  g05484(new_n5860_1, new_n5861);
not_1  g05485(new_n5629, new_n5862);
nand_1 g05486(new_n5862, new_n5621, new_n5863);
nand_1 g05487(new_n5646, new_n5630, new_n5864);
not_1  g05488(new_n5864, new_n5865);
nand_1 g05489(new_n5865, new_n5627, new_n5866);
nand_1 g05490(new_n5864, new_n5628, new_n5867);
nand_1 g05491(new_n5867, new_n5866, new_n5868);
nand_1 g05492(new_n5868, new_n5863, new_n5869);
xnor_1 g05493(new_n5869, new_n5861, new_n5870);
xnor_1 g05494(new_n5870, new_n5841, new_n5871);
xnor_1 g05495(new_n5871, new_n5839, new_n5872);
nand_1 g05496(new_n5724, new_n5653, new_n5873);
not_1  g05497(new_n5725, new_n5874);
nand_1 g05498(new_n5818, new_n5874, new_n5875);
nand_1 g05499(new_n5875, new_n5873, new_n5876);
xnor_1 g05500(new_n5876, new_n5872, new_n5877);
nor_1  g05501(new_n712, new_n5727, new_n5878);
nand_1 g05502(n6016, n2530, new_n5879);
not_1  g05503(n2347, new_n5880);
nor_1  g05504(new_n668, new_n5880, new_n5881);
xnor_1 g05505(new_n5881, new_n5879, new_n5882);
not_1  g05506(new_n5882, new_n5883);
nand_1 g05507(new_n5883, new_n5878, new_n5884);
nor_1  g05508(new_n5883, new_n5878, new_n5885);
not_1  g05509(new_n5885, new_n5886);
nand_1 g05510(new_n5886, new_n5884, new_n5887);
not_1  g05511(new_n5741, new_n5888);
nand_1 g05512(new_n5745, new_n5888, new_n5889);
nand_1 g05513(new_n5889, new_n5739, new_n5890);
nand_1 g05514(new_n5890, new_n5887, new_n5891);
not_1  g05515(new_n5887, new_n5892);
not_1  g05516(new_n5890, new_n5893);
nand_1 g05517(new_n5893, new_n5892, new_n5894);
nand_1 g05518(new_n5894, new_n5891, new_n5895);
not_1  g05519(new_n5895, new_n5896);
nand_1 g05520(n12648, n521, new_n5897);
xnor_1 g05521(new_n5897, new_n5735, new_n5898);
nor_1  g05522(new_n1048, new_n1235, new_n5899);
nand_1 g05523(n10545, n5579, new_n5900);
nand_1 g05524(n3616, n2558, new_n5901);
xnor_1 g05525(new_n5901, new_n5900, new_n5902);
xor_1  g05526(new_n5902, new_n5899, new_n5903);
xnor_1 g05527(new_n5903, new_n5898, new_n5904);
xnor_1 g05528(new_n5904, new_n5896, new_n5905);
not_1  g05529(new_n5754, new_n5906);
nand_1 g05530(new_n5906, new_n5746, new_n5907);
nand_1 g05531(new_n5759, new_n5755, new_n5908);
not_1  g05532(new_n5908, new_n5909);
nand_1 g05533(new_n5909, new_n5752, new_n5910);
nand_1 g05534(new_n5908, new_n5753, new_n5911);
nand_1 g05535(new_n5911, new_n5910, new_n5912);
nand_1 g05536(new_n5912, new_n5907, new_n5913);
xnor_1 g05537(new_n5913, new_n5905, new_n5914);
xnor_1 g05538(new_n5914, new_n5766, new_n5915);
nand_1 g05539(new_n5769, new_n5728, new_n5916);
not_1  g05540(new_n5726, new_n5917);
nand_1 g05541(new_n5770, new_n5917, new_n5918);
nand_1 g05542(new_n5918, new_n5916, new_n5919);
xnor_1 g05543(new_n5919, new_n5915, new_n5920);
not_1  g05544(new_n5782, new_n5921);
nand_1 g05545(new_n5786, new_n5921, new_n5922);
nand_1 g05546(new_n5922, new_n5780, new_n5923);
not_1  g05547(n5153, new_n5924);
nor_1  g05548(new_n696, new_n5924, new_n5925);
nand_1 g05549(n11892, n7270, new_n5926);
nand_1 g05550(n7965, n2507, new_n5927);
xnor_1 g05551(new_n5927, new_n5926, new_n5928);
xnor_1 g05552(new_n5928, new_n5925, new_n5929);
xnor_1 g05553(new_n5929, new_n5923, new_n5930);
not_1  g05554(new_n5930, new_n5931);
nor_1  g05555(new_n5777, new_n5776, new_n5932);
nor_1  g05556(new_n767, new_n1325, new_n5933);
xor_1  g05557(new_n5933, new_n5932, new_n5934_1);
nor_1  g05558(new_n1215, new_n1084, new_n5935);
nand_1 g05559(n5860, n3342, new_n5936);
nand_1 g05560(n9763, n5857, new_n5937);
xnor_1 g05561(new_n5937, new_n5936, new_n5938);
xor_1  g05562(new_n5938, new_n5935, new_n5939);
xnor_1 g05563(new_n5939, new_n5934_1, new_n5940);
not_1  g05564(new_n5940, new_n5941);
nand_1 g05565(new_n5941, new_n5931, new_n5942);
nand_1 g05566(new_n5940, new_n5930, new_n5943);
nand_1 g05567(new_n5943, new_n5942, new_n5944);
not_1  g05568(new_n5795, new_n5945);
nand_1 g05569(new_n5945, new_n5787, new_n5946);
nand_1 g05570(new_n5800, new_n5796, new_n5947);
not_1  g05571(new_n5947, new_n5948);
nand_1 g05572(new_n5948, new_n5793, new_n5949);
nand_1 g05573(new_n5947, new_n5794, new_n5950);
nand_1 g05574(new_n5950, new_n5949, new_n5951);
nand_1 g05575(new_n5951, new_n5946, new_n5952);
xnor_1 g05576(new_n5952, new_n5944, new_n5953);
xnor_1 g05577(new_n5953, new_n5808, new_n5954);
not_1  g05578(new_n5810, new_n5955);
nand_1 g05579(new_n5955, new_n5774, new_n5956);
nand_1 g05580(new_n5811, new_n5772, new_n5957);
nand_1 g05581(new_n5957, new_n5956, new_n5958);
xnor_1 g05582(new_n5958, new_n5954, new_n5959);
xnor_1 g05583(new_n5959, new_n5920, new_n5960);
not_1  g05584(new_n5771, new_n5961);
nand_1 g05585(new_n5812, new_n5961, new_n5962);
nand_1 g05586(new_n5817, new_n5813, new_n5963);
nand_1 g05587(new_n5963, new_n5962, new_n5964_1);
xnor_1 g05588(new_n5964_1, new_n5960, new_n5965);
xnor_1 g05589(new_n5965, new_n5877, new_n5966);
xnor_1 g05590(new_n5966, new_n5836, n1523);
nor_1  g05591(new_n378, new_n1121, new_n5968);
nand_1 g05592(n10223, n4189, new_n5969);
nor_1  g05593(new_n5969, new_n4611, new_n5970);
nand_1 g05594(n10223, n6687, new_n5971);
nand_1 g05595(n7265, n4189, new_n5972);
nand_1 g05596(new_n5972, new_n5971, new_n5973);
not_1  g05597(new_n5973, new_n5974);
nor_1  g05598(new_n1130, new_n1377, new_n5975);
not_1  g05599(new_n5975, new_n5976);
nor_1  g05600(new_n5976, new_n5974, new_n5977);
nor_1  g05601(new_n5977, new_n5970, new_n5978);
xnor_1 g05602(new_n5978, new_n5968, new_n5979);
nor_1  g05603(new_n1367, new_n1130, new_n5980);
nand_1 g05604(n10223, n2564, new_n5981);
nand_1 g05605(n7265, n6770, new_n5982);
xnor_1 g05606(new_n5982, new_n5981, new_n5983);
xnor_1 g05607(new_n5983, new_n5980, new_n5984);
xor_1  g05608(new_n5984, new_n5979, new_n5985);
nor_1  g05609(new_n5974, new_n5970, new_n5986);
not_1  g05610(new_n5986, new_n5987);
nor_1  g05611(new_n1142, new_n1377, new_n5988);
nor_1  g05612(new_n378, new_n1130, new_n5989);
and_1  g05613(new_n5989, new_n5988, new_n5990);
nand_1 g05614(new_n5990, new_n5987, new_n5991);
not_1  g05615(new_n5991, new_n5992);
nand_1 g05616(new_n5992, new_n5985, new_n5993);
not_1  g05617(new_n5993, new_n5994);
nor_1  g05618(new_n5516, new_n378, new_n5995);
nor_1  g05619(new_n1121, new_n1377, new_n5996);
nor_1  g05620(new_n4283, new_n1130, new_n5997);
not_1  g05621(new_n5997, new_n5998);
nand_1 g05622(n9920, n7265, new_n5999);
xnor_1 g05623(new_n5999, new_n5969, new_n6000);
xnor_1 g05624(new_n6000, new_n5998, new_n6001);
xnor_1 g05625(new_n6001, new_n5996, new_n6002);
nand_1 g05626(new_n5982, new_n5981, new_n6003);
not_1  g05627(new_n6003, new_n6004);
nor_1  g05628(new_n5983, new_n5980, new_n6005);
nor_1  g05629(new_n6005, new_n6004, new_n6006);
xor_1  g05630(new_n6006, new_n6002, new_n6007);
nand_1 g05631(new_n6007, new_n5995, new_n6008);
not_1  g05632(new_n6008, new_n6009);
nor_1  g05633(new_n6007, new_n5995, new_n6010);
nor_1  g05634(new_n6010, new_n6009, new_n6011);
not_1  g05635(new_n5968, new_n6012);
nor_1  g05636(new_n5978, new_n6012, new_n6013);
not_1  g05637(new_n6013, new_n6014);
nand_1 g05638(new_n5984, new_n5979, new_n6015);
nand_1 g05639(new_n6015, new_n6014, new_n6016_1);
nand_1 g05640(new_n6016_1, new_n6011, new_n6017);
not_1  g05641(new_n6017, new_n6018);
nor_1  g05642(new_n6016_1, new_n6011, new_n6019);
nor_1  g05643(new_n6019, new_n6018, new_n6020);
nand_1 g05644(new_n6020, new_n5994, new_n6021);
not_1  g05645(new_n6021, new_n6022);
nor_1  g05646(new_n6020, new_n5994, new_n6023);
nor_1  g05647(new_n6023, new_n6022, new_n6024);
nor_1  g05648(new_n382, new_n1278, new_n6025);
nand_1 g05649(n9189, n8336, new_n6026);
nand_1 g05650(n7946, n6986, new_n6027);
nand_1 g05651(new_n6027, new_n6026, new_n6028);
not_1  g05652(new_n6028, new_n6029);
nand_1 g05653(n9189, n6986, new_n6030);
nor_1  g05654(new_n6030, new_n4612, new_n6031);
nor_1  g05655(new_n1434, new_n1192, new_n6032);
nor_1  g05656(new_n6032, new_n6031, new_n6033);
nor_1  g05657(new_n6033, new_n6029, new_n6034);
xnor_1 g05658(new_n6034, new_n6025, new_n6035);
nor_1  g05659(new_n1508, new_n1192, new_n6036);
nor_1  g05660(new_n1434, new_n1199_1, new_n6037);
not_1  g05661(new_n6037, new_n6038_1);
nor_1  g05662(new_n1196, new_n4529, new_n6039);
not_1  g05663(new_n6039, new_n6040);
nand_1 g05664(new_n6040, new_n6038_1, new_n6041);
nor_1  g05665(new_n6040, new_n6038_1, new_n6042);
not_1  g05666(new_n6042, new_n6043);
nand_1 g05667(new_n6043, new_n6041, new_n6044);
xnor_1 g05668(new_n6044, new_n6036, new_n6045);
xnor_1 g05669(new_n6045, new_n6035, new_n6046);
not_1  g05670(new_n6032, new_n6047);
nor_1  g05671(new_n6047, new_n4613, new_n6048);
nor_1  g05672(new_n6031, new_n6029, new_n6049);
nor_1  g05673(new_n6049, new_n6048, new_n6050);
not_1  g05674(new_n6050, new_n6051);
nor_1  g05675(new_n6051, new_n6047, new_n6052);
nand_1 g05676(new_n6052, new_n6046, new_n6053);
nor_1  g05677(new_n5592, new_n382, new_n6054);
nand_1 g05678(n10928, n2522, new_n6055);
not_1  g05679(new_n6055, new_n6056);
not_1  g05680(new_n6041, new_n6057);
nor_1  g05681(new_n6042, new_n6036, new_n6058);
nor_1  g05682(new_n6058, new_n6057, new_n6059);
xnor_1 g05683(new_n6059, new_n6056, new_n6060);
nor_1  g05684(new_n4529, new_n1192, new_n6061);
not_1  g05685(new_n6061, new_n6062);
nand_1 g05686(n7946, n1094, new_n6063);
xnor_1 g05687(new_n6063, new_n6030, new_n6064);
xnor_1 g05688(new_n6064, new_n6062, new_n6065);
not_1  g05689(new_n6065, new_n6066);
xnor_1 g05690(new_n6066, new_n6060, new_n6067);
nand_1 g05691(new_n6067, new_n6054, new_n6068);
not_1  g05692(new_n6068, new_n6069);
nor_1  g05693(new_n6067, new_n6054, new_n6070);
nor_1  g05694(new_n6070, new_n6069, new_n6071);
nand_1 g05695(new_n6034, new_n6025, new_n6072);
not_1  g05696(new_n6035, new_n6073);
nand_1 g05697(new_n6045, new_n6073, new_n6074);
nand_1 g05698(new_n6074, new_n6072, new_n6075);
xnor_1 g05699(new_n6075, new_n6071, new_n6076);
xnor_1 g05700(new_n6076, new_n6053, new_n6077);
xnor_1 g05701(new_n6052, new_n6046, new_n6078);
not_1  g05702(new_n6078, new_n6079);
nor_1  g05703(new_n1533, new_n1310, new_n6080);
nand_1 g05704(n7891, n5579, new_n6081);
not_1  g05705(new_n6081, new_n6082);
nand_1 g05706(new_n6082, new_n4616, new_n6083);
nand_1 g05707(n12069, n5579, new_n6084);
nand_1 g05708(n7891, n2558, new_n6085);
nand_1 g05709(new_n6085, new_n6084, new_n6086);
nor_1  g05710(new_n1452, new_n1235, new_n6087);
nand_1 g05711(new_n6087, new_n6086, new_n6088);
nand_1 g05712(new_n6088, new_n6083, new_n6089_1);
nand_1 g05713(new_n6089_1, new_n6080, new_n6090);
not_1  g05714(new_n6090, new_n6091);
nor_1  g05715(new_n6089_1, new_n6080, new_n6092);
nor_1  g05716(new_n6092, new_n6091, new_n6093);
nor_1  g05717(new_n4386, new_n1235, new_n6094);
nand_1 g05718(n12391, n5579, new_n6095);
nand_1 g05719(n7160, n2558, new_n6096);
nand_1 g05720(new_n6096, new_n6095, new_n6097);
nor_1  g05721(new_n6096, new_n6095, new_n6098);
not_1  g05722(new_n6098, new_n6099);
nand_1 g05723(new_n6099, new_n6097, new_n6100);
xnor_1 g05724(new_n6100, new_n6094, new_n6101);
xnor_1 g05725(new_n6101, new_n6093, new_n6102);
nand_1 g05726(new_n6086, new_n6083, new_n6103);
nand_1 g05727(n12391, n2558, new_n6104);
nand_1 g05728(n12069, n2498, new_n6105);
nor_1  g05729(new_n6105, new_n6104, new_n6106);
nand_1 g05730(new_n6106, new_n6103, new_n6107);
not_1  g05731(new_n6107, new_n6108);
xnor_1 g05732(new_n6108, new_n6102, new_n6109);
nor_1  g05733(new_n385, new_n1325, new_n6110);
nand_1 g05734(n11222, n3342, new_n6111);
nand_1 g05735(n9763, n5314, new_n6112);
nand_1 g05736(new_n6112, new_n6111, new_n6113);
not_1  g05737(new_n6113, new_n6114);
nand_1 g05738(n5314, n3342, new_n6115);
nor_1  g05739(new_n6115, new_n4614, new_n6116);
nor_1  g05740(new_n1467, new_n1215, new_n6117);
nor_1  g05741(new_n6117, new_n6116, new_n6118);
nor_1  g05742(new_n6118, new_n6114, new_n6119);
nand_1 g05743(new_n6119, new_n6110, new_n6120);
not_1  g05744(new_n6120, new_n6121);
nor_1  g05745(new_n6119, new_n6110, new_n6122);
nor_1  g05746(new_n6122, new_n6121, new_n6123);
nor_1  g05747(new_n1215, new_n1562, new_n6124);
nand_1 g05748(n11153, n3342, new_n6125);
nand_1 g05749(n9763, n996, new_n6126_1);
nand_1 g05750(new_n6126_1, new_n6125, new_n6127);
nor_1  g05751(new_n6126_1, new_n6125, new_n6128);
not_1  g05752(new_n6128, new_n6129);
nand_1 g05753(new_n6129, new_n6127, new_n6130);
xnor_1 g05754(new_n6130, new_n6124, new_n6131);
xnor_1 g05755(new_n6131, new_n6123, new_n6132);
not_1  g05756(new_n6116, new_n6133);
nand_1 g05757(new_n6117, new_n4614, new_n6134);
nand_1 g05758(new_n6134, new_n6114, new_n6135);
nand_1 g05759(new_n6135, new_n6133, new_n6136);
nand_1 g05760(new_n6136, new_n6117, new_n6137);
not_1  g05761(new_n6137, new_n6138);
xnor_1 g05762(new_n6138, new_n6132, new_n6139);
nand_1 g05763(new_n6139, new_n6109, new_n6140);
nor_1  g05764(new_n6139, new_n6109, new_n6141);
not_1  g05765(new_n6141, new_n6142);
nand_1 g05766(new_n6142, new_n6140, new_n6143);
nor_1  g05767(new_n6134, new_n6114, new_n6144);
nor_1  g05768(new_n6144, new_n6136, new_n6145);
not_1  g05769(new_n6145, new_n6146);
xnor_1 g05770(new_n6105, new_n6104, new_n6147);
nand_1 g05771(new_n6147, new_n4619, new_n6148);
xnor_1 g05772(new_n6147, new_n4618, new_n6149);
nand_1 g05773(n11153, n9763, new_n6150);
nand_1 g05774(n11222, n9111, new_n6151);
xnor_1 g05775(new_n6151, new_n6150, new_n6152);
nand_1 g05776(new_n6152, new_n6149, new_n6153);
nand_1 g05777(new_n6153, new_n6148, new_n6154);
nand_1 g05778(new_n6154, new_n6146, new_n6155);
xnor_1 g05779(new_n6154, new_n6145, new_n6156);
nand_1 g05780(new_n6087, new_n4617, new_n6157);
nand_1 g05781(new_n6157, new_n6103, new_n6158);
not_1  g05782(new_n6157, new_n6159);
nand_1 g05783(new_n6159, new_n6086, new_n6160);
nand_1 g05784(new_n6160, new_n6158, new_n6161);
nand_1 g05785(new_n6161, new_n6156, new_n6162);
nand_1 g05786(new_n6162, new_n6155, new_n6163);
xnor_1 g05787(new_n6163, new_n6143, new_n6164);
not_1  g05788(new_n6164, new_n6165);
nand_1 g05789(new_n6165, new_n6079, new_n6166);
xnor_1 g05790(new_n6164, new_n6079, new_n6167);
nand_1 g05791(new_n6048, new_n6028, new_n6168);
nand_1 g05792(new_n6168, new_n6051, new_n6169);
not_1  g05793(new_n6161, new_n6170);
xnor_1 g05794(new_n6170, new_n6156, new_n6171);
nor_1  g05795(new_n6171, new_n6169, new_n6172);
not_1  g05796(new_n6172, new_n6173);
not_1  g05797(new_n6169, new_n6174);
xnor_1 g05798(new_n6171, new_n6174, new_n6175);
xnor_1 g05799(new_n6152, new_n6149, new_n6176);
nand_1 g05800(n10928, n7946, new_n6177);
nand_1 g05801(n8336, n2024, new_n6178);
xnor_1 g05802(new_n6178, new_n6177, new_n6179);
not_1  g05803(new_n6179, new_n6180);
nand_1 g05804(new_n6180, new_n6176, new_n6181);
nor_1  g05805(new_n4621, new_n4612, new_n6182);
xnor_1 g05806(new_n6179, new_n6176, new_n6183);
nand_1 g05807(new_n6183, new_n6182, new_n6184);
nand_1 g05808(new_n6184, new_n6181, new_n6185);
nand_1 g05809(new_n6185, new_n6175, new_n6186);
nand_1 g05810(new_n6186, new_n6173, new_n6187);
nand_1 g05811(new_n6187, new_n6167, new_n6188);
nand_1 g05812(new_n6188, new_n6166, new_n6189);
xnor_1 g05813(new_n6189, new_n6077, new_n6190);
nor_1  g05814(new_n6107, new_n6102, new_n6191);
nor_1  g05815(new_n1533, new_n5658, new_n6192_1);
not_1  g05816(new_n6192_1, new_n6193);
nor_1  g05817(new_n1452, new_n1310, new_n6194);
not_1  g05818(new_n6097, new_n6195);
nor_1  g05819(new_n6098, new_n6094, new_n6196);
nor_1  g05820(new_n6196, new_n6195, new_n6197);
nand_1 g05821(new_n6197, new_n6194, new_n6198);
not_1  g05822(new_n6198, new_n6199);
nor_1  g05823(new_n6197, new_n6194, new_n6200);
nor_1  g05824(new_n6200, new_n6199, new_n6201);
nor_1  g05825(new_n1538, new_n1235, new_n6202);
not_1  g05826(new_n6202, new_n6203);
nand_1 g05827(n4828, n2558, new_n6204);
xnor_1 g05828(new_n6204, new_n6081, new_n6205);
xnor_1 g05829(new_n6205, new_n6203, new_n6206);
not_1  g05830(new_n6206, new_n6207);
xnor_1 g05831(new_n6207, new_n6201, new_n6208);
xnor_1 g05832(new_n6208, new_n6193, new_n6209);
nand_1 g05833(new_n6101, new_n6093, new_n6210);
nand_1 g05834(new_n6210, new_n6090, new_n6211);
xnor_1 g05835(new_n6211, new_n6209, new_n6212);
xnor_1 g05836(new_n6212, new_n6191, new_n6213);
not_1  g05837(new_n6213, new_n6214);
nor_1  g05838(new_n6137, new_n6132, new_n6215);
nor_1  g05839(new_n385, new_n5685, new_n6216);
nor_1  g05840(new_n1467, new_n1325, new_n6217);
not_1  g05841(new_n6127, new_n6218);
nor_1  g05842(new_n6128, new_n6124, new_n6219);
nor_1  g05843(new_n6219, new_n6218, new_n6220);
xnor_1 g05844(new_n6220, new_n6217, new_n6221);
nor_1  g05845(new_n1215, new_n4542, new_n6222);
nand_1 g05846(n9763, n5767, new_n6223);
nand_1 g05847(new_n6223, new_n6115, new_n6224);
nor_1  g05848(new_n6223, new_n6115, new_n6225);
not_1  g05849(new_n6225, new_n6226);
nand_1 g05850(new_n6226, new_n6224, new_n6227);
xnor_1 g05851(new_n6227, new_n6222, new_n6228);
xnor_1 g05852(new_n6228, new_n6221, new_n6229);
nand_1 g05853(new_n6229, new_n6216, new_n6230);
not_1  g05854(new_n6230, new_n6231);
nor_1  g05855(new_n6229, new_n6216, new_n6232);
nor_1  g05856(new_n6232, new_n6231, new_n6233);
nand_1 g05857(new_n6131, new_n6123, new_n6234);
nand_1 g05858(new_n6234, new_n6120, new_n6235);
nor_1  g05859(new_n6235, new_n6233, new_n6236);
nand_1 g05860(new_n6235, new_n6233, new_n6237);
not_1  g05861(new_n6237, new_n6238);
nor_1  g05862(new_n6238, new_n6236, new_n6239);
nand_1 g05863(new_n6239, new_n6215, new_n6240);
not_1  g05864(new_n6240, new_n6241);
nor_1  g05865(new_n6239, new_n6215, new_n6242);
nor_1  g05866(new_n6242, new_n6241, new_n6243);
xnor_1 g05867(new_n6243, new_n6214, new_n6244);
not_1  g05868(new_n6143, new_n6245);
nand_1 g05869(new_n6163, new_n6245, new_n6246);
nand_1 g05870(new_n6246, new_n6142, new_n6247);
xnor_1 g05871(new_n6247, new_n6244, new_n6248);
not_1  g05872(new_n6248, new_n6249);
xnor_1 g05873(new_n6249, new_n6190, new_n6250);
xnor_1 g05874(new_n6250, new_n6024, new_n6251);
xnor_1 g05875(new_n5992, new_n5985, new_n6252);
xnor_1 g05876(new_n6187, new_n6167, new_n6253);
nand_1 g05877(new_n6253, new_n6252, new_n6254_1);
xnor_1 g05878(new_n6185, new_n6175, new_n6255);
nor_1  g05879(new_n5976, new_n4610, new_n6256);
nor_1  g05880(new_n6256, new_n5986, new_n6257);
nand_1 g05881(new_n6256, new_n5973, new_n6258);
not_1  g05882(new_n6258, new_n6259);
nor_1  g05883(new_n6259, new_n6257, new_n6260);
not_1  g05884(new_n6260, new_n6261);
nand_1 g05885(new_n6261, new_n6255, new_n6262);
xnor_1 g05886(new_n6260, new_n6255, new_n6263);
nand_1 g05887(new_n4622, new_n4610, new_n6264);
xnor_1 g05888(new_n5989, new_n5988, new_n6265);
nand_1 g05889(new_n6265, new_n6264, new_n6266);
xnor_1 g05890(new_n6183, new_n6182, new_n6267);
xor_1  g05891(new_n6265, new_n6264, new_n6268);
nand_1 g05892(new_n6268, new_n6267, new_n6269);
nand_1 g05893(new_n6269, new_n6266, new_n6270);
nand_1 g05894(new_n6270, new_n6263, new_n6271);
nand_1 g05895(new_n6271, new_n6262, new_n6272);
not_1  g05896(new_n6253, new_n6273_1);
xnor_1 g05897(new_n6273_1, new_n6252, new_n6274);
nand_1 g05898(new_n6274, new_n6272, new_n6275);
nand_1 g05899(new_n6275, new_n6254_1, new_n6276);
xnor_1 g05900(new_n6276, new_n6251, n1658);
nor_1  g05901(new_n1348, new_n1121, new_n6278);
nand_1 g05902(n10223, n7862, new_n6279);
nand_1 g05903(n7265, n3172, new_n6280);
nand_1 g05904(new_n6280, new_n6279, new_n6281);
not_1  g05905(new_n6281, new_n6282);
nor_1  g05906(new_n1348, new_n1142, new_n6283);
not_1  g05907(new_n6283, new_n6284);
nor_1  g05908(new_n1139, new_n1600, new_n6285);
not_1  g05909(new_n6285, new_n6286);
nor_1  g05910(new_n6286, new_n6284, new_n6287);
nor_1  g05911(new_n1130, new_n1590, new_n6288);
nor_1  g05912(new_n6288, new_n6287, new_n6289);
nor_1  g05913(new_n6289, new_n6282, new_n6290);
nand_1 g05914(new_n6290, new_n6278, new_n6291);
not_1  g05915(new_n6291, new_n6292);
nor_1  g05916(new_n6290, new_n6278, new_n6293);
nor_1  g05917(new_n6293, new_n6292, new_n6294_1);
nor_1  g05918(new_n1600, new_n1130, new_n6295);
nand_1 g05919(n10223, n1333, new_n6296);
nand_1 g05920(n11757, n7265, new_n6297);
nand_1 g05921(new_n6297, new_n6296, new_n6298);
nor_1  g05922(new_n6297, new_n6296, new_n6299);
not_1  g05923(new_n6299, new_n6300);
nand_1 g05924(new_n6300, new_n6298, new_n6301);
xnor_1 g05925(new_n6301, new_n6295, new_n6302);
nand_1 g05926(new_n6302, new_n6294_1, new_n6303);
not_1  g05927(new_n6303, new_n6304);
nor_1  g05928(new_n6302, new_n6294_1, new_n6305);
nor_1  g05929(new_n6305, new_n6304, new_n6306);
not_1  g05930(new_n6288, new_n6307);
nor_1  g05931(new_n6307, new_n6283, new_n6308);
nor_1  g05932(new_n6308, new_n6281, new_n6309);
nor_1  g05933(new_n6309, new_n6287, new_n6310);
nor_1  g05934(new_n6310, new_n6307, new_n6311);
xor_1  g05935(new_n6311, new_n6306, new_n6312);
nor_1  g05936(new_n1350, new_n1278, new_n6313);
not_1  g05937(new_n6313, new_n6314);
nor_1  g05938(new_n1729, new_n1192, new_n6315);
nand_1 g05939(n9400, n9189, new_n6316);
nand_1 g05940(n11311, n7946, new_n6317);
xnor_1 g05941(new_n6317, new_n6316, new_n6318);
nand_1 g05942(new_n6318, new_n6315, new_n6319);
nor_1  g05943(new_n6318, new_n6315, new_n6320);
not_1  g05944(new_n6320, new_n6321);
nand_1 g05945(new_n6321, new_n6319, new_n6322);
not_1  g05946(new_n6322, new_n6323);
nor_1  g05947(new_n6323, new_n6314, new_n6324);
nor_1  g05948(new_n6322, new_n6313, new_n6325);
nor_1  g05949(new_n6325, new_n6324, new_n6326);
nand_1 g05950(n9189, n6877, new_n6327);
nand_1 g05951(n7946, n2464, new_n6328);
nand_1 g05952(new_n6328, new_n6327, new_n6329);
not_1  g05953(new_n6329, new_n6330);
nor_1  g05954(new_n1196, new_n1350, new_n6331);
not_1  g05955(new_n6331, new_n6332);
nor_1  g05956(new_n1199_1, new_n1729, new_n6333);
not_1  g05957(new_n6333, new_n6334);
nor_1  g05958(new_n6334, new_n6332, new_n6335);
nor_1  g05959(new_n1735, new_n1192, new_n6336);
nor_1  g05960(new_n6336, new_n6335, new_n6337);
nor_1  g05961(new_n6337, new_n6330, new_n6338);
xnor_1 g05962(new_n6338, new_n6326, new_n6339);
not_1  g05963(new_n6339, new_n6340);
not_1  g05964(new_n6336, new_n6341);
nor_1  g05965(new_n6341, new_n6331, new_n6342);
nor_1  g05966(new_n6335, new_n6330, new_n6343);
nor_1  g05967(new_n6343, new_n6342, new_n6344);
not_1  g05968(new_n6344, new_n6345);
nor_1  g05969(new_n6345, new_n6341, new_n6346);
nor_1  g05970(new_n6346, new_n6340, new_n6347);
nand_1 g05971(new_n6346, new_n6340, new_n6348);
not_1  g05972(new_n6348, new_n6349);
nor_1  g05973(new_n6349, new_n6347, new_n6350);
nand_1 g05974(new_n6342, new_n6329, new_n6351);
nand_1 g05975(new_n6351, new_n6345, new_n6352);
not_1  g05976(new_n6352, new_n6353);
nand_1 g05977(n4805, n2558, new_n6354);
nand_1 g05978(n9763, n7236, new_n6355);
nor_1  g05979(new_n6355, new_n6354, new_n6356);
not_1  g05980(new_n6356, new_n6357);
nand_1 g05981(new_n6355, new_n6354, new_n6358_1);
nand_1 g05982(new_n6358_1, new_n6357, new_n6359_1);
nor_1  g05983(new_n6359_1, new_n6332, new_n6360);
nand_1 g05984(n9400, n7946, new_n6361);
nand_1 g05985(n6877, n2024, new_n6362);
xnor_1 g05986(new_n6362, new_n6361, new_n6363);
not_1  g05987(new_n6363, new_n6364);
nand_1 g05988(new_n6364, new_n6360, new_n6365);
nand_1 g05989(n9111, n7236, new_n6366);
nand_1 g05990(n9763, n3992, new_n6367);
nand_1 g05991(new_n6367, new_n6366, new_n6368);
nor_1  g05992(new_n6367, new_n6366, new_n6369);
not_1  g05993(new_n6369, new_n6370);
nand_1 g05994(new_n6370, new_n6368, new_n6371);
xnor_1 g05995(new_n6371, new_n6356, new_n6372);
nand_1 g05996(n4805, n2498, new_n6373);
nand_1 g05997(n11478, n2558, new_n6374);
xnor_1 g05998(new_n6374, new_n6373, new_n6375);
xnor_1 g05999(new_n6375, new_n6372, new_n6376);
xnor_1 g06000(new_n6363, new_n6360, new_n6377);
nand_1 g06001(new_n6377, new_n6376, new_n6378);
nand_1 g06002(new_n6378, new_n6365, new_n6379);
nor_1  g06003(new_n6379, new_n6353, new_n6380);
not_1  g06004(new_n6380, new_n6381);
nand_1 g06005(new_n6371, new_n6357, new_n6382);
nand_1 g06006(new_n6375, new_n6372, new_n6383);
nand_1 g06007(new_n6383, new_n6382, new_n6384);
nor_1  g06008(new_n1931, new_n1235, new_n6385);
nand_1 g06009(new_n6385, new_n6354, new_n6386);
not_1  g06010(new_n6386, new_n6387);
nand_1 g06011(n5283, n2558, new_n6388);
nand_1 g06012(n5579, n4805, new_n6389);
nand_1 g06013(new_n6389, new_n6388, new_n6390);
not_1  g06014(new_n6390, new_n6391);
nor_1  g06015(new_n6389, new_n6388, new_n6392);
nor_1  g06016(new_n6392, new_n6391, new_n6393);
nor_1  g06017(new_n6393, new_n6387, new_n6394);
nor_1  g06018(new_n6391, new_n6386, new_n6395);
nor_1  g06019(new_n6395, new_n6394, new_n6396);
xnor_1 g06020(new_n6396, new_n6384, new_n6397);
nor_1  g06021(new_n1215, new_n1835_1, new_n6398);
nand_1 g06022(new_n6398, new_n6355, new_n6399);
nand_1 g06023(n9763, n8384, new_n6400);
nand_1 g06024(n7236, n3342, new_n6401);
nand_1 g06025(new_n6401, new_n6400, new_n6402);
nor_1  g06026(new_n6402, new_n6399, new_n6403);
not_1  g06027(new_n6403, new_n6404);
not_1  g06028(new_n6402, new_n6405);
nor_1  g06029(new_n6401, new_n6400, new_n6406);
nor_1  g06030(new_n6406, new_n6405, new_n6407);
nand_1 g06031(new_n6407, new_n6399, new_n6408);
nand_1 g06032(new_n6408, new_n6404, new_n6409);
xnor_1 g06033(new_n6409, new_n6397, new_n6410);
xnor_1 g06034(new_n6379, new_n6352, new_n6411);
nand_1 g06035(new_n6411, new_n6410, new_n6412);
nand_1 g06036(new_n6412, new_n6381, new_n6413);
xnor_1 g06037(new_n6413, new_n6350, new_n6414);
nor_1  g06038(new_n1925, new_n1310, new_n6415);
nor_1  g06039(new_n6392, new_n6385, new_n6416);
nor_1  g06040(new_n6416, new_n6391, new_n6417);
nand_1 g06041(new_n6417, new_n6415, new_n6418);
not_1  g06042(new_n6418, new_n6419);
nor_1  g06043(new_n6417, new_n6415, new_n6420);
nor_1  g06044(new_n6420, new_n6419, new_n6421);
nor_1  g06045(new_n1923, new_n1235, new_n6422);
nand_1 g06046(n2558, n137, new_n6423);
nand_1 g06047(n11478, n5579, new_n6424);
nand_1 g06048(new_n6424, new_n6423, new_n6425);
nor_1  g06049(new_n6424, new_n6423, new_n6426);
not_1  g06050(new_n6426, new_n6427);
nand_1 g06051(new_n6427, new_n6425, new_n6428);
xnor_1 g06052(new_n6428, new_n6422, new_n6429_1);
xnor_1 g06053(new_n6429_1, new_n6421, new_n6430);
nand_1 g06054(new_n6394, new_n6385, new_n6431_1);
nor_1  g06055(new_n6431_1, new_n6430, new_n6432);
not_1  g06056(new_n6432, new_n6433);
nand_1 g06057(new_n6431_1, new_n6430, new_n6434);
nand_1 g06058(new_n6434, new_n6433, new_n6435);
nor_1  g06059(new_n1833, new_n1325, new_n6436);
not_1  g06060(new_n6406, new_n6437);
nand_1 g06061(new_n6402, new_n6398, new_n6438);
nand_1 g06062(new_n6438, new_n6437, new_n6439);
nand_1 g06063(new_n6439, new_n6436, new_n6440);
not_1  g06064(new_n6440, new_n6441_1);
nor_1  g06065(new_n6439, new_n6436, new_n6442);
nor_1  g06066(new_n6442, new_n6441_1, new_n6443);
nor_1  g06067(new_n1215, new_n1837, new_n6444);
nand_1 g06068(n9763, n6358, new_n6445_1);
nand_1 g06069(n3992, n3342, new_n6446);
nand_1 g06070(new_n6446, new_n6445_1, new_n6447);
nor_1  g06071(new_n6446, new_n6445_1, new_n6448);
not_1  g06072(new_n6448, new_n6449);
nand_1 g06073(new_n6449, new_n6447, new_n6450);
xnor_1 g06074(new_n6450, new_n6444, new_n6451);
xnor_1 g06075(new_n6451, new_n6443, new_n6452);
not_1  g06076(new_n6452, new_n6453);
nor_1  g06077(new_n6407, new_n6370, new_n6454);
nand_1 g06078(new_n6454, new_n6453, new_n6455);
not_1  g06079(new_n6455, new_n6456);
nor_1  g06080(new_n6454, new_n6453, new_n6457);
nor_1  g06081(new_n6457, new_n6456, new_n6458);
xnor_1 g06082(new_n6458, new_n6435, new_n6459);
not_1  g06083(new_n6396, new_n6460);
nand_1 g06084(new_n6460, new_n6384, new_n6461);
not_1  g06085(new_n6409, new_n6462);
nand_1 g06086(new_n6462, new_n6397, new_n6463);
nand_1 g06087(new_n6463, new_n6461, new_n6464);
xnor_1 g06088(new_n6464, new_n6459, new_n6465);
nor_1  g06089(new_n6465, new_n6414, new_n6466);
nand_1 g06090(new_n6465, new_n6414, new_n6467);
not_1  g06091(new_n6467, new_n6468);
nor_1  g06092(new_n6468, new_n6466, new_n6469);
nand_1 g06093(new_n6469, new_n6312, new_n6470);
not_1  g06094(new_n6312, new_n6471);
not_1  g06095(new_n6469, new_n6472);
nand_1 g06096(new_n6472, new_n6471, new_n6473);
nand_1 g06097(new_n6473, new_n6470, new_n6474);
nand_1 g06098(new_n6308, new_n6281, new_n6475);
nand_1 g06099(new_n6475, new_n6310, new_n6476);
not_1  g06100(new_n6412, new_n6477);
nor_1  g06101(new_n6411, new_n6410, new_n6478);
nor_1  g06102(new_n6478, new_n6477, new_n6479);
nor_1  g06103(new_n6479, new_n6476, new_n6480);
xnor_1 g06104(new_n6359_1, new_n6331, new_n6481);
nand_1 g06105(new_n6481, new_n6283, new_n6482);
nand_1 g06106(n7265, n1333, new_n6483);
nor_1  g06107(new_n1348, new_n1130, new_n6484);
xnor_1 g06108(new_n6484, new_n6483, new_n6485);
not_1  g06109(new_n6485, new_n6486);
nand_1 g06110(new_n6486, new_n6482, new_n6487);
not_1  g06111(new_n6487, new_n6488);
xnor_1 g06112(new_n6377, new_n6376, new_n6489);
nor_1  g06113(new_n6486, new_n6482, new_n6490);
nor_1  g06114(new_n6490, new_n6488, new_n6491);
and_1  g06115(new_n6491, new_n6489, new_n6492);
nor_1  g06116(new_n6492, new_n6488, new_n6493);
not_1  g06117(new_n6493, new_n6494);
xnor_1 g06118(new_n6479, new_n6476, new_n6495);
nor_1  g06119(new_n6495, new_n6494, new_n6496);
nor_1  g06120(new_n6496, new_n6480, new_n6497);
xor_1  g06121(new_n6497, new_n6474, n1847);
nor_1  g06122(new_n456, new_n4682, new_n6499);
nor_1  g06123(new_n552, new_n4085, new_n6500);
nand_1 g06124(n5645, n5331, new_n6501);
nand_1 g06125(n11876, n7965, new_n6502);
nor_1  g06126(new_n6502, new_n6501, new_n6503);
not_1  g06127(new_n6503, new_n6504);
nand_1 g06128(new_n6502, new_n6501, new_n6505);
nand_1 g06129(new_n6505, new_n6504, new_n6506);
xnor_1 g06130(new_n6506, new_n6500, new_n6507);
nand_1 g06131(new_n6507, new_n6499, new_n6508);
nor_1  g06132(new_n456, new_n4053, new_n6509);
not_1  g06133(new_n6509, new_n6510);
nor_1  g06134(new_n424, new_n4682, new_n6511);
xnor_1 g06135(new_n6511, new_n6510, new_n6512);
not_1  g06136(new_n6512, new_n6513);
xnor_1 g06137(new_n6513, new_n6508, new_n6514);
not_1  g06138(new_n6514, new_n6515);
not_1  g06139(new_n6500, new_n6516);
nor_1  g06140(new_n6506, new_n6516, new_n6517);
not_1  g06141(new_n6517, new_n6518);
nand_1 g06142(n9640, n8759, new_n6519);
nand_1 g06143(n6776, n6703, new_n6520);
xnor_1 g06144(new_n6520, new_n6519, new_n6521);
xnor_1 g06145(new_n6521, new_n6518, new_n6522);
not_1  g06146(new_n6522, new_n6523);
nand_1 g06147(n10898, n7965, new_n6524);
nand_1 g06148(n11876, n7388, new_n6525);
xnor_1 g06149(new_n6525, new_n6524, new_n6526);
xnor_1 g06150(new_n6526, new_n6503, new_n6527);
nand_1 g06151(n5331, n1067, new_n6528);
nand_1 g06152(n8476, n5645, new_n6529);
nand_1 g06153(new_n6529, new_n6528, new_n6530);
nor_1  g06154(new_n6529, new_n6528, new_n6531);
not_1  g06155(new_n6531, new_n6532);
nand_1 g06156(new_n6532, new_n6530, new_n6533);
not_1  g06157(new_n6533, new_n6534);
nor_1  g06158(new_n6534, new_n6527, new_n6535);
nand_1 g06159(new_n6534, new_n6527, new_n6536);
not_1  g06160(new_n6536, new_n6537);
nor_1  g06161(new_n6537, new_n6535, new_n6538);
nand_1 g06162(new_n6538, new_n6523, new_n6539);
not_1  g06163(new_n6539, new_n6540);
nor_1  g06164(new_n6538, new_n6523, new_n6541);
nor_1  g06165(new_n6541, new_n6540, new_n6542);
nand_1 g06166(new_n6542, new_n6515, new_n6543);
not_1  g06167(new_n6543, new_n6544);
nor_1  g06168(new_n6542, new_n6515, new_n6545);
nor_1  g06169(new_n6545, new_n6544, n2096);
and_1  g06170(new_n3899, new_n3896, new_n6547);
nor_1  g06171(new_n6547, new_n3900, n2131);
nor_1  g06172(new_n4044, new_n1377, new_n6549);
nor_1  g06173(new_n4067, new_n4061, new_n6550);
nor_1  g06174(new_n6550, new_n4066, new_n6551);
nand_1 g06175(new_n6551, new_n6549, new_n6552);
not_1  g06176(new_n6549, new_n6553);
xnor_1 g06177(new_n6551, new_n6553, new_n6554);
nor_1  g06178(new_n4283, new_n4053, new_n6555);
not_1  g06179(new_n6555, new_n6556);
nand_1 g06180(n9920, n1798, new_n6557);
nand_1 g06181(new_n6557, new_n4051, new_n6558);
not_1  g06182(new_n6558, new_n6559);
nor_1  g06183(new_n6557, new_n4051, new_n6560);
nor_1  g06184(new_n6560, new_n6559, new_n6561);
xnor_1 g06185(new_n6561, new_n6556, new_n6562);
nand_1 g06186(new_n6562, new_n6554, new_n6563);
nand_1 g06187(new_n6563, new_n6552, new_n6564);
nor_1  g06188(new_n4665, new_n1377, new_n6565);
not_1  g06189(new_n6565, new_n6566);
nor_1  g06190(new_n4044, new_n1367, new_n6567);
not_1  g06191(new_n6567, new_n6568);
nand_1 g06192(new_n6568, new_n6566, new_n6569);
nor_1  g06193(new_n6568, new_n6566, new_n6570);
not_1  g06194(new_n6570, new_n6571);
nand_1 g06195(new_n6571, new_n6569, new_n6572);
xnor_1 g06196(new_n6572, new_n6564, new_n6573);
nor_1  g06197(new_n4627, new_n4283, new_n6574);
nand_1 g06198(n3627, n1798, new_n6575);
nand_1 g06199(n9920, n3932, new_n6576);
nand_1 g06200(new_n6576, new_n6575, new_n6577);
not_1  g06201(new_n6577, new_n6578_1);
nor_1  g06202(new_n6576, new_n6575, new_n6579);
nor_1  g06203(new_n6579, new_n6578_1, new_n6580);
nand_1 g06204(new_n6580, new_n6574, new_n6581);
not_1  g06205(new_n6581, new_n6582);
nor_1  g06206(new_n6580, new_n6574, new_n6583);
nor_1  g06207(new_n6583, new_n6582, new_n6584);
nor_1  g06208(new_n6560, new_n6555, new_n6585);
nor_1  g06209(new_n6585, new_n6559, new_n6586);
nand_1 g06210(new_n6586, new_n6584, new_n6587);
not_1  g06211(new_n6587, new_n6588);
nor_1  g06212(new_n6586, new_n6584, new_n6589);
nor_1  g06213(new_n6589, new_n6588, new_n6590);
nand_1 g06214(new_n6590, new_n6573, new_n6591);
not_1  g06215(new_n6591, new_n6592);
nor_1  g06216(new_n6590, new_n6573, new_n6593);
nor_1  g06217(new_n6593, new_n6592, new_n6594);
nor_1  g06218(new_n4665, new_n378, new_n6595);
nand_1 g06219(new_n4070, new_n4057, new_n6596);
nor_1  g06220(new_n6596, new_n6595, new_n6597);
not_1  g06221(new_n6597, new_n6598);
xnor_1 g06222(new_n6562, new_n6554, new_n6599);
not_1  g06223(new_n6595, new_n6600);
xnor_1 g06224(new_n6596, new_n6600, new_n6601);
nand_1 g06225(new_n6601, new_n6599, new_n6602);
nand_1 g06226(new_n6602, new_n6598, new_n6603);
not_1  g06227(new_n6603, new_n6604_1);
nand_1 g06228(new_n6604_1, new_n6594, new_n6605);
nand_1 g06229(new_n6587, new_n6581, new_n6606);
nor_1  g06230(new_n4709, new_n1377, new_n6607);
nand_1 g06231(n11662, n4189, new_n6608);
nand_1 g06232(n9583, n6687, new_n6609);
xnor_1 g06233(new_n6609, new_n6608, new_n6610);
and_1  g06234(new_n6610, new_n6607, new_n6611_1);
nor_1  g06235(new_n6610, new_n6607, new_n6612);
nor_1  g06236(new_n6612, new_n6611_1, new_n6613);
xnor_1 g06237(new_n6613, new_n6606, new_n6614);
nand_1 g06238(n7456, n6770, new_n6615);
xnor_1 g06239(new_n6615, new_n6579, new_n6616);
not_1  g06240(n3627, new_n6617);
nor_1  g06241(new_n4053, new_n6617, new_n6618);
not_1  g06242(new_n6618, new_n6619);
nand_1 g06243(n12591, n9920, new_n6620);
nand_1 g06244(n4516, n1798, new_n6621);
nand_1 g06245(new_n6621, new_n6620, new_n6622);
not_1  g06246(new_n6620, new_n6623);
not_1  g06247(new_n6621, new_n6624);
nand_1 g06248(new_n6624, new_n6623, new_n6625);
nand_1 g06249(new_n6625, new_n6622, new_n6626);
xnor_1 g06250(new_n6626, new_n6619, new_n6627);
xnor_1 g06251(new_n6627, new_n6616, new_n6628);
xnor_1 g06252(new_n6628, new_n6614, new_n6629);
not_1  g06253(new_n6572, new_n6630);
nand_1 g06254(new_n6630, new_n6564, new_n6631);
nand_1 g06255(new_n6592, new_n6570, new_n6632);
nand_1 g06256(new_n6591, new_n6571, new_n6633);
nand_1 g06257(new_n6633, new_n6632, new_n6634);
nand_1 g06258(new_n6634, new_n6631, new_n6635);
xnor_1 g06259(new_n6635, new_n6629, new_n6636);
xnor_1 g06260(new_n6636, new_n6605, new_n6637);
nor_1  g06261(new_n4709, new_n378, new_n6638);
not_1  g06262(new_n6605, new_n6639);
nor_1  g06263(new_n6604_1, new_n6594, new_n6640);
nor_1  g06264(new_n6640, new_n6639, new_n6641);
nand_1 g06265(new_n6641, new_n6638, new_n6642);
nand_1 g06266(new_n4080, new_n4073, new_n6643);
not_1  g06267(new_n6602, new_n6644);
nor_1  g06268(new_n6601, new_n6599, new_n6645_1);
nor_1  g06269(new_n6645_1, new_n6644, new_n6646);
nor_1  g06270(new_n6646, new_n6643, new_n6647);
not_1  g06271(new_n6638, new_n6648);
xnor_1 g06272(new_n6641, new_n6648, new_n6649);
nand_1 g06273(new_n6649, new_n6647, new_n6650);
nand_1 g06274(new_n6650, new_n6642, new_n6651);
xor_1  g06275(new_n6651, new_n6637, new_n6652);
not_1  g06276(new_n6652, new_n6653);
nor_1  g06277(new_n4761, new_n4529, new_n6654);
nand_1 g06278(n9640, n1094, new_n6655);
nand_1 g06279(n10678, n6703, new_n6656);
nand_1 g06280(new_n6656, new_n6655, new_n6657);
not_1  g06281(new_n6657, new_n6658);
nor_1  g06282(new_n6656, new_n6655, new_n6659);
nor_1  g06283(new_n6659, new_n6658, new_n6660);
nand_1 g06284(new_n6660, new_n6654, new_n6661);
not_1  g06285(new_n6661, new_n6662);
nor_1  g06286(new_n6660, new_n6654, new_n6663);
nor_1  g06287(new_n6663, new_n6662, new_n6664);
nand_1 g06288(n6703, n1094, new_n6665);
nand_1 g06289(new_n6665, new_n4124, new_n6666);
not_1  g06290(new_n6666, new_n6667);
nor_1  g06291(new_n6665, new_n4124, new_n6668);
nor_1  g06292(new_n4116, new_n4529, new_n6669);
nor_1  g06293(new_n6669, new_n6668, new_n6670);
nor_1  g06294(new_n6670, new_n6667, new_n6671);
nand_1 g06295(new_n6671, new_n6664, new_n6672);
not_1  g06296(new_n6672, new_n6673);
nor_1  g06297(new_n6671, new_n6664, new_n6674);
nor_1  g06298(new_n6674, new_n6673, new_n6675);
nand_1 g06299(n10928, n10451, new_n6676);
nand_1 g06300(n11023, n6986, new_n6677);
nand_1 g06301(new_n6677, new_n6676, new_n6678);
nor_1  g06302(new_n6677, new_n6676, new_n6679);
not_1  g06303(new_n6679, new_n6680);
nand_1 g06304(new_n6680, new_n6678, new_n6681);
xnor_1 g06305(new_n6681, new_n6675, new_n6682);
nor_1  g06306(new_n4232, new_n1434, new_n6683);
not_1  g06307(new_n4240, new_n6684);
nor_1  g06308(new_n4241, new_n4237, new_n6685);
nor_1  g06309(new_n6685, new_n6684, new_n6686);
nand_1 g06310(new_n6686, new_n6683, new_n6687_1);
not_1  g06311(new_n6687_1, new_n6688);
nor_1  g06312(new_n6686, new_n6683, new_n6689_1);
nor_1  g06313(new_n6689_1, new_n6688, new_n6690);
not_1  g06314(new_n6669, new_n6691);
not_1  g06315(new_n6668, new_n6692);
nand_1 g06316(new_n6692, new_n6666, new_n6693);
xnor_1 g06317(new_n6693, new_n6691, new_n6694);
not_1  g06318(new_n6694, new_n6695);
nand_1 g06319(new_n6695, new_n6690, new_n6696);
nand_1 g06320(new_n6696, new_n6687_1, new_n6697);
xnor_1 g06321(new_n6697, new_n6682, new_n6698);
not_1  g06322(new_n6698, new_n6699);
nor_1  g06323(new_n4815, new_n382, new_n6700);
xnor_1 g06324(new_n6694, new_n6690, new_n6701);
nand_1 g06325(new_n6701, new_n6700, new_n6702);
nand_1 g06326(new_n4235, new_n4233, new_n6703_1);
not_1  g06327(new_n4236, new_n6704);
nand_1 g06328(new_n4244, new_n6704, new_n6705);
nand_1 g06329(new_n6705, new_n6703_1, new_n6706);
not_1  g06330(new_n6702, new_n6707);
nor_1  g06331(new_n6701, new_n6700, new_n6708);
nor_1  g06332(new_n6708, new_n6707, new_n6709);
nand_1 g06333(new_n6709, new_n6706, new_n6710);
nand_1 g06334(new_n6710, new_n6702, new_n6711);
nand_1 g06335(new_n6711, new_n6699, new_n6712);
nand_1 g06336(new_n6672, new_n6661, new_n6713);
nor_1  g06337(new_n1434, new_n4852, new_n6714);
nand_1 g06338(n10451, n6986, new_n6715);
nand_1 g06339(n11423, n8336, new_n6716);
xnor_1 g06340(new_n6716, new_n6715, new_n6717);
and_1  g06341(new_n6717, new_n6714, new_n6718);
nor_1  g06342(new_n6717, new_n6714, new_n6719);
nor_1  g06343(new_n6719, new_n6718, new_n6720);
xnor_1 g06344(new_n6720, new_n6713, new_n6721);
nor_1  g06345(new_n4232, new_n4529, new_n6722);
xnor_1 g06346(new_n6722, new_n6659, new_n6723);
not_1  g06347(new_n6723, new_n6724);
not_1  g06348(n10678, new_n6725);
nor_1  g06349(new_n6725, new_n4116, new_n6726);
not_1  g06350(new_n6726, new_n6727);
nand_1 g06351(n3022, n1094, new_n6728);
nand_1 g06352(n7320, n6703, new_n6729);
xnor_1 g06353(new_n6729, new_n6728, new_n6730);
xnor_1 g06354(new_n6730, new_n6727, new_n6731);
xnor_1 g06355(new_n6731, new_n6724, new_n6732);
xnor_1 g06356(new_n6732, new_n6721, new_n6733);
not_1  g06357(new_n6681, new_n6734);
nand_1 g06358(new_n6734, new_n6675, new_n6735);
nand_1 g06359(new_n6697, new_n6682, new_n6736);
xnor_1 g06360(new_n6736, new_n6680, new_n6737);
nand_1 g06361(new_n6737, new_n6735, new_n6738);
xnor_1 g06362(new_n6738, new_n6733, new_n6739);
not_1  g06363(new_n6739, new_n6740);
xnor_1 g06364(new_n6740, new_n6712, new_n6741);
nand_1 g06365(n10278, n8336, new_n6742_1);
xnor_1 g06366(new_n6711, new_n6698, new_n6743);
not_1  g06367(new_n6743, new_n6744);
nand_1 g06368(new_n6744, new_n6742_1, new_n6745);
not_1  g06369(new_n6710, new_n6746);
nor_1  g06370(new_n6709, new_n6706, new_n6747);
nor_1  g06371(new_n6747, new_n6746, new_n6748);
nand_1 g06372(new_n6748, new_n4249, new_n6749);
xnor_1 g06373(new_n6743, new_n6742_1, new_n6750);
nand_1 g06374(new_n6750, new_n6749, new_n6751);
nand_1 g06375(new_n6751, new_n6745, new_n6752);
xnor_1 g06376(new_n6752, new_n6741, new_n6753);
nor_1  g06377(new_n4132, new_n1538, new_n6754);
not_1  g06378(new_n6754, new_n6755);
nand_1 g06379(n4828, n1067, new_n6756);
nand_1 g06380(n5645, n2515, new_n6757);
xnor_1 g06381(new_n6757, new_n6756, new_n6758);
nor_1  g06382(new_n6758, new_n6755, new_n6759);
not_1  g06383(new_n6759, new_n6760);
nand_1 g06384(new_n6758, new_n6755, new_n6761);
nand_1 g06385(new_n6761, new_n6760, new_n6762);
not_1  g06386(new_n6762, new_n6763);
nand_1 g06387(n5645, n4828, new_n6764);
nand_1 g06388(n8665, n7891, new_n6765);
nand_1 g06389(new_n6765, new_n6764, new_n6766);
not_1  g06390(new_n6766, new_n6767);
nor_1  g06391(new_n1538, new_n4919, new_n6768);
xnor_1 g06392(new_n6765, new_n6764, new_n6769);
nor_1  g06393(new_n6769, new_n6768, new_n6770_1);
nor_1  g06394(new_n6770_1, new_n6767, new_n6771);
nand_1 g06395(new_n6771, new_n6763, new_n6772);
not_1  g06396(new_n6772, new_n6773);
nor_1  g06397(new_n6771, new_n6763, new_n6774);
nor_1  g06398(new_n6774, new_n6773, new_n6775);
nor_1  g06399(new_n1452, new_n4951, new_n6776_1);
not_1  g06400(new_n6776_1, new_n6777);
nor_1  g06401(new_n4187_1, new_n4386, new_n6778);
not_1  g06402(new_n6778, new_n6779);
nand_1 g06403(new_n6779, new_n6777, new_n6780);
nor_1  g06404(new_n6779, new_n6777, new_n6781);
not_1  g06405(new_n6781, new_n6782);
nand_1 g06406(new_n6782, new_n6780, new_n6783);
xnor_1 g06407(new_n6783, new_n6775, new_n6784);
nor_1  g06408(new_n1452, new_n4187_1, new_n6785);
nand_1 g06409(new_n4199, new_n4198, new_n6786);
not_1  g06410(new_n6786, new_n6787);
nor_1  g06411(new_n4200, new_n4196, new_n6788);
nor_1  g06412(new_n6788, new_n6787, new_n6789);
nand_1 g06413(new_n6789, new_n6785, new_n6790);
xnor_1 g06414(new_n6769, new_n6768, new_n6791);
not_1  g06415(new_n6785, new_n6792);
xnor_1 g06416(new_n6789, new_n6792, new_n6793);
nand_1 g06417(new_n6793, new_n6791, new_n6794);
nand_1 g06418(new_n6794, new_n6790, new_n6795);
xnor_1 g06419(new_n6795, new_n6784, new_n6796);
not_1  g06420(new_n6796, new_n6797_1);
nor_1  g06421(new_n1533, new_n4951, new_n6798);
xnor_1 g06422(new_n6793, new_n6791, new_n6799);
not_1  g06423(new_n6799, new_n6800);
nand_1 g06424(new_n6800, new_n6798, new_n6801);
not_1  g06425(new_n6798, new_n6802);
nand_1 g06426(new_n6799, new_n6802, new_n6803);
nand_1 g06427(new_n4193, new_n4188, new_n6804);
not_1  g06428(new_n4201, new_n6805);
nand_1 g06429(new_n6805, new_n4194, new_n6806_1);
nand_1 g06430(new_n6806_1, new_n6804, new_n6807);
nand_1 g06431(new_n6807, new_n6803, new_n6808);
nand_1 g06432(new_n6808, new_n6801, new_n6809_1);
nand_1 g06433(new_n6809_1, new_n6797_1, new_n6810);
nand_1 g06434(new_n6772, new_n6760, new_n6811);
nor_1  g06435(new_n4908, new_n1452, new_n6812);
nand_1 g06436(n7891, n2551, new_n6813);
nand_1 g06437(n12069, n4094, new_n6814);
xnor_1 g06438(new_n6814, new_n6813, new_n6815);
xnor_1 g06439(new_n6815, new_n6812, new_n6816);
not_1  g06440(new_n6816, new_n6817);
xnor_1 g06441(new_n6817, new_n6811, new_n6818);
nor_1  g06442(new_n6757, new_n6756, new_n6819);
nor_1  g06443(new_n4187_1, new_n1538, new_n6820);
xnor_1 g06444(new_n6820, new_n6819, new_n6821);
not_1  g06445(new_n6821, new_n6822_1);
not_1  g06446(n2515, new_n6823);
nor_1  g06447(new_n6823, new_n4919, new_n6824);
not_1  g06448(n4828, new_n6825);
nor_1  g06449(new_n4132, new_n6825, new_n6826_1);
not_1  g06450(new_n6826_1, new_n6827);
not_1  g06451(n1199, new_n6828);
nor_1  g06452(new_n4195, new_n6828, new_n6829);
not_1  g06453(new_n6829, new_n6830);
nand_1 g06454(new_n6830, new_n6827, new_n6831);
nand_1 g06455(new_n6829, new_n6826_1, new_n6832);
nand_1 g06456(new_n6832, new_n6831, new_n6833);
xnor_1 g06457(new_n6833, new_n6824, new_n6834);
xnor_1 g06458(new_n6834, new_n6822_1, new_n6835);
xnor_1 g06459(new_n6835, new_n6818, new_n6836);
not_1  g06460(new_n6775, new_n6837);
nor_1  g06461(new_n6783, new_n6837, new_n6838);
not_1  g06462(new_n6838, new_n6839);
nand_1 g06463(new_n6795, new_n6784, new_n6840);
xnor_1 g06464(new_n6840, new_n6782, new_n6841);
nand_1 g06465(new_n6841, new_n6839, new_n6842);
xnor_1 g06466(new_n6842, new_n6836, new_n6843);
xnor_1 g06467(new_n6843, new_n6810, new_n6844);
nor_1  g06468(new_n4908, new_n1533, new_n6845);
not_1  g06469(new_n6845, new_n6846);
xnor_1 g06470(new_n6809_1, new_n6796, new_n6847);
not_1  g06471(new_n6847, new_n6848);
nand_1 g06472(new_n6848, new_n6846, new_n6849);
nand_1 g06473(new_n4202, new_n4186, new_n6850);
not_1  g06474(new_n6850, new_n6851);
nand_1 g06475(new_n6803, new_n6801, new_n6852);
xnor_1 g06476(new_n6852, new_n6807, new_n6853);
nand_1 g06477(new_n6853, new_n6851, new_n6854);
nand_1 g06478(new_n6847, new_n6845, new_n6855);
nand_1 g06479(new_n6855, new_n6849, new_n6856);
not_1  g06480(new_n6856, new_n6857);
nand_1 g06481(new_n6857, new_n6854, new_n6858);
nand_1 g06482(new_n6858, new_n6849, new_n6859);
xnor_1 g06483(new_n6859, new_n6844, new_n6860_1);
nor_1  g06484(new_n5052, new_n4542, new_n6861);
nand_1 g06485(n10898, n5767, new_n6862);
nand_1 g06486(n11876, n5319, new_n6863);
xnor_1 g06487(new_n6863, new_n6862, new_n6864);
xnor_1 g06488(new_n6864, new_n6861, new_n6865);
nand_1 g06489(n10898, n996, new_n6866);
nand_1 g06490(new_n6866, new_n4151, new_n6867);
not_1  g06491(new_n6867, new_n6868);
not_1  g06492(n5767, new_n6869);
nor_1  g06493(new_n4088_1, new_n6869, new_n6870);
xnor_1 g06494(new_n6866, new_n4151, new_n6871);
nor_1  g06495(new_n6871, new_n6870, new_n6872);
nor_1  g06496(new_n6872, new_n6868, new_n6873);
nand_1 g06497(new_n6873, new_n6865, new_n6874);
not_1  g06498(new_n6874, new_n6875);
nor_1  g06499(new_n6873, new_n6865, new_n6876);
nor_1  g06500(new_n6876, new_n6875, new_n6877_1);
nor_1  g06501(new_n1467, new_n5065, new_n6878);
not_1  g06502(new_n6878, new_n6879);
nor_1  g06503(new_n1562, new_n4204, new_n6880);
not_1  g06504(new_n6880, new_n6881);
nand_1 g06505(new_n6881, new_n6879, new_n6882);
nor_1  g06506(new_n6881, new_n6879, new_n6883);
not_1  g06507(new_n6883, new_n6884);
nand_1 g06508(new_n6884, new_n6882, new_n6885);
xnor_1 g06509(new_n6885, new_n6877_1, new_n6886);
nor_1  g06510(new_n1467, new_n4204, new_n6887);
nand_1 g06511(new_n4215, new_n4214, new_n6888);
not_1  g06512(new_n6888, new_n6889);
nor_1  g06513(new_n4216, new_n4212, new_n6890);
nor_1  g06514(new_n6890, new_n6889, new_n6891);
nand_1 g06515(new_n6891, new_n6887, new_n6892);
not_1  g06516(new_n6892, new_n6893);
nor_1  g06517(new_n6891, new_n6887, new_n6894);
nor_1  g06518(new_n6894, new_n6893, new_n6895);
not_1  g06519(new_n6870, new_n6896);
xnor_1 g06520(new_n6871, new_n6896, new_n6897);
not_1  g06521(new_n6897, new_n6898);
nand_1 g06522(new_n6898, new_n6895, new_n6899);
nand_1 g06523(new_n6899, new_n6892, new_n6900);
nand_1 g06524(new_n6900, new_n6886, new_n6901);
not_1  g06525(new_n6901, new_n6902);
nor_1  g06526(new_n6900, new_n6886, new_n6903);
nor_1  g06527(new_n6903, new_n6902, new_n6904);
nor_1  g06528(new_n385, new_n5065, new_n6905);
xnor_1 g06529(new_n6898, new_n6895, new_n6906);
not_1  g06530(new_n6906, new_n6907);
nand_1 g06531(new_n6907, new_n6905, new_n6908);
not_1  g06532(new_n6905, new_n6909);
nand_1 g06533(new_n6906, new_n6909, new_n6910);
nand_1 g06534(new_n4218, new_n4211, new_n6911);
nand_1 g06535(new_n6911, new_n4208, new_n6912);
nand_1 g06536(new_n6912, new_n6910, new_n6913);
nand_1 g06537(new_n6913, new_n6908, new_n6914);
nand_1 g06538(new_n6914, new_n6904, new_n6915);
not_1  g06539(new_n6885, new_n6916);
nand_1 g06540(new_n6916, new_n6877_1, new_n6917);
nand_1 g06541(new_n6902, new_n6883, new_n6918);
nand_1 g06542(new_n6901, new_n6884, new_n6919);
nand_1 g06543(new_n6919, new_n6918, new_n6920);
nand_1 g06544(new_n6920, new_n6917, new_n6921);
not_1  g06545(new_n6861, new_n6922);
nor_1  g06546(new_n6864, new_n6922, new_n6923);
nor_1  g06547(new_n6875, new_n6923, new_n6924);
nor_1  g06548(new_n1467, new_n5107, new_n6925);
nand_1 g06549(n5314, n159, new_n6926);
nand_1 g06550(n12247, n11222, new_n6927);
xnor_1 g06551(new_n6927, new_n6926, new_n6928);
xnor_1 g06552(new_n6928, new_n6925, new_n6929);
xnor_1 g06553(new_n6929, new_n6924, new_n6930);
not_1  g06554(new_n6930, new_n6931);
nor_1  g06555(new_n6863, new_n6862, new_n6932);
nor_1  g06556(new_n4204, new_n4542, new_n6933);
xnor_1 g06557(new_n6933, new_n6932, new_n6934);
not_1  g06558(n5319, new_n6935);
nor_1  g06559(new_n4143, new_n6935, new_n6936);
nand_1 g06560(n11876, n9457, new_n6937);
nand_1 g06561(n5767, n3754, new_n6938);
xnor_1 g06562(new_n6938, new_n6937, new_n6939);
xnor_1 g06563(new_n6939, new_n6936, new_n6940);
not_1  g06564(new_n6940, new_n6941);
nand_1 g06565(new_n6941, new_n6934, new_n6942);
not_1  g06566(new_n6934, new_n6943);
nand_1 g06567(new_n6940, new_n6943, new_n6944);
and_1  g06568(new_n6944, new_n6942, new_n6945);
not_1  g06569(new_n6945, new_n6946);
nor_1  g06570(new_n6946, new_n6931, new_n6947);
nor_1  g06571(new_n6945, new_n6930, new_n6948);
nor_1  g06572(new_n6948, new_n6947, new_n6949);
not_1  g06573(new_n6949, new_n6950);
xnor_1 g06574(new_n6950, new_n6921, new_n6951);
xnor_1 g06575(new_n6951, new_n6915, new_n6952);
nor_1  g06576(new_n385, new_n5107, new_n6953);
not_1  g06577(new_n6915, new_n6954);
nor_1  g06578(new_n6914, new_n6904, new_n6955);
nor_1  g06579(new_n6955, new_n6954, new_n6956);
nor_1  g06580(new_n6956, new_n6953, new_n6957);
nor_1  g06581(new_n4220, new_n4219, new_n6958);
nand_1 g06582(new_n6910, new_n6908, new_n6959);
xnor_1 g06583(new_n6959, new_n6912, new_n6960);
nand_1 g06584(new_n6960, new_n6958, new_n6961);
not_1  g06585(new_n6961, new_n6962);
xnor_1 g06586(new_n6956, new_n6953, new_n6963);
nor_1  g06587(new_n6963, new_n6962, new_n6964);
nor_1  g06588(new_n6964, new_n6957, new_n6965);
xnor_1 g06589(new_n6965, new_n6952, new_n6966);
xnor_1 g06590(new_n6963, new_n6962, new_n6967);
xnor_1 g06591(new_n6856, new_n6854, new_n6968);
not_1  g06592(new_n6968, new_n6969);
nand_1 g06593(new_n6969, new_n6967, new_n6970);
not_1  g06594(new_n6967, new_n6971);
nand_1 g06595(new_n6968, new_n6971, new_n6972);
xnor_1 g06596(new_n6853, new_n6851, new_n6973);
not_1  g06597(new_n4222, new_n6974);
nand_1 g06598(new_n6974, new_n4203_1, new_n6975);
nand_1 g06599(new_n4227, new_n6975, new_n6976);
nand_1 g06600(new_n6976, new_n6973, new_n6977);
not_1  g06601(new_n6977, new_n6978);
nor_1  g06602(new_n6960, new_n6958, new_n6979);
nor_1  g06603(new_n6979, new_n6962, new_n6980);
xnor_1 g06604(new_n6976, new_n6973, new_n6981);
nor_1  g06605(new_n6981, new_n6980, new_n6982);
nor_1  g06606(new_n6982, new_n6978, new_n6983);
nand_1 g06607(new_n6983, new_n6972, new_n6984);
nand_1 g06608(new_n6984, new_n6970, new_n6985);
xnor_1 g06609(new_n6985, new_n6966, new_n6986_1);
xnor_1 g06610(new_n6986_1, new_n6860_1, new_n6987);
xnor_1 g06611(new_n6987, new_n6753, new_n6988);
xnor_1 g06612(new_n6750, new_n6749, new_n6989);
xnor_1 g06613(new_n6748, new_n4248, new_n6990);
not_1  g06614(new_n6990, new_n6991);
not_1  g06615(new_n6980, new_n6992);
xnor_1 g06616(new_n6981, new_n6992, new_n6993);
nor_1  g06617(new_n6993, new_n6991, new_n6994);
not_1  g06618(new_n6994, new_n6995);
nor_1  g06619(new_n4261, new_n4256, new_n6996);
not_1  g06620(new_n6996, new_n6997);
xnor_1 g06621(new_n6993, new_n6990, new_n6998);
nand_1 g06622(new_n6998, new_n6997, new_n6999);
nand_1 g06623(new_n6999, new_n6995, new_n7000);
nand_1 g06624(new_n7000, new_n6989, new_n7001);
xnor_1 g06625(new_n7000, new_n6989, new_n7002);
nand_1 g06626(new_n6972, new_n6970, new_n7003);
xnor_1 g06627(new_n7003, new_n6983, new_n7004);
not_1  g06628(new_n7004, new_n7005);
nor_1  g06629(new_n7005, new_n7002, new_n7006);
not_1  g06630(new_n7006, new_n7007);
nand_1 g06631(new_n7007, new_n7001, new_n7008);
xnor_1 g06632(new_n7008, new_n6988, new_n7009);
nor_1  g06633(new_n7009, new_n6653, new_n7010);
not_1  g06634(new_n7009, new_n7011);
nor_1  g06635(new_n7011, new_n6652, new_n7012);
nor_1  g06636(new_n7012, new_n7010, new_n7013);
xor_1  g06637(new_n6649, new_n6647, new_n7014);
not_1  g06638(new_n7014, new_n7015);
nand_1 g06639(new_n7005, new_n7002, new_n7016);
nand_1 g06640(new_n7016, new_n7007, new_n7017);
nor_1  g06641(new_n7017, new_n7015, new_n7018);
not_1  g06642(new_n7017, new_n7019);
nor_1  g06643(new_n7019, new_n7014, new_n7020);
xor_1  g06644(new_n6646, new_n6643, new_n7021);
xnor_1 g06645(new_n6998, new_n6996, new_n7022);
nor_1  g06646(new_n7022, new_n7021, new_n7023);
not_1  g06647(new_n7023, new_n7024);
nor_1  g06648(new_n4184, new_n4082, new_n7025);
not_1  g06649(new_n4262, new_n7026);
nor_1  g06650(new_n7026, new_n4185, new_n7027);
nor_1  g06651(new_n7027, new_n7025, new_n7028);
not_1  g06652(new_n7021, new_n7029);
xnor_1 g06653(new_n7022, new_n7029, new_n7030);
nand_1 g06654(new_n7030, new_n7028, new_n7031);
nand_1 g06655(new_n7031, new_n7024, new_n7032);
nor_1  g06656(new_n7032, new_n7020, new_n7033);
nor_1  g06657(new_n7033, new_n7018, new_n7034);
xnor_1 g06658(new_n7034, new_n7013, n2301);
xnor_1 g06659(new_n4182, new_n4180, n2316);
nand_1 g06660(n4634, n1333, new_n7037);
not_1  g06661(new_n7037, new_n7038);
not_1  g06662(new_n6298, new_n7039);
nor_1  g06663(new_n6299, new_n6295, new_n7040);
nor_1  g06664(new_n7040, new_n7039, new_n7041);
nand_1 g06665(new_n7041, new_n7038, new_n7042);
xnor_1 g06666(new_n7041, new_n7037, new_n7043);
nor_1  g06667(new_n1592, new_n1130, new_n7044);
nor_1  g06668(new_n1142, new_n4720, new_n7045);
not_1  g06669(new_n7045, new_n7046);
nand_1 g06670(new_n7046, new_n6286, new_n7047);
nand_1 g06671(new_n7045, new_n6285, new_n7048);
nand_1 g06672(new_n7048, new_n7047, new_n7049);
xnor_1 g06673(new_n7049, new_n7044, new_n7050);
nand_1 g06674(new_n7050, new_n7043, new_n7051);
nand_1 g06675(new_n7051, new_n7042, new_n7052);
nor_1  g06676(new_n1121, new_n1600, new_n7053);
not_1  g06677(new_n7053, new_n7054);
nor_1  g06678(new_n5516, new_n1590, new_n7055);
not_1  g06679(new_n7055, new_n7056);
nor_1  g06680(new_n7056, new_n7054, new_n7057);
not_1  g06681(new_n7057, new_n7058);
nand_1 g06682(new_n7056, new_n7054, new_n7059);
nand_1 g06683(new_n7059, new_n7058, new_n7060);
xnor_1 g06684(new_n7060, new_n7052, new_n7061);
nand_1 g06685(n11757, n10223, new_n7062);
nand_1 g06686(n5240, n2879, new_n7063);
nand_1 g06687(n11821, n7265, new_n7064);
nand_1 g06688(new_n7064, new_n7063, new_n7065);
nor_1  g06689(new_n7064, new_n7063, new_n7066);
not_1  g06690(new_n7066, new_n7067);
nand_1 g06691(new_n7067, new_n7065, new_n7068);
xnor_1 g06692(new_n7068, new_n7062, new_n7069);
not_1  g06693(new_n7069, new_n7070);
not_1  g06694(new_n7047, new_n7071);
not_1  g06695(new_n7048, new_n7072);
nor_1  g06696(new_n7072, new_n7044, new_n7073);
nor_1  g06697(new_n7073, new_n7071, new_n7074);
not_1  g06698(new_n7074, new_n7075);
nand_1 g06699(new_n7075, new_n7070, new_n7076);
nand_1 g06700(new_n7074, new_n7069, new_n7077);
nand_1 g06701(new_n7077, new_n7076, new_n7078);
xnor_1 g06702(new_n7078, new_n7061, new_n7079);
not_1  g06703(new_n7079, new_n7080);
nor_1  g06704(new_n5516, new_n1348, new_n7081);
not_1  g06705(new_n7051, new_n7082);
nor_1  g06706(new_n7050, new_n7043, new_n7083);
nor_1  g06707(new_n7083, new_n7082, new_n7084);
nand_1 g06708(new_n7084, new_n7081, new_n7085);
nand_1 g06709(new_n6303, new_n6291, new_n7086);
not_1  g06710(new_n7085, new_n7087);
nor_1  g06711(new_n7084, new_n7081, new_n7088);
nor_1  g06712(new_n7088, new_n7087, new_n7089);
nand_1 g06713(new_n7089, new_n7086, new_n7090);
nand_1 g06714(new_n7090, new_n7085, new_n7091);
nand_1 g06715(new_n7091, new_n7080, new_n7092);
nand_1 g06716(new_n7068, new_n7062, new_n7093);
nand_1 g06717(new_n7076, new_n7093, new_n7094);
nor_1  g06718(new_n5550, new_n1590, new_n7095);
nand_1 g06719(n9195, n3172, new_n7096);
nand_1 g06720(n7862, n3865, new_n7097);
nor_1  g06721(new_n7097, new_n7096, new_n7098);
nand_1 g06722(new_n7097, new_n7096, new_n7099);
not_1  g06723(new_n7099, new_n7100);
nor_1  g06724(new_n7100, new_n7098, new_n7101);
xnor_1 g06725(new_n7101, new_n7095, new_n7102);
xnor_1 g06726(new_n7102, new_n7094, new_n7103);
nor_1  g06727(new_n1592, new_n1121, new_n7104);
not_1  g06728(new_n7104, new_n7105);
nand_1 g06729(new_n7105, new_n7067, new_n7106);
nand_1 g06730(new_n7104, new_n7066, new_n7107);
and_1  g06731(new_n7107, new_n7106, new_n7108);
not_1  g06732(new_n7108, new_n7109);
nor_1  g06733(new_n1682, new_n1130, new_n7110);
nand_1 g06734(n10223, n5240, new_n7111);
nand_1 g06735(n9080, n7265, new_n7112);
xnor_1 g06736(new_n7112, new_n7111, new_n7113);
xor_1  g06737(new_n7113, new_n7110, new_n7114);
xnor_1 g06738(new_n7114, new_n7109, new_n7115);
xnor_1 g06739(new_n7115, new_n7103, new_n7116);
not_1  g06740(new_n7052, new_n7117);
nor_1  g06741(new_n7060, new_n7117, new_n7118);
nand_1 g06742(new_n7078, new_n7061, new_n7119);
xnor_1 g06743(new_n7119, new_n7057, new_n7120);
nor_1  g06744(new_n7120, new_n7118, new_n7121);
nor_1  g06745(new_n7121, new_n7116, new_n7122);
and_1  g06746(new_n7121, new_n7116, new_n7123);
nor_1  g06747(new_n7123, new_n7122, new_n7124);
xnor_1 g06748(new_n7124, new_n7092, new_n7125);
nor_1  g06749(new_n1348, new_n5550, new_n7126);
not_1  g06750(new_n7092, new_n7127);
nor_1  g06751(new_n7091, new_n7080, new_n7128);
nor_1  g06752(new_n7128, new_n7127, new_n7129);
nand_1 g06753(new_n7129, new_n7126, new_n7130);
nand_1 g06754(new_n6311, new_n6306, new_n7131);
xnor_1 g06755(new_n7089, new_n7086, new_n7132);
nor_1  g06756(new_n7132, new_n7131, new_n7133);
not_1  g06757(new_n7126, new_n7134);
xnor_1 g06758(new_n7129, new_n7134, new_n7135);
nand_1 g06759(new_n7135, new_n7133, new_n7136);
nand_1 g06760(new_n7136, new_n7130, new_n7137);
xnor_1 g06761(new_n7137, new_n7125, new_n7138);
xnor_1 g06762(new_n7135, new_n7133, new_n7139);
xnor_1 g06763(new_n7132, new_n7131, new_n7140);
nor_1  g06764(new_n5592, new_n1350, new_n7141);
nand_1 g06765(n9400, n2522, new_n7142);
nor_1  g06766(new_n1747, new_n1192, new_n7143);
nor_1  g06767(new_n1196, new_n4769, new_n7144);
not_1  g06768(new_n7144, new_n7145);
nand_1 g06769(new_n7145, new_n6334, new_n7146);
nand_1 g06770(new_n7144, new_n6333, new_n7147);
nand_1 g06771(new_n7147, new_n7146, new_n7148);
xnor_1 g06772(new_n7148, new_n7143, new_n7149);
xnor_1 g06773(new_n7149, new_n7142, new_n7150);
nand_1 g06774(new_n6317, new_n6316, new_n7151);
not_1  g06775(new_n7151, new_n7152);
nor_1  g06776(new_n6320, new_n7152, new_n7153);
xnor_1 g06777(new_n7153, new_n7150, new_n7154);
xnor_1 g06778(new_n7154, new_n7141, new_n7155);
nand_1 g06779(new_n6338, new_n6326, new_n7156);
not_1  g06780(new_n7156, new_n7157);
nor_1  g06781(new_n7157, new_n6324, new_n7158);
xnor_1 g06782(new_n7158, new_n7155, new_n7159_1);
nand_1 g06783(new_n7159_1, new_n6349, new_n7160_1);
not_1  g06784(new_n7160_1, new_n7161);
nor_1  g06785(new_n7159_1, new_n6349, new_n7162);
nor_1  g06786(new_n7162, new_n7161, new_n7163);
not_1  g06787(new_n7163, new_n7164);
not_1  g06788(new_n6413, new_n7165);
nand_1 g06789(new_n7165, new_n6350, new_n7166);
nand_1 g06790(new_n6467, new_n7166, new_n7167);
xnor_1 g06791(new_n7167, new_n7164, new_n7168);
nor_1  g06792(new_n1931, new_n1310, new_n7169);
not_1  g06793(new_n6425, new_n7170);
nor_1  g06794(new_n6426, new_n6422, new_n7171);
nor_1  g06795(new_n7171, new_n7170, new_n7172);
nand_1 g06796(new_n7172, new_n7169, new_n7173);
not_1  g06797(new_n7173, new_n7174);
nor_1  g06798(new_n7172, new_n7169, new_n7175);
nor_1  g06799(new_n7175, new_n7174, new_n7176);
nor_1  g06800(new_n1235, new_n1959, new_n7177);
nor_1  g06801(new_n1244, new_n1923, new_n7178);
not_1  g06802(new_n7178, new_n7179);
nor_1  g06803(new_n3966, new_n4615, new_n7180);
not_1  g06804(new_n7180, new_n7181);
nand_1 g06805(new_n7181, new_n7179, new_n7182);
nor_1  g06806(new_n7181, new_n7179, new_n7183);
not_1  g06807(new_n7183, new_n7184);
nand_1 g06808(new_n7184, new_n7182, new_n7185);
xnor_1 g06809(new_n7185, new_n7177, new_n7186);
xnor_1 g06810(new_n7186, new_n7176, new_n7187);
nor_1  g06811(new_n5658, new_n1925, new_n7188);
not_1  g06812(new_n7188, new_n7189);
nand_1 g06813(new_n6429_1, new_n6421, new_n7190);
nand_1 g06814(new_n7190, new_n6418, new_n7191);
xnor_1 g06815(new_n7191, new_n7189, new_n7192);
nand_1 g06816(new_n7192, new_n7187, new_n7193_1);
not_1  g06817(new_n7193_1, new_n7194);
nor_1  g06818(new_n7192, new_n7187, new_n7195);
nor_1  g06819(new_n7195, new_n7194, new_n7196);
xnor_1 g06820(new_n7196, new_n6432, new_n7197);
nor_1  g06821(new_n5685, new_n1833, new_n7198);
not_1  g06822(new_n7198, new_n7199);
nand_1 g06823(new_n6451, new_n6443, new_n7200);
nand_1 g06824(new_n7200, new_n6440, new_n7201);
xnor_1 g06825(new_n7201, new_n7199, new_n7202);
nor_1  g06826(new_n1835_1, new_n1325, new_n7203);
not_1  g06827(new_n6447, new_n7204);
nor_1  g06828(new_n6448, new_n6444, new_n7205);
nor_1  g06829(new_n7205, new_n7204, new_n7206);
nand_1 g06830(new_n7206, new_n7203, new_n7207);
not_1  g06831(new_n7207, new_n7208);
nor_1  g06832(new_n7206, new_n7203, new_n7209);
nor_1  g06833(new_n7209, new_n7208, new_n7210);
nor_1  g06834(new_n1215, new_n1866, new_n7211);
nand_1 g06835(n8384, n3342, new_n7212);
nand_1 g06836(n9763, n5198, new_n7213);
xnor_1 g06837(new_n7213, new_n7212, new_n7214);
nor_1  g06838(new_n7214, new_n7211, new_n7215);
not_1  g06839(new_n7215, new_n7216);
nand_1 g06840(new_n7214, new_n7211, new_n7217);
nand_1 g06841(new_n7217, new_n7216, new_n7218);
nand_1 g06842(new_n7218, new_n7210, new_n7219);
not_1  g06843(new_n7219, new_n7220);
nor_1  g06844(new_n7218, new_n7210, new_n7221);
nor_1  g06845(new_n7221, new_n7220, new_n7222);
not_1  g06846(new_n7222, new_n7223);
xnor_1 g06847(new_n7223, new_n7202, new_n7224);
not_1  g06848(new_n7224, new_n7225);
nor_1  g06849(new_n7225, new_n6455, new_n7226);
nor_1  g06850(new_n7224, new_n6456, new_n7227);
nor_1  g06851(new_n7227, new_n7226, new_n7228);
not_1  g06852(new_n7228, new_n7229);
xnor_1 g06853(new_n7229, new_n7197, new_n7230);
not_1  g06854(new_n6458, new_n7231);
nand_1 g06855(new_n7231, new_n6435, new_n7232);
nand_1 g06856(new_n6464, new_n6459, new_n7233);
nand_1 g06857(new_n7233, new_n7232, new_n7234);
nand_1 g06858(new_n7234, new_n7230, new_n7235);
not_1  g06859(new_n7235, new_n7236_1);
nor_1  g06860(new_n7234, new_n7230, new_n7237);
nor_1  g06861(new_n7237, new_n7236_1, new_n7238);
nand_1 g06862(new_n7238, new_n7168, new_n7239);
not_1  g06863(new_n7239, new_n7240);
nor_1  g06864(new_n7238, new_n7168, new_n7241);
nor_1  g06865(new_n7241, new_n7240, new_n7242);
nand_1 g06866(new_n7242, new_n7140, new_n7243);
not_1  g06867(new_n7140, new_n7244);
xnor_1 g06868(new_n7242, new_n7244, new_n7245);
nand_1 g06869(new_n6497, new_n6470, new_n7246);
nand_1 g06870(new_n7246, new_n6473, new_n7247);
nand_1 g06871(new_n7247, new_n7245, new_n7248);
nand_1 g06872(new_n7248, new_n7243, new_n7249);
nand_1 g06873(new_n7249, new_n7139, new_n7250);
nor_1  g06874(new_n7167, new_n7163, new_n7251);
not_1  g06875(new_n7251, new_n7252);
nand_1 g06876(new_n7239, new_n7252, new_n7253);
nor_1  g06877(new_n5615, new_n1350, new_n7254);
not_1  g06878(new_n7254, new_n7255);
not_1  g06879(new_n7141, new_n7256);
nor_1  g06880(new_n7154, new_n7256, new_n7257);
not_1  g06881(new_n7155, new_n7258);
nor_1  g06882(new_n7158, new_n7258, new_n7259);
nor_1  g06883(new_n7259, new_n7257, new_n7260);
not_1  g06884(new_n7260, new_n7261);
not_1  g06885(new_n7149, new_n7262);
nand_1 g06886(new_n7262, new_n7142, new_n7263);
not_1  g06887(new_n7153, new_n7264);
nand_1 g06888(new_n7264, new_n7150, new_n7265_1);
nand_1 g06889(new_n7265_1, new_n7263, new_n7266);
nand_1 g06890(n11311, n9189, new_n7267);
nand_1 g06891(n7946, n4203, new_n7268);
nand_1 g06892(n4187, n2024, new_n7269);
xnor_1 g06893(new_n7269, new_n7268, new_n7270_1);
xnor_1 g06894(new_n7270_1, new_n7267, new_n7271);
not_1  g06895(new_n7271, new_n7272);
not_1  g06896(new_n7147, new_n7273);
nor_1  g06897(new_n7273, new_n7143, new_n7274);
not_1  g06898(new_n7274, new_n7275);
and_1  g06899(new_n7275, new_n7146, new_n7276);
not_1  g06900(new_n7276, new_n7277);
nand_1 g06901(new_n7277, new_n7272, new_n7278);
nand_1 g06902(new_n7276, new_n7271, new_n7279);
nand_1 g06903(new_n7279, new_n7278, new_n7280);
not_1  g06904(new_n7280, new_n7281);
nand_1 g06905(n12145, n9400, new_n7282);
nand_1 g06906(n2522, n2464, new_n7283);
xor_1  g06907(new_n7283, new_n7282, new_n7284);
not_1  g06908(new_n7284, new_n7285);
nand_1 g06909(new_n7285, new_n7281, new_n7286);
nand_1 g06910(new_n7284, new_n7280, new_n7287);
nand_1 g06911(new_n7287, new_n7286, new_n7288);
xnor_1 g06912(new_n7288, new_n7266, new_n7289);
xnor_1 g06913(new_n7289, new_n7261, new_n7290);
xnor_1 g06914(new_n7290, new_n7255, new_n7291);
xnor_1 g06915(new_n7291, new_n7160_1, new_n7292);
xnor_1 g06916(new_n7292, new_n7253, new_n7293);
nor_1  g06917(new_n1833, new_n5924, new_n7294_1);
not_1  g06918(new_n7294_1, new_n7295);
nor_1  g06919(new_n1866, new_n1219, new_n7296);
not_1  g06920(new_n7296, new_n7297);
nand_1 g06921(n9111, n5198, new_n7298);
nand_1 g06922(n9763, n1471, new_n7299);
xnor_1 g06923(new_n7299, new_n7298, new_n7300);
xnor_1 g06924(new_n7300, new_n7297, new_n7301);
not_1  g06925(new_n7301, new_n7302);
nand_1 g06926(new_n7213, new_n7212, new_n7303);
nand_1 g06927(new_n7216, new_n7303, new_n7304);
xnor_1 g06928(new_n7304, new_n7302, new_n7305);
nand_1 g06929(n7270, n3992, new_n7306);
nand_1 g06930(n8384, n806, new_n7307);
nand_1 g06931(new_n7307, new_n7306, new_n7308);
nor_1  g06932(new_n7307, new_n7306, new_n7309);
not_1  g06933(new_n7309, new_n7310);
nand_1 g06934(new_n7310, new_n7308, new_n7311);
xnor_1 g06935(new_n7311, new_n7305, new_n7312);
nor_1  g06936(new_n7220, new_n7208, new_n7313);
not_1  g06937(new_n7313, new_n7314);
xnor_1 g06938(new_n7314, new_n7312, new_n7315);
nor_1  g06939(new_n7201, new_n7198, new_n7316);
not_1  g06940(new_n7316, new_n7317);
nand_1 g06941(new_n7223, new_n7202, new_n7318);
nand_1 g06942(new_n7318, new_n7317, new_n7319);
nor_1  g06943(new_n7319, new_n7315, new_n7320_1);
not_1  g06944(new_n7320_1, new_n7321);
nand_1 g06945(new_n7319, new_n7315, new_n7322);
nand_1 g06946(new_n7322, new_n7321, new_n7323);
xnor_1 g06947(new_n7323, new_n7295, new_n7324);
xnor_1 g06948(new_n7324, new_n7226, new_n7325);
nor_1  g06949(new_n7196, new_n6433, new_n7326);
not_1  g06950(new_n7326, new_n7327);
nor_1  g06951(new_n5727, new_n1925, new_n7328);
not_1  g06952(new_n7328, new_n7329);
nor_1  g06953(new_n1244, new_n1959, new_n7330);
not_1  g06954(new_n7330, new_n7331);
nand_1 g06955(n6797, n2558, new_n7332);
nand_1 g06956(n6294, n2498, new_n7333);
xnor_1 g06957(new_n7333, new_n7332, new_n7334);
xnor_1 g06958(new_n7334, new_n7331, new_n7335);
not_1  g06959(new_n7335, new_n7336);
not_1  g06960(new_n7182, new_n7337);
nor_1  g06961(new_n7183, new_n7177, new_n7338);
nor_1  g06962(new_n7338, new_n7337, new_n7339);
nand_1 g06963(new_n7339, new_n7336, new_n7340);
not_1  g06964(new_n7340, new_n7341);
nor_1  g06965(new_n7339, new_n7336, new_n7342);
nor_1  g06966(new_n7342, new_n7341, new_n7343);
nand_1 g06967(n11478, n6016, new_n7344);
nand_1 g06968(n5283, n521, new_n7345);
nor_1  g06969(new_n7345, new_n7344, new_n7346);
not_1  g06970(new_n7346, new_n7347);
nand_1 g06971(new_n7345, new_n7344, new_n7348);
nand_1 g06972(new_n7348, new_n7347, new_n7349);
xnor_1 g06973(new_n7349, new_n7343, new_n7350);
nand_1 g06974(new_n7186, new_n7176, new_n7351);
nand_1 g06975(new_n7351, new_n7173, new_n7352);
xnor_1 g06976(new_n7352, new_n7350, new_n7353);
nor_1  g06977(new_n7191, new_n7188, new_n7354_1);
not_1  g06978(new_n7354_1, new_n7355);
nand_1 g06979(new_n7193_1, new_n7355, new_n7356);
xnor_1 g06980(new_n7356, new_n7353, new_n7357);
nand_1 g06981(new_n7357, new_n7329, new_n7358);
not_1  g06982(new_n7357, new_n7359);
nand_1 g06983(new_n7359, new_n7328, new_n7360);
nand_1 g06984(new_n7360, new_n7358, new_n7361);
xnor_1 g06985(new_n7361, new_n7327, new_n7362);
xnor_1 g06986(new_n7362, new_n7325, new_n7363);
nor_1  g06987(new_n7228, new_n7197, new_n7364);
not_1  g06988(new_n7364, new_n7365);
nand_1 g06989(new_n7235, new_n7365, new_n7366);
xnor_1 g06990(new_n7366, new_n7363, new_n7367);
nand_1 g06991(new_n7367, new_n7293, new_n7368);
not_1  g06992(new_n7253, new_n7369);
xnor_1 g06993(new_n7292, new_n7369, new_n7370);
not_1  g06994(new_n7367, new_n7371);
nand_1 g06995(new_n7371, new_n7370, new_n7372);
nand_1 g06996(new_n7372, new_n7368, new_n7373);
not_1  g06997(new_n7139, new_n7374);
xnor_1 g06998(new_n7249, new_n7374, new_n7375);
nand_1 g06999(new_n7375, new_n7373, new_n7376);
nand_1 g07000(new_n7376, new_n7250, new_n7377);
nand_1 g07001(new_n7377, new_n7138, new_n7378);
not_1  g07002(new_n7138, new_n7379);
xnor_1 g07003(new_n7377, new_n7379, new_n7380);
nor_1  g07004(new_n7289, new_n7260, new_n7381);
nand_1 g07005(new_n7270_1, new_n7267, new_n7382);
nand_1 g07006(new_n7278, new_n7382, new_n7383);
nor_1  g07007(new_n5615, new_n1735, new_n7384);
nand_1 g07008(n12145, n2464, new_n7385);
nand_1 g07009(n10217, n6877, new_n7386);
xnor_1 g07010(new_n7386, new_n7385, new_n7387);
xor_1  g07011(new_n7387, new_n7384, new_n7388_1);
xnor_1 g07012(new_n7388_1, new_n7383, new_n7389);
nor_1  g07013(new_n7269, new_n7268, new_n7390);
nor_1  g07014(new_n1747, new_n1278, new_n7391);
xor_1  g07015(new_n7391, new_n7390, new_n7392);
nor_1  g07016(new_n2119, new_n1192, new_n7393);
nor_1  g07017(new_n1199_1, new_n4769, new_n7394);
not_1  g07018(new_n7394, new_n7395);
nor_1  g07019(new_n2450, new_n1196, new_n7396);
not_1  g07020(new_n7396, new_n7397);
nand_1 g07021(new_n7397, new_n7395, new_n7398);
nand_1 g07022(new_n7396, new_n7394, new_n7399);
nand_1 g07023(new_n7399, new_n7398, new_n7400);
xnor_1 g07024(new_n7400, new_n7393, new_n7401);
xnor_1 g07025(new_n7401, new_n7392, new_n7402);
xnor_1 g07026(new_n7402, new_n7389, new_n7403);
nor_1  g07027(new_n7283, new_n7282, new_n7404);
not_1  g07028(new_n7286, new_n7405);
nor_1  g07029(new_n7405, new_n7266, new_n7406);
xnor_1 g07030(new_n7406, new_n7404, new_n7407);
nand_1 g07031(new_n7407, new_n7287, new_n7408);
xnor_1 g07032(new_n7408, new_n7403, new_n7409);
xnor_1 g07033(new_n7409, new_n7381, new_n7410);
nand_1 g07034(new_n7290, new_n7254, new_n7411);
nand_1 g07035(new_n7291, new_n7161, new_n7412);
nand_1 g07036(new_n7412, new_n7411, new_n7413);
xnor_1 g07037(new_n7413, new_n7410, new_n7414);
not_1  g07038(new_n7414, new_n7415);
nor_1  g07039(new_n7356, new_n7353, new_n7416);
nor_1  g07040(new_n1925, new_n5880, new_n7417);
nand_1 g07041(n6016, n5283, new_n7418);
nand_1 g07042(n11478, n5798, new_n7419);
xnor_1 g07043(new_n7419, new_n7418, new_n7420);
xor_1  g07044(new_n7420, new_n7417, new_n7421);
nor_1  g07045(new_n7334, new_n7331, new_n7422);
nor_1  g07046(new_n7341, new_n7422, new_n7423);
not_1  g07047(new_n7423, new_n7424);
xnor_1 g07048(new_n7424, new_n7421, new_n7425);
nor_1  g07049(new_n7333, new_n7332, new_n7426);
nor_1  g07050(new_n1310, new_n1959, new_n7427);
xor_1  g07051(new_n7427, new_n7426, new_n7428);
nor_1  g07052(new_n2205, new_n1235, new_n7429);
nand_1 g07053(n6294, n5579, new_n7430);
nand_1 g07054(n3146, n2558, new_n7431);
xnor_1 g07055(new_n7431, new_n7430, new_n7432);
xor_1  g07056(new_n7432, new_n7429, new_n7433);
xnor_1 g07057(new_n7433, new_n7428, new_n7434);
xnor_1 g07058(new_n7434, new_n7425, new_n7435);
not_1  g07059(new_n7349, new_n7436_1);
nand_1 g07060(new_n7436_1, new_n7343, new_n7437);
nand_1 g07061(new_n7352, new_n7350, new_n7438);
xnor_1 g07062(new_n7438, new_n7347, new_n7439);
nand_1 g07063(new_n7439, new_n7437, new_n7440);
xnor_1 g07064(new_n7440, new_n7435, new_n7441);
xnor_1 g07065(new_n7441, new_n7416, new_n7442);
nand_1 g07066(new_n7358, new_n7326, new_n7443);
nand_1 g07067(new_n7443, new_n7360, new_n7444);
xnor_1 g07068(new_n7444, new_n7442, new_n7445);
not_1  g07069(new_n7445, new_n7446);
not_1  g07070(new_n7311, new_n7447);
nand_1 g07071(new_n7447, new_n7305, new_n7448);
nand_1 g07072(new_n7314, new_n7312, new_n7449);
not_1  g07073(new_n7449, new_n7450);
nand_1 g07074(new_n7450, new_n7309, new_n7451);
nand_1 g07075(new_n7449, new_n7310, new_n7452);
nand_1 g07076(new_n7452, new_n7451, new_n7453);
nand_1 g07077(new_n7453, new_n7448, new_n7454);
nor_1  g07078(new_n7299, new_n7298, new_n7455);
nor_1  g07079(new_n1866, new_n1325, new_n7456_1);
xor_1  g07080(new_n7456_1, new_n7455, new_n7457);
nor_1  g07081(new_n1215, new_n2154, new_n7458);
nor_1  g07082(new_n4006, new_n1219, new_n7459);
not_1  g07083(new_n7459, new_n7460);
nor_1  g07084(new_n5696, new_n4009, new_n7461);
not_1  g07085(new_n7461, new_n7462);
nand_1 g07086(new_n7462, new_n7460, new_n7463);
nand_1 g07087(new_n7461, new_n7459, new_n7464);
nand_1 g07088(new_n7464, new_n7463, new_n7465);
xor_1  g07089(new_n7465, new_n7458, new_n7466);
xnor_1 g07090(new_n7466, new_n7457, new_n7467);
nor_1  g07091(new_n7300, new_n7297, new_n7468);
nor_1  g07092(new_n7304, new_n7301, new_n7469);
nor_1  g07093(new_n7469, new_n7468, new_n7470);
not_1  g07094(new_n7470, new_n7471);
nor_1  g07095(new_n5924, new_n1835_1, new_n7472);
nand_1 g07096(n8384, n7270, new_n7473);
nand_1 g07097(n7236, n2507, new_n7474);
xnor_1 g07098(new_n7474, new_n7473, new_n7475);
xor_1  g07099(new_n7475, new_n7472, new_n7476);
xnor_1 g07100(new_n7476, new_n7471, new_n7477);
xnor_1 g07101(new_n7477, new_n7467, new_n7478);
xnor_1 g07102(new_n7478, new_n7454, new_n7479);
xnor_1 g07103(new_n7479, new_n7320_1, new_n7480);
nand_1 g07104(new_n7323, new_n7295, new_n7481);
not_1  g07105(new_n7481, new_n7482);
nor_1  g07106(new_n7323, new_n7295, new_n7483);
nor_1  g07107(new_n7483, new_n7226, new_n7484);
nor_1  g07108(new_n7484, new_n7482, new_n7485);
xnor_1 g07109(new_n7485, new_n7480, new_n7486);
xnor_1 g07110(new_n7486, new_n7446, new_n7487);
not_1  g07111(new_n7325, new_n7488);
nand_1 g07112(new_n7362, new_n7488, new_n7489);
nand_1 g07113(new_n7366, new_n7363, new_n7490);
nand_1 g07114(new_n7490, new_n7489, new_n7491);
xnor_1 g07115(new_n7491, new_n7487, new_n7492);
xnor_1 g07116(new_n7492, new_n7415, new_n7493);
nand_1 g07117(new_n7292, new_n7369, new_n7494);
nand_1 g07118(new_n7368, new_n7494, new_n7495);
xnor_1 g07119(new_n7495, new_n7493, new_n7496);
nand_1 g07120(new_n7496, new_n7380, new_n7497);
nand_1 g07121(new_n7497, new_n7378, new_n7498);
nand_1 g07122(new_n7492, new_n7414, new_n7499);
nand_1 g07123(new_n7495, new_n7493, new_n7500_1);
nand_1 g07124(new_n7500_1, new_n7499, new_n7501);
nand_1 g07125(n4805, n1576, new_n7502);
or_1   g07126(new_n7438, new_n7347, new_n7503);
not_1  g07127(new_n7435, new_n7504);
nand_1 g07128(new_n7440, new_n7504, new_n7505);
nand_1 g07129(new_n7505, new_n7503, new_n7506);
xnor_1 g07130(new_n7506, new_n7502, new_n7507);
xnor_1 g07131(new_n7507, new_n7501, new_n7508);
nand_1 g07132(new_n7409, new_n7381, new_n7509);
not_1  g07133(new_n7410, new_n7510);
nand_1 g07134(new_n7413, new_n7510, new_n7511);
nand_1 g07135(new_n7511, new_n7509, new_n7512);
nand_1 g07136(new_n7479, new_n7320_1, new_n7513);
not_1  g07137(new_n7480, new_n7514);
nand_1 g07138(new_n7485, new_n7514, new_n7515);
nand_1 g07139(new_n7515, new_n7513, new_n7516);
nand_1 g07140(new_n7388_1, new_n7383, new_n7517);
not_1  g07141(new_n7389, new_n7518);
nand_1 g07142(new_n7402, new_n7518, new_n7519);
nand_1 g07143(new_n7519, new_n7517, new_n7520);
nand_1 g07144(n9189, n4203, new_n7521);
nand_1 g07145(n4187, n2522, new_n7522);
xnor_1 g07146(new_n7522, new_n7521, new_n7523_1);
nand_1 g07147(n9763, n4722, new_n7524);
nand_1 g07148(n10217, n9400, new_n7525);
xnor_1 g07149(new_n7525, new_n7524, new_n7526);
xnor_1 g07150(new_n7526, new_n7523_1, new_n7527);
nand_1 g07151(n9111, n7646, new_n7528);
nand_1 g07152(n12221, n2464, new_n7529);
nand_1 g07153(n12145, n11311, new_n7530);
xnor_1 g07154(new_n7530, new_n7529, new_n7531);
xnor_1 g07155(new_n7531, new_n7528, new_n7532);
xnor_1 g07156(new_n7532, new_n7527, new_n7533);
xnor_1 g07157(new_n7533, new_n7520, new_n7534);
xnor_1 g07158(new_n7534, new_n7516, new_n7535);
xnor_1 g07159(new_n7535, new_n7512, new_n7536);
nand_1 g07160(new_n7406, new_n7404, new_n7537);
not_1  g07161(new_n7403, new_n7538);
nand_1 g07162(new_n7408, new_n7538, new_n7539);
nand_1 g07163(new_n7539, new_n7537, new_n7540);
not_1  g07164(new_n7478, new_n7541);
nand_1 g07165(new_n7541, new_n7454, new_n7542);
nand_1 g07166(new_n7542, new_n7451, new_n7543);
xnor_1 g07167(new_n7543, new_n7540, new_n7544);
nand_1 g07168(n11821, n10223, new_n7545);
nand_1 g07169(n9080, n2879, new_n7546_1);
xnor_1 g07170(new_n7546_1, new_n7545, new_n7547);
nand_1 g07171(n11757, n9195, new_n7548);
nand_1 g07172(n7862, n2512, new_n7549);
xnor_1 g07173(new_n7549, new_n7548, new_n7550);
xnor_1 g07174(new_n7550, new_n7547, new_n7551);
and_1  g07175(new_n7099, new_n7095, new_n7552);
nor_1  g07176(new_n7552, new_n7098, new_n7553);
xnor_1 g07177(new_n7553, new_n7551, new_n7554);
nor_1  g07178(new_n2450, new_n1192, new_n7555);
nand_1 g07179(n3865, n1333, new_n7556);
nand_1 g07180(n5240, n4634, new_n7557);
xnor_1 g07181(new_n7557, new_n7556, new_n7558);
xnor_1 g07182(new_n7558, new_n7555, new_n7559);
xnor_1 g07183(new_n7559, new_n7554, new_n7560);
xnor_1 g07184(new_n7560, new_n7544, new_n7561);
nor_1  g07185(new_n7119, new_n7058, new_n7562);
nor_1  g07186(new_n7122, new_n7562, new_n7563);
nand_1 g07187(new_n7102, new_n7094, new_n7564);
not_1  g07188(new_n7103, new_n7565);
nand_1 g07189(new_n7115, new_n7565, new_n7566);
nand_1 g07190(new_n7566, new_n7564, new_n7567);
nand_1 g07191(new_n7391, new_n7390, new_n7568_1);
nand_1 g07192(new_n7401, new_n7392, new_n7569);
nand_1 g07193(new_n7569, new_n7568_1, new_n7570);
nand_1 g07194(n8384, n5153, new_n7571);
nor_1  g07195(new_n5685, new_n1866, new_n7572);
xnor_1 g07196(new_n7572, new_n7571, new_n7573);
nand_1 g07197(new_n7398, new_n7393, new_n7574);
nand_1 g07198(new_n7574, new_n7399, new_n7575);
xnor_1 g07199(new_n7575, new_n7573, new_n7576);
xnor_1 g07200(new_n7576, new_n7570, new_n7577);
xnor_1 g07201(new_n7577, new_n7567, new_n7578);
nand_1 g07202(n5198, n806, new_n7579);
nand_1 g07203(n3992, n2507, new_n7580);
xnor_1 g07204(new_n7580, new_n7579, new_n7581);
nand_1 g07205(n7823, n6877, new_n7582);
nand_1 g07206(n3342, n1471, new_n7583);
xnor_1 g07207(new_n7583, new_n7582, new_n7584);
xnor_1 g07208(new_n7584, new_n7581, new_n7585);
nand_1 g07209(new_n7463, new_n7458, new_n7586);
nand_1 g07210(new_n7586, new_n7464, new_n7587);
xnor_1 g07211(new_n7587, new_n7585, new_n7588);
xnor_1 g07212(new_n7588, new_n7578, new_n7589);
nand_1 g07213(new_n7476, new_n7470, new_n7590);
not_1  g07214(new_n7467, new_n7591);
nand_1 g07215(new_n7477, new_n7591, new_n7592);
nand_1 g07216(new_n7592, new_n7590, new_n7593);
nand_1 g07217(new_n7386, new_n7385, new_n7594);
not_1  g07218(new_n7594, new_n7595);
nor_1  g07219(new_n7387, new_n7384, new_n7596);
nor_1  g07220(new_n7596, new_n7595, new_n7597);
nand_1 g07221(n7236, n6431, new_n7598);
nand_1 g07222(n10174, n7946, new_n7599);
xnor_1 g07223(new_n7599, new_n7598, new_n7600);
xnor_1 g07224(new_n7600, new_n7597, new_n7601);
xnor_1 g07225(new_n7601, new_n7593, new_n7602);
xnor_1 g07226(new_n7602, new_n7589, new_n7603);
xnor_1 g07227(new_n7603, new_n7563, new_n7604);
xnor_1 g07228(new_n7604, new_n7561, new_n7605);
xnor_1 g07229(new_n7605, new_n7536, new_n7606);
not_1  g07230(new_n7486, new_n7607);
nand_1 g07231(new_n7607, new_n7446, new_n7608);
nand_1 g07232(new_n7491, new_n7487, new_n7609);
nand_1 g07233(new_n7609, new_n7608, new_n7610_1);
nand_1 g07234(new_n7124, new_n7127, new_n7611);
nand_1 g07235(new_n7137, new_n7125, new_n7612);
nand_1 g07236(new_n7612, new_n7611, new_n7613);
nand_1 g07237(new_n7441, new_n7416, new_n7614);
not_1  g07238(new_n7442, new_n7615);
nand_1 g07239(new_n7444, new_n7615, new_n7616);
nand_1 g07240(new_n7616, new_n7614, new_n7617);
nand_1 g07241(new_n7456_1, new_n7455, new_n7618);
not_1  g07242(new_n7466, new_n7619);
nand_1 g07243(new_n7619, new_n7457, new_n7620);
nand_1 g07244(new_n7620, new_n7618, new_n7621);
nand_1 g07245(new_n7427, new_n7426, new_n7622);
not_1  g07246(new_n7433, new_n7623);
nand_1 g07247(new_n7623, new_n7428, new_n7624);
nand_1 g07248(new_n7624, new_n7622, new_n7625);
xnor_1 g07249(new_n7625, new_n7621, new_n7626);
nand_1 g07250(new_n7114, new_n7108, new_n7627);
nand_1 g07251(new_n7627, new_n7106, new_n7628);
nand_1 g07252(n3172, n2253, new_n7629);
nand_1 g07253(n6797, n5579, new_n7630);
nand_1 g07254(n5798, n5283, new_n7631);
xnor_1 g07255(new_n7631, new_n7630, new_n7632);
xnor_1 g07256(new_n7632, new_n7629, new_n7633);
xnor_1 g07257(new_n7633, new_n7628, new_n7634);
nand_1 g07258(new_n7419, new_n7418, new_n7635);
not_1  g07259(new_n7635, new_n7636);
nor_1  g07260(new_n7420, new_n7417, new_n7637);
nor_1  g07261(new_n7637, new_n7636, new_n7638);
nand_1 g07262(new_n7431, new_n7430, new_n7639);
not_1  g07263(new_n7639, new_n7640);
nor_1  g07264(new_n7432, new_n7429, new_n7641);
nor_1  g07265(new_n7641, new_n7640, new_n7642);
xnor_1 g07266(new_n7642, new_n7638, new_n7643);
nand_1 g07267(n11478, n2347, new_n7644);
nand_1 g07268(n3146, n2498, new_n7645);
xnor_1 g07269(new_n7645, new_n7644, new_n7646_1);
xnor_1 g07270(new_n7646_1, new_n7643, new_n7647);
xnor_1 g07271(new_n7647, new_n7634, new_n7648);
xnor_1 g07272(new_n7648, new_n7626, new_n7649);
nand_1 g07273(new_n7423, new_n7421, new_n7650);
not_1  g07274(new_n7434, new_n7651);
nand_1 g07275(new_n7651, new_n7425, new_n7652);
nand_1 g07276(new_n7652, new_n7650, new_n7653);
nand_1 g07277(new_n7112, new_n7111, new_n7654);
not_1  g07278(new_n7654, new_n7655);
nor_1  g07279(new_n7113, new_n7110, new_n7656);
nor_1  g07280(new_n7656, new_n7655, new_n7657);
nand_1 g07281(n6016, n137, new_n7658);
nand_1 g07282(n7265, n6826, new_n7659);
nand_1 g07283(n6294, n521, new_n7660);
xnor_1 g07284(new_n7660, new_n7659, new_n7661);
xnor_1 g07285(new_n7661, new_n7658, new_n7662);
xnor_1 g07286(new_n7662, new_n7657, new_n7663);
not_1  g07287(n4938, new_n7664);
nor_1  g07288(new_n7664, new_n4615, new_n7665);
nand_1 g07289(new_n7474, new_n7473, new_n7666);
not_1  g07290(new_n7666, new_n7667);
nor_1  g07291(new_n7475, new_n7472, new_n7668);
nor_1  g07292(new_n7668, new_n7667, new_n7669);
xnor_1 g07293(new_n7669, new_n7665, new_n7670);
xnor_1 g07294(new_n7670, new_n7663, new_n7671);
xnor_1 g07295(new_n7671, new_n7653, new_n7672);
xnor_1 g07296(new_n7672, new_n7649, new_n7673);
xnor_1 g07297(new_n7673, new_n7617, new_n7674);
xnor_1 g07298(new_n7674, new_n7613, new_n7675);
xnor_1 g07299(new_n7675, new_n7610_1, new_n7676_1);
xnor_1 g07300(new_n7676_1, new_n7606, new_n7677);
xnor_1 g07301(new_n7677, new_n7508, new_n7678);
xnor_1 g07302(new_n7678, new_n7498, n2383);
xnor_1 g07303(new_n6270, new_n6263, n2425);
not_1  g07304(new_n3106, new_n7681);
xnor_1 g07305(new_n3152, new_n7681, n2431);
xnor_1 g07306(new_n2271, new_n2270, n2434);
xnor_1 g07307(new_n5292, new_n5289, n2581);
nor_1  g07308(new_n7020, new_n7018, new_n7685);
xnor_1 g07309(new_n7685, new_n7032, n2624);
nor_1  g07310(new_n2462, new_n4283, new_n7687);
not_1  g07311(new_n7687, new_n7688);
nand_1 g07312(n9920, n4921, new_n7689);
nand_1 g07313(n9956, n3627, new_n7690_1);
nand_1 g07314(new_n7690_1, new_n7689, new_n7691);
nor_1  g07315(new_n7690_1, new_n7689, new_n7692);
not_1  g07316(new_n7692, new_n7693);
nand_1 g07317(new_n7693, new_n7691, new_n7694);
xnor_1 g07318(new_n7694, new_n7688, new_n7695);
nand_1 g07319(new_n4318, new_n4271, new_n7696);
not_1  g07320(new_n7696, new_n7697);
nor_1  g07321(new_n4319, new_n4317, new_n7698);
nor_1  g07322(new_n7698, new_n7697, new_n7699);
xnor_1 g07323(new_n7699, new_n7695, new_n7700);
nor_1  g07324(new_n2481, new_n1377, new_n7701);
not_1  g07325(new_n7701, new_n7702);
nor_1  g07326(new_n1367, new_n2484, new_n7703);
not_1  g07327(new_n7703, new_n7704);
nor_1  g07328(new_n7704, new_n7702, new_n7705);
not_1  g07329(new_n7705, new_n7706);
nand_1 g07330(new_n7704, new_n7702, new_n7707);
nand_1 g07331(new_n7707, new_n7706, new_n7708);
xnor_1 g07332(new_n7708, new_n7700, new_n7709);
not_1  g07333(new_n7709, new_n7710);
nor_1  g07334(new_n4322, new_n4314, new_n7711);
nor_1  g07335(new_n7711, new_n7710, new_n7712);
not_1  g07336(new_n7712, new_n7713);
nand_1 g07337(new_n7711, new_n7710, new_n7714);
nand_1 g07338(new_n7714, new_n7713, new_n7715);
not_1  g07339(new_n7715, new_n7716);
nand_1 g07340(new_n4325, new_n4305, new_n7717);
nand_1 g07341(new_n7717, new_n7716, new_n7718);
nand_1 g07342(n6770, n3842, new_n7719);
xnor_1 g07343(new_n7719, new_n7692, new_n7720);
nor_1  g07344(new_n2476, new_n6617, new_n7721);
not_1  g07345(new_n7721, new_n7722);
nand_1 g07346(n11917, n9920, new_n7723);
nand_1 g07347(n9956, n4516, new_n7724);
xnor_1 g07348(new_n7724, new_n7723, new_n7725);
xnor_1 g07349(new_n7725, new_n7722, new_n7726);
xor_1  g07350(new_n7726, new_n7720, new_n7727);
and_1  g07351(new_n7694, new_n7688, new_n7728);
nor_1  g07352(new_n7699, new_n7695, new_n7729);
nor_1  g07353(new_n7729, new_n7728, new_n7730_1);
nor_1  g07354(new_n2551_1, new_n1377, new_n7731);
nand_1 g07355(n4189, n2577, new_n7732);
nand_1 g07356(n6687, n1835, new_n7733_1);
xnor_1 g07357(new_n7733_1, new_n7732, new_n7734);
xor_1  g07358(new_n7734, new_n7731, new_n7735);
xnor_1 g07359(new_n7735, new_n7730_1, new_n7736);
xnor_1 g07360(new_n7736, new_n7727, new_n7737);
not_1  g07361(new_n7737, new_n7738);
not_1  g07362(new_n7708, new_n7739);
nand_1 g07363(new_n7739, new_n7700, new_n7740);
nand_1 g07364(new_n7712, new_n7705, new_n7741);
nand_1 g07365(new_n7713, new_n7706, new_n7742);
nand_1 g07366(new_n7742, new_n7741, new_n7743);
nand_1 g07367(new_n7743, new_n7740, new_n7744);
xnor_1 g07368(new_n7744, new_n7738, new_n7745);
xnor_1 g07369(new_n7745, new_n7718, new_n7746);
nor_1  g07370(new_n2551_1, new_n378, new_n7747);
not_1  g07371(new_n7718, new_n7748);
nor_1  g07372(new_n7717, new_n7716, new_n7749);
nor_1  g07373(new_n7749, new_n7748, new_n7750);
nand_1 g07374(new_n7750, new_n7747, new_n7751);
not_1  g07375(new_n7747, new_n7752);
xnor_1 g07376(new_n7750, new_n7752, new_n7753);
nand_1 g07377(new_n7753, new_n4330, new_n7754);
nand_1 g07378(new_n7754, new_n7751, new_n7755);
xor_1  g07379(new_n7755, new_n7746, new_n7756);
nor_1  g07380(new_n2725, new_n4529, new_n7757);
not_1  g07381(new_n7757, new_n7758);
nand_1 g07382(n3602, n1094, new_n7759);
nand_1 g07383(n10678, n3719, new_n7760);
xnor_1 g07384(new_n7760, new_n7759, new_n7761);
nand_1 g07385(new_n7761, new_n7758, new_n7762);
not_1  g07386(new_n7762, new_n7763);
nor_1  g07387(new_n7761, new_n7758, new_n7764);
nor_1  g07388(new_n7764, new_n7763, new_n7765);
nand_1 g07389(new_n4531, new_n4342, new_n7766);
not_1  g07390(new_n7766, new_n7767);
nor_1  g07391(new_n4534, new_n7767, new_n7768);
xnor_1 g07392(new_n7768, new_n7765, new_n7769);
not_1  g07393(new_n7769, new_n7770);
nor_1  g07394(new_n1434, new_n2623, new_n7771);
not_1  g07395(new_n7771, new_n7772);
nor_1  g07396(new_n2626, new_n1508, new_n7773);
not_1  g07397(new_n7773, new_n7774);
nand_1 g07398(new_n7774, new_n7772, new_n7775);
nor_1  g07399(new_n7774, new_n7772, new_n7776);
not_1  g07400(new_n7776, new_n7777);
nand_1 g07401(new_n7777, new_n7775, new_n7778);
not_1  g07402(new_n7778, new_n7779);
nand_1 g07403(new_n7779, new_n7770, new_n7780);
nand_1 g07404(new_n7778, new_n7769, new_n7781);
nand_1 g07405(new_n7781, new_n7780, new_n7782);
nand_1 g07406(new_n4527, new_n4523, new_n7783);
not_1  g07407(new_n7783, new_n7784);
not_1  g07408(new_n4536, new_n7785);
nor_1  g07409(new_n7785, new_n4528, new_n7786);
nor_1  g07410(new_n7786, new_n7784, new_n7787);
nor_1  g07411(new_n7787, new_n7782, new_n7788);
not_1  g07412(new_n7788, new_n7789);
nand_1 g07413(new_n7787, new_n7782, new_n7790);
nand_1 g07414(new_n7790, new_n7789, new_n7791);
not_1  g07415(new_n7791, new_n7792);
nand_1 g07416(new_n4537, new_n4522, new_n7793);
nand_1 g07417(new_n7793, new_n4519, new_n7794);
nand_1 g07418(new_n7794, new_n7792, new_n7795);
not_1  g07419(new_n7795, new_n7796);
not_1  g07420(new_n7765, new_n7797);
nor_1  g07421(new_n7768, new_n7797, new_n7798);
nor_1  g07422(new_n7798, new_n7763, new_n7799);
nor_1  g07423(new_n1434, new_n2603, new_n7800);
nand_1 g07424(n10439, n6986, new_n7801);
nand_1 g07425(n10391, n8336, new_n7802);
xnor_1 g07426(new_n7802, new_n7801, new_n7803);
xor_1  g07427(new_n7803, new_n7800, new_n7804);
xnor_1 g07428(new_n7804, new_n7799, new_n7805);
nor_1  g07429(new_n7760, new_n7759, new_n7806);
nor_1  g07430(new_n2626, new_n4529, new_n7807);
xor_1  g07431(new_n7807, new_n7806, new_n7808);
nor_1  g07432(new_n6725, new_n2618, new_n7809);
nand_1 g07433(n6126, n1094, new_n7810);
nand_1 g07434(n7320, n3719, new_n7811);
xnor_1 g07435(new_n7811, new_n7810, new_n7812);
xnor_1 g07436(new_n7812, new_n7809, new_n7813);
xnor_1 g07437(new_n7813, new_n7808, new_n7814);
not_1  g07438(new_n7814, new_n7815);
xnor_1 g07439(new_n7815, new_n7805, new_n7816);
nand_1 g07440(new_n7788, new_n7776, new_n7817);
nand_1 g07441(new_n7789, new_n7777, new_n7818);
nand_1 g07442(new_n7818, new_n7817, new_n7819);
nand_1 g07443(new_n7819, new_n7780, new_n7820);
xnor_1 g07444(new_n7820, new_n7816, new_n7821);
xnor_1 g07445(new_n7821, new_n7796, new_n7822);
nand_1 g07446(n8336, n8065, new_n7823_1);
nor_1  g07447(new_n7794, new_n7792, new_n7824);
nor_1  g07448(new_n7824, new_n7796, new_n7825);
not_1  g07449(new_n7825, new_n7826);
nand_1 g07450(new_n7826, new_n7823_1, new_n7827);
nand_1 g07451(new_n4538, new_n4372, new_n7828);
xnor_1 g07452(new_n7825, new_n7823_1, new_n7829);
nand_1 g07453(new_n7829, new_n7828, new_n7830);
nand_1 g07454(new_n7830, new_n7827, new_n7831);
xnor_1 g07455(new_n7831, new_n7822, new_n7832);
not_1  g07456(new_n7832, new_n7833);
nand_1 g07457(n7160, n4826, new_n7834);
nand_1 g07458(n7733, n4828, new_n7835);
nand_1 g07459(n12925, n2515, new_n7836);
xnor_1 g07460(new_n7836, new_n7835, new_n7837);
nor_1  g07461(new_n7837, new_n7834, new_n7838);
not_1  g07462(new_n7838, new_n7839);
nand_1 g07463(new_n7837, new_n7834, new_n7840);
nand_1 g07464(new_n7840, new_n7839, new_n7841);
nand_1 g07465(new_n4579, new_n4380, new_n7842);
not_1  g07466(new_n7842, new_n7843);
nor_1  g07467(new_n4580, new_n4578, new_n7844);
nor_1  g07468(new_n7844, new_n7843, new_n7845);
xnor_1 g07469(new_n7845, new_n7841, new_n7846);
nor_1  g07470(new_n1452, new_n2767, new_n7847);
not_1  g07471(new_n7847, new_n7848);
nor_1  g07472(new_n4386, new_n2770, new_n7849);
not_1  g07473(new_n7849, new_n7850);
nand_1 g07474(new_n7850, new_n7848, new_n7851);
nor_1  g07475(new_n7850, new_n7848, new_n7852);
not_1  g07476(new_n7852, new_n7853);
nand_1 g07477(new_n7853, new_n7851, new_n7854);
xnor_1 g07478(new_n7854, new_n7846, new_n7855);
not_1  g07479(new_n4571, new_n7856);
nand_1 g07480(new_n4575, new_n7856, new_n7857);
nand_1 g07481(new_n4581, new_n4576, new_n7858);
nand_1 g07482(new_n7858, new_n7857, new_n7859);
xnor_1 g07483(new_n7859, new_n7855, new_n7860);
nand_1 g07484(new_n4589, new_n4583, new_n7861);
not_1  g07485(new_n7861, new_n7862_1);
nor_1  g07486(new_n7862_1, new_n7860, new_n7863);
not_1  g07487(new_n7863, new_n7864);
not_1  g07488(new_n7841, new_n7865);
nand_1 g07489(new_n7845, new_n7865, new_n7866);
nand_1 g07490(new_n7866, new_n7839, new_n7867);
nor_1  g07491(new_n1452, new_n2846, new_n7868);
nand_1 g07492(n7891, n4970, new_n7869);
nand_1 g07493(n12069, n10965, new_n7870);
xnor_1 g07494(new_n7870, new_n7869, new_n7871);
xor_1  g07495(new_n7871, new_n7868, new_n7872);
xnor_1 g07496(new_n7872, new_n7867, new_n7873);
nor_1  g07497(new_n7836, new_n7835, new_n7874);
nor_1  g07498(new_n2770, new_n1538, new_n7875);
xor_1  g07499(new_n7875, new_n7874, new_n7876);
nor_1  g07500(new_n2761, new_n6823, new_n7877);
nand_1 g07501(n4828, n4826, new_n7878);
nand_1 g07502(n12925, n1199, new_n7879);
xnor_1 g07503(new_n7879, new_n7878, new_n7880);
xor_1  g07504(new_n7880, new_n7877, new_n7881);
xnor_1 g07505(new_n7881, new_n7876, new_n7882);
xnor_1 g07506(new_n7882, new_n7873, new_n7883);
not_1  g07507(new_n7854, new_n7884);
nand_1 g07508(new_n7884, new_n7846, new_n7885);
nand_1 g07509(new_n7859, new_n7855, new_n7886);
xnor_1 g07510(new_n7886, new_n7852, new_n7887);
not_1  g07511(new_n7887, new_n7888);
nand_1 g07512(new_n7888, new_n7885, new_n7889);
xnor_1 g07513(new_n7889, new_n7883, new_n7890);
xnor_1 g07514(new_n7890, new_n7864, new_n7891_1);
nor_1  g07515(new_n1533, new_n2846, new_n7892);
xnor_1 g07516(new_n7861, new_n7860, new_n7893);
nand_1 g07517(new_n7893, new_n7892, new_n7894);
not_1  g07518(new_n7892, new_n7895);
xnor_1 g07519(new_n7893, new_n7895, new_n7896);
nand_1 g07520(new_n7896, new_n4594, new_n7897);
nand_1 g07521(new_n7897, new_n7894, new_n7898);
xnor_1 g07522(new_n7898, new_n7891_1, new_n7899);
nor_1  g07523(new_n385, new_n2980, new_n7900);
nor_1  g07524(new_n3772, new_n4542, new_n7901);
not_1  g07525(new_n7901, new_n7902);
nand_1 g07526(n5767, n405, new_n7903);
nand_1 g07527(n8433, n5319, new_n7904);
xnor_1 g07528(new_n7904, new_n7903, new_n7905);
nor_1  g07529(new_n7905, new_n7902, new_n7906);
not_1  g07530(new_n7906, new_n7907);
nand_1 g07531(new_n7905, new_n7902, new_n7908);
nand_1 g07532(new_n7908, new_n7907, new_n7909);
nor_1  g07533(new_n4549, new_n4543, new_n7910);
nor_1  g07534(new_n7910, new_n4548, new_n7911);
xnor_1 g07535(new_n7911, new_n7909, new_n7912);
nor_1  g07536(new_n1467, new_n2895, new_n7913);
not_1  g07537(new_n7913, new_n7914);
nor_1  g07538(new_n1562, new_n2898, new_n7915);
not_1  g07539(new_n7915, new_n7916);
nand_1 g07540(new_n7916, new_n7914, new_n7917);
nor_1  g07541(new_n7916, new_n7914, new_n7918);
not_1  g07542(new_n7918, new_n7919);
nand_1 g07543(new_n7919, new_n7917, new_n7920);
xnor_1 g07544(new_n7920, new_n7912, new_n7921);
nand_1 g07545(new_n4551, new_n4541, new_n7922);
not_1  g07546(new_n4552, new_n7923);
nand_1 g07547(new_n4555, new_n7923, new_n7924);
nand_1 g07548(new_n7924, new_n7922, new_n7925);
xnor_1 g07549(new_n7925, new_n7921, new_n7926);
nand_1 g07550(new_n4562, new_n4560, new_n7927);
nand_1 g07551(new_n7927, new_n4557, new_n7928);
xnor_1 g07552(new_n7928, new_n7926, new_n7929);
nand_1 g07553(new_n7929, new_n7900, new_n7930);
not_1  g07554(new_n7900, new_n7931);
xnor_1 g07555(new_n7929, new_n7931, new_n7932);
nand_1 g07556(new_n7932, new_n4565, new_n7933);
nand_1 g07557(new_n7933, new_n7930, new_n7934);
not_1  g07558(new_n7928, new_n7935);
nor_1  g07559(new_n7935, new_n7926, new_n7936);
nor_1  g07560(new_n7904, new_n7903, new_n7937);
nor_1  g07561(new_n4542, new_n2898, new_n7938);
xor_1  g07562(new_n7938, new_n7937, new_n7939);
nor_1  g07563(new_n6935, new_n2889, new_n7940);
nand_1 g07564(n5767, n4086, new_n7941);
nand_1 g07565(n9457, n8433, new_n7942);
xnor_1 g07566(new_n7942, new_n7941, new_n7943);
xnor_1 g07567(new_n7943, new_n7940, new_n7944);
not_1  g07568(new_n7944, new_n7945);
xnor_1 g07569(new_n7945, new_n7939, new_n7946_1);
nor_1  g07570(new_n1467, new_n2980, new_n7947);
nor_1  g07571(new_n2895, new_n1562, new_n7948);
nand_1 g07572(n11296, n11222, new_n7949);
xnor_1 g07573(new_n7949, new_n7948, new_n7950);
xnor_1 g07574(new_n7950, new_n7947, new_n7951);
not_1  g07575(new_n7909, new_n7952);
nand_1 g07576(new_n7911, new_n7952, new_n7953);
nand_1 g07577(new_n7953, new_n7907, new_n7954);
xnor_1 g07578(new_n7954, new_n7951, new_n7955);
xnor_1 g07579(new_n7955, new_n7946_1, new_n7956);
not_1  g07580(new_n7920, new_n7957);
nand_1 g07581(new_n7957, new_n7912, new_n7958);
nand_1 g07582(new_n7925, new_n7921, new_n7959);
xnor_1 g07583(new_n7959, new_n7919, new_n7960);
nand_1 g07584(new_n7960, new_n7958, new_n7961);
xnor_1 g07585(new_n7961, new_n7956, new_n7962);
xnor_1 g07586(new_n7962, new_n7936, new_n7963);
xnor_1 g07587(new_n7963, new_n7934, new_n7964);
not_1  g07588(new_n7964, new_n7965_1);
xnor_1 g07589(new_n7965_1, new_n7899, new_n7966_1);
xnor_1 g07590(new_n7896, new_n4594, new_n7967);
xnor_1 g07591(new_n7932, new_n4566, new_n7968);
not_1  g07592(new_n7968, new_n7969);
nand_1 g07593(new_n7969, new_n7967, new_n7970);
not_1  g07594(new_n4596, new_n7971);
nand_1 g07595(new_n4599, new_n7971, new_n7972);
nand_1 g07596(new_n4600, new_n4567, new_n7973);
nand_1 g07597(new_n7973, new_n7972, new_n7974);
xnor_1 g07598(new_n7968, new_n7967, new_n7975);
nand_1 g07599(new_n7975, new_n7974, new_n7976);
nand_1 g07600(new_n7976, new_n7970, new_n7977);
xnor_1 g07601(new_n7977, new_n7966_1, new_n7978);
xnor_1 g07602(new_n7978, new_n7833, new_n7979);
xnor_1 g07603(new_n7829, new_n7828, new_n7980);
not_1  g07604(new_n7980, new_n7981_1);
xnor_1 g07605(new_n7969, new_n7967, new_n7982);
xnor_1 g07606(new_n7982, new_n7974, new_n7983);
nand_1 g07607(new_n7983, new_n7981_1, new_n7984);
xnor_1 g07608(new_n7983, new_n7980, new_n7985);
not_1  g07609(new_n4539, new_n7986);
nor_1  g07610(new_n4601, new_n7986, new_n7987);
not_1  g07611(new_n4602, new_n7988);
nor_1  g07612(new_n4607, new_n7988, new_n7989);
nor_1  g07613(new_n7989, new_n7987, new_n7990);
nand_1 g07614(new_n7990, new_n7985, new_n7991);
nand_1 g07615(new_n7991, new_n7984, new_n7992);
xnor_1 g07616(new_n7992, new_n7979, new_n7993);
nand_1 g07617(new_n7993, new_n7756, new_n7994);
xnor_1 g07618(new_n7753, new_n4329, new_n7995);
not_1  g07619(new_n4515, new_n7996);
nand_1 g07620(new_n7996, new_n4332, new_n7997);
nand_1 g07621(new_n4608, new_n4516_1, new_n7998);
nand_1 g07622(new_n7998, new_n7997, new_n7999);
nor_1  g07623(new_n7999, new_n7995, new_n8000);
xnor_1 g07624(new_n7990, new_n7985, new_n8001);
xnor_1 g07625(new_n7999, new_n7995, new_n8002);
nor_1  g07626(new_n8002, new_n8001, new_n8003);
nor_1  g07627(new_n8003, new_n8000, new_n8004);
not_1  g07628(new_n7756, new_n8005);
xnor_1 g07629(new_n7993, new_n8005, new_n8006);
nand_1 g07630(new_n8006, new_n8004, new_n8007);
nand_1 g07631(new_n8007, new_n7994, new_n8008);
nor_1  g07632(new_n7886, new_n7853, new_n8009);
not_1  g07633(new_n7889, new_n8010);
nor_1  g07634(new_n8010, new_n7883, new_n8011);
nor_1  g07635(new_n8011, new_n8009, new_n8012);
nand_1 g07636(new_n7875, new_n7874, new_n8013);
not_1  g07637(new_n7881, new_n8014);
nand_1 g07638(new_n8014, new_n7876, new_n8015);
nand_1 g07639(new_n8015, new_n8013, new_n8016);
nand_1 g07640(new_n7733_1, new_n7732, new_n8017);
not_1  g07641(new_n8017, new_n8018);
nor_1  g07642(new_n7734, new_n7731, new_n8019);
nor_1  g07643(new_n8019, new_n8018, new_n8020);
nor_1  g07644(new_n4283, new_n2481, new_n8021);
xnor_1 g07645(new_n8021, new_n8020, new_n8022);
nand_1 g07646(n9637, n4189, new_n8023);
nand_1 g07647(n11917, n3627, new_n8024);
xnor_1 g07648(new_n8024, new_n8023, new_n8025);
xnor_1 g07649(new_n8025, new_n8022, new_n8026);
nand_1 g07650(new_n7870, new_n7869, new_n8027);
not_1  g07651(new_n8027, new_n8028_1);
nor_1  g07652(new_n7871, new_n7868, new_n8029);
nor_1  g07653(new_n8029, new_n8028_1, new_n8030);
nand_1 g07654(new_n7719, new_n7693, new_n8031);
nand_1 g07655(new_n7726, new_n7720, new_n8032);
nand_1 g07656(new_n8032, new_n8031, new_n8033);
xnor_1 g07657(new_n8033, new_n8030, new_n8034);
xnor_1 g07658(new_n8034, new_n8026, new_n8035);
xnor_1 g07659(new_n8035, new_n8016, new_n8036);
not_1  g07660(new_n7867, new_n8037);
nand_1 g07661(new_n7872, new_n8037, new_n8038);
not_1  g07662(new_n7882, new_n8039);
nand_1 g07663(new_n8039, new_n7873, new_n8040);
nand_1 g07664(new_n8040, new_n8038, new_n8041);
nand_1 g07665(new_n7811, new_n7810, new_n8042);
not_1  g07666(new_n8042, new_n8043);
nor_1  g07667(new_n7812, new_n7809, new_n8044);
nor_1  g07668(new_n8044, new_n8043, new_n8045);
nand_1 g07669(n7523, n3719, new_n8046);
nand_1 g07670(n11222, n1357, new_n8047);
xnor_1 g07671(new_n8047, new_n8046, new_n8048);
nand_1 g07672(n8336, n4190, new_n8049);
nand_1 g07673(n7320, n3602, new_n8050);
xnor_1 g07674(new_n8050, new_n8049, new_n8051);
xnor_1 g07675(new_n8051, new_n8048, new_n8052);
xnor_1 g07676(new_n8052, new_n8045, new_n8053);
xnor_1 g07677(new_n8053, new_n8041, new_n8054);
xnor_1 g07678(new_n8054, new_n8036, new_n8055);
nand_1 g07679(new_n7744, new_n7737, new_n8056);
nand_1 g07680(new_n8056, new_n7741, new_n8057);
not_1  g07681(new_n7816, new_n8058);
nand_1 g07682(new_n7820, new_n8058, new_n8059);
nand_1 g07683(new_n8059, new_n7817, new_n8060);
xnor_1 g07684(new_n8060, new_n8057, new_n8061);
xnor_1 g07685(new_n8061, new_n8055, new_n8062);
xnor_1 g07686(new_n8062, new_n8012, new_n8063);
and_1  g07687(new_n7821, new_n7796, new_n8064);
nor_1  g07688(new_n7831, new_n7822, new_n8065_1);
nor_1  g07689(new_n8065_1, new_n8064, new_n8066);
nand_1 g07690(new_n7802, new_n7801, new_n8067);
not_1  g07691(new_n8067, new_n8068);
nor_1  g07692(new_n7803, new_n7800, new_n8069);
nor_1  g07693(new_n8069, new_n8068, new_n8070);
nand_1 g07694(n5319, n4086, new_n8071);
nor_1  g07695(new_n1434, new_n3287_1, new_n8072);
xnor_1 g07696(new_n8072, new_n8071, new_n8073);
xnor_1 g07697(new_n8073, new_n8070, new_n8074);
xnor_1 g07698(new_n8074, new_n8066, new_n8075);
xnor_1 g07699(new_n8075, new_n8063, new_n8076);
nand_1 g07700(new_n7890, new_n7863, new_n8077);
nand_1 g07701(new_n7898, new_n7891_1, new_n8078);
nand_1 g07702(new_n8078, new_n8077, new_n8079);
and_1  g07703(new_n7962, new_n7936, new_n8080);
not_1  g07704(new_n7934, new_n8081);
nor_1  g07705(new_n7963, new_n8081, new_n8082);
nor_1  g07706(new_n8082, new_n8080, new_n8083);
xnor_1 g07707(new_n8083, new_n8079, new_n8084);
xnor_1 g07708(new_n8084, new_n8076, new_n8085);
nand_1 g07709(n4826, n2515, new_n8086);
not_1  g07710(n6578, new_n8087);
nor_1  g07711(new_n3969, new_n8087, new_n8088);
xnor_1 g07712(new_n8088, new_n8086, new_n8089);
nand_1 g07713(n6359, n5314, new_n8090);
nand_1 g07714(n12069, n7546, new_n8091);
xnor_1 g07715(new_n8091, new_n8090, new_n8092);
xnor_1 g07716(new_n8092, new_n8089, new_n8093);
nand_1 g07717(new_n7942, new_n7941, new_n8094);
not_1  g07718(new_n8094, new_n8095);
nor_1  g07719(new_n7943, new_n7940, new_n8096);
nor_1  g07720(new_n8096, new_n8095, new_n8097);
not_1  g07721(new_n7948, new_n8098);
not_1  g07722(new_n7950, new_n8099);
nor_1  g07723(new_n8099, new_n7947, new_n8100_1);
nor_1  g07724(new_n8100_1, new_n8098, new_n8101);
nor_1  g07725(new_n2969, new_n1467, new_n8102);
nand_1 g07726(new_n8102, new_n8101, new_n8103);
not_1  g07727(new_n8101, new_n8104);
nand_1 g07728(new_n8102, new_n7931, new_n8105);
nand_1 g07729(new_n8105, new_n8104, new_n8106);
nand_1 g07730(new_n8106, new_n8103, new_n8107);
xnor_1 g07731(new_n8107, new_n8097, new_n8108);
xnor_1 g07732(new_n8108, new_n8093, new_n8109);
xnor_1 g07733(new_n8109, new_n8085, new_n8110);
nand_1 g07734(new_n7978, new_n7832, new_n8111);
nand_1 g07735(new_n7992, new_n7979, new_n8112);
nand_1 g07736(new_n8112, new_n8111, new_n8113);
nand_1 g07737(new_n7965_1, new_n7899, new_n8114);
xnor_1 g07738(new_n7964, new_n7899, new_n8115);
nand_1 g07739(new_n7977, new_n8115, new_n8116);
nand_1 g07740(new_n8116, new_n8114, new_n8117);
nand_1 g07741(new_n7745, new_n7748, new_n8118);
nand_1 g07742(new_n7755, new_n7746, new_n8119);
nand_1 g07743(new_n8119, new_n8118, new_n8120);
nor_1  g07744(new_n7959, new_n7919, new_n8121);
not_1  g07745(new_n7961, new_n8122);
nor_1  g07746(new_n8122, new_n7956, new_n8123);
nor_1  g07747(new_n8123, new_n8121, new_n8124);
not_1  g07748(new_n7735, new_n8125);
nand_1 g07749(new_n8125, new_n7730_1, new_n8126);
not_1  g07750(new_n7727, new_n8127);
nand_1 g07751(new_n7736, new_n8127, new_n8128);
nand_1 g07752(new_n8128, new_n8126, new_n8129);
not_1  g07753(new_n7799, new_n8130);
nand_1 g07754(new_n7804, new_n8130, new_n8131);
nand_1 g07755(new_n7814, new_n7805, new_n8132);
nand_1 g07756(new_n8132, new_n8131, new_n8133);
xnor_1 g07757(new_n8133, new_n8129, new_n8134);
nand_1 g07758(new_n7938, new_n7937, new_n8135);
nand_1 g07759(new_n7944, new_n7939, new_n8136);
nand_1 g07760(new_n8136, new_n8135, new_n8137);
not_1  g07761(n1094, new_n8138_1);
nor_1  g07762(new_n2626, new_n8138_1, new_n8139);
nand_1 g07763(n2564, n1835, new_n8140);
xnor_1 g07764(new_n8140, new_n8139, new_n8141);
xnor_1 g07765(new_n8141, new_n8137, new_n8142);
nand_1 g07766(new_n7879, new_n7878, new_n8143);
not_1  g07767(new_n8143, new_n8144);
nor_1  g07768(new_n7880, new_n7877, new_n8145);
nor_1  g07769(new_n8145, new_n8144, new_n8146);
nand_1 g07770(n12391, n10965, new_n8147);
nand_1 g07771(n7891, n503, new_n8148);
nand_1 g07772(n9457, n405, new_n8149);
xnor_1 g07773(new_n8149, new_n8148, new_n8150);
xnor_1 g07774(new_n8150, new_n8147, new_n8151);
xnor_1 g07775(new_n8151, new_n8146, new_n8152);
nand_1 g07776(n8065, n6986, new_n8153);
nand_1 g07777(n10439, n2226, new_n8154);
xnor_1 g07778(new_n8154, new_n8153, new_n8155);
xnor_1 g07779(new_n8155, new_n8152, new_n8156);
xnor_1 g07780(new_n8156, new_n8142, new_n8157);
nand_1 g07781(new_n7724, new_n7723, new_n8158);
not_1  g07782(new_n8158, new_n8159);
nor_1  g07783(new_n7725, new_n7721, new_n8160);
nor_1  g07784(new_n8160, new_n8159, new_n8161);
nand_1 g07785(n11536, n6687, new_n8162);
nand_1 g07786(n6611, n996, new_n8163);
xnor_1 g07787(new_n8163, new_n8162, new_n8164);
nand_1 g07788(n4921, n4516, new_n8165);
nand_1 g07789(n9920, n3842, new_n8166);
xnor_1 g07790(new_n8166, new_n8165, new_n8167);
xnor_1 g07791(new_n8167, new_n8164, new_n8168);
xnor_1 g07792(new_n8168, new_n8161, new_n8169);
nand_1 g07793(n9956, n2087, new_n8170);
nand_1 g07794(n7733, n1199, new_n8171);
nand_1 g07795(n5767, n217, new_n8172);
xnor_1 g07796(new_n8172, new_n8171, new_n8173);
nand_1 g07797(n7160, n4970, new_n8174);
nand_1 g07798(n7610, n4828, new_n8175);
xnor_1 g07799(new_n8175, new_n8174, new_n8176);
xnor_1 g07800(new_n8176, new_n8173, new_n8177);
xnor_1 g07801(new_n8177, new_n8170, new_n8178);
xnor_1 g07802(new_n8178, new_n8169, new_n8179);
nand_1 g07803(new_n7807, new_n7806, new_n8180);
nand_1 g07804(new_n7813, new_n7808, new_n8181);
nand_1 g07805(new_n8181, new_n8180, new_n8182);
nand_1 g07806(n8433, n4817, new_n8183);
nor_1  g07807(new_n6725, new_n2725, new_n8184);
xnor_1 g07808(new_n8184, new_n8183, new_n8185);
xnor_1 g07809(new_n8185, new_n8182, new_n8186);
xnor_1 g07810(new_n8186, new_n8179, new_n8187);
xnor_1 g07811(new_n8187, new_n8157, new_n8188);
xnor_1 g07812(new_n8188, new_n8134, new_n8189);
xnor_1 g07813(new_n8189, new_n8124, new_n8190);
xnor_1 g07814(new_n8190, new_n8120, new_n8191);
xnor_1 g07815(new_n8191, new_n8117, new_n8192);
not_1  g07816(new_n7954, new_n8193);
nand_1 g07817(new_n8193, new_n7951, new_n8194);
not_1  g07818(new_n7946_1, new_n8195);
nand_1 g07819(new_n7955, new_n8195, new_n8196);
nand_1 g07820(new_n8196, new_n8194, new_n8197);
xnor_1 g07821(new_n8197, new_n8192, new_n8198);
xnor_1 g07822(new_n8198, new_n8113, new_n8199);
xnor_1 g07823(new_n8199, new_n8110, new_n8200);
xnor_1 g07824(new_n8200, new_n8008, n2679);
nor_1  g07825(new_n378, new_n5550, new_n8202_1);
nand_1 g07826(n10223, n6770, new_n8203);
nand_1 g07827(n9920, n2879, new_n8204);
nand_1 g07828(n7265, n3627, new_n8205);
nand_1 g07829(new_n8205, new_n8204, new_n8206);
nor_1  g07830(new_n8205, new_n8204, new_n8207);
not_1  g07831(new_n8207, new_n8208);
nand_1 g07832(new_n8208, new_n8206, new_n8209);
nor_1  g07833(new_n8209, new_n8203, new_n8210);
not_1  g07834(new_n8210, new_n8211);
nand_1 g07835(new_n8209, new_n8203, new_n8212);
nand_1 g07836(new_n8212, new_n8211, new_n8213);
nand_1 g07837(new_n5999, new_n5969, new_n8214);
not_1  g07838(new_n8214, new_n8215);
nor_1  g07839(new_n6000, new_n5997, new_n8216);
nor_1  g07840(new_n8216, new_n8215, new_n8217);
xnor_1 g07841(new_n8217, new_n8213, new_n8218);
nor_1  g07842(new_n5516, new_n1377, new_n8219);
not_1  g07843(new_n8219, new_n8220);
nor_1  g07844(new_n1121, new_n1367, new_n8221);
not_1  g07845(new_n8221, new_n8222);
nand_1 g07846(new_n8222, new_n8220, new_n8223);
nor_1  g07847(new_n8222, new_n8220, new_n8224);
not_1  g07848(new_n8224, new_n8225);
nand_1 g07849(new_n8225, new_n8223, new_n8226);
xnor_1 g07850(new_n8226, new_n8218, new_n8227);
not_1  g07851(new_n5996, new_n8228);
nor_1  g07852(new_n6001, new_n8228, new_n8229);
not_1  g07853(new_n8229, new_n8230);
nand_1 g07854(new_n6006, new_n6002, new_n8231);
nand_1 g07855(new_n8231, new_n8230, new_n8232);
xnor_1 g07856(new_n8232, new_n8227, new_n8233);
nand_1 g07857(new_n6017, new_n6008, new_n8234);
xnor_1 g07858(new_n8234, new_n8233, new_n8235);
xnor_1 g07859(new_n8235, new_n8202_1, new_n8236_1);
xnor_1 g07860(new_n8236_1, new_n6021, new_n8237);
not_1  g07861(new_n6024, new_n8238);
nand_1 g07862(new_n6250, new_n8238, new_n8239);
nand_1 g07863(new_n6276, new_n6251, new_n8240);
nand_1 g07864(new_n8240, new_n8239, new_n8241);
xnor_1 g07865(new_n8241, new_n8237, new_n8242);
nor_1  g07866(new_n6076, new_n6053, new_n8243);
nor_1  g07867(new_n5615, new_n382, new_n8244);
not_1  g07868(new_n8244, new_n8245);
nor_1  g07869(new_n1199_1, new_n4529, new_n8246);
nand_1 g07870(n2024, n1094, new_n8247);
nand_1 g07871(n10678, n7946, new_n8248);
nand_1 g07872(new_n8248, new_n8247, new_n8249);
nor_1  g07873(new_n8248, new_n8247, new_n8250);
not_1  g07874(new_n8250, new_n8251);
nand_1 g07875(new_n8251, new_n8249, new_n8252);
xnor_1 g07876(new_n8252, new_n8246, new_n8253);
nand_1 g07877(new_n6063, new_n6030, new_n8254);
not_1  g07878(new_n8254, new_n8255);
nor_1  g07879(new_n6064, new_n6061, new_n8256);
nor_1  g07880(new_n8256, new_n8255, new_n8257);
xnor_1 g07881(new_n8257, new_n8253, new_n8258);
nor_1  g07882(new_n5592, new_n1434, new_n8259);
not_1  g07883(new_n8259, new_n8260);
nor_1  g07884(new_n1508, new_n1278, new_n8261);
not_1  g07885(new_n8261, new_n8262);
nand_1 g07886(new_n8262, new_n8260, new_n8263);
nor_1  g07887(new_n8262, new_n8260, new_n8264);
not_1  g07888(new_n8264, new_n8265);
nand_1 g07889(new_n8265, new_n8263, new_n8266);
not_1  g07890(new_n8266, new_n8267);
xnor_1 g07891(new_n8267, new_n8258, new_n8268);
nand_1 g07892(new_n6059, new_n6056, new_n8269);
not_1  g07893(new_n8269, new_n8270);
nor_1  g07894(new_n6065, new_n6060, new_n8271);
nor_1  g07895(new_n8271, new_n8270, new_n8272);
not_1  g07896(new_n8272, new_n8273);
xnor_1 g07897(new_n8273, new_n8268, new_n8274);
not_1  g07898(new_n8274, new_n8275);
nand_1 g07899(new_n6075, new_n6071, new_n8276_1);
nand_1 g07900(new_n8276_1, new_n6068, new_n8277);
nand_1 g07901(new_n8277, new_n8275, new_n8278);
not_1  g07902(new_n8278, new_n8279);
nor_1  g07903(new_n8277, new_n8275, new_n8280);
nor_1  g07904(new_n8280, new_n8279, new_n8281);
xnor_1 g07905(new_n8281, new_n8245, new_n8282);
xnor_1 g07906(new_n8282, new_n8243, new_n8283);
not_1  g07907(new_n8283, new_n8284);
not_1  g07908(new_n6077, new_n8285);
nand_1 g07909(new_n6189, new_n8285, new_n8286);
nand_1 g07910(new_n6249, new_n6190, new_n8287);
nand_1 g07911(new_n8287, new_n8286, new_n8288);
xnor_1 g07912(new_n8288, new_n8284, new_n8289);
nand_1 g07913(new_n6212, new_n6191, new_n8290);
nor_1  g07914(new_n1533, new_n5727, new_n8291);
not_1  g07915(new_n8291, new_n8292);
nor_1  g07916(new_n1538, new_n1244, new_n8293);
nor_1  g07917(new_n6205, new_n6202, new_n8294);
nor_1  g07918(new_n8294, new_n6204, new_n8295);
nor_1  g07919(new_n8295, new_n8293, new_n8296);
not_1  g07920(new_n8293, new_n8297);
nor_1  g07921(new_n8295, new_n6094, new_n8298);
nor_1  g07922(new_n8298, new_n8297, new_n8299);
nor_1  g07923(new_n8299, new_n8296, new_n8300);
nand_1 g07924(n4828, n2498, new_n8301);
nand_1 g07925(n2558, n2515, new_n8302);
xnor_1 g07926(new_n8302, new_n8301, new_n8303_1);
xnor_1 g07927(new_n8303_1, new_n8300, new_n8304);
nor_1  g07928(new_n1452, new_n5658, new_n8305);
not_1  g07929(new_n8305, new_n8306);
nor_1  g07930(new_n4386, new_n1310, new_n8307);
not_1  g07931(new_n8307, new_n8308);
nand_1 g07932(new_n8308, new_n8306, new_n8309);
nor_1  g07933(new_n8308, new_n8306, new_n8310);
not_1  g07934(new_n8310, new_n8311);
nand_1 g07935(new_n8311, new_n8309, new_n8312);
xnor_1 g07936(new_n8312, new_n8304, new_n8313);
nand_1 g07937(new_n6207, new_n6201, new_n8314);
nand_1 g07938(new_n8314, new_n6198, new_n8315);
nand_1 g07939(new_n8315, new_n8313, new_n8316);
not_1  g07940(new_n8316, new_n8317);
nor_1  g07941(new_n8315, new_n8313, new_n8318);
nor_1  g07942(new_n8318, new_n8317, new_n8319);
nor_1  g07943(new_n6208, new_n6193, new_n8320);
not_1  g07944(new_n6211, new_n8321);
nor_1  g07945(new_n8321, new_n6209, new_n8322);
nor_1  g07946(new_n8322, new_n8320, new_n8323);
xnor_1 g07947(new_n8323, new_n8319, new_n8324);
xnor_1 g07948(new_n8324, new_n8292, new_n8325);
xnor_1 g07949(new_n8325, new_n8290, new_n8326);
nor_1  g07950(new_n385, new_n5924, new_n8327);
nor_1  g07951(new_n1219, new_n4542, new_n8328);
nand_1 g07952(n9111, n5767, new_n8329);
nand_1 g07953(n9763, n5319, new_n8330);
xnor_1 g07954(new_n8330, new_n8329, new_n8331);
xnor_1 g07955(new_n8331, new_n8328, new_n8332);
not_1  g07956(new_n6224, new_n8333);
nor_1  g07957(new_n6225, new_n6222, new_n8334);
nor_1  g07958(new_n8334, new_n8333, new_n8335);
nand_1 g07959(new_n8335, new_n8332, new_n8336_1);
not_1  g07960(new_n8336_1, new_n8337);
nor_1  g07961(new_n8335, new_n8332, new_n8338);
nor_1  g07962(new_n8338, new_n8337, new_n8339);
nand_1 g07963(n11153, n7270, new_n8340);
nand_1 g07964(n5314, n806, new_n8341);
nand_1 g07965(new_n8341, new_n8340, new_n8342);
nor_1  g07966(new_n8341, new_n8340, new_n8343);
not_1  g07967(new_n8343, new_n8344);
nand_1 g07968(new_n8344, new_n8342, new_n8345);
xnor_1 g07969(new_n8345, new_n8339, new_n8346);
nand_1 g07970(new_n6220, new_n6217, new_n8347);
not_1  g07971(new_n6221, new_n8348);
nand_1 g07972(new_n6228, new_n8348, new_n8349);
nand_1 g07973(new_n8349, new_n8347, new_n8350);
xnor_1 g07974(new_n8350, new_n8346, new_n8351);
not_1  g07975(new_n8351, new_n8352);
nand_1 g07976(new_n6237, new_n6230, new_n8353);
xnor_1 g07977(new_n8353, new_n8352, new_n8354);
xnor_1 g07978(new_n8354, new_n8327, new_n8355);
xnor_1 g07979(new_n8355, new_n6241, new_n8356);
xnor_1 g07980(new_n8356, new_n8326, new_n8357);
nor_1  g07981(new_n6243, new_n6214, new_n8358);
not_1  g07982(new_n6247, new_n8359);
nor_1  g07983(new_n8359, new_n6244, new_n8360);
nor_1  g07984(new_n8360, new_n8358, new_n8361);
nand_1 g07985(new_n8361, new_n8357, new_n8362);
not_1  g07986(new_n8357, new_n8363);
not_1  g07987(new_n8361, new_n8364);
nand_1 g07988(new_n8364, new_n8363, new_n8365);
nand_1 g07989(new_n8365, new_n8362, new_n8366);
nor_1  g07990(new_n8366, new_n8289, new_n8367);
not_1  g07991(new_n8367, new_n8368);
nand_1 g07992(new_n8366, new_n8289, new_n8369);
nand_1 g07993(new_n8369, new_n8368, new_n8370);
nor_1  g07994(new_n8370, new_n8242, new_n8371);
and_1  g07995(new_n8370, new_n8242, new_n8372);
nor_1  g07996(new_n8372, new_n8371, n2708);
xnor_1 g07997(new_n987, new_n984, n2818);
xnor_1 g07998(new_n2273, new_n2249, n2902);
nor_1  g07999(new_n1368, new_n456, new_n8376);
nor_1  g08000(new_n1402, new_n552, new_n8377);
nand_1 g08001(n12489, n5331, new_n8378);
nand_1 g08002(n10990, n7965, new_n8379);
nor_1  g08003(new_n8379, new_n8378, new_n8380);
not_1  g08004(new_n8380, new_n8381);
nand_1 g08005(new_n8379, new_n8378, new_n8382);
nand_1 g08006(new_n8382, new_n8381, new_n8383);
xnor_1 g08007(new_n8383, new_n8377, new_n8384_1);
nand_1 g08008(new_n8384_1, new_n8376, new_n8385);
not_1  g08009(new_n8385, new_n8386);
nor_1  g08010(new_n8384_1, new_n8376, new_n8387);
nor_1  g08011(new_n8387, new_n8386, n3071);
xnor_1 g08012(new_n3145, new_n3144, n3124);
nand_1 g08013(n11407, n5964, new_n8390);
nor_1  g08014(new_n456, new_n1378, new_n8391);
xnor_1 g08015(new_n8391, new_n8390, new_n8392);
not_1  g08016(new_n8392, new_n8393);
nand_1 g08017(new_n8393, new_n8385, new_n8394);
not_1  g08018(new_n8377, new_n8395);
nor_1  g08019(new_n8383, new_n8395, new_n8396);
nand_1 g08020(n11728, n8759, new_n8397);
nand_1 g08021(n12709, n6776, new_n8398_1);
xnor_1 g08022(new_n8398_1, new_n8397, new_n8399);
xnor_1 g08023(new_n8399, new_n8396, new_n8400);
nand_1 g08024(n7159, n5331, new_n8401);
nand_1 g08025(n12489, n8476, new_n8402);
xnor_1 g08026(new_n8402, new_n8401, new_n8403);
xnor_1 g08027(new_n8403, new_n8380, new_n8404);
nand_1 g08028(n7965, n5760, new_n8405);
nand_1 g08029(n10990, n7388, new_n8406);
xnor_1 g08030(new_n8406, new_n8405, new_n8407);
xnor_1 g08031(new_n8407, new_n8404, new_n8408);
xnor_1 g08032(new_n8408, new_n8400, new_n8409);
xnor_1 g08033(new_n8392, new_n8385, new_n8410);
nand_1 g08034(new_n8410, new_n8409, new_n8411);
nand_1 g08035(new_n8411, new_n8394, new_n8412);
nor_1  g08036(new_n424, new_n1378, new_n8413);
not_1  g08037(new_n8413, new_n8414);
nor_1  g08038(new_n8414, new_n8376, new_n8415);
nor_1  g08039(new_n1368, new_n419, new_n8416);
not_1  g08040(new_n8416, new_n8417);
nor_1  g08041(new_n1371, new_n456, new_n8418);
not_1  g08042(new_n8418, new_n8419);
nand_1 g08043(new_n8419, new_n8417, new_n8420);
not_1  g08044(new_n8420, new_n8421);
nor_1  g08045(new_n8419, new_n8417, new_n8422);
nor_1  g08046(new_n8422, new_n8421, new_n8423);
nor_1  g08047(new_n8423, new_n8415, new_n8424);
not_1  g08048(new_n8424, new_n8425);
nand_1 g08049(new_n8420, new_n8415, new_n8426);
nand_1 g08050(new_n8426, new_n8425, new_n8427);
xnor_1 g08051(new_n8427, new_n8412, new_n8428);
not_1  g08052(new_n8396, new_n8429);
nor_1  g08053(new_n8399, new_n8429, new_n8430);
not_1  g08054(new_n8430, new_n8431);
nand_1 g08055(new_n8408, new_n8400, new_n8432);
nand_1 g08056(new_n8432, new_n8431, new_n8433_1);
not_1  g08057(new_n8433_1, new_n8434);
nor_1  g08058(new_n1435, new_n563, new_n8435);
not_1  g08059(new_n8435, new_n8436);
nor_1  g08060(new_n8436, new_n8377, new_n8437);
nand_1 g08061(n12709, n12299, new_n8438);
nand_1 g08062(n8759, n6429, new_n8439);
nand_1 g08063(new_n8439, new_n8438, new_n8440);
not_1  g08064(new_n8440, new_n8441);
nor_1  g08065(new_n8439, new_n8438, new_n8442);
nor_1  g08066(new_n8442, new_n8441, new_n8443);
nor_1  g08067(new_n8443, new_n8437, new_n8444);
not_1  g08068(new_n8444, new_n8445);
nand_1 g08069(new_n8440, new_n8437, new_n8446);
nand_1 g08070(new_n8446, new_n8445, new_n8447);
xnor_1 g08071(new_n8447, new_n8434, new_n8448);
nand_1 g08072(n8476, n7159, new_n8449);
not_1  g08073(new_n8449, new_n8450);
nand_1 g08074(new_n8450, new_n8378, new_n8451);
not_1  g08075(new_n8451, new_n8452);
nand_1 g08076(n12489, n2530, new_n8453);
nand_1 g08077(n12777, n5331, new_n8454);
nand_1 g08078(new_n8454, new_n8453, new_n8455);
not_1  g08079(new_n8455, new_n8456);
nand_1 g08080(n12777, n2530, new_n8457);
nor_1  g08081(new_n8457, new_n8378, new_n8458);
nor_1  g08082(new_n8458, new_n8456, new_n8459);
nor_1  g08083(new_n8459, new_n8452, new_n8460);
nor_1  g08084(new_n8456, new_n8451, new_n8461);
nor_1  g08085(new_n8461, new_n8460, new_n8462);
nand_1 g08086(n7388, n5760, new_n8463);
not_1  g08087(new_n8463, new_n8464);
nand_1 g08088(new_n8464, new_n8379, new_n8465);
not_1  g08089(n10990, new_n8466);
nor_1  g08090(new_n762, new_n8466, new_n8467);
not_1  g08091(new_n8467, new_n8468);
not_1  g08092(n1478, new_n8469);
nor_1  g08093(new_n754, new_n8469, new_n8470);
not_1  g08094(new_n8470, new_n8471);
nand_1 g08095(new_n8471, new_n8468, new_n8472);
nor_1  g08096(new_n8471, new_n8468, new_n8473);
not_1  g08097(new_n8473, new_n8474);
nand_1 g08098(new_n8474, new_n8472, new_n8475);
nand_1 g08099(new_n8475, new_n8465, new_n8476_1);
not_1  g08100(new_n8465, new_n8477);
nand_1 g08101(new_n8472, new_n8477, new_n8478);
nand_1 g08102(new_n8478, new_n8476_1, new_n8479);
xnor_1 g08103(new_n8479, new_n8462, new_n8480);
nand_1 g08104(new_n8403, new_n8381, new_n8481);
nand_1 g08105(new_n8407, new_n8404, new_n8482);
nand_1 g08106(new_n8482, new_n8481, new_n8483);
xnor_1 g08107(new_n8483, new_n8480, new_n8484);
xnor_1 g08108(new_n8484, new_n8448, new_n8485);
xnor_1 g08109(new_n8485, new_n8428, n3214);
xnor_1 g08110(new_n5831, new_n5830, n3230);
not_1  g08111(new_n5254, new_n8488);
xnor_1 g08112(new_n5304, new_n8488, n3272);
nor_1  g08113(new_n424, new_n1365, new_n8490);
nand_1 g08114(n11407, n4312, new_n8491);
nand_1 g08115(n11877, n5964, new_n8492);
nand_1 g08116(new_n8492, new_n8491, new_n8493);
not_1  g08117(new_n8493, new_n8494);
nor_1  g08118(new_n8492, new_n8491, new_n8495);
nor_1  g08119(new_n1378, new_n419, new_n8496);
nor_1  g08120(new_n8496, new_n8495, new_n8497);
nor_1  g08121(new_n8497, new_n8494, new_n8498);
nand_1 g08122(new_n8498, new_n8490, new_n8499);
xnor_1 g08123(new_n8498, new_n8490, new_n8500);
not_1  g08124(new_n8500, new_n8501);
nor_1  g08125(new_n1378, new_n395, new_n8502);
nor_1  g08126(new_n1371, new_n419, new_n8503);
not_1  g08127(new_n8503, new_n8504);
not_1  g08128(n12705, new_n8505);
nor_1  g08129(new_n8505, new_n1368, new_n8506);
not_1  g08130(new_n8506, new_n8507);
nand_1 g08131(new_n8507, new_n8504, new_n8508);
nor_1  g08132(new_n8507, new_n8504, new_n8509);
not_1  g08133(new_n8509, new_n8510);
nand_1 g08134(new_n8510, new_n8508, new_n8511);
xnor_1 g08135(new_n8511, new_n8502, new_n8512);
nand_1 g08136(new_n8512, new_n8501, new_n8513);
nand_1 g08137(new_n8513, new_n8499, new_n8514);
not_1  g08138(n5320, new_n8515);
nor_1  g08139(new_n424, new_n8515, new_n8516);
not_1  g08140(new_n8516, new_n8517);
nor_1  g08141(new_n1365, new_n419, new_n8518);
xnor_1 g08142(new_n8518, new_n8517, new_n8519);
xnor_1 g08143(new_n8519, new_n8514, new_n8520);
nor_1  g08144(new_n1371, new_n395, new_n8521);
nand_1 g08145(n12705, n5212, new_n8522);
nand_1 g08146(n12025, n11407, new_n8523);
xnor_1 g08147(new_n8523, new_n8522, new_n8524);
xnor_1 g08148(new_n8524, new_n8521, new_n8525);
not_1  g08149(new_n8508, new_n8526);
nor_1  g08150(new_n8509, new_n8502, new_n8527);
nor_1  g08151(new_n8527, new_n8526, new_n8528);
xnor_1 g08152(new_n8528, new_n8525, new_n8529);
nor_1  g08153(new_n8529, new_n8520, new_n8530);
not_1  g08154(new_n8530, new_n8531);
nand_1 g08155(new_n8529, new_n8520, new_n8532);
nand_1 g08156(new_n8532, new_n8531, new_n8533);
nor_1  g08157(new_n8515, new_n456, new_n8534);
xnor_1 g08158(new_n8512, new_n8500, new_n8535);
nor_1  g08159(new_n8535, new_n8534, new_n8536);
not_1  g08160(new_n8536, new_n8537);
nand_1 g08161(new_n8535, new_n8534, new_n8538);
nand_1 g08162(new_n8538, new_n8537, new_n8539);
not_1  g08163(new_n8539, new_n8540);
nor_1  g08164(new_n456, new_n1365, new_n8541);
nor_1  g08165(new_n8422, new_n8413, new_n8542);
nor_1  g08166(new_n8542, new_n8421, new_n8543);
nand_1 g08167(new_n8543, new_n8541, new_n8544);
not_1  g08168(new_n8544, new_n8545);
nor_1  g08169(new_n8543, new_n8541, new_n8546);
nor_1  g08170(new_n8546, new_n8545, new_n8547);
not_1  g08171(new_n8547, new_n8548);
nor_1  g08172(new_n8495, new_n8494, new_n8549);
xnor_1 g08173(new_n8549, new_n8496, new_n8550);
nor_1  g08174(new_n8550, new_n8548, new_n8551);
nor_1  g08175(new_n8551, new_n8545, new_n8552);
nand_1 g08176(new_n8552, new_n8540, new_n8553);
nand_1 g08177(new_n8553, new_n8537, new_n8554);
nor_1  g08178(new_n8554, new_n8533, new_n8555);
not_1  g08179(new_n8521, new_n8556);
nand_1 g08180(new_n8524, new_n8556, new_n8557);
not_1  g08181(new_n8528, new_n8558);
nand_1 g08182(new_n8558, new_n8525, new_n8559);
nand_1 g08183(new_n8559, new_n8557, new_n8560);
not_1  g08184(n12000, new_n8561);
nor_1  g08185(new_n8561, new_n424, new_n8562);
nand_1 g08186(n5320, n1097, new_n8563);
nand_1 g08187(n9725, n5305, new_n8564);
xnor_1 g08188(new_n8564, new_n8563, new_n8565);
xnor_1 g08189(new_n8565, new_n8562, new_n8566);
xnor_1 g08190(new_n8566, new_n8560, new_n8567);
nor_1  g08191(new_n8523, new_n8522, new_n8568);
nor_1  g08192(new_n1365, new_n395, new_n8569);
xnor_1 g08193(new_n8569, new_n8568, new_n8570);
nor_1  g08194(new_n511, new_n1378, new_n8571);
nand_1 g08195(n12705, n11877, new_n8572);
nand_1 g08196(n11407, n11257, new_n8573);
xnor_1 g08197(new_n8573, new_n8572, new_n8574);
xor_1  g08198(new_n8574, new_n8571, new_n8575);
xnor_1 g08199(new_n8575, new_n8570, new_n8576);
xnor_1 g08200(new_n8576, new_n8567, new_n8577);
not_1  g08201(new_n8577, new_n8578);
nand_1 g08202(new_n8519, new_n8514, new_n8579);
not_1  g08203(new_n8518, new_n8580);
nor_1  g08204(new_n8580, new_n8517, new_n8581);
xnor_1 g08205(new_n8530, new_n8581, new_n8582);
nand_1 g08206(new_n8582, new_n8579, new_n8583);
xnor_1 g08207(new_n8583, new_n8578, new_n8584);
xnor_1 g08208(new_n8584, new_n8555, new_n8585);
nor_1  g08209(new_n8561, new_n456, new_n8586);
not_1  g08210(new_n8533, new_n8587);
xnor_1 g08211(new_n8554, new_n8587, new_n8588);
nand_1 g08212(new_n8588, new_n8586, new_n8589);
xnor_1 g08213(new_n8550, new_n8547, new_n8590);
nor_1  g08214(new_n8425, new_n8414, new_n8591);
and_1  g08215(new_n8591, new_n8590, new_n8592);
xnor_1 g08216(new_n8552, new_n8539, new_n8593);
not_1  g08217(new_n8593, new_n8594);
nand_1 g08218(new_n8594, new_n8592, new_n8595_1);
not_1  g08219(new_n8595_1, new_n8596);
not_1  g08220(new_n8586, new_n8597);
xnor_1 g08221(new_n8588, new_n8597, new_n8598);
nand_1 g08222(new_n8598, new_n8596, new_n8599);
nand_1 g08223(new_n8599, new_n8589, new_n8600);
xnor_1 g08224(new_n8600, new_n8585, new_n8601);
not_1  g08225(n8717, new_n8602);
nor_1  g08226(new_n552, new_n8602, new_n8603);
nand_1 g08227(n7436, n6429, new_n8604);
nand_1 g08228(n12709, n9241, new_n8605);
nand_1 g08229(n11728, n8276, new_n8606);
xnor_1 g08230(new_n8606, new_n8605, new_n8607);
xnor_1 g08231(new_n8607, new_n8604, new_n8608);
not_1  g08232(new_n8608, new_n8609);
nand_1 g08233(n12299, n6429, new_n8610);
nand_1 g08234(n12709, n8276, new_n8611);
nand_1 g08235(new_n8611, new_n8610, new_n8612);
not_1  g08236(new_n8612, new_n8613);
nor_1  g08237(new_n8611, new_n8610, new_n8614);
nor_1  g08238(new_n1435, new_n599, new_n8615);
nor_1  g08239(new_n8615, new_n8614, new_n8616);
nor_1  g08240(new_n8616, new_n8613, new_n8617);
not_1  g08241(new_n8617, new_n8618);
nand_1 g08242(new_n8618, new_n8609, new_n8619);
nand_1 g08243(new_n8617, new_n8608, new_n8620);
nand_1 g08244(new_n8620, new_n8619, new_n8621);
not_1  g08245(n2433, new_n8622);
nor_1  g08246(new_n563, new_n8622, new_n8623);
not_1  g08247(new_n8623, new_n8624);
nor_1  g08248(new_n554, new_n1506, new_n8625);
not_1  g08249(new_n8625, new_n8626);
nor_1  g08250(new_n8626, new_n8624, new_n8627);
not_1  g08251(new_n8627, new_n8628);
nand_1 g08252(new_n8626, new_n8624, new_n8629);
nand_1 g08253(new_n8629, new_n8628, new_n8630);
xnor_1 g08254(new_n8630, new_n8621, new_n8631);
nand_1 g08255(n8819, n6776, new_n8632);
not_1  g08256(new_n8632, new_n8633);
nand_1 g08257(n12709, n7436, new_n8634);
nand_1 g08258(n6776, n6429, new_n8635);
nand_1 g08259(new_n8635, new_n8634, new_n8636);
not_1  g08260(new_n8636, new_n8637);
nor_1  g08261(new_n8635, new_n8634, new_n8638);
nor_1  g08262(new_n554, new_n1435, new_n8639);
nor_1  g08263(new_n8639, new_n8638, new_n8640);
nor_1  g08264(new_n8640, new_n8637, new_n8641);
nand_1 g08265(new_n8641, new_n8633, new_n8642);
not_1  g08266(new_n8642, new_n8643);
xnor_1 g08267(new_n8641, new_n8633, new_n8644);
not_1  g08268(new_n8615, new_n8645);
xnor_1 g08269(new_n8611, new_n8610, new_n8646);
xnor_1 g08270(new_n8646, new_n8645, new_n8647);
nor_1  g08271(new_n8647, new_n8644, new_n8648);
nor_1  g08272(new_n8648, new_n8643, new_n8649);
not_1  g08273(new_n8649, new_n8650);
nand_1 g08274(new_n8650, new_n8631, new_n8651);
not_1  g08275(new_n8651, new_n8652);
nor_1  g08276(new_n8650, new_n8631, new_n8653);
nor_1  g08277(new_n8653, new_n8652, new_n8654);
nor_1  g08278(new_n552, new_n8622, new_n8655);
not_1  g08279(new_n8655, new_n8656);
xnor_1 g08280(new_n8647, new_n8644, new_n8657);
nand_1 g08281(new_n8657, new_n8656, new_n8658);
xnor_1 g08282(new_n8657, new_n8655, new_n8659);
nor_1  g08283(new_n1506, new_n552, new_n8660);
nor_1  g08284(new_n8442, new_n8435, new_n8661);
nor_1  g08285(new_n8661, new_n8441, new_n8662);
nand_1 g08286(new_n8662, new_n8660, new_n8663);
not_1  g08287(new_n8663, new_n8664);
xnor_1 g08288(new_n8662, new_n8660, new_n8665_1);
nor_1  g08289(new_n8638, new_n8637, new_n8666);
xnor_1 g08290(new_n8666, new_n8639, new_n8667);
nor_1  g08291(new_n8667, new_n8665_1, new_n8668);
nor_1  g08292(new_n8668, new_n8664, new_n8669);
nand_1 g08293(new_n8669, new_n8659, new_n8670);
nand_1 g08294(new_n8670, new_n8658, new_n8671);
not_1  g08295(new_n8671, new_n8672);
nand_1 g08296(new_n8672, new_n8654, new_n8673);
not_1  g08297(new_n8673, new_n8674);
nor_1  g08298(new_n8672, new_n8654, new_n8675);
nor_1  g08299(new_n8675, new_n8674, new_n8676);
nand_1 g08300(new_n8676, new_n8603, new_n8677);
xnor_1 g08301(new_n8667, new_n8665_1, new_n8678);
nor_1  g08302(new_n8445, new_n8436, new_n8679);
not_1  g08303(new_n8679, new_n8680);
nor_1  g08304(new_n8680, new_n8678, new_n8681);
xnor_1 g08305(new_n8669, new_n8659, new_n8682);
nand_1 g08306(new_n8682, new_n8681, new_n8683);
not_1  g08307(new_n8683, new_n8684);
not_1  g08308(new_n8603, new_n8685);
xnor_1 g08309(new_n8676, new_n8685, new_n8686);
nand_1 g08310(new_n8686, new_n8684, new_n8687);
nand_1 g08311(new_n8687, new_n8677, new_n8688);
nand_1 g08312(new_n8607, new_n8604, new_n8689);
nand_1 g08313(new_n8619, new_n8689, new_n8690);
nor_1  g08314(new_n8602, new_n563, new_n8691);
nor_1  g08315(new_n554, new_n8622, new_n8692);
nand_1 g08316(n8759, n7730, new_n8693);
not_1  g08317(new_n8693, new_n8694);
nand_1 g08318(new_n8694, new_n8692, new_n8695);
not_1  g08319(new_n8692, new_n8696);
nand_1 g08320(new_n8693, new_n8696, new_n8697);
nand_1 g08321(new_n8697, new_n8695, new_n8698);
xnor_1 g08322(new_n8698, new_n8691, new_n8699);
xnor_1 g08323(new_n8699, new_n8690, new_n8700);
nor_1  g08324(new_n8606, new_n8605, new_n8701);
nor_1  g08325(new_n1506, new_n599, new_n8702);
xor_1  g08326(new_n8702, new_n8701, new_n8703);
nor_1  g08327(new_n1435, new_n2723, new_n8704);
nand_1 g08328(n8276, n6429, new_n8705);
nand_1 g08329(n12709, n10510, new_n8706);
xnor_1 g08330(new_n8706, new_n8705, new_n8707);
xor_1  g08331(new_n8707, new_n8704, new_n8708);
xnor_1 g08332(new_n8708, new_n8703, new_n8709);
xnor_1 g08333(new_n8709, new_n8700, new_n8710);
not_1  g08334(new_n8630, new_n8711);
nand_1 g08335(new_n8711, new_n8621, new_n8712);
nand_1 g08336(new_n8652, new_n8627, new_n8713);
nand_1 g08337(new_n8651, new_n8628, new_n8714);
nand_1 g08338(new_n8714, new_n8713, new_n8715);
nand_1 g08339(new_n8715, new_n8712, new_n8716);
xnor_1 g08340(new_n8716, new_n8710, new_n8717_1);
xnor_1 g08341(new_n8717_1, new_n8673, new_n8718);
xnor_1 g08342(new_n8718, new_n8688, new_n8719);
nor_1  g08343(new_n767, new_n8469, new_n8720);
not_1  g08344(new_n8720, new_n8721);
nand_1 g08345(n5860, n5760, new_n8722);
nand_1 g08346(n10990, n3986, new_n8723);
xnor_1 g08347(new_n8723, new_n8722, new_n8724);
xnor_1 g08348(new_n8724, new_n8721, new_n8725);
not_1  g08349(new_n8725, new_n8726);
nor_1  g08350(new_n762, new_n8469, new_n8727);
not_1  g08351(new_n8727, new_n8728);
nor_1  g08352(new_n8466, new_n802, new_n8729);
not_1  g08353(new_n8729, new_n8730);
nand_1 g08354(new_n8730, new_n8728, new_n8731);
not_1  g08355(new_n8731, new_n8732);
nor_1  g08356(new_n8730, new_n8728, new_n8733);
nor_1  g08357(new_n1466, new_n767, new_n8734);
nor_1  g08358(new_n8734, new_n8733, new_n8735);
nor_1  g08359(new_n8735, new_n8732, new_n8736);
nand_1 g08360(new_n8736, new_n8726, new_n8737);
not_1  g08361(new_n8737, new_n8738);
nor_1  g08362(new_n8736, new_n8726, new_n8739);
nor_1  g08363(new_n8739, new_n8738, new_n8740);
nand_1 g08364(n12947, n7388, new_n8741);
nand_1 g08365(n11892, n11791, new_n8742);
nand_1 g08366(new_n8742, new_n8741, new_n8743);
nor_1  g08367(new_n8742, new_n8741, new_n8744);
not_1  g08368(new_n8744, new_n8745);
nand_1 g08369(new_n8745, new_n8743, new_n8746);
xnor_1 g08370(new_n8746, new_n8740, new_n8747);
not_1  g08371(n11791, new_n8748);
nor_1  g08372(new_n8748, new_n696, new_n8749);
nand_1 g08373(n10990, n2393, new_n8750);
nand_1 g08374(n7388, n1478, new_n8751);
nand_1 g08375(new_n8751, new_n8750, new_n8752);
not_1  g08376(new_n8752, new_n8753);
nor_1  g08377(new_n8751, new_n8750, new_n8754);
nor_1  g08378(new_n762, new_n1466, new_n8755);
nor_1  g08379(new_n8755, new_n8754, new_n8756);
nor_1  g08380(new_n8756, new_n8753, new_n8757);
nand_1 g08381(new_n8757, new_n8749, new_n8758);
not_1  g08382(new_n8758, new_n8759_1);
nor_1  g08383(new_n8757, new_n8749, new_n8760);
nor_1  g08384(new_n8760, new_n8759_1, new_n8761);
not_1  g08385(new_n8733, new_n8762);
nand_1 g08386(new_n8762, new_n8731, new_n8763);
xnor_1 g08387(new_n8763, new_n8734, new_n8764);
nand_1 g08388(new_n8764, new_n8761, new_n8765);
nand_1 g08389(new_n8765, new_n8758, new_n8766);
xnor_1 g08390(new_n8766, new_n8747, new_n8767);
not_1  g08391(n12947, new_n8768);
nor_1  g08392(new_n8768, new_n754, new_n8769);
nor_1  g08393(new_n8748, new_n754, new_n8770);
not_1  g08394(new_n8472, new_n8771);
nor_1  g08395(new_n8473, new_n8464, new_n8772);
nor_1  g08396(new_n8772, new_n8771, new_n8773);
nand_1 g08397(new_n8773, new_n8770, new_n8774);
not_1  g08398(new_n8774, new_n8775);
nor_1  g08399(new_n8773, new_n8770, new_n8776);
nor_1  g08400(new_n8776, new_n8775, new_n8777);
not_1  g08401(new_n8754, new_n8778);
nand_1 g08402(new_n8778, new_n8752, new_n8779);
xnor_1 g08403(new_n8779, new_n8755, new_n8780);
nand_1 g08404(new_n8780, new_n8777, new_n8781);
nand_1 g08405(new_n8781, new_n8774, new_n8782);
nor_1  g08406(new_n8782, new_n8769, new_n8783);
not_1  g08407(new_n8783, new_n8784);
xnor_1 g08408(new_n8764, new_n8761, new_n8785);
not_1  g08409(new_n8769, new_n8786);
xnor_1 g08410(new_n8782, new_n8786, new_n8787);
nand_1 g08411(new_n8787, new_n8785, new_n8788);
nand_1 g08412(new_n8788, new_n8784, new_n8789);
nor_1  g08413(new_n8789, new_n8767, new_n8790);
nor_1  g08414(new_n8723, new_n8722, new_n8791);
nor_1  g08415(new_n8748, new_n767, new_n8792);
xnor_1 g08416(new_n8792, new_n8791, new_n8793);
nor_1  g08417(new_n1466, new_n1084, new_n8794);
nand_1 g08418(n5860, n1478, new_n8795);
nand_1 g08419(n10990, n5857, new_n8796);
nand_1 g08420(new_n8796, new_n8795, new_n8797);
not_1  g08421(new_n8797, new_n8798);
nor_1  g08422(new_n8796, new_n8795, new_n8799);
nor_1  g08423(new_n8799, new_n8798, new_n8800);
xnor_1 g08424(new_n8800, new_n8794, new_n8801);
xnor_1 g08425(new_n8801, new_n8793, new_n8802);
not_1  g08426(new_n8802, new_n8803);
not_1  g08427(n6441, new_n8804);
nor_1  g08428(new_n696, new_n8804, new_n8805);
nand_1 g08429(n12947, n11892, new_n8806);
not_1  g08430(new_n8806, new_n8807);
nand_1 g08431(n11999, n7965, new_n8808);
xnor_1 g08432(new_n8808, new_n8807, new_n8809);
xnor_1 g08433(new_n8809, new_n8805, new_n8810);
nor_1  g08434(new_n8724, new_n8721, new_n8811);
nor_1  g08435(new_n8738, new_n8811, new_n8812);
not_1  g08436(new_n8812, new_n8813);
xnor_1 g08437(new_n8813, new_n8810, new_n8814);
xnor_1 g08438(new_n8814, new_n8803, new_n8815);
not_1  g08439(new_n8746, new_n8816);
nand_1 g08440(new_n8816, new_n8740, new_n8817);
nand_1 g08441(new_n8766, new_n8747, new_n8818);
not_1  g08442(new_n8818, new_n8819_1);
nand_1 g08443(new_n8819_1, new_n8744, new_n8820);
nand_1 g08444(new_n8818, new_n8745, new_n8821);
nand_1 g08445(new_n8821, new_n8820, new_n8822);
nand_1 g08446(new_n8822, new_n8817, new_n8823);
xnor_1 g08447(new_n8823, new_n8815, new_n8824);
xnor_1 g08448(new_n8824, new_n8790, new_n8825);
nor_1  g08449(new_n754, new_n8804, new_n8826);
xnor_1 g08450(new_n8789, new_n8767, new_n8827);
not_1  g08451(new_n8827, new_n8828);
nand_1 g08452(new_n8828, new_n8826, new_n8829);
not_1  g08453(new_n8826, new_n8830);
nand_1 g08454(new_n8827, new_n8830, new_n8831);
xnor_1 g08455(new_n8780, new_n8777, new_n8832);
nor_1  g08456(new_n8476_1, new_n8463, new_n8833);
not_1  g08457(new_n8833, new_n8834);
nor_1  g08458(new_n8834, new_n8832, new_n8835);
xnor_1 g08459(new_n8787, new_n8785, new_n8836);
nand_1 g08460(new_n8836, new_n8835, new_n8837);
not_1  g08461(new_n8837, new_n8838);
nand_1 g08462(new_n8838, new_n8831, new_n8839);
nand_1 g08463(new_n8839, new_n8829, new_n8840);
xnor_1 g08464(new_n8840, new_n8825, new_n8841);
not_1  g08465(new_n8841, new_n8842);
not_1  g08466(n12777, new_n8843);
nor_1  g08467(new_n8843, new_n829, new_n8844);
not_1  g08468(new_n8844, new_n8845);
nand_1 g08469(n10545, n7159, new_n8846);
nand_1 g08470(n12489, n7690, new_n8847);
xnor_1 g08471(new_n8847, new_n8846, new_n8848);
xnor_1 g08472(new_n8848, new_n8845, new_n8849);
not_1  g08473(new_n8849, new_n8850);
nand_1 g08474(n12489, n10545, new_n8851);
nand_1 g08475(new_n8851, new_n8457, new_n8852);
not_1  g08476(new_n8852, new_n8853);
nor_1  g08477(new_n8851, new_n8457, new_n8854);
nor_1  g08478(new_n829, new_n1451, new_n8855);
nor_1  g08479(new_n8855, new_n8854, new_n8856);
nor_1  g08480(new_n8856, new_n8853, new_n8857);
nand_1 g08481(new_n8857, new_n8850, new_n8858);
not_1  g08482(new_n8858, new_n8859);
nor_1  g08483(new_n8857, new_n8850, new_n8860);
nor_1  g08484(new_n8860, new_n8859, new_n8861);
nand_1 g08485(n6254, n2530, new_n8862);
nand_1 g08486(n11967, n8476, new_n8863);
nand_1 g08487(new_n8863, new_n8862, new_n8864);
nor_1  g08488(new_n8863, new_n8862, new_n8865);
not_1  g08489(new_n8865, new_n8866);
nand_1 g08490(new_n8866, new_n8864, new_n8867);
xnor_1 g08491(new_n8867, new_n8861, new_n8868);
nor_1  g08492(new_n712, new_n1532, new_n8869);
nand_1 g08493(n12648, n12489, new_n8870);
nand_1 g08494(n12777, n8476, new_n8871);
nand_1 g08495(new_n8871, new_n8870, new_n8872);
not_1  g08496(new_n8872, new_n8873);
nor_1  g08497(new_n8871, new_n8870, new_n8874);
nor_1  g08498(new_n1451, new_n740, new_n8875);
nor_1  g08499(new_n8875, new_n8874, new_n8876);
nor_1  g08500(new_n8876, new_n8873, new_n8877);
nand_1 g08501(new_n8877, new_n8869, new_n8878);
not_1  g08502(new_n8878, new_n8879);
nor_1  g08503(new_n8877, new_n8869, new_n8880);
nor_1  g08504(new_n8880, new_n8879, new_n8881);
not_1  g08505(new_n8854, new_n8882);
nand_1 g08506(new_n8882, new_n8852, new_n8883);
xnor_1 g08507(new_n8883, new_n8855, new_n8884);
nand_1 g08508(new_n8884, new_n8881, new_n8885);
nand_1 g08509(new_n8885, new_n8878, new_n8886);
xnor_1 g08510(new_n8886, new_n8868, new_n8887);
not_1  g08511(n11967, new_n8888);
nor_1  g08512(new_n8888, new_n668, new_n8889);
not_1  g08513(new_n8889, new_n8890);
xnor_1 g08514(new_n8884, new_n8881, new_n8891);
nand_1 g08515(new_n8891, new_n8890, new_n8892);
xnor_1 g08516(new_n8891, new_n8889, new_n8893);
nor_1  g08517(new_n1532, new_n668, new_n8894);
nor_1  g08518(new_n8458, new_n8450, new_n8895);
nor_1  g08519(new_n8895, new_n8456, new_n8896);
nand_1 g08520(new_n8896, new_n8894, new_n8897);
not_1  g08521(new_n8897, new_n8898);
nor_1  g08522(new_n8896, new_n8894, new_n8899);
nor_1  g08523(new_n8899, new_n8898, new_n8900);
not_1  g08524(new_n8900, new_n8901);
not_1  g08525(new_n8874, new_n8902);
nand_1 g08526(new_n8902, new_n8872, new_n8903);
xnor_1 g08527(new_n8903, new_n8875, new_n8904);
not_1  g08528(new_n8904, new_n8905);
nor_1  g08529(new_n8905, new_n8901, new_n8906);
nor_1  g08530(new_n8906, new_n8898, new_n8907);
nand_1 g08531(new_n8907, new_n8893, new_n8908);
nand_1 g08532(new_n8908, new_n8892, new_n8909);
nor_1  g08533(new_n8909, new_n8887, new_n8910);
not_1  g08534(n1353, new_n8911);
nor_1  g08535(new_n668, new_n8911, new_n8912);
nand_1 g08536(n11967, n2530, new_n8913);
nand_1 g08537(n8476, n447, new_n8914);
xnor_1 g08538(new_n8914, new_n8913, new_n8915);
xor_1  g08539(new_n8915, new_n8912, new_n8916);
nor_1  g08540(new_n8848, new_n8845, new_n8917);
nor_1  g08541(new_n8859, new_n8917, new_n8918);
not_1  g08542(new_n8918, new_n8919);
xnor_1 g08543(new_n8919, new_n8916, new_n8920);
nor_1  g08544(new_n8847, new_n8846, new_n8921);
nor_1  g08545(new_n829, new_n1532, new_n8922);
xor_1  g08546(new_n8922, new_n8921, new_n8923);
nor_1  g08547(new_n1048, new_n1451, new_n8924);
nand_1 g08548(n12777, n10545, new_n8925);
nand_1 g08549(n12489, n3616, new_n8926);
xnor_1 g08550(new_n8926, new_n8925, new_n8927);
xnor_1 g08551(new_n8927, new_n8924, new_n8928);
not_1  g08552(new_n8928, new_n8929);
xnor_1 g08553(new_n8929, new_n8923, new_n8930);
xnor_1 g08554(new_n8930, new_n8920, new_n8931);
not_1  g08555(new_n8867, new_n8932);
nand_1 g08556(new_n8932, new_n8861, new_n8933);
nand_1 g08557(new_n8886, new_n8868, new_n8934);
not_1  g08558(new_n8934, new_n8935);
nand_1 g08559(new_n8935, new_n8865, new_n8936);
nand_1 g08560(new_n8934, new_n8866, new_n8937);
nand_1 g08561(new_n8937, new_n8936, new_n8938);
nand_1 g08562(new_n8938, new_n8933, new_n8939);
xnor_1 g08563(new_n8939, new_n8931, new_n8940);
xnor_1 g08564(new_n8940, new_n8910, new_n8941);
not_1  g08565(n447, new_n8942);
nor_1  g08566(new_n668, new_n8942, new_n8943);
xnor_1 g08567(new_n8909, new_n8887, new_n8944);
not_1  g08568(new_n8944, new_n8945);
nand_1 g08569(new_n8945, new_n8943, new_n8946);
not_1  g08570(new_n8943, new_n8947);
nand_1 g08571(new_n8944, new_n8947, new_n8948);
nor_1  g08572(new_n8904, new_n8900, new_n8949);
nor_1  g08573(new_n8949, new_n8906, new_n8950);
not_1  g08574(new_n8950, new_n8951);
nand_1 g08575(new_n8460, new_n8450, new_n8952);
nor_1  g08576(new_n8952, new_n8951, new_n8953);
not_1  g08577(new_n8953, new_n8954);
xnor_1 g08578(new_n8907, new_n8893, new_n8955);
not_1  g08579(new_n8955, new_n8956);
nor_1  g08580(new_n8956, new_n8954, new_n8957);
nand_1 g08581(new_n8957, new_n8948, new_n8958);
nand_1 g08582(new_n8958, new_n8946, new_n8959);
xnor_1 g08583(new_n8959, new_n8941, new_n8960);
not_1  g08584(new_n8960, new_n8961);
nand_1 g08585(new_n8961, new_n8842, new_n8962);
nand_1 g08586(new_n8960, new_n8841, new_n8963);
nand_1 g08587(new_n8963, new_n8962, new_n8964);
nand_1 g08588(new_n8831, new_n8829, new_n8965);
xnor_1 g08589(new_n8965, new_n8837, new_n8966);
nand_1 g08590(new_n8948, new_n8946, new_n8967);
xnor_1 g08591(new_n8967, new_n8957, new_n8968);
not_1  g08592(new_n8968, new_n8969);
nand_1 g08593(new_n8969, new_n8966, new_n8970);
xnor_1 g08594(new_n8955, new_n8953, new_n8971);
nor_1  g08595(new_n8836, new_n8835, new_n8972);
nor_1  g08596(new_n8972, new_n8838, new_n8973);
not_1  g08597(new_n8973, new_n8974);
nand_1 g08598(new_n8974, new_n8971, new_n8975);
xnor_1 g08599(new_n8973, new_n8971, new_n8976);
xnor_1 g08600(new_n8952, new_n8950, new_n8977);
xnor_1 g08601(new_n8833, new_n8832, new_n8978);
and_1  g08602(new_n8978, new_n8977, new_n8979);
not_1  g08603(new_n8462, new_n8980);
nor_1  g08604(new_n8479, new_n8980, new_n8981);
not_1  g08605(new_n8480, new_n8982);
nor_1  g08606(new_n8483, new_n8982, new_n8983);
nor_1  g08607(new_n8983, new_n8981, new_n8984);
xnor_1 g08608(new_n8978, new_n8977, new_n8985);
nor_1  g08609(new_n8985, new_n8984, new_n8986);
nor_1  g08610(new_n8986, new_n8979, new_n8987);
nand_1 g08611(new_n8987, new_n8976, new_n8988);
nand_1 g08612(new_n8988, new_n8975, new_n8989);
xnor_1 g08613(new_n8968, new_n8966, new_n8990);
nand_1 g08614(new_n8990, new_n8989, new_n8991);
nand_1 g08615(new_n8991, new_n8970, new_n8992);
xnor_1 g08616(new_n8992, new_n8964, new_n8993);
xnor_1 g08617(new_n8993, new_n8719, new_n8994);
xnor_1 g08618(new_n8686, new_n8683, new_n8995);
not_1  g08619(new_n8995, new_n8996);
not_1  g08620(new_n8990, new_n8997);
xnor_1 g08621(new_n8997, new_n8989, new_n8998);
nand_1 g08622(new_n8998, new_n8996, new_n8999);
xnor_1 g08623(new_n8998, new_n8995, new_n9000);
nor_1  g08624(new_n8682, new_n8681, new_n9001);
nor_1  g08625(new_n9001, new_n8684, new_n9002);
not_1  g08626(new_n9002, new_n9003);
not_1  g08627(new_n8976, new_n9004);
xnor_1 g08628(new_n8987, new_n9004, new_n9005);
nor_1  g08629(new_n9005, new_n9003, new_n9006);
xnor_1 g08630(new_n8679, new_n8678, new_n9007);
not_1  g08631(new_n9007, new_n9008);
xnor_1 g08632(new_n8985, new_n8984, new_n9009);
nor_1  g08633(new_n9009, new_n9008, new_n9010);
xnor_1 g08634(new_n9009, new_n9007, new_n9011);
not_1  g08635(new_n9011, new_n9012);
nor_1  g08636(new_n8447, new_n8434, new_n9013);
not_1  g08637(new_n8484, new_n9014);
nor_1  g08638(new_n9014, new_n8448, new_n9015);
nor_1  g08639(new_n9015, new_n9013, new_n9016);
nor_1  g08640(new_n9016, new_n9012, new_n9017);
nor_1  g08641(new_n9017, new_n9010, new_n9018);
xnor_1 g08642(new_n9005, new_n9002, new_n9019);
not_1  g08643(new_n9019, new_n9020);
nor_1  g08644(new_n9020, new_n9018, new_n9021);
nor_1  g08645(new_n9021, new_n9006, new_n9022);
nand_1 g08646(new_n9022, new_n9000, new_n9023);
nand_1 g08647(new_n9023, new_n8999, new_n9024);
xnor_1 g08648(new_n9024, new_n8994, new_n9025);
not_1  g08649(new_n9025, new_n9026);
nand_1 g08650(new_n9026, new_n8601, new_n9027);
xnor_1 g08651(new_n9025, new_n8601, new_n9028);
xnor_1 g08652(new_n8598, new_n8595_1, new_n9029);
not_1  g08653(new_n9029, new_n9030);
xnor_1 g08654(new_n8998, new_n8996, new_n9031);
xnor_1 g08655(new_n9022, new_n9031, new_n9032);
nand_1 g08656(new_n9032, new_n9030, new_n9033);
not_1  g08657(new_n9033, new_n9034);
xnor_1 g08658(new_n9032, new_n9030, new_n9035);
nor_1  g08659(new_n8594, new_n8592, new_n9036);
nor_1  g08660(new_n9036, new_n8596, new_n9037);
xnor_1 g08661(new_n9019, new_n9018, new_n9038);
nor_1  g08662(new_n9038, new_n9037, new_n9039);
xnor_1 g08663(new_n9038, new_n9037, new_n9040);
nor_1  g08664(new_n8591, new_n8590, new_n9041);
nor_1  g08665(new_n9041, new_n8592, new_n9042);
xnor_1 g08666(new_n9016, new_n9011, new_n9043);
nor_1  g08667(new_n9043, new_n9042, new_n9044);
nor_1  g08668(new_n8427, new_n8412, new_n9045);
not_1  g08669(new_n8485, new_n9046);
nor_1  g08670(new_n9046, new_n8428, new_n9047);
nor_1  g08671(new_n9047, new_n9045, new_n9048);
not_1  g08672(new_n9048, new_n9049);
xnor_1 g08673(new_n9043, new_n9042, new_n9050);
nor_1  g08674(new_n9050, new_n9049, new_n9051);
nor_1  g08675(new_n9051, new_n9044, new_n9052);
nor_1  g08676(new_n9052, new_n9040, new_n9053);
nor_1  g08677(new_n9053, new_n9039, new_n9054);
nor_1  g08678(new_n9054, new_n9035, new_n9055);
nor_1  g08679(new_n9055, new_n9034, new_n9056);
nand_1 g08680(new_n9056, new_n9028, new_n9057);
nand_1 g08681(new_n9057, new_n9027, new_n9058);
nand_1 g08682(new_n8993, new_n8719, new_n9059);
not_1  g08683(new_n8994, new_n9060);
nand_1 g08684(new_n9024, new_n9060, new_n9061);
nand_1 g08685(new_n9061, new_n9059, new_n9062);
nand_1 g08686(new_n8584, new_n8555, new_n9063);
not_1  g08687(new_n8585, new_n9064);
nand_1 g08688(new_n8600, new_n9064, new_n9065);
nand_1 g08689(new_n9065, new_n9063, new_n9066);
nand_1 g08690(new_n8573, new_n8572, new_n9067);
not_1  g08691(new_n9067, new_n9068);
nor_1  g08692(new_n8574, new_n8571, new_n9069);
nor_1  g08693(new_n9069, new_n9068, new_n9070);
nand_1 g08694(new_n8564, new_n8563, new_n9071);
not_1  g08695(new_n9071, new_n9072);
nor_1  g08696(new_n8565, new_n8562, new_n9073);
nor_1  g08697(new_n9073, new_n9072, new_n9074);
not_1  g08698(n9725, new_n9075);
nor_1  g08699(new_n9075, new_n424, new_n9076);
xnor_1 g08700(new_n9076, new_n9074, new_n9077);
xnor_1 g08701(new_n9077, new_n9070, new_n9078);
xnor_1 g08702(new_n9078, new_n9066, new_n9079);
nand_1 g08703(new_n8717_1, new_n8674, new_n9080_1);
nand_1 g08704(new_n8718, new_n8688, new_n9081);
nand_1 g08705(new_n9081, new_n9080_1, new_n9082);
nand_1 g08706(new_n8940, new_n8910, new_n9083);
not_1  g08707(new_n8941, new_n9084);
nand_1 g08708(new_n8959, new_n9084, new_n9085);
nand_1 g08709(new_n9085, new_n9083, new_n9086);
xnor_1 g08710(new_n9086, new_n9082, new_n9087);
nand_1 g08711(new_n8824, new_n8790, new_n9088);
not_1  g08712(new_n8825, new_n9089);
nand_1 g08713(new_n8840, new_n9089, new_n9090);
nand_1 g08714(new_n9090, new_n9088, new_n9091);
nand_1 g08715(new_n8918, new_n8916, new_n9092);
not_1  g08716(new_n8930, new_n9093);
nand_1 g08717(new_n9093, new_n8920, new_n9094);
nand_1 g08718(new_n9094, new_n9092, new_n9095);
nand_1 g08719(new_n8697, new_n8691, new_n9096);
nand_1 g08720(new_n9096, new_n8695, new_n9097);
nand_1 g08721(n3986, n1478, new_n9098);
nand_1 g08722(n9241, n6429, new_n9099);
nand_1 g08723(n10022, n7965, new_n9100);
xnor_1 g08724(new_n9100, new_n9099, new_n9101);
xnor_1 g08725(new_n9101, new_n9098, new_n9102);
xnor_1 g08726(new_n9102, new_n9097, new_n9103);
xnor_1 g08727(new_n9103, new_n9095, new_n9104);
nand_1 g08728(new_n8926, new_n8925, new_n9105);
not_1  g08729(new_n9105, new_n9106);
nor_1  g08730(new_n8927, new_n8924, new_n9107);
nor_1  g08731(new_n9107, new_n9106, new_n9108);
not_1  g08732(new_n8809, new_n9109);
nor_1  g08733(new_n9109, new_n8805, new_n9110);
nor_1  g08734(new_n9110, new_n8806, new_n9111_1);
and_1  g08735(n11999, n7388, new_n9112);
nand_1 g08736(new_n9112, new_n9111_1, new_n9113);
not_1  g08737(new_n9111_1, new_n9114);
nand_1 g08738(new_n9112, new_n8830, new_n9115);
nand_1 g08739(new_n9115, new_n9114, new_n9116);
nand_1 g08740(new_n9116, new_n9113, new_n9117);
xnor_1 g08741(new_n9117, new_n9108, new_n9118);
nand_1 g08742(new_n8922, new_n8921, new_n9119);
nand_1 g08743(new_n8928, new_n8923, new_n9120);
nand_1 g08744(new_n9120, new_n9119, new_n9121);
and_1  g08745(new_n8797, new_n8794, new_n9122);
nor_1  g08746(new_n9122, new_n8799, new_n9123);
nand_1 g08747(n2530, n447, new_n9124);
nand_1 g08748(n12777, n7690, new_n9125);
nand_1 g08749(n8476, n1353, new_n9126);
xnor_1 g08750(new_n9126, new_n9125, new_n9127);
xnor_1 g08751(new_n9127, new_n9124, new_n9128);
xnor_1 g08752(new_n9128, new_n9123, new_n9129);
xnor_1 g08753(new_n9129, new_n9121, new_n9130);
xnor_1 g08754(new_n9130, new_n9118, new_n9131);
nand_1 g08755(n8759, n1198, new_n9132);
nand_1 g08756(n11728, n10510, new_n9133);
xnor_1 g08757(new_n9133, new_n9132, new_n9134);
nand_1 g08758(n12489, n4499, new_n9135);
nand_1 g08759(n10545, n6254, new_n9136);
xnor_1 g08760(new_n9136, new_n9135, new_n9137_1);
nand_1 g08761(n5331, n4436, new_n9138);
nand_1 g08762(n12947, n2393, new_n9139);
xnor_1 g08763(new_n9139, new_n9138, new_n9140);
xnor_1 g08764(new_n9140, new_n9137_1, new_n9141);
xnor_1 g08765(new_n9141, new_n9134, new_n9142);
nor_1  g08766(new_n829, new_n8888, new_n9143);
nand_1 g08767(n7159, n3616, new_n9144);
nand_1 g08768(n12709, n10644, new_n9145);
xnor_1 g08769(new_n9145, new_n9144, new_n9146);
xnor_1 g08770(new_n9146, new_n9143, new_n9147);
nand_1 g08771(n8819, n8276, new_n9148);
nand_1 g08772(n7730, n6776, new_n9149);
xnor_1 g08773(new_n9149, new_n9148, new_n9150);
xnor_1 g08774(new_n9150, new_n9147, new_n9151);
xnor_1 g08775(new_n9151, new_n9142, new_n9152);
xnor_1 g08776(new_n9152, new_n9131, new_n9153);
xnor_1 g08777(new_n9153, new_n9104, new_n9154);
not_1  g08778(new_n8815, new_n9155);
nand_1 g08779(new_n8823, new_n9155, new_n9156);
nand_1 g08780(new_n9156, new_n8820, new_n9157);
nand_1 g08781(n12705, n4370, new_n9158);
not_1  g08782(new_n8566, new_n9159);
nand_1 g08783(new_n9159, new_n8560, new_n9160);
nand_1 g08784(new_n8576, new_n8567, new_n9161);
nand_1 g08785(new_n9161, new_n9160, new_n9162);
nand_1 g08786(new_n8812, new_n8810, new_n9163);
nand_1 g08787(new_n8814, new_n8802, new_n9164);
nand_1 g08788(new_n9164, new_n9163, new_n9165);
xnor_1 g08789(new_n9165, new_n9162, new_n9166);
xnor_1 g08790(new_n9166, new_n9158, new_n9167);
xnor_1 g08791(new_n9167, new_n9157, new_n9168);
xnor_1 g08792(new_n9168, new_n9154, new_n9169);
xnor_1 g08793(new_n9169, new_n9091, new_n9170);
xnor_1 g08794(new_n9170, new_n9087, new_n9171);
xnor_1 g08795(new_n9171, new_n9079, new_n9172);
not_1  g08796(new_n8964, new_n9173);
nand_1 g08797(new_n8992, new_n9173, new_n9174);
nand_1 g08798(new_n9174, new_n8962, new_n9175);
not_1  g08799(new_n8710, new_n9176);
nand_1 g08800(new_n8716, new_n9176, new_n9177);
nand_1 g08801(new_n9177, new_n8713, new_n9178);
nand_1 g08802(n11407, n10547, new_n9179);
nor_1  g08803(new_n8515, new_n395, new_n9180);
xnor_1 g08804(new_n9180, new_n9179, new_n9181);
nand_1 g08805(n12299, n8717, new_n9182);
nand_1 g08806(n5857, n5760, new_n9183);
xnor_1 g08807(new_n9183, new_n9182, new_n9184);
nand_1 g08808(n12025, n11877, new_n9185);
nand_1 g08809(n12000, n1097, new_n9186);
xnor_1 g08810(new_n9186, new_n9185, new_n9187);
xnor_1 g08811(new_n9187, new_n9184, new_n9188);
xnor_1 g08812(new_n9188, new_n9181, new_n9189_1);
nand_1 g08813(new_n8706, new_n8705, new_n9190);
not_1  g08814(new_n9190, new_n9191);
nor_1  g08815(new_n8707, new_n8704, new_n9192);
nor_1  g08816(new_n9192, new_n9191, new_n9193);
nand_1 g08817(n10990, n45, new_n9194);
xnor_1 g08818(new_n9194, new_n9193, new_n9195_1);
xnor_1 g08819(new_n9195_1, new_n9189_1, new_n9196);
nand_1 g08820(new_n8702, new_n8701, new_n9197);
not_1  g08821(new_n8708, new_n9198);
nand_1 g08822(new_n9198, new_n8703, new_n9199);
nand_1 g08823(new_n9199, new_n9197, new_n9200);
nor_1  g08824(new_n599, new_n8622, new_n9201);
xnor_1 g08825(new_n9201, new_n9200, new_n9202);
xnor_1 g08826(new_n9202, new_n9196, new_n9203);
nand_1 g08827(new_n8914, new_n8913, new_n9204);
not_1  g08828(new_n9204, new_n9205);
nor_1  g08829(new_n8915, new_n8912, new_n9206);
nor_1  g08830(new_n9206, new_n9205, new_n9207);
not_1  g08831(new_n8699, new_n9208);
nand_1 g08832(new_n9208, new_n8690, new_n9209);
not_1  g08833(new_n8709, new_n9210);
nand_1 g08834(new_n9210, new_n8700, new_n9211);
nand_1 g08835(new_n9211, new_n9209, new_n9212);
xnor_1 g08836(new_n9212, new_n9207, new_n9213);
xnor_1 g08837(new_n9213, new_n9203, new_n9214);
xnor_1 g08838(new_n9214, new_n9178, new_n9215);
not_1  g08839(new_n8931, new_n9216);
nand_1 g08840(new_n8939, new_n9216, new_n9217);
nand_1 g08841(new_n9217, new_n8936, new_n9218);
nand_1 g08842(new_n8792, new_n8791, new_n9219);
or_1   g08843(new_n8801, new_n8793, new_n9220);
nand_1 g08844(new_n9220, new_n9219, new_n9221);
nand_1 g08845(n11892, n6441, new_n9222);
nand_1 g08846(n11791, n5860, new_n9223);
xnor_1 g08847(new_n9223, new_n9222, new_n9224);
nand_1 g08848(n11257, n5212, new_n9225);
nand_1 g08849(n6604, n5305, new_n9226);
xnor_1 g08850(new_n9226, new_n9225, new_n9227);
xnor_1 g08851(new_n9227, new_n9224, new_n9228);
xnor_1 g08852(new_n9228, new_n9221, new_n9229);
xnor_1 g08853(new_n9229, new_n9218, new_n9230);
xnor_1 g08854(new_n9230, new_n9215, new_n9231);
nor_1  g08855(new_n8569, new_n8568, new_n9232);
not_1  g08856(new_n8575, new_n9233);
nor_1  g08857(new_n9233, new_n8570, new_n9234);
nor_1  g08858(new_n9234, new_n9232, new_n9235);
nand_1 g08859(new_n8530, new_n8581, new_n9236);
nand_1 g08860(new_n8583, new_n8577, new_n9237);
nand_1 g08861(new_n9237, new_n9236, new_n9238);
xnor_1 g08862(new_n9238, new_n9235, new_n9239);
xnor_1 g08863(new_n9239, new_n9231, new_n9240);
xnor_1 g08864(new_n9240, new_n9175, new_n9241_1);
xnor_1 g08865(new_n9241_1, new_n9172, new_n9242);
xnor_1 g08866(new_n9242, new_n9062, new_n9243);
xnor_1 g08867(new_n9243, new_n9058, n3287);
xnor_1 g08868(new_n9054, new_n9035, n3339);
xnor_1 g08869(new_n4178, new_n4175, n3456);
nor_1  g08870(new_n378, new_n492, new_n9247);
nor_1  g08871(new_n396, new_n4283, new_n9248);
not_1  g08872(new_n9248, new_n9249);
nand_1 g08873(n9920, n2509, new_n9250);
nand_1 g08874(n6038, n3627, new_n9251);
nand_1 g08875(new_n9251, new_n9250, new_n9252);
nor_1  g08876(new_n9251, new_n9250, new_n9253);
not_1  g08877(new_n9253, new_n9254);
nand_1 g08878(new_n9254, new_n9252, new_n9255);
nand_1 g08879(new_n9255, new_n9249, new_n9256);
not_1  g08880(new_n9256, new_n9257);
nor_1  g08881(new_n9255, new_n9249, new_n9258);
nor_1  g08882(new_n9258, new_n9257, new_n9259);
not_1  g08883(new_n9259, new_n9260);
nand_1 g08884(n9920, n6038, new_n9261);
nand_1 g08885(n12720, n4189, new_n9262);
nand_1 g08886(new_n9262, new_n9261, new_n9263);
not_1  g08887(new_n9263, new_n9264);
nor_1  g08888(new_n4283, new_n413, new_n9265);
nor_1  g08889(new_n9262, new_n9261, new_n9266);
nor_1  g08890(new_n9266, new_n9264, new_n9267);
not_1  g08891(new_n9267, new_n9268);
nor_1  g08892(new_n9268, new_n9265, new_n9269);
nor_1  g08893(new_n9269, new_n9264, new_n9270);
xnor_1 g08894(new_n9270, new_n9260, new_n9271);
nor_1  g08895(new_n1377, new_n420, new_n9272);
nand_1 g08896(n6770, n6038, new_n9273);
nand_1 g08897(n4189, n2509, new_n9274);
nand_1 g08898(new_n9274, new_n9273, new_n9275);
not_1  g08899(new_n9275, new_n9276);
nor_1  g08900(new_n396, new_n1377, new_n9277);
xnor_1 g08901(new_n9274, new_n9273, new_n9278);
nor_1  g08902(new_n9278, new_n9277, new_n9279);
nor_1  g08903(new_n9279, new_n9276, new_n9280);
nand_1 g08904(new_n9280, new_n9272, new_n9281);
xnor_1 g08905(new_n9268, new_n9265, new_n9282);
not_1  g08906(new_n9281, new_n9283);
nor_1  g08907(new_n9280, new_n9272, new_n9284);
nor_1  g08908(new_n9284, new_n9283, new_n9285);
nand_1 g08909(new_n9285, new_n9282, new_n9286);
nand_1 g08910(new_n9286, new_n9281, new_n9287);
nor_1  g08911(new_n423, new_n1377, new_n9288);
not_1  g08912(new_n9288, new_n9289);
nor_1  g08913(new_n1367, new_n420, new_n9290);
not_1  g08914(new_n9290, new_n9291);
nor_1  g08915(new_n9291, new_n9289, new_n9292);
not_1  g08916(new_n9292, new_n9293);
nand_1 g08917(new_n9291, new_n9289, new_n9294);
nand_1 g08918(new_n9294, new_n9293, new_n9295);
xnor_1 g08919(new_n9295, new_n9287, new_n9296);
xnor_1 g08920(new_n9296, new_n9271, new_n9297);
not_1  g08921(new_n9297, new_n9298);
nor_1  g08922(new_n378, new_n423, new_n9299);
nor_1  g08923(new_n378, new_n420, new_n9300);
not_1  g08924(new_n9262, new_n9301);
nand_1 g08925(new_n9301, new_n379, new_n9302);
nand_1 g08926(n6038, n4189, new_n9303);
nand_1 g08927(n12720, n6687, new_n9304);
nand_1 g08928(new_n9304, new_n9303, new_n9305);
nor_1  g08929(new_n1377, new_n413, new_n9306);
nand_1 g08930(new_n9306, new_n9305, new_n9307);
nand_1 g08931(new_n9307, new_n9302, new_n9308);
nand_1 g08932(new_n9308, new_n9300, new_n9309);
not_1  g08933(new_n9309, new_n9310);
nor_1  g08934(new_n9308, new_n9300, new_n9311);
nor_1  g08935(new_n9311, new_n9310, new_n9312);
xnor_1 g08936(new_n9278, new_n9277, new_n9313);
nand_1 g08937(new_n9313, new_n9312, new_n9314);
nand_1 g08938(new_n9314, new_n9309, new_n9315);
nor_1  g08939(new_n9315, new_n9299, new_n9316);
xnor_1 g08940(new_n9285, new_n9282, new_n9317);
not_1  g08941(new_n9317, new_n9318);
xnor_1 g08942(new_n9315, new_n9299, new_n9319);
nor_1  g08943(new_n9319, new_n9318, new_n9320);
nor_1  g08944(new_n9320, new_n9316, new_n9321);
nand_1 g08945(new_n9321, new_n9298, new_n9322);
not_1  g08946(new_n9322, new_n9323);
nor_1  g08947(new_n9321, new_n9298, new_n9324);
nor_1  g08948(new_n9324, new_n9323, new_n9325);
nand_1 g08949(new_n9325, new_n9247, new_n9326);
xor_1  g08950(new_n9313, new_n9312, new_n9327);
nand_1 g08951(new_n9305, new_n9302, new_n9328);
not_1  g08952(new_n9328, new_n9329);
nor_1  g08953(new_n378, new_n413, new_n9330);
nor_1  g08954(new_n377, new_n1377, new_n9331);
nand_1 g08955(new_n9331, new_n9330, new_n9332);
nor_1  g08956(new_n9332, new_n9329, new_n9333);
nand_1 g08957(new_n9333, new_n9327, new_n9334);
xnor_1 g08958(new_n9319, new_n9317, new_n9335);
nor_1  g08959(new_n9335, new_n9334, new_n9336);
not_1  g08960(new_n9247, new_n9337);
xnor_1 g08961(new_n9325, new_n9337, new_n9338);
nand_1 g08962(new_n9338, new_n9336, new_n9339);
nand_1 g08963(new_n9339, new_n9326, new_n9340);
nor_1  g08964(new_n9270, new_n9260, new_n9341);
nor_1  g08965(new_n9341, new_n9257, new_n9342);
not_1  g08966(new_n9342, new_n9343);
nor_1  g08967(new_n492, new_n1377, new_n9344);
nand_1 g08968(n4189, n2585, new_n9345);
nand_1 g08969(n12706, n6687, new_n9346);
xnor_1 g08970(new_n9346, new_n9345, new_n9347);
xnor_1 g08971(new_n9347, new_n9344, new_n9348);
not_1  g08972(new_n9348, new_n9349);
nand_1 g08973(new_n9349, new_n9343, new_n9350);
nand_1 g08974(new_n9348, new_n9342, new_n9351);
nand_1 g08975(new_n9351, new_n9350, new_n9352);
nand_1 g08976(n6770, n2508, new_n9353);
xnor_1 g08977(new_n9353, new_n9253, new_n9354);
not_1  g08978(new_n9354, new_n9355);
nand_1 g08979(n3627, n2509, new_n9356);
nand_1 g08980(n12720, n9920, new_n9357);
nand_1 g08981(n6038, n4516, new_n9358);
nor_1  g08982(new_n9358, new_n9357, new_n9359);
nand_1 g08983(new_n9358, new_n9357, new_n9360);
not_1  g08984(new_n9360, new_n9361);
nor_1  g08985(new_n9361, new_n9359, new_n9362);
xor_1  g08986(new_n9362, new_n9356, new_n9363);
xnor_1 g08987(new_n9363, new_n9355, new_n9364);
xnor_1 g08988(new_n9364, new_n9352, new_n9365);
not_1  g08989(new_n9295, new_n9366);
nand_1 g08990(new_n9366, new_n9287, new_n9367);
nand_1 g08991(new_n9296, new_n9271, new_n9368);
xnor_1 g08992(new_n9368, new_n9293, new_n9369);
nand_1 g08993(new_n9369, new_n9367, new_n9370);
xnor_1 g08994(new_n9370, new_n9365, new_n9371);
xnor_1 g08995(new_n9371, new_n9322, new_n9372);
xor_1  g08996(new_n9372, new_n9340, new_n9373);
not_1  g08997(new_n9373, new_n9374);
nor_1  g08998(new_n382, new_n551, new_n9375);
nor_1  g08999(new_n1434, new_n564, new_n9376);
nand_1 g09000(n8336, n1209, new_n9377);
nand_1 g09001(n7354, n6986, new_n9378);
nand_1 g09002(new_n9378, new_n9377, new_n9379);
nand_1 g09003(new_n9379, new_n9376, new_n9380);
not_1  g09004(new_n9377, new_n9381);
not_1  g09005(new_n9378, new_n9382);
nand_1 g09006(new_n9382, new_n9381, new_n9383);
nand_1 g09007(new_n9383, new_n9380, new_n9384);
nand_1 g09008(new_n9384, new_n9375, new_n9385);
not_1  g09009(new_n9385, new_n9386);
nor_1  g09010(new_n9384, new_n9375, new_n9387_1);
nor_1  g09011(new_n9387_1, new_n9386, new_n9388);
nor_1  g09012(new_n564, new_n1508, new_n9389);
nand_1 g09013(n7354, n2226, new_n9390);
nand_1 g09014(n10928, n1209, new_n9391);
nand_1 g09015(new_n9391, new_n9390, new_n9392);
not_1  g09016(new_n9390, new_n9393);
not_1  g09017(new_n9391, new_n9394);
nand_1 g09018(new_n9394, new_n9393, new_n9395);
nand_1 g09019(new_n9395, new_n9392, new_n9396);
xnor_1 g09020(new_n9396, new_n9389, new_n9397);
nand_1 g09021(new_n9397, new_n9388, new_n9398);
not_1  g09022(new_n9398, new_n9399);
nor_1  g09023(new_n9397, new_n9388, new_n9400_1);
nor_1  g09024(new_n9400_1, new_n9399, new_n9401);
nand_1 g09025(new_n9383, new_n9379, new_n9402);
nor_1  g09026(new_n1434, new_n381_1, new_n9403);
nor_1  g09027(new_n382, new_n564, new_n9404);
and_1  g09028(new_n9404, new_n9403, new_n9405);
nand_1 g09029(new_n9405, new_n9402, new_n9406);
not_1  g09030(new_n9406, new_n9407);
and_1  g09031(new_n9407, new_n9401, new_n9408);
nor_1  g09032(new_n382, new_n588, new_n9409);
nand_1 g09033(new_n9398, new_n9385, new_n9410);
xnor_1 g09034(new_n9410, new_n9409, new_n9411);
nor_1  g09035(new_n1434, new_n551, new_n9412);
not_1  g09036(new_n9392, new_n9413);
not_1  g09037(new_n9395, new_n9414);
nor_1  g09038(new_n9414, new_n9389, new_n9415);
nor_1  g09039(new_n9415, new_n9413, new_n9416);
nand_1 g09040(new_n9416, new_n9412, new_n9417);
not_1  g09041(new_n9417, new_n9418);
nor_1  g09042(new_n9416, new_n9412, new_n9419);
nor_1  g09043(new_n9419, new_n9418, new_n9420);
nor_1  g09044(new_n1508, new_n557, new_n9421);
nand_1 g09045(n7354, n1094, new_n9422);
nand_1 g09046(n7500, n2226, new_n9423);
xnor_1 g09047(new_n9423, new_n9422, new_n9424);
nor_1  g09048(new_n9424, new_n9421, new_n9425);
not_1  g09049(new_n9425, new_n9426);
nand_1 g09050(new_n9424, new_n9421, new_n9427);
nand_1 g09051(new_n9427, new_n9426, new_n9428);
nand_1 g09052(new_n9428, new_n9420, new_n9429);
not_1  g09053(new_n9429, new_n9430);
nor_1  g09054(new_n9428, new_n9420, new_n9431);
nor_1  g09055(new_n9431, new_n9430, new_n9432);
xnor_1 g09056(new_n9432, new_n9411, new_n9433);
nand_1 g09057(new_n9433, new_n9408, new_n9434);
nor_1  g09058(new_n382, new_n621, new_n9435);
not_1  g09059(new_n9435, new_n9436);
nor_1  g09060(new_n4529, new_n557, new_n9437);
nand_1 g09061(new_n9423, new_n9422, new_n9438);
not_1  g09062(new_n9438, new_n9439);
nor_1  g09063(new_n9425, new_n9439, new_n9440);
nand_1 g09064(new_n9440, new_n9437, new_n9441);
not_1  g09065(new_n9441, new_n9442);
nor_1  g09066(new_n9440, new_n9437, new_n9443);
nor_1  g09067(new_n9443, new_n9442, new_n9444);
nand_1 g09068(n7500, n1094, new_n9445);
nand_1 g09069(n10678, n7354, new_n9446);
nand_1 g09070(new_n9446, new_n9445, new_n9447);
nor_1  g09071(new_n9446, new_n9445, new_n9448);
not_1  g09072(new_n9448, new_n9449);
nand_1 g09073(new_n9449, new_n9447, new_n9450);
xnor_1 g09074(new_n9450, new_n9444, new_n9451);
nand_1 g09075(n10928, n4141, new_n9452);
nand_1 g09076(n6986, n5105, new_n9453);
nand_1 g09077(new_n9453, new_n9452, new_n9454);
nor_1  g09078(new_n9453, new_n9452, new_n9455);
not_1  g09079(new_n9455, new_n9456);
nand_1 g09080(new_n9456, new_n9454, new_n9457_1);
xnor_1 g09081(new_n9457_1, new_n9451, new_n9458);
nor_1  g09082(new_n9430, new_n9418, new_n9459);
not_1  g09083(new_n9459, new_n9460);
nand_1 g09084(new_n9460, new_n9458, new_n9461);
not_1  g09085(new_n9461, new_n9462);
nor_1  g09086(new_n9460, new_n9458, new_n9463);
nor_1  g09087(new_n9463, new_n9462, new_n9464);
nor_1  g09088(new_n9410, new_n9409, new_n9465);
nor_1  g09089(new_n9432, new_n9411, new_n9466);
nor_1  g09090(new_n9466, new_n9465, new_n9467);
nand_1 g09091(new_n9467, new_n9464, new_n9468);
not_1  g09092(new_n9468, new_n9469);
nor_1  g09093(new_n9467, new_n9464, new_n9470);
nor_1  g09094(new_n9470, new_n9469, new_n9471);
xnor_1 g09095(new_n9471, new_n9436, new_n9472);
nand_1 g09096(new_n9472, new_n9434, new_n9473);
not_1  g09097(new_n9473, new_n9474);
nor_1  g09098(new_n9472, new_n9434, new_n9475);
nor_1  g09099(new_n9475, new_n9474, new_n9476);
nor_1  g09100(new_n385, new_n753_1, new_n9477);
nand_1 g09101(n11222, n1980, new_n9478);
nand_1 g09102(n8028, n5314, new_n9479);
nor_1  g09103(new_n9479, new_n9478, new_n9480);
not_1  g09104(new_n9480, new_n9481);
nand_1 g09105(new_n9479, new_n9478, new_n9482);
nor_1  g09106(new_n1467, new_n697, new_n9483);
nand_1 g09107(new_n9483, new_n9482, new_n9484);
nand_1 g09108(new_n9484, new_n9481, new_n9485);
xnor_1 g09109(new_n9485, new_n9477, new_n9486);
nor_1  g09110(new_n697, new_n1562, new_n9487);
nand_1 g09111(n8028, n996, new_n9488);
nand_1 g09112(n11153, n1980, new_n9489);
nor_1  g09113(new_n9489, new_n9488, new_n9490);
not_1  g09114(new_n9490, new_n9491);
nand_1 g09115(new_n9489, new_n9488, new_n9492);
nand_1 g09116(new_n9492, new_n9491, new_n9493);
xnor_1 g09117(new_n9493, new_n9487, new_n9494);
not_1  g09118(new_n9494, new_n9495);
nor_1  g09119(new_n9495, new_n9486, new_n9496);
not_1  g09120(new_n9496, new_n9497);
nand_1 g09121(new_n9495, new_n9486, new_n9498);
nand_1 g09122(new_n9498, new_n9497, new_n9499);
not_1  g09123(new_n9499, new_n9500);
not_1  g09124(new_n9482, new_n9501);
nor_1  g09125(new_n9501, new_n9480, new_n9502);
not_1  g09126(new_n9502, new_n9503);
nand_1 g09127(n11153, n8028, new_n9504);
nand_1 g09128(n11222, n10848, new_n9505);
nor_1  g09129(new_n9505, new_n9504, new_n9506);
and_1  g09130(new_n9506, new_n9503, new_n9507);
nand_1 g09131(new_n9507, new_n9500, new_n9508);
nand_1 g09132(new_n9485, new_n9477, new_n9509);
not_1  g09133(new_n9509, new_n9510);
nor_1  g09134(new_n9496, new_n9510, new_n9511);
nor_1  g09135(new_n790, new_n385, new_n9512);
not_1  g09136(new_n9512, new_n9513);
nor_1  g09137(new_n1467, new_n753_1, new_n9514);
not_1  g09138(new_n9492, new_n9515);
nor_1  g09139(new_n9490, new_n9487, new_n9516);
nor_1  g09140(new_n9516, new_n9515, new_n9517);
nand_1 g09141(new_n9517, new_n9514, new_n9518);
not_1  g09142(new_n9518, new_n9519);
nor_1  g09143(new_n9517, new_n9514, new_n9520);
nor_1  g09144(new_n9520, new_n9519, new_n9521);
nor_1  g09145(new_n697, new_n4542, new_n9522);
nor_1  g09146(new_n1562, new_n764, new_n9523);
not_1  g09147(new_n9523, new_n9524);
nor_1  g09148(new_n384, new_n6869, new_n9525);
not_1  g09149(new_n9525, new_n9526);
nor_1  g09150(new_n9526, new_n9524, new_n9527);
nand_1 g09151(new_n9526, new_n9524, new_n9528);
not_1  g09152(new_n9528, new_n9529);
nor_1  g09153(new_n9529, new_n9527, new_n9530);
xnor_1 g09154(new_n9530, new_n9522, new_n9531);
xnor_1 g09155(new_n9531, new_n9521, new_n9532);
xnor_1 g09156(new_n9532, new_n9513, new_n9533);
nand_1 g09157(new_n9533, new_n9511, new_n9534);
not_1  g09158(new_n9534, new_n9535);
nor_1  g09159(new_n9533, new_n9511, new_n9536);
nor_1  g09160(new_n9536, new_n9535, new_n9537);
nor_1  g09161(new_n9537, new_n9508, new_n9538);
nor_1  g09162(new_n385, new_n915, new_n9539);
not_1  g09163(new_n9539, new_n9540);
nand_1 g09164(n1980, n996, new_n9541);
nand_1 g09165(n8028, n5319, new_n9542);
nand_1 g09166(n10848, n5767, new_n9543);
xnor_1 g09167(new_n9543, new_n9542, new_n9544);
nor_1  g09168(new_n9544, new_n9541, new_n9545);
not_1  g09169(new_n9545, new_n9546);
nand_1 g09170(new_n9544, new_n9541, new_n9547);
nand_1 g09171(new_n9547, new_n9546, new_n9548);
nor_1  g09172(new_n9527, new_n9522, new_n9549);
nor_1  g09173(new_n9549, new_n9529, new_n9550);
xnor_1 g09174(new_n9550, new_n9548, new_n9551);
nor_1  g09175(new_n790, new_n1467, new_n9552);
not_1  g09176(new_n9552, new_n9553);
nor_1  g09177(new_n753_1, new_n1562, new_n9554);
not_1  g09178(new_n9554, new_n9555);
nand_1 g09179(new_n9555, new_n9553, new_n9556);
nor_1  g09180(new_n9555, new_n9553, new_n9557);
not_1  g09181(new_n9557, new_n9558);
nand_1 g09182(new_n9558, new_n9556, new_n9559);
xnor_1 g09183(new_n9559, new_n9551, new_n9560);
not_1  g09184(new_n9521, new_n9561);
nor_1  g09185(new_n9531, new_n9561, new_n9562);
nor_1  g09186(new_n9562, new_n9519, new_n9563);
not_1  g09187(new_n9563, new_n9564);
nand_1 g09188(new_n9564, new_n9560, new_n9565);
not_1  g09189(new_n9565, new_n9566);
nor_1  g09190(new_n9564, new_n9560, new_n9567);
nor_1  g09191(new_n9567, new_n9566, new_n9568);
not_1  g09192(new_n9532, new_n9569);
nand_1 g09193(new_n9569, new_n9513, new_n9570);
nand_1 g09194(new_n9534, new_n9570, new_n9571_1);
xnor_1 g09195(new_n9571_1, new_n9568, new_n9572);
xnor_1 g09196(new_n9572, new_n9540, new_n9573);
xnor_1 g09197(new_n9573, new_n9538, new_n9574);
not_1  g09198(new_n9574, new_n9575);
nor_1  g09199(new_n1533, new_n735, new_n9576);
nor_1  g09200(new_n4386, new_n667, new_n9577);
not_1  g09201(new_n9577, new_n9578_1);
nor_1  g09202(new_n1533, new_n869, new_n9579);
not_1  g09203(new_n9579, new_n9580);
nand_1 g09204(new_n9580, new_n9578_1, new_n9581);
nor_1  g09205(new_n1452, new_n711, new_n9582);
nand_1 g09206(new_n9582, new_n9581, new_n9583_1);
nand_1 g09207(new_n9579, new_n9577, new_n9584);
nand_1 g09208(new_n9584, new_n9583_1, new_n9585);
xnor_1 g09209(new_n9585, new_n9576, new_n9586);
nor_1  g09210(new_n4386, new_n711, new_n9587);
not_1  g09211(new_n9587, new_n9588);
nand_1 g09212(n7160, n1564, new_n9589);
nand_1 g09213(n12391, n533, new_n9590);
xnor_1 g09214(new_n9590, new_n9589, new_n9591);
xnor_1 g09215(new_n9591, new_n9588, new_n9592);
xnor_1 g09216(new_n9592, new_n9586, new_n9593);
nand_1 g09217(new_n9584, new_n9581, new_n9594);
nand_1 g09218(n12391, n1564, new_n9595);
nand_1 g09219(n12069, n1512, new_n9596);
nor_1  g09220(new_n9596, new_n9595, new_n9597);
nand_1 g09221(new_n9597, new_n9594, new_n9598);
nor_1  g09222(new_n9598, new_n9593, new_n9599);
not_1  g09223(new_n9599, new_n9600);
nor_1  g09224(new_n1533, new_n820, new_n9601);
not_1  g09225(new_n9601, new_n9602);
nand_1 g09226(n12391, n2802, new_n9603);
nand_1 g09227(new_n9590, new_n9589, new_n9604);
not_1  g09228(new_n9604, new_n9605);
nor_1  g09229(new_n9591, new_n9587, new_n9606);
nor_1  g09230(new_n9606, new_n9605, new_n9607);
xnor_1 g09231(new_n9607, new_n9603, new_n9608);
nand_1 g09232(n7891, n533, new_n9609);
nand_1 g09233(n4828, n1564, new_n9610);
nand_1 g09234(n7160, n1512, new_n9611);
xnor_1 g09235(new_n9611, new_n9610, new_n9612);
xnor_1 g09236(new_n9612, new_n9609, new_n9613);
xnor_1 g09237(new_n9613, new_n9608, new_n9614);
xnor_1 g09238(new_n9614, new_n9602, new_n9615);
nand_1 g09239(new_n9585, new_n9576, new_n9616);
not_1  g09240(new_n9616, new_n9617);
nor_1  g09241(new_n9592, new_n9586, new_n9618);
nor_1  g09242(new_n9618, new_n9617, new_n9619);
nand_1 g09243(new_n9619, new_n9615, new_n9620);
not_1  g09244(new_n9620, new_n9621);
nor_1  g09245(new_n9619, new_n9615, new_n9622);
nor_1  g09246(new_n9622, new_n9621, new_n9623);
nor_1  g09247(new_n9623, new_n9600, new_n9624);
not_1  g09248(new_n9624, new_n9625);
nor_1  g09249(new_n1533, new_n867, new_n9626);
not_1  g09250(new_n9626, new_n9627);
nand_1 g09251(n7160, n533, new_n9628);
not_1  g09252(new_n9628, new_n9629);
nand_1 g09253(n2515, n1564, new_n9630);
nand_1 g09254(n4828, n1512, new_n9631);
xnor_1 g09255(new_n9631, new_n9630, new_n9632);
xnor_1 g09256(new_n9632, new_n9629, new_n9633);
nand_1 g09257(new_n9611, new_n9610, new_n9634);
not_1  g09258(new_n9634, new_n9635);
not_1  g09259(new_n9609, new_n9636);
nor_1  g09260(new_n9612, new_n9636, new_n9637_1);
nor_1  g09261(new_n9637_1, new_n9635, new_n9638);
nand_1 g09262(new_n9638, new_n9633, new_n9639);
not_1  g09263(new_n9639, new_n9640_1);
nor_1  g09264(new_n9638, new_n9633, new_n9641);
nor_1  g09265(new_n9641, new_n9640_1, new_n9642);
nor_1  g09266(new_n4386, new_n735, new_n9643);
not_1  g09267(new_n9643, new_n9644);
nor_1  g09268(new_n1452, new_n820, new_n9645);
not_1  g09269(new_n9645, new_n9646);
nor_1  g09270(new_n9646, new_n9644, new_n9647);
not_1  g09271(new_n9647, new_n9648);
nand_1 g09272(new_n9646, new_n9644, new_n9649);
nand_1 g09273(new_n9649, new_n9648, new_n9650);
xnor_1 g09274(new_n9650, new_n9642, new_n9651);
not_1  g09275(new_n9603, new_n9652);
nand_1 g09276(new_n9607, new_n9652, new_n9653);
not_1  g09277(new_n9613, new_n9654);
nand_1 g09278(new_n9654, new_n9608, new_n9655);
nand_1 g09279(new_n9655, new_n9653, new_n9656);
nand_1 g09280(new_n9656, new_n9651, new_n9657);
not_1  g09281(new_n9657, new_n9658);
nor_1  g09282(new_n9656, new_n9651, new_n9659);
nor_1  g09283(new_n9659, new_n9658, new_n9660);
not_1  g09284(new_n9660, new_n9661);
not_1  g09285(new_n9614, new_n9662);
nand_1 g09286(new_n9662, new_n9602, new_n9663);
nand_1 g09287(new_n9620, new_n9663, new_n9664);
xnor_1 g09288(new_n9664, new_n9661, new_n9665);
nand_1 g09289(new_n9665, new_n9627, new_n9666);
xnor_1 g09290(new_n9664, new_n9660, new_n9667);
nand_1 g09291(new_n9667, new_n9626, new_n9668);
nand_1 g09292(new_n9668, new_n9666, new_n9669);
xnor_1 g09293(new_n9669, new_n9625, new_n9670);
xnor_1 g09294(new_n9670, new_n9575, new_n9671);
xnor_1 g09295(new_n9537, new_n9508, new_n9672);
not_1  g09296(new_n9598, new_n9673);
xnor_1 g09297(new_n9673, new_n9593, new_n9674);
xnor_1 g09298(new_n9507, new_n9499, new_n9675);
nor_1  g09299(new_n9675, new_n9674, new_n9676);
not_1  g09300(new_n9676, new_n9677);
nand_1 g09301(new_n9582, new_n388, new_n9678);
nand_1 g09302(new_n9678, new_n9594, new_n9679);
not_1  g09303(new_n9583_1, new_n9680);
nand_1 g09304(new_n9680, new_n388, new_n9681);
nand_1 g09305(new_n9681, new_n9679, new_n9682);
not_1  g09306(new_n9682, new_n9683);
nand_1 g09307(new_n9483, new_n387, new_n9684);
not_1  g09308(new_n9684, new_n9685);
nor_1  g09309(new_n9685, new_n9502, new_n9686);
nor_1  g09310(new_n9684, new_n9501, new_n9687);
nor_1  g09311(new_n9687, new_n9686, new_n9688);
nand_1 g09312(new_n9688, new_n9683, new_n9689);
xnor_1 g09313(new_n9505, new_n9504, new_n9690);
nand_1 g09314(new_n9690, new_n390, new_n9691);
xnor_1 g09315(new_n9690, new_n389, new_n9692);
xnor_1 g09316(new_n9596, new_n9595, new_n9693);
nand_1 g09317(new_n9693, new_n9692, new_n9694);
nand_1 g09318(new_n9694, new_n9691, new_n9695);
not_1  g09319(new_n9695, new_n9696);
not_1  g09320(new_n9689, new_n9697);
nor_1  g09321(new_n9688, new_n9683, new_n9698);
nor_1  g09322(new_n9698, new_n9697, new_n9699);
nand_1 g09323(new_n9699, new_n9696, new_n9700);
nand_1 g09324(new_n9700, new_n9689, new_n9701);
not_1  g09325(new_n9701, new_n9702);
not_1  g09326(new_n9674, new_n9703);
xnor_1 g09327(new_n9675, new_n9703, new_n9704);
nand_1 g09328(new_n9704, new_n9702, new_n9705);
nand_1 g09329(new_n9705, new_n9677, new_n9706_1);
nand_1 g09330(new_n9706_1, new_n9672, new_n9707);
xnor_1 g09331(new_n9623, new_n9599, new_n9708);
not_1  g09332(new_n9708, new_n9709);
not_1  g09333(new_n9672, new_n9710);
xnor_1 g09334(new_n9706_1, new_n9710, new_n9711);
nand_1 g09335(new_n9711, new_n9709, new_n9712);
nand_1 g09336(new_n9712, new_n9707, new_n9713);
nand_1 g09337(new_n9713, new_n9671, new_n9714);
not_1  g09338(new_n9714, new_n9715);
nor_1  g09339(new_n9713, new_n9671, new_n9716);
nor_1  g09340(new_n9716, new_n9715, new_n9717);
nor_1  g09341(new_n9717, new_n9476, new_n9718);
xnor_1 g09342(new_n9717, new_n9476, new_n9719);
xnor_1 g09343(new_n9433, new_n9408, new_n9720);
xnor_1 g09344(new_n9711, new_n9708, new_n9721);
nor_1  g09345(new_n9721, new_n9720, new_n9722);
xnor_1 g09346(new_n9721, new_n9720, new_n9723);
nor_1  g09347(new_n9407, new_n9401, new_n9724);
nor_1  g09348(new_n9724, new_n9408, new_n9725_1);
not_1  g09349(new_n9725_1, new_n9726);
xnor_1 g09350(new_n9704, new_n9701, new_n9727);
nor_1  g09351(new_n9727, new_n9726, new_n9728);
xnor_1 g09352(new_n9727, new_n9725_1, new_n9729);
not_1  g09353(new_n9729, new_n9730);
not_1  g09354(new_n9699, new_n9731);
nand_1 g09355(new_n9731, new_n9695, new_n9732);
nand_1 g09356(new_n9732, new_n9700, new_n9733);
not_1  g09357(new_n9733, new_n9734);
not_1  g09358(new_n383, new_n9735);
nand_1 g09359(new_n9376, new_n9735, new_n9736);
nor_1  g09360(new_n9736, new_n9379, new_n9737);
not_1  g09361(new_n9736, new_n9738);
nor_1  g09362(new_n9738, new_n9402, new_n9739);
nor_1  g09363(new_n9739, new_n9737, new_n9740);
not_1  g09364(new_n9740, new_n9741);
nor_1  g09365(new_n9741, new_n9734, new_n9742);
nor_1  g09366(new_n9740, new_n9733, new_n9743);
nor_1  g09367(new_n9743, new_n9742, new_n9744);
not_1  g09368(new_n9744, new_n9745);
xnor_1 g09369(new_n9693, new_n9692, new_n9746);
xor_1  g09370(new_n9404, new_n9403, new_n9747);
nand_1 g09371(new_n9747, new_n9746, new_n9748);
nor_1  g09372(new_n392, new_n9735, new_n9749);
not_1  g09373(new_n9748, new_n9750);
nor_1  g09374(new_n9747, new_n9746, new_n9751);
nor_1  g09375(new_n9751, new_n9750, new_n9752);
nand_1 g09376(new_n9752, new_n9749, new_n9753);
nand_1 g09377(new_n9753, new_n9748, new_n9754);
nor_1  g09378(new_n9754, new_n9745, new_n9755);
nor_1  g09379(new_n9755, new_n9742, new_n9756_1);
not_1  g09380(new_n9756_1, new_n9757);
nor_1  g09381(new_n9757, new_n9730, new_n9758);
nor_1  g09382(new_n9758, new_n9728, new_n9759);
nor_1  g09383(new_n9759, new_n9723, new_n9760);
nor_1  g09384(new_n9760, new_n9722, new_n9761);
nor_1  g09385(new_n9761, new_n9719, new_n9762);
nor_1  g09386(new_n9762, new_n9718, new_n9763_1);
not_1  g09387(new_n9450, new_n9764);
nand_1 g09388(new_n9764, new_n9444, new_n9765);
nand_1 g09389(new_n9765, new_n9441, new_n9766);
nor_1  g09390(new_n1434, new_n621, new_n9767_1);
nand_1 g09391(n6986, n4141, new_n9768);
nand_1 g09392(n8336, n8236, new_n9769);
xnor_1 g09393(new_n9769, new_n9768, new_n9770);
xor_1  g09394(new_n9770, new_n9767_1, new_n9771);
xnor_1 g09395(new_n9771, new_n9766, new_n9772);
nand_1 g09396(n5105, n2226, new_n9773);
xnor_1 g09397(new_n9773, new_n9448, new_n9774);
nor_1  g09398(new_n6725, new_n564, new_n9775);
nand_1 g09399(n7354, n7320, new_n9776);
nand_1 g09400(n1209, n1094, new_n9777);
xnor_1 g09401(new_n9777, new_n9776, new_n9778);
xor_1  g09402(new_n9778, new_n9775, new_n9779);
xnor_1 g09403(new_n9779, new_n9774, new_n9780);
xnor_1 g09404(new_n9780, new_n9772, new_n9781);
not_1  g09405(new_n9457_1, new_n9782);
nand_1 g09406(new_n9782, new_n9451, new_n9783);
nand_1 g09407(new_n9462, new_n9455, new_n9784);
nand_1 g09408(new_n9461, new_n9456, new_n9785);
nand_1 g09409(new_n9785, new_n9784, new_n9786);
nand_1 g09410(new_n9786, new_n9783, new_n9787);
xnor_1 g09411(new_n9787, new_n9781, new_n9788);
xnor_1 g09412(new_n9788, new_n9468, new_n9789);
not_1  g09413(new_n9471, new_n9790);
nand_1 g09414(new_n9790, new_n9436, new_n9791);
nand_1 g09415(new_n9473, new_n9791, new_n9792);
xnor_1 g09416(new_n9792, new_n9789, new_n9793);
not_1  g09417(new_n9793, new_n9794);
not_1  g09418(new_n9571_1, new_n9795);
nand_1 g09419(new_n9795, new_n9568, new_n9796);
not_1  g09420(new_n9548, new_n9797);
nand_1 g09421(new_n9550, new_n9797, new_n9798);
nand_1 g09422(new_n9798, new_n9546, new_n9799);
nor_1  g09423(new_n1467, new_n915, new_n9800);
nand_1 g09424(n12704, n5314, new_n9801);
nand_1 g09425(n11222, n4903, new_n9802);
xnor_1 g09426(new_n9802, new_n9801, new_n9803);
xnor_1 g09427(new_n9803, new_n9800, new_n9804);
xnor_1 g09428(new_n9804, new_n9799, new_n9805);
not_1  g09429(new_n9805, new_n9806);
nor_1  g09430(new_n9543, new_n9542, new_n9807);
nor_1  g09431(new_n753_1, new_n4542, new_n9808);
xor_1  g09432(new_n9808, new_n9807, new_n9809);
nor_1  g09433(new_n697, new_n6935, new_n9810);
nand_1 g09434(n5767, n1980, new_n9811);
nand_1 g09435(n9457, n8028, new_n9812);
xnor_1 g09436(new_n9812, new_n9811, new_n9813);
xor_1  g09437(new_n9813, new_n9810, new_n9814);
xnor_1 g09438(new_n9814, new_n9809, new_n9815);
not_1  g09439(new_n9815, new_n9816);
nand_1 g09440(new_n9816, new_n9806, new_n9817);
nand_1 g09441(new_n9815, new_n9805, new_n9818);
nand_1 g09442(new_n9818, new_n9817, new_n9819);
not_1  g09443(new_n9819, new_n9820_1);
not_1  g09444(new_n9559, new_n9821);
nand_1 g09445(new_n9821, new_n9551, new_n9822);
nand_1 g09446(new_n9566, new_n9557, new_n9823);
nand_1 g09447(new_n9565, new_n9558, new_n9824);
nand_1 g09448(new_n9824, new_n9823, new_n9825);
nand_1 g09449(new_n9825, new_n9822, new_n9826);
xnor_1 g09450(new_n9826, new_n9820_1, new_n9827);
xnor_1 g09451(new_n9827, new_n9796, new_n9828);
not_1  g09452(new_n9828, new_n9829);
nand_1 g09453(new_n9572, new_n9539, new_n9830);
nand_1 g09454(new_n9573, new_n9538, new_n9831);
nand_1 g09455(new_n9831, new_n9830, new_n9832);
xnor_1 g09456(new_n9832, new_n9829, new_n9833);
nor_1  g09457(new_n9664, new_n9661, new_n9834);
not_1  g09458(new_n9650, new_n9835);
nand_1 g09459(new_n9835, new_n9642, new_n9836);
nand_1 g09460(new_n9658, new_n9647, new_n9837);
nand_1 g09461(new_n9657, new_n9648, new_n9838);
nand_1 g09462(new_n9838, new_n9837, new_n9839);
nand_1 g09463(new_n9839, new_n9836, new_n9840);
nor_1  g09464(new_n9631, new_n9630, new_n9841);
nor_1  g09465(new_n1538, new_n735, new_n9842);
xor_1  g09466(new_n9842, new_n9841, new_n9843);
nor_1  g09467(new_n6823, new_n711, new_n9844);
nor_1  g09468(new_n667, new_n6828, new_n9845);
not_1  g09469(new_n9845, new_n9846);
nor_1  g09470(new_n6825, new_n869, new_n9847);
not_1  g09471(new_n9847, new_n9848);
nand_1 g09472(new_n9848, new_n9846, new_n9849);
nand_1 g09473(new_n9847, new_n9845, new_n9850);
nand_1 g09474(new_n9850, new_n9849, new_n9851);
xor_1  g09475(new_n9851, new_n9844, new_n9852);
xnor_1 g09476(new_n9852, new_n9843, new_n9853);
nor_1  g09477(new_n9632, new_n9628, new_n9854);
nor_1  g09478(new_n9640_1, new_n9854, new_n9855);
not_1  g09479(new_n9855, new_n9856);
nor_1  g09480(new_n1452, new_n867, new_n9857);
nand_1 g09481(n7891, n6806, new_n9858);
nand_1 g09482(n12069, n12044, new_n9859);
xnor_1 g09483(new_n9859, new_n9858, new_n9860);
xor_1  g09484(new_n9860, new_n9857, new_n9861);
xnor_1 g09485(new_n9861, new_n9856, new_n9862);
xnor_1 g09486(new_n9862, new_n9853, new_n9863);
xnor_1 g09487(new_n9863, new_n9840, new_n9864);
xnor_1 g09488(new_n9864, new_n9834, new_n9865);
nand_1 g09489(new_n9666, new_n9624, new_n9866);
nand_1 g09490(new_n9866, new_n9668, new_n9867);
xnor_1 g09491(new_n9867, new_n9865, new_n9868);
nand_1 g09492(new_n9670, new_n9574, new_n9869);
nand_1 g09493(new_n9714, new_n9869, new_n9870);
xnor_1 g09494(new_n9870, new_n9868, new_n9871);
xnor_1 g09495(new_n9871, new_n9833, new_n9872);
xnor_1 g09496(new_n9872, new_n9794, new_n9873);
xnor_1 g09497(new_n9873, new_n9763_1, new_n9874);
nand_1 g09498(new_n9874, new_n9374, new_n9875);
xor_1  g09499(new_n9338, new_n9336, new_n9876);
not_1  g09500(new_n9876, new_n9877);
xor_1  g09501(new_n9335, new_n9334, new_n9878);
not_1  g09502(new_n9878, new_n9879);
xnor_1 g09503(new_n9759, new_n9723, new_n9880);
nand_1 g09504(new_n9880, new_n9879, new_n9881);
xnor_1 g09505(new_n9333, new_n9327, new_n9882);
nor_1  g09506(new_n9756_1, new_n9729, new_n9883);
nor_1  g09507(new_n9883, new_n9758, new_n9884);
not_1  g09508(new_n9884, new_n9885);
nand_1 g09509(new_n9885, new_n9882, new_n9886);
xnor_1 g09510(new_n9884, new_n9882, new_n9887);
not_1  g09511(new_n9754, new_n9888);
nor_1  g09512(new_n9888, new_n9744, new_n9889);
nor_1  g09513(new_n9889, new_n9755, new_n9890);
nand_1 g09514(new_n9306, new_n380, new_n9891);
nand_1 g09515(new_n9891, new_n9328, new_n9892);
not_1  g09516(new_n9891, new_n9893);
nand_1 g09517(new_n9893, new_n9305, new_n9894);
nand_1 g09518(new_n9894, new_n9892, new_n9895);
nand_1 g09519(new_n9895, new_n9890, new_n9896);
not_1  g09520(new_n9890, new_n9897);
xnor_1 g09521(new_n9895, new_n9897, new_n9898);
nand_1 g09522(new_n393, new_n379, new_n9899);
xnor_1 g09523(new_n9331, new_n9330, new_n9900);
nand_1 g09524(new_n9900, new_n9899, new_n9901);
xnor_1 g09525(new_n9752, new_n9749, new_n9902);
xor_1  g09526(new_n9900, new_n9899, new_n9903);
nand_1 g09527(new_n9903, new_n9902, new_n9904);
nand_1 g09528(new_n9904, new_n9901, new_n9905);
nand_1 g09529(new_n9905, new_n9898, new_n9906);
nand_1 g09530(new_n9906, new_n9896, new_n9907);
nand_1 g09531(new_n9907, new_n9887, new_n9908);
nand_1 g09532(new_n9908, new_n9886, new_n9909);
xnor_1 g09533(new_n9880, new_n9878, new_n9910);
nand_1 g09534(new_n9910, new_n9909, new_n9911);
nand_1 g09535(new_n9911, new_n9881, new_n9912);
nand_1 g09536(new_n9912, new_n9877, new_n9913);
xnor_1 g09537(new_n9761, new_n9719, new_n9914);
xnor_1 g09538(new_n9912, new_n9876, new_n9915);
nand_1 g09539(new_n9915, new_n9914, new_n9916);
nand_1 g09540(new_n9916, new_n9913, new_n9917);
xnor_1 g09541(new_n9874, new_n9373, new_n9918);
nand_1 g09542(new_n9918, new_n9917, new_n9919);
nand_1 g09543(new_n9919, new_n9875, new_n9920_1);
not_1  g09544(new_n9870, new_n9921);
nor_1  g09545(new_n9921, new_n9868, new_n9922);
not_1  g09546(new_n9871, new_n9923);
nor_1  g09547(new_n9923, new_n9833, new_n9924);
nor_1  g09548(new_n9924, new_n9922, new_n9925);
nand_1 g09549(new_n9872, new_n9794, new_n9926);
xnor_1 g09550(new_n9872, new_n9793, new_n9927);
nand_1 g09551(new_n9927, new_n9763_1, new_n9928);
nand_1 g09552(new_n9928, new_n9926, new_n9929);
xnor_1 g09553(new_n9929, new_n9925, new_n9930);
nand_1 g09554(new_n9788, new_n9469, new_n9931);
not_1  g09555(new_n9792, new_n9932);
nand_1 g09556(new_n9932, new_n9789, new_n9933);
nand_1 g09557(new_n9933, new_n9931, new_n9934);
not_1  g09558(new_n9863, new_n9935);
nand_1 g09559(new_n9935, new_n9840, new_n9936);
nand_1 g09560(new_n9936, new_n9837, new_n9937);
nand_1 g09561(new_n9808, new_n9807, new_n9938_1);
not_1  g09562(new_n9814, new_n9939);
nand_1 g09563(new_n9939, new_n9809, new_n9940);
nand_1 g09564(new_n9940, new_n9938_1, new_n9941);
nand_1 g09565(new_n9849, new_n9844, new_n9942);
nand_1 g09566(new_n9942, new_n9850, new_n9943);
xnor_1 g09567(new_n9943, new_n9941, new_n9944);
nand_1 g09568(n8028, n4817, new_n9945);
not_1  g09569(n7523, new_n9946);
nor_1  g09570(new_n9946, new_n381_1, new_n9947);
xnor_1 g09571(new_n9947, new_n9945, new_n9948);
nand_1 g09572(n10848, n9457, new_n9949);
nand_1 g09573(n11222, n1906, new_n9950);
xnor_1 g09574(new_n9950, new_n9949, new_n9951);
nand_1 g09575(n6986, n4928, new_n9952);
nand_1 g09576(n4141, n2226, new_n9953);
xnor_1 g09577(new_n9953, new_n9952, new_n9954);
xnor_1 g09578(new_n9954, new_n9951, new_n9955);
xnor_1 g09579(new_n9955, new_n9948, new_n9956_1);
nor_1  g09580(new_n9361, new_n9356, new_n9957);
nor_1  g09581(new_n9957, new_n9359, new_n9958);
nand_1 g09582(n4516, n2509, new_n9959);
nand_1 g09583(n12704, n996, new_n9960);
nand_1 g09584(n12720, n3627, new_n9961);
xnor_1 g09585(new_n9961, new_n9960, new_n9962);
xnor_1 g09586(new_n9962, new_n9959, new_n9963);
xnor_1 g09587(new_n9963, new_n9958, new_n9964);
xnor_1 g09588(new_n9964, new_n9956_1, new_n9965);
nand_1 g09589(n2515, n533, new_n9966);
nand_1 g09590(n1512, n1199, new_n9967);
nand_1 g09591(n12391, n12044, new_n9968);
xnor_1 g09592(new_n9968, new_n9967, new_n9969);
xnor_1 g09593(new_n9969, new_n9966, new_n9970);
xnor_1 g09594(new_n9970, new_n9965, new_n9971);
xnor_1 g09595(new_n9971, new_n9944, new_n9972);
or_1   g09596(new_n9804, new_n9799, new_n9973);
nand_1 g09597(new_n9817, new_n9973, new_n9974);
nand_1 g09598(new_n9812, new_n9811, new_n9975);
not_1  g09599(new_n9975, new_n9976);
nor_1  g09600(new_n9813, new_n9810, new_n9977);
nor_1  g09601(new_n9977, new_n9976, new_n9978);
nand_1 g09602(n12069, n5694, new_n9979);
nand_1 g09603(n11153, n4903, new_n9980);
xnor_1 g09604(new_n9980, new_n9979, new_n9981);
nand_1 g09605(n7294, n5767, new_n9982);
nand_1 g09606(n8336, n783, new_n9983);
xnor_1 g09607(new_n9983, new_n9982, new_n9984);
xnor_1 g09608(new_n9984, new_n9981, new_n9985);
xnor_1 g09609(new_n9985, new_n9978, new_n9986);
nand_1 g09610(n4189, n4005, new_n9987);
nor_1  g09611(new_n915, new_n1562, new_n9988);
xnor_1 g09612(new_n9988, new_n9987, new_n9989);
xnor_1 g09613(new_n9989, new_n9986, new_n9990);
xnor_1 g09614(new_n9990, new_n9974, new_n9991);
xnor_1 g09615(new_n9991, new_n9972, new_n9992);
xnor_1 g09616(new_n9992, new_n9937, new_n9993);
xnor_1 g09617(new_n9993, new_n9934, new_n9994);
nand_1 g09618(new_n9864, new_n9834, new_n9995);
not_1  g09619(new_n9865, new_n9996);
nand_1 g09620(new_n9867, new_n9996, new_n9997);
nand_1 g09621(new_n9997, new_n9995, new_n9998);
not_1  g09622(new_n9796, new_n9999);
nand_1 g09623(new_n9827, new_n9999, new_n10000);
nand_1 g09624(new_n9832, new_n9828, new_n10001);
nand_1 g09625(new_n10001, new_n10000, new_n10002);
not_1  g09626(new_n9352, new_n10003);
nand_1 g09627(new_n9364, new_n10003, new_n10004);
nand_1 g09628(new_n10004, new_n9350, new_n10005);
nand_1 g09629(new_n9346, new_n9345, new_n10006);
not_1  g09630(new_n10006, new_n10007);
nor_1  g09631(new_n9347, new_n9344, new_n10008);
nor_1  g09632(new_n10008, new_n10007, new_n10009);
xnor_1 g09633(new_n10009, new_n10005, new_n10010);
nand_1 g09634(new_n9802, new_n9801, new_n10011);
not_1  g09635(new_n10011, new_n10012);
nor_1  g09636(new_n9803, new_n9800, new_n10013);
nor_1  g09637(new_n10013, new_n10012, new_n10014);
nand_1 g09638(new_n9859, new_n9858, new_n10015);
not_1  g09639(new_n10015, new_n10016);
nor_1  g09640(new_n9860, new_n9857, new_n10017);
nor_1  g09641(new_n10017, new_n10016, new_n10018);
xnor_1 g09642(new_n10018, new_n10014, new_n10019);
xnor_1 g09643(new_n10019, new_n10010, new_n10020);
xnor_1 g09644(new_n10020, new_n10002, new_n10021);
nand_1 g09645(new_n9371, new_n9323, new_n10022_1);
nand_1 g09646(new_n9372, new_n9340, new_n10023);
nand_1 g09647(new_n10023, new_n10022_1, new_n10024);
nand_1 g09648(new_n9861, new_n9855, new_n10025);
not_1  g09649(new_n9853, new_n10026);
nand_1 g09650(new_n9862, new_n10026, new_n10027);
nand_1 g09651(new_n10027, new_n10025, new_n10028);
nor_1  g09652(new_n8087, new_n667, new_n10029);
xnor_1 g09653(new_n10029, new_n10028, new_n10030);
xnor_1 g09654(new_n10030, new_n10024, new_n10031);
xnor_1 g09655(new_n10031, new_n10021, new_n10032);
nand_1 g09656(new_n9826, new_n9819, new_n10033);
nand_1 g09657(new_n10033, new_n9823, new_n10034);
nor_1  g09658(new_n9773, new_n9449, new_n10035);
not_1  g09659(new_n9774, new_n10036);
nor_1  g09660(new_n9779, new_n10036, new_n10037);
nor_1  g09661(new_n10037, new_n10035, new_n10038);
nand_1 g09662(new_n9769, new_n9768, new_n10039);
not_1  g09663(new_n10039, new_n10040);
nor_1  g09664(new_n9770, new_n9767_1, new_n10041);
nor_1  g09665(new_n10041, new_n10040, new_n10042);
nand_1 g09666(n5319, n1980, new_n10043);
nand_1 g09667(n9920, n2508, new_n10044);
nand_1 g09668(n10678, n1209, new_n10045);
xnor_1 g09669(new_n10045, new_n10044, new_n10046);
xnor_1 g09670(new_n10046, new_n10043, new_n10047);
xnor_1 g09671(new_n10047, new_n10042, new_n10048);
xnor_1 g09672(new_n10048, new_n10038, new_n10049);
xnor_1 g09673(new_n10049, new_n10034, new_n10050);
not_1  g09674(new_n9766, new_n10051);
nand_1 g09675(new_n9771, new_n10051, new_n10052);
not_1  g09676(new_n9780, new_n10053);
nand_1 g09677(new_n10053, new_n9772, new_n10054);
nand_1 g09678(new_n10054, new_n10052, new_n10055);
nand_1 g09679(new_n9777, new_n9776, new_n10056);
not_1  g09680(new_n10056, new_n10057);
nor_1  g09681(new_n9778, new_n9775, new_n10058);
nor_1  g09682(new_n10058, new_n10057, new_n10059);
nand_1 g09683(n4828, n2802, new_n10060);
nand_1 g09684(n10928, n8236, new_n10061);
nand_1 g09685(n5105, n1094, new_n10062);
xnor_1 g09686(new_n10062, new_n10061, new_n10063);
xnor_1 g09687(new_n10063, new_n10060, new_n10064);
xnor_1 g09688(new_n10064, new_n10059, new_n10065);
xnor_1 g09689(new_n10065, new_n10055, new_n10066);
xnor_1 g09690(new_n10066, new_n10050, new_n10067);
nand_1 g09691(new_n9842, new_n9841, new_n10068);
not_1  g09692(new_n9852, new_n10069);
nand_1 g09693(new_n10069, new_n9843, new_n10070);
nand_1 g09694(new_n10070, new_n10068, new_n10071);
nand_1 g09695(n7891, n5069, new_n10072);
not_1  g09696(n2087, new_n10073);
nor_1  g09697(new_n377, new_n10073, new_n10074);
xnor_1 g09698(new_n10074, new_n10072, new_n10075);
xnor_1 g09699(new_n10075, new_n10071, new_n10076);
nand_1 g09700(n7160, n6806, new_n10077);
nand_1 g09701(n6687, n615, new_n10078);
xnor_1 g09702(new_n10078, new_n10077, new_n10079);
xnor_1 g09703(new_n10079, new_n10076, new_n10080);
xnor_1 g09704(new_n10080, new_n10067, new_n10081);
nor_1  g09705(new_n9368, new_n9293, new_n10082);
not_1  g09706(new_n9370, new_n10083);
nor_1  g09707(new_n10083, new_n9365, new_n10084);
nor_1  g09708(new_n10084, new_n10082, new_n10085);
not_1  g09709(new_n9781, new_n10086);
nand_1 g09710(new_n9787, new_n10086, new_n10087);
nand_1 g09711(new_n10087, new_n9784, new_n10088);
nand_1 g09712(new_n9353, new_n9254, new_n10089);
nand_1 g09713(new_n9363, new_n9354, new_n10090);
nand_1 g09714(new_n10090, new_n10089, new_n10091);
nand_1 g09715(n7500, n7320, new_n10092);
nand_1 g09716(n12706, n2564, new_n10093);
nand_1 g09717(n6770, n2585, new_n10094);
xnor_1 g09718(new_n10094, new_n10093, new_n10095);
xnor_1 g09719(new_n10095, new_n10092, new_n10096);
xnor_1 g09720(new_n10096, new_n10091, new_n10097);
xnor_1 g09721(new_n10097, new_n10088, new_n10098);
xnor_1 g09722(new_n10098, new_n10085, new_n10099);
xnor_1 g09723(new_n10099, new_n10081, new_n10100);
xnor_1 g09724(new_n10100, new_n10032, new_n10101);
xnor_1 g09725(new_n10101, new_n9998, new_n10102);
xnor_1 g09726(new_n10102, new_n9994, new_n10103);
xnor_1 g09727(new_n10103, new_n9930, new_n10104);
xnor_1 g09728(new_n10104, new_n9920_1, n3654);
xnor_1 g09729(new_n9915, new_n9914, n3661);
nor_1  g09730(new_n4044, new_n456, new_n10107);
nor_1  g09731(new_n424, new_n4053, new_n10108);
nand_1 g09732(n1798, n1097, new_n10109);
nand_1 g09733(n12591, n5305, new_n10110);
nand_1 g09734(new_n10110, new_n10109, new_n10111);
nand_1 g09735(new_n10111, new_n10108, new_n10112);
nor_1  g09736(new_n10110, new_n10109, new_n10113);
not_1  g09737(new_n10113, new_n10114);
nand_1 g09738(new_n10114, new_n10112, new_n10115);
xnor_1 g09739(new_n10115, new_n10107, new_n10116);
nor_1  g09740(new_n4053, new_n419, new_n10117);
nand_1 g09741(n4312, n1798, new_n10118);
nand_1 g09742(n12591, n5964, new_n10119);
xnor_1 g09743(new_n10119, new_n10118, new_n10120);
xnor_1 g09744(new_n10120, new_n10117, new_n10121);
xnor_1 g09745(new_n10121, new_n10116, new_n10122);
not_1  g09746(new_n6511, new_n10123);
nor_1  g09747(new_n10123, new_n6510, new_n10124);
not_1  g09748(new_n10124, new_n10125);
and_1  g09749(new_n10114, new_n10111, new_n10126);
nor_1  g09750(new_n10126, new_n10125, new_n10127);
nand_1 g09751(new_n10127, new_n10122, new_n10128);
nor_1  g09752(new_n4665, new_n456, new_n10129);
not_1  g09753(new_n10129, new_n10130);
nor_1  g09754(new_n4044, new_n424, new_n10131);
nor_1  g09755(new_n395, new_n4053, new_n10132);
not_1  g09756(new_n10132, new_n10133);
nand_1 g09757(n12591, n1097, new_n10134);
nand_1 g09758(n12705, n1798, new_n10135);
xnor_1 g09759(new_n10135, new_n10134, new_n10136);
xnor_1 g09760(new_n10136, new_n10133, new_n10137);
xnor_1 g09761(new_n10137, new_n10131, new_n10138);
nand_1 g09762(new_n10119, new_n10118, new_n10139);
not_1  g09763(new_n10139, new_n10140);
nor_1  g09764(new_n10120, new_n10117, new_n10141);
nor_1  g09765(new_n10141, new_n10140, new_n10142);
xnor_1 g09766(new_n10142, new_n10138, new_n10143);
xnor_1 g09767(new_n10143, new_n10130, new_n10144);
nand_1 g09768(new_n10115, new_n10107, new_n10145);
not_1  g09769(new_n10145, new_n10146);
not_1  g09770(new_n10121, new_n10147);
nor_1  g09771(new_n10147, new_n10116, new_n10148);
nor_1  g09772(new_n10148, new_n10146, new_n10149);
xnor_1 g09773(new_n10149, new_n10144, new_n10150);
xor_1  g09774(new_n10150, new_n10128, new_n10151);
not_1  g09775(new_n10151, new_n10152);
xnor_1 g09776(new_n10127, new_n10122, new_n10153);
not_1  g09777(new_n10153, new_n10154);
nor_1  g09778(new_n4232, new_n552, new_n10155);
nand_1 g09779(n8759, n3022, new_n10156);
nand_1 g09780(n12299, n6703, new_n10157);
nand_1 g09781(new_n10157, new_n10156, new_n10158);
not_1  g09782(new_n10158, new_n10159);
nand_1 g09783(n12299, n3022, new_n10160);
nor_1  g09784(new_n10160, new_n6516, new_n10161);
nor_1  g09785(new_n4116, new_n563, new_n10162);
nor_1  g09786(new_n10162, new_n10161, new_n10163);
nor_1  g09787(new_n10163, new_n10159, new_n10164);
nand_1 g09788(new_n10164, new_n10155, new_n10165);
not_1  g09789(new_n10165, new_n10166);
nor_1  g09790(new_n10164, new_n10155, new_n10167);
nor_1  g09791(new_n10167, new_n10166, new_n10168);
nor_1  g09792(new_n554, new_n4116, new_n10169);
nand_1 g09793(n6776, n3022, new_n10170);
nand_1 g09794(n7436, n6703, new_n10171);
nand_1 g09795(new_n10171, new_n10170, new_n10172);
not_1  g09796(new_n10172, new_n10173);
nor_1  g09797(new_n10171, new_n10170, new_n10174_1);
nor_1  g09798(new_n10174_1, new_n10173, new_n10175);
xor_1  g09799(new_n10175, new_n10169, new_n10176);
nand_1 g09800(new_n10176, new_n10168, new_n10177);
not_1  g09801(new_n10177, new_n10178);
nor_1  g09802(new_n10176, new_n10168, new_n10179);
nor_1  g09803(new_n10179, new_n10178, new_n10180);
not_1  g09804(new_n10162, new_n10181);
nor_1  g09805(new_n10181, new_n6500, new_n10182);
nor_1  g09806(new_n10161, new_n10159, new_n10183);
nor_1  g09807(new_n10183, new_n10182, new_n10184);
not_1  g09808(new_n10184, new_n10185);
nor_1  g09809(new_n10185, new_n10181, new_n10186);
nor_1  g09810(new_n10186, new_n10180, new_n10187);
nand_1 g09811(new_n10186, new_n10180, new_n10188);
not_1  g09812(new_n10188, new_n10189);
nor_1  g09813(new_n10189, new_n10187, new_n10190);
nor_1  g09814(new_n4187_1, new_n668, new_n10191);
nor_1  g09815(new_n740, new_n4919, new_n10192);
nand_1 g09816(n8665, n8476, new_n10193);
nand_1 g09817(n12648, n5645, new_n10194);
nand_1 g09818(new_n10194, new_n10193, new_n10195);
nor_1  g09819(new_n10194, new_n10193, new_n10196);
not_1  g09820(new_n10196, new_n10197);
nand_1 g09821(new_n10197, new_n10195, new_n10198);
xnor_1 g09822(new_n10198, new_n10192, new_n10199);
xnor_1 g09823(new_n10199, new_n10191, new_n10200);
nand_1 g09824(n8665, n5331, new_n10201);
nand_1 g09825(n5645, n2530, new_n10202);
nand_1 g09826(new_n10202, new_n10201, new_n10203);
not_1  g09827(new_n10203, new_n10204);
nor_1  g09828(new_n712, new_n4919, new_n10205);
nor_1  g09829(new_n4132, new_n740, new_n10206);
not_1  g09830(new_n10206, new_n10207);
nor_1  g09831(new_n10207, new_n6501, new_n10208);
nor_1  g09832(new_n10208, new_n10205, new_n10209);
nor_1  g09833(new_n10209, new_n10204, new_n10210);
xnor_1 g09834(new_n10210, new_n10200, new_n10211);
nor_1  g09835(new_n10208, new_n10204, new_n10212);
nor_1  g09836(new_n10212, new_n6532, new_n10213);
nor_1  g09837(new_n10213, new_n10211, new_n10214);
nand_1 g09838(new_n10213, new_n10211, new_n10215);
not_1  g09839(new_n10215, new_n10216);
nor_1  g09840(new_n10216, new_n10214, new_n10217_1);
nor_1  g09841(new_n754, new_n4204, new_n10218);
nand_1 g09842(n7965, n3754, new_n10219);
nand_1 g09843(n11892, n11876, new_n10220);
nand_1 g09844(new_n10220, new_n10219, new_n10221);
not_1  g09845(new_n10221, new_n10222);
nor_1  g09846(new_n762, new_n5052, new_n10223_1);
not_1  g09847(new_n10223_1, new_n10224);
nor_1  g09848(new_n10224, new_n6502, new_n10225);
nor_1  g09849(new_n4143, new_n696, new_n10226);
nor_1  g09850(new_n10226, new_n10225, new_n10227);
nor_1  g09851(new_n10227, new_n10222, new_n10228);
nand_1 g09852(new_n10228, new_n10218, new_n10229);
not_1  g09853(new_n10229, new_n10230);
nor_1  g09854(new_n10228, new_n10218, new_n10231);
nor_1  g09855(new_n10231, new_n10230, new_n10232);
nor_1  g09856(new_n762, new_n4143, new_n10233);
nand_1 g09857(n7388, n3754, new_n10234);
nand_1 g09858(n11876, n2393, new_n10235);
xnor_1 g09859(new_n10235, new_n10234, new_n10236);
xnor_1 g09860(new_n10236, new_n10233, new_n10237);
xnor_1 g09861(new_n10237, new_n10232, new_n10238);
nand_1 g09862(new_n10226, new_n6502, new_n10239);
not_1  g09863(new_n10239, new_n10240);
nor_1  g09864(new_n10225, new_n10222, new_n10241);
nor_1  g09865(new_n10241, new_n10240, new_n10242);
nand_1 g09866(new_n10242, new_n10226, new_n10243);
nor_1  g09867(new_n10243, new_n10238, new_n10244);
not_1  g09868(new_n10244, new_n10245);
nand_1 g09869(new_n10243, new_n10238, new_n10246);
nand_1 g09870(new_n10246, new_n10245, new_n10247);
xnor_1 g09871(new_n10247, new_n10217_1, new_n10248);
not_1  g09872(new_n10248, new_n10249);
not_1  g09873(new_n10242, new_n10250);
nand_1 g09874(new_n10240, new_n10221, new_n10251);
nand_1 g09875(new_n10251, new_n10250, new_n10252);
nor_1  g09876(new_n6526, new_n6504, new_n10253);
nor_1  g09877(new_n6537, new_n10253, new_n10254);
nand_1 g09878(new_n10254, new_n10252, new_n10255);
xnor_1 g09879(new_n10254, new_n10252, new_n10256);
not_1  g09880(new_n10256, new_n10257);
nand_1 g09881(new_n10205, new_n6501, new_n10258);
nor_1  g09882(new_n10258, new_n10203, new_n10259);
and_1  g09883(new_n10258, new_n10212, new_n10260);
nor_1  g09884(new_n10260, new_n10259, new_n10261);
nand_1 g09885(new_n10261, new_n10257, new_n10262);
nand_1 g09886(new_n10262, new_n10255, new_n10263);
xnor_1 g09887(new_n10263, new_n10249, new_n10264);
xnor_1 g09888(new_n10264, new_n10190, new_n10265);
nand_1 g09889(new_n10182, new_n10158, new_n10266);
nand_1 g09890(new_n10266, new_n10185, new_n10267);
nor_1  g09891(new_n6521, new_n6518, new_n10268);
nor_1  g09892(new_n6540, new_n10268, new_n10269);
nand_1 g09893(new_n10269, new_n10267, new_n10270);
xnor_1 g09894(new_n10261, new_n10256, new_n10271);
not_1  g09895(new_n10269, new_n10272);
xnor_1 g09896(new_n10272, new_n10267, new_n10273);
nand_1 g09897(new_n10273, new_n10271, new_n10274);
nand_1 g09898(new_n10274, new_n10270, new_n10275);
xnor_1 g09899(new_n10275, new_n10265, new_n10276);
nand_1 g09900(new_n10276, new_n10154, new_n10277);
not_1  g09901(new_n10277, new_n10278_1);
xnor_1 g09902(new_n10276, new_n10154, new_n10279);
xnor_1 g09903(new_n10273, new_n10271, new_n10280);
not_1  g09904(new_n6499, new_n10281);
nand_1 g09905(new_n10108, new_n10281, new_n10282);
nor_1  g09906(new_n10282, new_n10111, new_n10283);
nand_1 g09907(new_n10282, new_n10126, new_n10284);
not_1  g09908(new_n10284, new_n10285);
nor_1  g09909(new_n10285, new_n10283, new_n10286);
not_1  g09910(new_n10286, new_n10287);
nor_1  g09911(new_n10287, new_n10280, new_n10288);
nor_1  g09912(new_n6513, new_n6508, new_n10289);
nor_1  g09913(new_n6544, new_n10289, new_n10290);
not_1  g09914(new_n10290, new_n10291);
xnor_1 g09915(new_n10287, new_n10280, new_n10292);
nor_1  g09916(new_n10292, new_n10291, new_n10293);
nor_1  g09917(new_n10293, new_n10288, new_n10294);
not_1  g09918(new_n10294, new_n10295);
nor_1  g09919(new_n10295, new_n10279, new_n10296);
nor_1  g09920(new_n10296, new_n10278_1, new_n10297);
xnor_1 g09921(new_n10297, new_n10152, new_n10298);
nor_1  g09922(new_n4815, new_n552, new_n10299);
not_1  g09923(new_n10299, new_n10300);
nand_1 g09924(n11023, n6776, new_n10301);
nor_1  g09925(new_n10174_1, new_n10169, new_n10302);
nor_1  g09926(new_n10302, new_n10173, new_n10303);
xnor_1 g09927(new_n10303, new_n10301, new_n10304);
nor_1  g09928(new_n4116, new_n599, new_n10305);
nand_1 g09929(n8276, n6703, new_n10306);
nand_1 g09930(new_n10306, new_n10160, new_n10307);
not_1  g09931(new_n10160, new_n10308);
not_1  g09932(new_n10306, new_n10309);
nand_1 g09933(new_n10309, new_n10308, new_n10310);
nand_1 g09934(new_n10310, new_n10307, new_n10311);
xnor_1 g09935(new_n10311, new_n10305, new_n10312);
xor_1  g09936(new_n10312, new_n10304, new_n10313);
xnor_1 g09937(new_n10313, new_n10300, new_n10314);
nor_1  g09938(new_n10178, new_n10166, new_n10315);
not_1  g09939(new_n10315, new_n10316);
nor_1  g09940(new_n10316, new_n10314, new_n10317);
nand_1 g09941(new_n10316, new_n10314, new_n10318);
not_1  g09942(new_n10318, new_n10319);
nor_1  g09943(new_n10319, new_n10317, new_n10320);
nand_1 g09944(new_n10320, new_n10189, new_n10321);
not_1  g09945(new_n10320, new_n10322);
nand_1 g09946(new_n10322, new_n10188, new_n10323);
nand_1 g09947(new_n10323, new_n10321, new_n10324);
nor_1  g09948(new_n754, new_n5065, new_n10325);
nand_1 g09949(new_n10237, new_n10232, new_n10326);
nand_1 g09950(new_n10326, new_n10229, new_n10327_1);
xnor_1 g09951(new_n10327_1, new_n10325, new_n10328);
nor_1  g09952(new_n696, new_n4204, new_n10329);
nand_1 g09953(new_n10235, new_n10234, new_n10330);
not_1  g09954(new_n10330, new_n10331);
nor_1  g09955(new_n10236, new_n10233, new_n10332);
nor_1  g09956(new_n10332, new_n10331, new_n10333);
xnor_1 g09957(new_n10333, new_n10329, new_n10334);
not_1  g09958(new_n10334, new_n10335);
nand_1 g09959(n11876, n5860, new_n10336);
nand_1 g09960(n10898, n2393, new_n10337);
xnor_1 g09961(new_n10337, new_n10336, new_n10338);
nand_1 g09962(new_n10338, new_n10223_1, new_n10339);
nor_1  g09963(new_n10338, new_n10223_1, new_n10340);
not_1  g09964(new_n10340, new_n10341);
nand_1 g09965(new_n10341, new_n10339, new_n10342);
nand_1 g09966(new_n10342, new_n10335, new_n10343);
not_1  g09967(new_n10342, new_n10344);
nand_1 g09968(new_n10344, new_n10334, new_n10345);
nand_1 g09969(new_n10345, new_n10343, new_n10346);
not_1  g09970(new_n10346, new_n10347);
xnor_1 g09971(new_n10347, new_n10328, new_n10348);
nand_1 g09972(new_n10348, new_n10244, new_n10349);
not_1  g09973(new_n10349, new_n10350);
nor_1  g09974(new_n10348, new_n10244, new_n10351);
nor_1  g09975(new_n10351, new_n10350, new_n10352);
nor_1  g09976(new_n668, new_n4951, new_n10353);
nor_1  g09977(new_n4187_1, new_n712, new_n10354);
not_1  g09978(new_n10195, new_n10355);
nor_1  g09979(new_n10196, new_n10192, new_n10356);
nor_1  g09980(new_n10356, new_n10355, new_n10357);
nand_1 g09981(new_n10357, new_n10354, new_n10358);
not_1  g09982(new_n10358, new_n10359);
nor_1  g09983(new_n10357, new_n10354, new_n10360);
nor_1  g09984(new_n10360, new_n10359, new_n10361);
nor_1  g09985(new_n829, new_n4919, new_n10362);
nor_1  g09986(new_n5668, new_n4195, new_n10363);
not_1  g09987(new_n10363, new_n10364);
nand_1 g09988(new_n10364, new_n10207, new_n10365);
nor_1  g09989(new_n10364, new_n10207, new_n10366);
not_1  g09990(new_n10366, new_n10367);
nand_1 g09991(new_n10367, new_n10365, new_n10368);
xnor_1 g09992(new_n10368, new_n10362, new_n10369);
nand_1 g09993(new_n10369, new_n10361, new_n10370);
not_1  g09994(new_n10370, new_n10371);
nor_1  g09995(new_n10369, new_n10361, new_n10372);
nor_1  g09996(new_n10372, new_n10371, new_n10373);
nand_1 g09997(new_n10373, new_n10353, new_n10374);
not_1  g09998(new_n10374, new_n10375);
nor_1  g09999(new_n10373, new_n10353, new_n10376);
nor_1  g10000(new_n10376, new_n10375, new_n10377);
not_1  g10001(new_n10191, new_n10378);
not_1  g10002(new_n10199, new_n10379);
nor_1  g10003(new_n10379, new_n10378, new_n10380);
not_1  g10004(new_n10210, new_n10381);
nor_1  g10005(new_n10381, new_n10200, new_n10382);
nor_1  g10006(new_n10382, new_n10380, new_n10383);
xnor_1 g10007(new_n10383, new_n10377, new_n10384);
nand_1 g10008(new_n10384, new_n10216, new_n10385);
not_1  g10009(new_n10385, new_n10386);
nor_1  g10010(new_n10384, new_n10216, new_n10387);
nor_1  g10011(new_n10387, new_n10386, new_n10388);
nand_1 g10012(new_n10388, new_n10352, new_n10389);
not_1  g10013(new_n10352, new_n10390);
not_1  g10014(new_n10388, new_n10391_1);
nand_1 g10015(new_n10391_1, new_n10390, new_n10392);
nand_1 g10016(new_n10392, new_n10389, new_n10393);
not_1  g10017(new_n10217_1, new_n10394);
nand_1 g10018(new_n10247, new_n10394, new_n10395);
nand_1 g10019(new_n10263, new_n10248, new_n10396);
nand_1 g10020(new_n10396, new_n10395, new_n10397);
xnor_1 g10021(new_n10397, new_n10393, new_n10398);
xnor_1 g10022(new_n10398, new_n10324, new_n10399);
not_1  g10023(new_n10190, new_n10400);
nand_1 g10024(new_n10264, new_n10400, new_n10401);
nand_1 g10025(new_n10275, new_n10265, new_n10402);
nand_1 g10026(new_n10402, new_n10401, new_n10403);
xnor_1 g10027(new_n10403, new_n10399, new_n10404);
xor_1  g10028(new_n10404, new_n10298, n3677);
xnor_1 g10029(new_n9050, new_n9049, n3849);
xnor_1 g10030(new_n6495, new_n6493, n4088);
xnor_1 g10031(new_n1259, new_n1127, n4155);
not_1  g10032(new_n3150, new_n10409);
xnor_1 g10033(new_n10409, new_n3149, n4159);
xnor_1 g10034(new_n6481, new_n6284, n4226);
nor_1  g10035(new_n4627, new_n395, new_n10412);
not_1  g10036(new_n10412, new_n10413);
nand_1 g10037(new_n10135, new_n10134, new_n10414);
not_1  g10038(new_n10414, new_n10415);
nor_1  g10039(new_n10136, new_n10132, new_n10416);
nor_1  g10040(new_n10416, new_n10415, new_n10417);
xnor_1 g10041(new_n10417, new_n10413, new_n10418);
nor_1  g10042(new_n8505, new_n4053, new_n10419);
not_1  g10043(new_n10419, new_n10420);
nor_1  g10044(new_n511, new_n4682, new_n10421);
not_1  g10045(new_n10421, new_n10422);
nand_1 g10046(new_n10422, new_n10420, new_n10423);
nor_1  g10047(new_n10422, new_n10420, new_n10424);
not_1  g10048(new_n10424, new_n10425);
nand_1 g10049(new_n10425, new_n10423, new_n10426);
xnor_1 g10050(new_n10426, new_n10418, new_n10427);
nor_1  g10051(new_n4665, new_n424, new_n10428);
not_1  g10052(new_n10428, new_n10429);
nor_1  g10053(new_n4044, new_n419, new_n10430);
not_1  g10054(new_n10430, new_n10431);
nor_1  g10055(new_n10431, new_n10429, new_n10432);
not_1  g10056(new_n10432, new_n10433);
nand_1 g10057(new_n10431, new_n10429, new_n10434);
nand_1 g10058(new_n10434, new_n10433, new_n10435);
xnor_1 g10059(new_n10435, new_n10427, new_n10436);
not_1  g10060(new_n10131, new_n10437);
nor_1  g10061(new_n10137, new_n10437, new_n10438);
not_1  g10062(new_n10438, new_n10439_1);
nand_1 g10063(new_n10142, new_n10138, new_n10440);
nand_1 g10064(new_n10440, new_n10439_1, new_n10441);
nand_1 g10065(new_n10441, new_n10436, new_n10442);
not_1  g10066(new_n10442, new_n10443);
nor_1  g10067(new_n10441, new_n10436, new_n10444);
nor_1  g10068(new_n10444, new_n10443, new_n10445);
nor_1  g10069(new_n10143, new_n10130, new_n10446);
nor_1  g10070(new_n10149, new_n10144, new_n10447);
nor_1  g10071(new_n10447, new_n10446, new_n10448);
not_1  g10072(new_n10448, new_n10449);
nand_1 g10073(new_n10449, new_n10445, new_n10450);
not_1  g10074(new_n10417, new_n10451_1);
nand_1 g10075(new_n10451_1, new_n10413, new_n10452);
nand_1 g10076(new_n10426, new_n10418, new_n10453);
nand_1 g10077(new_n10453, new_n10452, new_n10454);
nor_1  g10078(new_n4709, new_n424, new_n10455);
nand_1 g10079(n11662, n1097, new_n10456);
nand_1 g10080(n9583, n5305, new_n10457);
xnor_1 g10081(new_n10457, new_n10456, new_n10458);
xnor_1 g10082(new_n10458, new_n10455, new_n10459);
xnor_1 g10083(new_n10459, new_n10454, new_n10460);
nor_1  g10084(new_n4044, new_n395, new_n10461);
not_1  g10085(new_n10461, new_n10462);
nand_1 g10086(new_n10462, new_n10425, new_n10463);
nand_1 g10087(new_n10461, new_n10424, new_n10464);
nand_1 g10088(new_n10464, new_n10463, new_n10465);
nor_1  g10089(new_n511, new_n4053, new_n10466);
nand_1 g10090(n12705, n12591, new_n10467);
nand_1 g10091(n11257, n1798, new_n10468);
xnor_1 g10092(new_n10468, new_n10467, new_n10469);
xor_1  g10093(new_n10469, new_n10466, new_n10470);
xnor_1 g10094(new_n10470, new_n10465, new_n10471);
xnor_1 g10095(new_n10471, new_n10460, new_n10472);
not_1  g10096(new_n10472, new_n10473);
not_1  g10097(new_n10435, new_n10474);
nand_1 g10098(new_n10474, new_n10427, new_n10475);
nand_1 g10099(new_n10443, new_n10432, new_n10476_1);
nand_1 g10100(new_n10442, new_n10433, new_n10477);
nand_1 g10101(new_n10477, new_n10476_1, new_n10478);
nand_1 g10102(new_n10478, new_n10475, new_n10479);
xnor_1 g10103(new_n10479, new_n10473, new_n10480);
xnor_1 g10104(new_n10480, new_n10450, new_n10481);
nor_1  g10105(new_n4709, new_n456, new_n10482);
not_1  g10106(new_n10450, new_n10483);
nor_1  g10107(new_n10449, new_n10445, new_n10484);
nor_1  g10108(new_n10484, new_n10483, new_n10485);
nor_1  g10109(new_n10485, new_n10482, new_n10486);
nor_1  g10110(new_n10150, new_n10128, new_n10487);
xnor_1 g10111(new_n10485, new_n10482, new_n10488);
nor_1  g10112(new_n10488, new_n10487, new_n10489);
nor_1  g10113(new_n10489, new_n10486, new_n10490);
xor_1  g10114(new_n10490, new_n10481, new_n10491);
not_1  g10115(new_n10491, new_n10492);
not_1  g10116(new_n10301, new_n10493);
nand_1 g10117(new_n10303, new_n10493, new_n10494);
nand_1 g10118(new_n10312, new_n10304, new_n10495);
nand_1 g10119(new_n10495, new_n10494, new_n10496);
nor_1  g10120(new_n4815, new_n563, new_n10497);
not_1  g10121(new_n10497, new_n10498);
nor_1  g10122(new_n554, new_n4232, new_n10499);
not_1  g10123(new_n10499, new_n10500);
nor_1  g10124(new_n10500, new_n10498, new_n10501);
not_1  g10125(new_n10501, new_n10502);
nand_1 g10126(new_n10500, new_n10498, new_n10503);
nand_1 g10127(new_n10503, new_n10502, new_n10504);
xnor_1 g10128(new_n10504, new_n10496, new_n10505);
nor_1  g10129(new_n599, new_n4761, new_n10506);
nand_1 g10130(n9640, n8276, new_n10507);
nand_1 g10131(n9241, n6703, new_n10508);
xnor_1 g10132(new_n10508, new_n10507, new_n10509);
xnor_1 g10133(new_n10509, new_n10506, new_n10510_1);
not_1  g10134(new_n10307, new_n10511);
not_1  g10135(new_n10310, new_n10512);
nor_1  g10136(new_n10512, new_n10305, new_n10513);
nor_1  g10137(new_n10513, new_n10511, new_n10514);
xnor_1 g10138(new_n10514, new_n10510_1, new_n10515);
not_1  g10139(new_n10515, new_n10516);
nand_1 g10140(new_n10516, new_n10505, new_n10517);
not_1  g10141(new_n10517, new_n10518);
nor_1  g10142(new_n10516, new_n10505, new_n10519);
nor_1  g10143(new_n10519, new_n10518, new_n10520);
nand_1 g10144(new_n10313, new_n10299, new_n10521);
nand_1 g10145(new_n10318, new_n10521, new_n10522);
nand_1 g10146(new_n10522, new_n10520, new_n10523);
not_1  g10147(new_n10506, new_n10524);
nand_1 g10148(new_n10509, new_n10524, new_n10525);
not_1  g10149(new_n10514, new_n10526);
nand_1 g10150(new_n10526, new_n10510_1, new_n10527);
nand_1 g10151(new_n10527, new_n10525, new_n10528);
nor_1  g10152(new_n4852, new_n563, new_n10529);
nand_1 g10153(n12299, n10451, new_n10530);
nand_1 g10154(n11423, n8759, new_n10531);
xnor_1 g10155(new_n10531, new_n10530, new_n10532);
xor_1  g10156(new_n10532, new_n10529, new_n10533);
xnor_1 g10157(new_n10533, new_n10528, new_n10534);
not_1  g10158(new_n10534, new_n10535);
nor_1  g10159(new_n10508, new_n10507, new_n10536);
nor_1  g10160(new_n4232, new_n599, new_n10537);
xor_1  g10161(new_n10537, new_n10536, new_n10538);
nor_1  g10162(new_n4116, new_n2723, new_n10539);
nand_1 g10163(n8276, n3022, new_n10540);
nand_1 g10164(n10510, n6703, new_n10541);
xnor_1 g10165(new_n10541, new_n10540, new_n10542);
xor_1  g10166(new_n10542, new_n10539, new_n10543);
xnor_1 g10167(new_n10543, new_n10538, new_n10544);
not_1  g10168(new_n10544, new_n10545_1);
nand_1 g10169(new_n10545_1, new_n10535, new_n10546);
nand_1 g10170(new_n10544, new_n10534, new_n10547_1);
nand_1 g10171(new_n10547_1, new_n10546, new_n10548);
not_1  g10172(new_n10504, new_n10549);
nand_1 g10173(new_n10549, new_n10496, new_n10550);
nand_1 g10174(new_n10518, new_n10501, new_n10551);
nand_1 g10175(new_n10517, new_n10502, new_n10552);
nand_1 g10176(new_n10552, new_n10551, new_n10553);
nand_1 g10177(new_n10553, new_n10550, new_n10554);
xnor_1 g10178(new_n10554, new_n10548, new_n10555);
not_1  g10179(new_n10555, new_n10556);
xnor_1 g10180(new_n10556, new_n10523, new_n10557);
nor_1  g10181(new_n4852, new_n552, new_n10558);
not_1  g10182(new_n10520, new_n10559);
xnor_1 g10183(new_n10522, new_n10559, new_n10560);
nand_1 g10184(new_n10560, new_n10558, new_n10561);
not_1  g10185(new_n10321, new_n10562);
not_1  g10186(new_n10558, new_n10563);
xnor_1 g10187(new_n10560, new_n10563, new_n10564);
nand_1 g10188(new_n10564, new_n10562, new_n10565);
nand_1 g10189(new_n10565, new_n10561, new_n10566);
xnor_1 g10190(new_n10566, new_n10557, new_n10567);
nand_1 g10191(n12648, n8665, new_n10568);
not_1  g10192(new_n10568, new_n10569);
nand_1 g10193(n10545, n1067, new_n10570);
nand_1 g10194(n7690, n5645, new_n10571);
xnor_1 g10195(new_n10571, new_n10570, new_n10572);
xnor_1 g10196(new_n10572, new_n10569, new_n10573);
not_1  g10197(new_n10365, new_n10574);
nor_1  g10198(new_n10366, new_n10362, new_n10575);
nor_1  g10199(new_n10575, new_n10574, new_n10576);
nand_1 g10200(new_n10576, new_n10573, new_n10577);
not_1  g10201(new_n10577, new_n10578);
nor_1  g10202(new_n10576, new_n10573, new_n10579);
nor_1  g10203(new_n10579, new_n10578, new_n10580);
nand_1 g10204(n8476, n2551, new_n10581);
nand_1 g10205(n11922, n2530, new_n10582);
nor_1  g10206(new_n10582, new_n10581, new_n10583);
not_1  g10207(new_n10583, new_n10584);
nand_1 g10208(new_n10582, new_n10581, new_n10585);
nand_1 g10209(new_n10585, new_n10584, new_n10586);
xnor_1 g10210(new_n10586, new_n10580, new_n10587);
nand_1 g10211(new_n10370, new_n10358, new_n10588);
xnor_1 g10212(new_n10588, new_n10587, new_n10589_1);
not_1  g10213(new_n10589_1, new_n10590);
not_1  g10214(new_n10383, new_n10591);
nand_1 g10215(new_n10591, new_n10377, new_n10592);
nand_1 g10216(new_n10592, new_n10374, new_n10593);
nand_1 g10217(new_n10593, new_n10590, new_n10594);
not_1  g10218(new_n10594, new_n10595);
nor_1  g10219(new_n10571, new_n10570, new_n10596);
nor_1  g10220(new_n829, new_n4187_1, new_n10597);
xnor_1 g10221(new_n10597, new_n10596, new_n10598);
not_1  g10222(new_n10598, new_n10599);
nor_1  g10223(new_n1048, new_n4919, new_n10600);
nand_1 g10224(n10545, n8665, new_n10601);
nand_1 g10225(n5645, n3616, new_n10602);
xnor_1 g10226(new_n10602, new_n10601, new_n10603);
xnor_1 g10227(new_n10603, new_n10600, new_n10604);
xnor_1 g10228(new_n10604, new_n10599, new_n10605);
nor_1  g10229(new_n10572, new_n10568, new_n10606);
not_1  g10230(new_n10606, new_n10607);
nand_1 g10231(new_n10577, new_n10607, new_n10608);
nor_1  g10232(new_n4908, new_n712, new_n10609);
not_1  g10233(new_n10609, new_n10610);
nand_1 g10234(n2551, n2530, new_n10611);
nand_1 g10235(n5331, n4094, new_n10612);
xnor_1 g10236(new_n10612, new_n10611, new_n10613);
xnor_1 g10237(new_n10613, new_n10610, new_n10614);
xnor_1 g10238(new_n10614, new_n10608, new_n10615);
xnor_1 g10239(new_n10615, new_n10605, new_n10616);
not_1  g10240(new_n10616, new_n10617);
not_1  g10241(new_n10586, new_n10618);
nand_1 g10242(new_n10618, new_n10580, new_n10619);
nand_1 g10243(new_n10588, new_n10587, new_n10620);
not_1  g10244(new_n10620, new_n10621);
nand_1 g10245(new_n10621, new_n10583, new_n10622);
nand_1 g10246(new_n10620, new_n10584, new_n10623);
nand_1 g10247(new_n10623, new_n10622, new_n10624);
nand_1 g10248(new_n10624, new_n10619, new_n10625);
xnor_1 g10249(new_n10625, new_n10617, new_n10626);
xnor_1 g10250(new_n10626, new_n10595, new_n10627);
nand_1 g10251(n12826, n5331, new_n10628);
nor_1  g10252(new_n10593, new_n10590, new_n10629);
nor_1  g10253(new_n10629, new_n10595, new_n10630);
not_1  g10254(new_n10630, new_n10631);
nand_1 g10255(new_n10631, new_n10628, new_n10632);
xnor_1 g10256(new_n10630, new_n10628, new_n10633);
nand_1 g10257(new_n10633, new_n10385, new_n10634);
nand_1 g10258(new_n10634, new_n10632, new_n10635);
xnor_1 g10259(new_n10635, new_n10627, new_n10636);
nor_1  g10260(new_n754, new_n5107, new_n10637);
nand_1 g10261(new_n10333, new_n10329, new_n10638);
nand_1 g10262(new_n10343, new_n10638, new_n10639);
nand_1 g10263(n7388, n159, new_n10640);
nand_1 g10264(n11892, n2749, new_n10641);
xnor_1 g10265(new_n10641, new_n10640, new_n10642);
xnor_1 g10266(new_n10642, new_n10639, new_n10643);
nor_1  g10267(new_n5052, new_n767, new_n10644_1);
nand_1 g10268(n10898, n5860, new_n10645);
nand_1 g10269(n11876, n3986, new_n10646);
nand_1 g10270(new_n10646, new_n10645, new_n10647);
not_1  g10271(new_n10647, new_n10648);
nor_1  g10272(new_n10646, new_n10645, new_n10649);
nor_1  g10273(new_n10649, new_n10648, new_n10650);
nand_1 g10274(new_n10650, new_n10644_1, new_n10651);
not_1  g10275(new_n10651, new_n10652);
nor_1  g10276(new_n10650, new_n10644_1, new_n10653);
nor_1  g10277(new_n10653, new_n10652, new_n10654);
nand_1 g10278(new_n10337, new_n10336, new_n10655);
not_1  g10279(new_n10655, new_n10656);
nor_1  g10280(new_n10340, new_n10656, new_n10657);
xnor_1 g10281(new_n10657, new_n10654, new_n10658);
xnor_1 g10282(new_n10658, new_n10643, new_n10659);
nand_1 g10283(new_n10327_1, new_n10325, new_n10660);
not_1  g10284(new_n10660, new_n10661);
nor_1  g10285(new_n10346, new_n10328, new_n10662);
nor_1  g10286(new_n10662, new_n10661, new_n10663);
xnor_1 g10287(new_n10663, new_n10659, new_n10664);
nand_1 g10288(new_n10664, new_n10637, new_n10665);
not_1  g10289(new_n10637, new_n10666);
xnor_1 g10290(new_n10664, new_n10666, new_n10667);
nand_1 g10291(new_n10667, new_n10350, new_n10668);
nand_1 g10292(new_n10668, new_n10665, new_n10669);
not_1  g10293(new_n10659, new_n10670);
nor_1  g10294(new_n10663, new_n10670, new_n10671);
nor_1  g10295(new_n10641, new_n10640, new_n10672);
not_1  g10296(new_n10639, new_n10673);
nand_1 g10297(new_n10642, new_n10673, new_n10674);
nand_1 g10298(new_n10658, new_n10643, new_n10675);
nand_1 g10299(new_n10675, new_n10674, new_n10676);
xnor_1 g10300(new_n10676, new_n10672, new_n10677);
nor_1  g10301(new_n696, new_n5107, new_n10678_1);
nand_1 g10302(n11892, n159, new_n10679);
nand_1 g10303(n12247, n7965, new_n10680);
xnor_1 g10304(new_n10680, new_n10679, new_n10681);
nor_1  g10305(new_n10681, new_n10678_1, new_n10682);
and_1  g10306(new_n10681, new_n10678_1, new_n10683);
nor_1  g10307(new_n10683, new_n10682, new_n10684);
nand_1 g10308(new_n10657, new_n10654, new_n10685_1);
nand_1 g10309(new_n10685_1, new_n10651, new_n10686);
xnor_1 g10310(new_n10686, new_n10684, new_n10687);
nand_1 g10311(n2749, n2393, new_n10688);
xnor_1 g10312(new_n10688, new_n10649, new_n10689);
nor_1  g10313(new_n4143, new_n1084, new_n10690);
nand_1 g10314(n11876, n5857, new_n10691);
nand_1 g10315(n5860, n3754, new_n10692);
xnor_1 g10316(new_n10692, new_n10691, new_n10693);
and_1  g10317(new_n10693, new_n10690, new_n10694);
nor_1  g10318(new_n10693, new_n10690, new_n10695_1);
nor_1  g10319(new_n10695_1, new_n10694, new_n10696);
xnor_1 g10320(new_n10696, new_n10689, new_n10697);
xnor_1 g10321(new_n10697, new_n10687, new_n10698);
xnor_1 g10322(new_n10698, new_n10677, new_n10699);
xnor_1 g10323(new_n10699, new_n10671, new_n10700);
xnor_1 g10324(new_n10700, new_n10669, new_n10701);
not_1  g10325(new_n10701, new_n10702);
xnor_1 g10326(new_n10702, new_n10636, new_n10703);
xnor_1 g10327(new_n10667, new_n10349, new_n10704);
not_1  g10328(new_n10704, new_n10705);
xnor_1 g10329(new_n10633, new_n10386, new_n10706);
nand_1 g10330(new_n10706, new_n10705, new_n10707);
not_1  g10331(new_n10393, new_n10708);
nand_1 g10332(new_n10397, new_n10708, new_n10709);
nand_1 g10333(new_n10709, new_n10392, new_n10710);
xnor_1 g10334(new_n10706, new_n10704, new_n10711);
nand_1 g10335(new_n10711, new_n10710, new_n10712);
nand_1 g10336(new_n10712, new_n10707, new_n10713);
xnor_1 g10337(new_n10713, new_n10703, new_n10714);
xnor_1 g10338(new_n10714, new_n10567, new_n10715);
xnor_1 g10339(new_n10564, new_n10562, new_n10716);
xnor_1 g10340(new_n10706, new_n10705, new_n10717);
xnor_1 g10341(new_n10717, new_n10710, new_n10718);
nand_1 g10342(new_n10718, new_n10716, new_n10719);
nor_1  g10343(new_n10398, new_n10324, new_n10720);
nor_1  g10344(new_n10403, new_n10399, new_n10721);
nor_1  g10345(new_n10721, new_n10720, new_n10722);
xnor_1 g10346(new_n10564, new_n10321, new_n10723);
xnor_1 g10347(new_n10718, new_n10723, new_n10724);
nand_1 g10348(new_n10724, new_n10722, new_n10725);
nand_1 g10349(new_n10725, new_n10719, new_n10726);
xnor_1 g10350(new_n10726, new_n10715, new_n10727);
nand_1 g10351(new_n10727, new_n10492, new_n10728);
xnor_1 g10352(new_n10727, new_n10491, new_n10729);
not_1  g10353(new_n10487, new_n10730);
xnor_1 g10354(new_n10488, new_n10730, new_n10731);
xnor_1 g10355(new_n10718, new_n10716, new_n10732);
xnor_1 g10356(new_n10732, new_n10722, new_n10733);
nand_1 g10357(new_n10733, new_n10731, new_n10734);
not_1  g10358(new_n10731, new_n10735);
xnor_1 g10359(new_n10733, new_n10735, new_n10736);
nor_1  g10360(new_n10297, new_n10152, new_n10737);
nor_1  g10361(new_n10404, new_n10298, new_n10738);
nor_1  g10362(new_n10738, new_n10737, new_n10739);
nand_1 g10363(new_n10739, new_n10736, new_n10740);
nand_1 g10364(new_n10740, new_n10734, new_n10741);
nand_1 g10365(new_n10741, new_n10729, new_n10742);
nand_1 g10366(new_n10742, new_n10728, new_n10743);
nor_1  g10367(new_n10555, new_n10523, new_n10744);
and_1  g10368(new_n10566, new_n10557, new_n10745);
nor_1  g10369(new_n10745, new_n10744, new_n10746);
nand_1 g10370(new_n10714, new_n10567, new_n10747);
xnor_1 g10371(new_n10701, new_n10636, new_n10748);
xnor_1 g10372(new_n10713, new_n10748, new_n10749);
xnor_1 g10373(new_n10749, new_n10567, new_n10750);
nand_1 g10374(new_n10726, new_n10750, new_n10751);
nand_1 g10375(new_n10751, new_n10747, new_n10752);
not_1  g10376(new_n10465, new_n10753);
nand_1 g10377(new_n10470, new_n10753, new_n10754);
nand_1 g10378(new_n10754, new_n10463, new_n10755);
nand_1 g10379(n11662, n4312, new_n10756);
xnor_1 g10380(new_n10756, new_n10755, new_n10757);
nand_1 g10381(new_n10537, new_n10536, new_n10758);
not_1  g10382(new_n10543, new_n10759);
nand_1 g10383(new_n10759, new_n10538, new_n10760);
nand_1 g10384(new_n10760, new_n10758, new_n10761);
nand_1 g10385(n12299, n10278, new_n10762);
xnor_1 g10386(new_n10762, new_n10761, new_n10763);
nand_1 g10387(new_n10531, new_n10530, new_n10764);
not_1  g10388(new_n10764, new_n10765);
nor_1  g10389(new_n10532, new_n10529, new_n10766);
nor_1  g10390(new_n10766, new_n10765, new_n10767);
nand_1 g10391(n10451, n7436, new_n10768);
nand_1 g10392(n9241, n3022, new_n10769);
xnor_1 g10393(new_n10769, new_n10768, new_n10770);
nand_1 g10394(n11257, n3932, new_n10771);
nand_1 g10395(n10327, n1097, new_n10772);
xnor_1 g10396(new_n10772, new_n10771, new_n10773);
xnor_1 g10397(new_n10773, new_n10770, new_n10774);
xnor_1 g10398(new_n10774, new_n10767, new_n10775);
nand_1 g10399(new_n10692, new_n10691, new_n10776);
not_1  g10400(new_n10776, new_n10777);
nor_1  g10401(new_n10695_1, new_n10777, new_n10778);
nand_1 g10402(n2393, n159, new_n10779);
nand_1 g10403(n5860, n2749, new_n10780);
xnor_1 g10404(new_n10780, new_n10779, new_n10781);
xnor_1 g10405(new_n10781, new_n10778, new_n10782);
xnor_1 g10406(new_n10782, new_n10775, new_n10783);
xnor_1 g10407(new_n10783, new_n10763, new_n10784);
xnor_1 g10408(new_n10784, new_n10757, new_n10785);
and_1  g10409(new_n10626, new_n10595, new_n10786);
nor_1  g10410(new_n10635, new_n10627, new_n10787);
nor_1  g10411(new_n10787, new_n10786, new_n10788);
xnor_1 g10412(new_n10788, new_n10785, new_n10789_1);
not_1  g10413(new_n10676, new_n10790);
nand_1 g10414(new_n10790, new_n10672, new_n10791);
not_1  g10415(new_n10698, new_n10792);
nand_1 g10416(new_n10792, new_n10677, new_n10793);
nand_1 g10417(new_n10793, new_n10791, new_n10794);
nor_1  g10418(new_n10682, new_n10679, new_n10795);
and_1  g10419(n12247, n7388, new_n10796);
nand_1 g10420(new_n10796, new_n10795, new_n10797);
not_1  g10421(new_n10795, new_n10798);
nand_1 g10422(new_n10796, new_n10666, new_n10799);
nand_1 g10423(new_n10799, new_n10798, new_n10800);
nand_1 g10424(new_n10800, new_n10797, new_n10801);
nor_1  g10425(new_n4143, new_n3280, new_n10802);
nand_1 g10426(n12591, n12025, new_n10803);
nand_1 g10427(n11876, n45, new_n10804);
xnor_1 g10428(new_n10804, new_n10803, new_n10805);
xnor_1 g10429(new_n10805, new_n10802, new_n10806);
xnor_1 g10430(new_n10806, new_n10801, new_n10807);
xnor_1 g10431(new_n10807, new_n10794, new_n10808);
nand_1 g10432(new_n10541, new_n10540, new_n10809);
not_1  g10433(new_n10809, new_n10810);
nor_1  g10434(new_n10542, new_n10539, new_n10811);
nor_1  g10435(new_n10811, new_n10810, new_n10812);
nand_1 g10436(n12705, n7456, new_n10813);
nand_1 g10437(n11023, n8276, new_n10814);
xnor_1 g10438(new_n10814, new_n10813, new_n10815);
xnor_1 g10439(new_n10815, new_n10812, new_n10816);
nand_1 g10440(n9583, n5964, new_n10817);
nand_1 g10441(n12511, n7965, new_n10818);
xnor_1 g10442(new_n10818, new_n10817, new_n10819);
xnor_1 g10443(new_n10819, new_n10816, new_n10820);
nand_1 g10444(new_n10554, new_n10548, new_n10821);
nand_1 g10445(new_n10821, new_n10551, new_n10822);
nand_1 g10446(new_n10533, new_n10528, new_n10823);
nand_1 g10447(new_n10546, new_n10823, new_n10824);
xnor_1 g10448(new_n10824, new_n10822, new_n10825);
xnor_1 g10449(new_n10825, new_n10820, new_n10826);
xnor_1 g10450(new_n10826, new_n10808, new_n10827);
nand_1 g10451(new_n10699, new_n10671, new_n10828);
not_1  g10452(new_n10700, new_n10829);
nand_1 g10453(new_n10829, new_n10669, new_n10830);
nand_1 g10454(new_n10830, new_n10828, new_n10831);
nand_1 g10455(new_n10625, new_n10616, new_n10832);
nand_1 g10456(new_n10832, new_n10622, new_n10833);
not_1  g10457(new_n10459, new_n10834);
nand_1 g10458(new_n10834, new_n10454, new_n10835);
nand_1 g10459(new_n10471, new_n10460, new_n10836);
nand_1 g10460(new_n10836, new_n10835, new_n10837);
xnor_1 g10461(new_n10837, new_n10833, new_n10838);
nand_1 g10462(n3986, n3754, new_n10839);
nand_1 g10463(n11423, n6776, new_n10840);
xnor_1 g10464(new_n10840, new_n10839, new_n10841);
nand_1 g10465(n8759, n2278, new_n10842);
nand_1 g10466(n10510, n9640, new_n10843);
xnor_1 g10467(new_n10843, new_n10842, new_n10844);
xnor_1 g10468(new_n10844, new_n10841, new_n10845);
nand_1 g10469(n8476, n4094, new_n10846);
nand_1 g10470(n5305, n753, new_n10847);
xnor_1 g10471(new_n10847, new_n10846, new_n10848_1);
nand_1 g10472(n3616, n1067, new_n10849);
nand_1 g10473(n10644, n6703, new_n10850);
xnor_1 g10474(new_n10850, new_n10849, new_n10851_1);
xnor_1 g10475(new_n10851_1, new_n10848_1, new_n10852);
xnor_1 g10476(new_n10852, new_n10845, new_n10853);
nand_1 g10477(new_n10457, new_n10456, new_n10854);
not_1  g10478(new_n10854, new_n10855);
nor_1  g10479(new_n10458, new_n10455, new_n10856);
nor_1  g10480(new_n10856, new_n10855, new_n10857);
nand_1 g10481(new_n10468, new_n10467, new_n10858);
not_1  g10482(new_n10858, new_n10859);
nor_1  g10483(new_n10469, new_n10466, new_n10860);
nor_1  g10484(new_n10860, new_n10859, new_n10861);
xnor_1 g10485(new_n10861, new_n10857, new_n10862);
xnor_1 g10486(new_n10862, new_n10853, new_n10863);
xnor_1 g10487(new_n10863, new_n10838, new_n10864);
nand_1 g10488(new_n10479, new_n10472, new_n10865);
nand_1 g10489(new_n10865, new_n10476_1, new_n10866);
not_1  g10490(new_n10686, new_n10867);
nand_1 g10491(new_n10867, new_n10684, new_n10868);
not_1  g10492(new_n10697, new_n10869);
nand_1 g10493(new_n10869, new_n10687, new_n10870);
nand_1 g10494(new_n10870, new_n10868, new_n10871);
not_1  g10495(new_n10649, new_n10872);
nor_1  g10496(new_n10688, new_n10872, new_n10873);
not_1  g10497(new_n10689, new_n10874);
nor_1  g10498(new_n10696, new_n10874, new_n10875);
nor_1  g10499(new_n10875, new_n10873, new_n10876);
nand_1 g10500(new_n10602, new_n10601, new_n10877);
not_1  g10501(new_n10877, new_n10878);
nor_1  g10502(new_n10603, new_n10600, new_n10879);
nor_1  g10503(new_n10879, new_n10878, new_n10880);
nand_1 g10504(n10547, n1798, new_n10881);
nand_1 g10505(n8665, n7690, new_n10882);
xnor_1 g10506(new_n10882, new_n10881, new_n10883);
nand_1 g10507(n12826, n2530, new_n10884);
nand_1 g10508(n11892, n1510, new_n10885);
xnor_1 g10509(new_n10885, new_n10884, new_n10886);
xnor_1 g10510(new_n10886, new_n10883, new_n10887);
xnor_1 g10511(new_n10887, new_n10880, new_n10888);
xnor_1 g10512(new_n10888, new_n10876, new_n10889);
xnor_1 g10513(new_n10889, new_n10871, new_n10890);
nor_1  g10514(new_n4187_1, new_n5668, new_n10891);
not_1  g10515(new_n10608, new_n10892);
nand_1 g10516(new_n10614, new_n10892, new_n10893);
nand_1 g10517(new_n10615, new_n10605, new_n10894);
nand_1 g10518(new_n10894, new_n10893, new_n10895);
xnor_1 g10519(new_n10895, new_n10891, new_n10896);
nand_1 g10520(new_n10597, new_n10596, new_n10897);
nand_1 g10521(new_n10604, new_n10599, new_n10898_1);
nand_1 g10522(new_n10898_1, new_n10897, new_n10899);
nand_1 g10523(new_n10612, new_n10611, new_n10900);
not_1  g10524(new_n10900, new_n10901);
nor_1  g10525(new_n10613, new_n10609, new_n10902);
nor_1  g10526(new_n10902, new_n10901, new_n10903);
xnor_1 g10527(new_n10903, new_n10899, new_n10904);
nand_1 g10528(n12648, n2551, new_n10905);
nand_1 g10529(n10685, n5331, new_n10906);
nand_1 g10530(n5645, n4499, new_n10907);
xnor_1 g10531(new_n10907, new_n10906, new_n10908);
xnor_1 g10532(new_n10908, new_n10905, new_n10909);
xnor_1 g10533(new_n10909, new_n10904, new_n10910);
xnor_1 g10534(new_n10910, new_n10896, new_n10911);
xnor_1 g10535(new_n10911, new_n10890, new_n10912);
xnor_1 g10536(new_n10912, new_n10866, new_n10913_1);
xnor_1 g10537(new_n10913_1, new_n10864, new_n10914);
xnor_1 g10538(new_n10914, new_n10831, new_n10915);
xnor_1 g10539(new_n10915, new_n10827, new_n10916);
xnor_1 g10540(new_n10916, new_n10789_1, new_n10917);
nand_1 g10541(new_n10480, new_n10483, new_n10918);
nand_1 g10542(new_n10490, new_n10481, new_n10919);
nand_1 g10543(new_n10919, new_n10918, new_n10920);
nand_1 g10544(new_n10702, new_n10636, new_n10921);
nand_1 g10545(new_n10713, new_n10748, new_n10922);
nand_1 g10546(new_n10922, new_n10921, new_n10923);
xnor_1 g10547(new_n10923, new_n10920, new_n10924);
xnor_1 g10548(new_n10924, new_n10917, new_n10925);
xnor_1 g10549(new_n10925, new_n10752, new_n10926);
xnor_1 g10550(new_n10926, new_n10746, new_n10927);
xnor_1 g10551(new_n10927, new_n10743, n4230);
xnor_1 g10552(new_n6274, new_n6272, n4300);
xnor_1 g10553(new_n3889, new_n3888, n4326);
nand_1 g10554(new_n1400, new_n1394, new_n10931);
nor_1  g10555(new_n378, new_n8515, new_n10932);
nand_1 g10556(new_n1391, new_n1382, new_n10933);
xnor_1 g10557(new_n10933, new_n10932, new_n10934);
nor_1  g10558(new_n1365, new_n1377, new_n10935);
nand_1 g10559(new_n1388, new_n1387, new_n10936);
not_1  g10560(new_n10936, new_n10937);
nor_1  g10561(new_n1389, new_n1386, new_n10938);
nor_1  g10562(new_n10938, new_n10937, new_n10939);
xnor_1 g10563(new_n10939, new_n10935, new_n10940);
not_1  g10564(new_n10940, new_n10941);
nor_1  g10565(new_n4283, new_n1378, new_n10942);
nand_1 g10566(n11877, n4189, new_n10943);
nand_1 g10567(n11407, n9920, new_n10944);
xnor_1 g10568(new_n10944, new_n10943, new_n10945);
nand_1 g10569(new_n10945, new_n10942, new_n10946);
nor_1  g10570(new_n10945, new_n10942, new_n10947);
not_1  g10571(new_n10947, new_n10948);
nand_1 g10572(new_n10948, new_n10946, new_n10949_1);
nand_1 g10573(new_n10949_1, new_n10941, new_n10950);
not_1  g10574(new_n10949_1, new_n10951);
nand_1 g10575(new_n10951, new_n10940, new_n10952);
nand_1 g10576(new_n10952, new_n10950, new_n10953);
not_1  g10577(new_n10953, new_n10954);
xnor_1 g10578(new_n10954, new_n10934, new_n10955);
xnor_1 g10579(new_n10955, new_n10931, new_n10956);
nor_1  g10580(new_n382, new_n8622, new_n10957);
nor_1  g10581(new_n1434, new_n1506, new_n10958);
not_1  g10582(new_n1512_1, new_n10959);
nor_1  g10583(new_n1513, new_n1509, new_n10960);
nor_1  g10584(new_n10960, new_n10959, new_n10961);
xnor_1 g10585(new_n10961, new_n10958, new_n10962);
nor_1  g10586(new_n1435, new_n4529, new_n10963);
nand_1 g10587(n12709, n1094, new_n10964);
nand_1 g10588(new_n10964, new_n1439, new_n10965_1);
not_1  g10589(new_n1439, new_n10966);
not_1  g10590(new_n10964, new_n10967);
nand_1 g10591(new_n10967, new_n10966, new_n10968);
nand_1 g10592(new_n10968, new_n10965_1, new_n10969);
xnor_1 g10593(new_n10969, new_n10963, new_n10970);
xnor_1 g10594(new_n10970, new_n10962, new_n10971);
nand_1 g10595(new_n10971, new_n10957, new_n10972);
not_1  g10596(new_n10972, new_n10973);
nor_1  g10597(new_n10971, new_n10957, new_n10974);
nor_1  g10598(new_n10974, new_n10973, new_n10975);
nand_1 g10599(new_n1523_1, new_n1520, new_n10976);
nand_1 g10600(new_n10976, new_n1517, new_n10977);
nor_1  g10601(new_n10977, new_n10975, new_n10978);
nand_1 g10602(new_n10977, new_n10975, new_n10979);
not_1  g10603(new_n10979, new_n10980);
nor_1  g10604(new_n10980, new_n10978, new_n10981);
xnor_1 g10605(new_n10981, new_n1529, new_n10982);
nand_1 g10606(new_n1578, new_n1530, new_n10983);
nand_1 g10607(new_n1584, new_n10983, new_n10984);
xnor_1 g10608(new_n10984, new_n10982, new_n10985);
nor_1  g10609(new_n1533, new_n8888, new_n10986);
not_1  g10610(new_n10986, new_n10987);
nor_1  g10611(new_n1452, new_n1532, new_n10988);
nand_1 g10612(new_n1543, new_n1542, new_n10989);
not_1  g10613(new_n10989, new_n10990_1);
nor_1  g10614(new_n1544, new_n1540, new_n10991);
nor_1  g10615(new_n10991, new_n10990_1, new_n10992);
nand_1 g10616(new_n10992, new_n10988, new_n10993);
not_1  g10617(new_n10993, new_n10994);
nor_1  g10618(new_n10992, new_n10988, new_n10995);
nor_1  g10619(new_n10995, new_n10994, new_n10996);
nor_1  g10620(new_n1538, new_n1451, new_n10997);
nor_1  g10621(new_n8843, new_n4386, new_n10998);
not_1  g10622(new_n10998, new_n10999);
nor_1  g10623(new_n1539, new_n6825, new_n11000);
not_1  g10624(new_n11000, new_n11001);
nand_1 g10625(new_n11001, new_n10999, new_n11002);
nor_1  g10626(new_n11001, new_n10999, new_n11003);
not_1  g10627(new_n11003, new_n11004);
nand_1 g10628(new_n11004, new_n11002, new_n11005);
xnor_1 g10629(new_n11005, new_n10997, new_n11006);
nand_1 g10630(new_n11006, new_n10996, new_n11007);
not_1  g10631(new_n11007, new_n11008);
nor_1  g10632(new_n11006, new_n10996, new_n11009);
nor_1  g10633(new_n11009, new_n11008, new_n11010);
xnor_1 g10634(new_n11010, new_n10987, new_n11011);
nand_1 g10635(new_n1536, new_n1534, new_n11012);
nor_1  g10636(new_n1545, new_n1537, new_n11013);
not_1  g10637(new_n11013, new_n11014);
nand_1 g10638(new_n11014, new_n11012, new_n11015);
nand_1 g10639(new_n11015, new_n11011, new_n11016);
not_1  g10640(new_n11016, new_n11017);
nor_1  g10641(new_n11015, new_n11011, new_n11018);
nor_1  g10642(new_n11018, new_n11017, new_n11019);
xnor_1 g10643(new_n11019, new_n1551, new_n11020);
not_1  g10644(new_n11020, new_n11021);
not_1  g10645(new_n1569, new_n11022);
nor_1  g10646(new_n1570, new_n11022, new_n11023_1);
nor_1  g10647(new_n8768, new_n385, new_n11024);
nor_1  g10648(new_n8748, new_n1467, new_n11025);
not_1  g10649(new_n11025, new_n11026);
nand_1 g10650(new_n1566, new_n1565, new_n11027);
not_1  g10651(new_n11027, new_n11028);
nor_1  g10652(new_n1567, new_n1563, new_n11029);
nor_1  g10653(new_n11029, new_n11028, new_n11030);
xnor_1 g10654(new_n11030, new_n11026, new_n11031);
nor_1  g10655(new_n1466, new_n4542, new_n11032);
nor_1  g10656(new_n1562, new_n8469, new_n11033);
not_1  g10657(new_n11033, new_n11034);
nor_1  g10658(new_n8466, new_n6869, new_n11035);
not_1  g10659(new_n11035, new_n11036);
nand_1 g10660(new_n11036, new_n11034, new_n11037);
nand_1 g10661(new_n11035, new_n11033, new_n11038);
nand_1 g10662(new_n11038, new_n11037, new_n11039);
xnor_1 g10663(new_n11039, new_n11032, new_n11040);
nand_1 g10664(new_n11040, new_n11031, new_n11041);
not_1  g10665(new_n11041, new_n11042);
nor_1  g10666(new_n11040, new_n11031, new_n11043);
nor_1  g10667(new_n11043, new_n11042, new_n11044);
nand_1 g10668(new_n11044, new_n11024, new_n11045);
not_1  g10669(new_n11045, new_n11046);
nor_1  g10670(new_n11044, new_n11024, new_n11047);
nor_1  g10671(new_n11047, new_n11046, new_n11048);
not_1  g10672(new_n1561, new_n11049);
nor_1  g10673(new_n1568, new_n11049, new_n11050);
nor_1  g10674(new_n11050, new_n1559, new_n11051);
not_1  g10675(new_n11051, new_n11052);
xnor_1 g10676(new_n11052, new_n11048, new_n11053);
xnor_1 g10677(new_n11053, new_n11023_1, new_n11054);
nor_1  g10678(new_n1571, new_n1553, new_n11055);
not_1  g10679(new_n11055, new_n11056);
nand_1 g10680(new_n1577, new_n1573, new_n11057);
nand_1 g10681(new_n11057, new_n11056, new_n11058);
xnor_1 g10682(new_n11058, new_n11054, new_n11059);
xnor_1 g10683(new_n11059, new_n11021, new_n11060);
nand_1 g10684(new_n11060, new_n10985, new_n11061);
not_1  g10685(new_n11061, new_n11062);
nor_1  g10686(new_n11060, new_n10985, new_n11063);
nor_1  g10687(new_n11063, new_n11062, new_n11064);
nor_1  g10688(new_n11064, new_n10956, new_n11065);
nand_1 g10689(new_n11064, new_n10956, new_n11066);
not_1  g10690(new_n11066, new_n11067);
nor_1  g10691(new_n11067, new_n11065, new_n11068);
not_1  g10692(new_n1401, new_n11069);
nor_1  g10693(new_n1504, new_n11069, new_n11070);
not_1  g10694(new_n11070, new_n11071);
nand_1 g10695(new_n1587, new_n1505, new_n11072);
nand_1 g10696(new_n11072, new_n11071, new_n11073);
xor_1  g10697(new_n11073, new_n11068, n4333);
nor_1  g10698(new_n1371, new_n1592, new_n11075);
not_1  g10699(new_n11075, new_n11076);
nand_1 g10700(n5240, n5212, new_n11077);
nand_1 g10701(n11821, n11407, new_n11078);
nor_1  g10702(new_n11078, new_n11077, new_n11079);
not_1  g10703(new_n11079, new_n11080);
nand_1 g10704(new_n11078, new_n11077, new_n11081);
nand_1 g10705(new_n11081, new_n11080, new_n11082);
xnor_1 g10706(new_n11082, new_n11076, new_n11083);
nand_1 g10707(n11407, n5240, new_n11084);
nand_1 g10708(n11877, n3172, new_n11085);
nand_1 g10709(new_n11085, new_n11084, new_n11086);
not_1  g10710(new_n11086, new_n11087);
nor_1  g10711(new_n1592, new_n1378, new_n11088);
xnor_1 g10712(new_n11085, new_n11084, new_n11089);
nor_1  g10713(new_n11089, new_n11088, new_n11090);
nor_1  g10714(new_n11090, new_n11087, new_n11091);
nor_1  g10715(new_n11091, new_n11083, new_n11092);
not_1  g10716(new_n11092, new_n11093);
nand_1 g10717(new_n11091, new_n11083, new_n11094);
nand_1 g10718(new_n11094, new_n11093, new_n11095);
nor_1  g10719(new_n8515, new_n1590, new_n11096);
not_1  g10720(new_n11096, new_n11097);
nor_1  g10721(new_n1365, new_n1600, new_n11098);
not_1  g10722(new_n11098, new_n11099);
nand_1 g10723(new_n11099, new_n11097, new_n11100);
nor_1  g10724(new_n11099, new_n11097, new_n11101);
not_1  g10725(new_n11101, new_n11102);
nand_1 g10726(new_n11102, new_n11100, new_n11103);
xnor_1 g10727(new_n11103, new_n11095, new_n11104);
nor_1  g10728(new_n1365, new_n1590, new_n11105);
nand_1 g10729(n11877, n1333, new_n11106);
nand_1 g10730(n11757, n11407, new_n11107);
nand_1 g10731(new_n11107, new_n11106, new_n11108);
not_1  g10732(new_n11108, new_n11109);
nor_1  g10733(new_n1378, new_n1600, new_n11110);
xnor_1 g10734(new_n11107, new_n11106, new_n11111);
nor_1  g10735(new_n11111, new_n11110, new_n11112);
nor_1  g10736(new_n11112, new_n11109, new_n11113);
nand_1 g10737(new_n11113, new_n11105, new_n11114);
not_1  g10738(new_n11114, new_n11115);
nor_1  g10739(new_n11113, new_n11105, new_n11116);
nor_1  g10740(new_n11116, new_n11115, new_n11117);
xnor_1 g10741(new_n11089, new_n11088, new_n11118);
nand_1 g10742(new_n11118, new_n11117, new_n11119);
nand_1 g10743(new_n11119, new_n11114, new_n11120);
nand_1 g10744(new_n11120, new_n11104, new_n11121);
not_1  g10745(new_n11121, new_n11122);
nor_1  g10746(new_n11120, new_n11104, new_n11123);
nor_1  g10747(new_n11123, new_n11122, new_n11124);
not_1  g10748(new_n11124, new_n11125);
nor_1  g10749(new_n1348, new_n8515, new_n11126);
not_1  g10750(new_n11119, new_n11127);
nor_1  g10751(new_n11118, new_n11117, new_n11128);
nor_1  g10752(new_n11128, new_n11127, new_n11129);
nor_1  g10753(new_n11129, new_n11126, new_n11130);
not_1  g10754(new_n11130, new_n11131);
nand_1 g10755(new_n11129, new_n11126, new_n11132);
nand_1 g10756(new_n11132, new_n11131, new_n11133);
not_1  g10757(new_n11133, new_n11134);
nor_1  g10758(new_n1348, new_n1365, new_n11135);
nand_1 g10759(n11407, n3172, new_n11136);
nand_1 g10760(n11877, n7862, new_n11137);
nand_1 g10761(new_n11137, new_n11136, new_n11138);
not_1  g10762(new_n11138, new_n11139);
nor_1  g10763(new_n1368, new_n1348, new_n11140);
not_1  g10764(new_n11140, new_n11141);
nor_1  g10765(new_n11141, new_n11085, new_n11142);
nor_1  g10766(new_n1378, new_n1590, new_n11143);
nor_1  g10767(new_n11143, new_n11142, new_n11144);
nor_1  g10768(new_n11144, new_n11139, new_n11145);
nand_1 g10769(new_n11145, new_n11135, new_n11146);
not_1  g10770(new_n11146, new_n11147);
xnor_1 g10771(new_n11145, new_n11135, new_n11148);
xnor_1 g10772(new_n11111, new_n11110, new_n11149);
not_1  g10773(new_n11149, new_n11150);
nor_1  g10774(new_n11150, new_n11148, new_n11151);
nor_1  g10775(new_n11151, new_n11147, new_n11152);
nand_1 g10776(new_n11152, new_n11134, new_n11153_1);
nand_1 g10777(new_n11153_1, new_n11131, new_n11154);
nor_1  g10778(new_n11154, new_n11125, new_n11155);
not_1  g10779(new_n11155, new_n11156);
not_1  g10780(new_n11103, new_n11157);
nand_1 g10781(new_n11157, new_n11095, new_n11158);
nand_1 g10782(new_n11122, new_n11101, new_n11159);
nand_1 g10783(new_n11121, new_n11102, new_n11160);
nand_1 g10784(new_n11160, new_n11159, new_n11161);
nand_1 g10785(new_n11161, new_n11158, new_n11162);
nand_1 g10786(n11757, n4370, new_n11163);
xnor_1 g10787(new_n11163, new_n11079, new_n11164);
nand_1 g10788(n11821, n5212, new_n11165);
nand_1 g10789(n11877, n5240, new_n11166);
nand_1 g10790(n11407, n9080, new_n11167);
xnor_1 g10791(new_n11167, new_n11166, new_n11168);
xnor_1 g10792(new_n11168, new_n11165, new_n11169);
xor_1  g10793(new_n11169, new_n11164, new_n11170);
nand_1 g10794(new_n11082, new_n11076, new_n11171);
nand_1 g10795(new_n11093, new_n11171, new_n11172);
not_1  g10796(new_n11172, new_n11173);
nor_1  g10797(new_n8561, new_n1590, new_n11174);
nand_1 g10798(n5320, n3172, new_n11175);
nand_1 g10799(n9725, n7862, new_n11176);
xnor_1 g10800(new_n11176, new_n11175, new_n11177);
xor_1  g10801(new_n11177, new_n11174, new_n11178);
xnor_1 g10802(new_n11178, new_n11173, new_n11179);
xnor_1 g10803(new_n11179, new_n11170, new_n11180);
xor_1  g10804(new_n11180, new_n11162, new_n11181);
xnor_1 g10805(new_n11181, new_n11156, new_n11182);
nor_1  g10806(new_n8561, new_n1348, new_n11183);
nand_1 g10807(new_n11154, new_n11125, new_n11184);
nand_1 g10808(new_n11184, new_n11156, new_n11185);
not_1  g10809(new_n11185, new_n11186);
nor_1  g10810(new_n11186, new_n11183, new_n11187);
xnor_1 g10811(new_n11149, new_n11148, new_n11188);
nor_1  g10812(new_n11142, new_n11139, new_n11189);
nor_1  g10813(new_n1368, new_n1590, new_n11190);
nor_1  g10814(new_n1348, new_n1378, new_n11191);
nand_1 g10815(new_n11191, new_n11190, new_n11192);
nor_1  g10816(new_n11192, new_n11189, new_n11193);
nand_1 g10817(new_n11193, new_n11188, new_n11194);
xnor_1 g10818(new_n11152, new_n11133, new_n11195);
nor_1  g10819(new_n11195, new_n11194, new_n11196);
not_1  g10820(new_n11187, new_n11197);
nand_1 g10821(new_n11186, new_n11183, new_n11198);
nand_1 g10822(new_n11198, new_n11197, new_n11199);
nor_1  g10823(new_n11199, new_n11196, new_n11200);
nor_1  g10824(new_n11200, new_n11187, new_n11201);
not_1  g10825(new_n11201, new_n11202);
xnor_1 g10826(new_n11202, new_n11182, new_n11203);
not_1  g10827(new_n11203, new_n11204);
nor_1  g10828(new_n1506, new_n1350, new_n11205);
nor_1  g10829(new_n1402, new_n1729, new_n11206);
not_1  g10830(new_n11206, new_n11207);
not_1  g10831(n6429, new_n11208);
nor_1  g10832(new_n1350, new_n11208, new_n11209);
not_1  g10833(new_n11209, new_n11210);
nor_1  g10834(new_n11210, new_n11207, new_n11211);
not_1  g10835(new_n11211, new_n11212);
nand_1 g10836(new_n11210, new_n11207, new_n11213);
nor_1  g10837(new_n1435, new_n1735, new_n11214);
nand_1 g10838(new_n11214, new_n11213, new_n11215);
nand_1 g10839(new_n11215, new_n11212, new_n11216_1);
xnor_1 g10840(new_n11216_1, new_n11205, new_n11217);
nor_1  g10841(new_n1435, new_n1729, new_n11218);
nor_1  g10842(new_n1402, new_n1747, new_n11219);
not_1  g10843(new_n11219, new_n11220);
nor_1  g10844(new_n1735, new_n11208, new_n11221);
not_1  g10845(new_n11221, new_n11222_1);
nand_1 g10846(new_n11222_1, new_n11220, new_n11223);
nand_1 g10847(new_n11221, new_n11219, new_n11224);
nand_1 g10848(new_n11224, new_n11223, new_n11225);
xnor_1 g10849(new_n11225, new_n11218, new_n11226);
xnor_1 g10850(new_n11226, new_n11217, new_n11227);
not_1  g10851(new_n11213, new_n11228);
nor_1  g10852(new_n11228, new_n11211, new_n11229);
nor_1  g10853(new_n1402, new_n1735, new_n11230);
nor_1  g10854(new_n1435, new_n1350, new_n11231);
nand_1 g10855(new_n11231, new_n11230, new_n11232);
nor_1  g10856(new_n11232, new_n11229, new_n11233);
nand_1 g10857(new_n11233, new_n11227, new_n11234);
nor_1  g10858(new_n1350, new_n8622, new_n11235);
nor_1  g10859(new_n1735, new_n1506, new_n11236);
not_1  g10860(new_n11236, new_n11237);
not_1  g10861(new_n11223, new_n11238);
not_1  g10862(new_n11218, new_n11239);
and_1  g10863(new_n11224, new_n11239, new_n11240);
nor_1  g10864(new_n11240, new_n11238, new_n11241);
xnor_1 g10865(new_n11241, new_n11237, new_n11242);
nor_1  g10866(new_n1435, new_n1747, new_n11243);
nand_1 g10867(n6429, n2464, new_n11244);
nand_1 g10868(n12709, n4187, new_n11245);
xnor_1 g10869(new_n11245, new_n11244, new_n11246);
xor_1  g10870(new_n11246, new_n11243, new_n11247);
xnor_1 g10871(new_n11247, new_n11242, new_n11248);
nand_1 g10872(new_n11248, new_n11235, new_n11249);
not_1  g10873(new_n11249, new_n11250);
nor_1  g10874(new_n11248, new_n11235, new_n11251);
nor_1  g10875(new_n11251, new_n11250, new_n11252);
nand_1 g10876(new_n11216_1, new_n11205, new_n11253);
not_1  g10877(new_n11226, new_n11254);
nor_1  g10878(new_n11254, new_n11217, new_n11255);
not_1  g10879(new_n11255, new_n11256);
nand_1 g10880(new_n11256, new_n11253, new_n11257_1);
xnor_1 g10881(new_n11257_1, new_n11252, new_n11258);
nor_1  g10882(new_n11258, new_n11234, new_n11259);
nor_1  g10883(new_n8602, new_n1350, new_n11260);
nor_1  g10884(new_n1747, new_n11208, new_n11261);
nand_1 g10885(n12709, n4203, new_n11262);
nand_1 g10886(n11728, n4187, new_n11263);
nand_1 g10887(new_n11263, new_n11262, new_n11264);
nor_1  g10888(new_n11263, new_n11262, new_n11265);
not_1  g10889(new_n11265, new_n11266);
nand_1 g10890(new_n11266, new_n11264, new_n11267);
xnor_1 g10891(new_n11267, new_n11261, new_n11268);
nand_1 g10892(new_n11245, new_n11244, new_n11269);
not_1  g10893(new_n11269, new_n11270);
nor_1  g10894(new_n11246, new_n11243, new_n11271);
nor_1  g10895(new_n11271, new_n11270, new_n11272);
xnor_1 g10896(new_n11272, new_n11268, new_n11273);
not_1  g10897(new_n11273, new_n11274);
nor_1  g10898(new_n1735, new_n8622, new_n11275);
not_1  g10899(new_n11275, new_n11276);
nor_1  g10900(new_n1506, new_n1729, new_n11277);
not_1  g10901(new_n11277, new_n11278);
nor_1  g10902(new_n11278, new_n11276, new_n11279);
not_1  g10903(new_n11279, new_n11280);
nand_1 g10904(new_n11278, new_n11276, new_n11281);
and_1  g10905(new_n11281, new_n11280, new_n11282);
nand_1 g10906(new_n11282, new_n11274, new_n11283);
not_1  g10907(new_n11282, new_n11284);
nand_1 g10908(new_n11284, new_n11273, new_n11285);
nand_1 g10909(new_n11285, new_n11283, new_n11286);
not_1  g10910(new_n11286, new_n11287);
nand_1 g10911(new_n11241, new_n11236, new_n11288);
not_1  g10912(new_n11288, new_n11289);
xnor_1 g10913(new_n11241, new_n11236, new_n11290);
nor_1  g10914(new_n11247, new_n11290, new_n11291);
nor_1  g10915(new_n11291, new_n11289, new_n11292);
not_1  g10916(new_n11292, new_n11293);
nand_1 g10917(new_n11293, new_n11287, new_n11294);
nand_1 g10918(new_n11292, new_n11286, new_n11295);
nand_1 g10919(new_n11295, new_n11294, new_n11296_1);
nand_1 g10920(new_n11257_1, new_n11252, new_n11297);
nand_1 g10921(new_n11297, new_n11249, new_n11298);
xnor_1 g10922(new_n11298, new_n11296_1, new_n11299);
xnor_1 g10923(new_n11299, new_n11260, new_n11300);
xnor_1 g10924(new_n11300, new_n11259, new_n11301);
not_1  g10925(new_n11301, new_n11302);
xnor_1 g10926(new_n11258, new_n11234, new_n11303);
xnor_1 g10927(new_n11233, new_n11227, new_n11304);
nand_1 g10928(n12489, n4805, new_n11305);
nand_1 g10929(n10990, n7236, new_n11306);
nor_1  g10930(new_n11306, new_n11305, new_n11307);
not_1  g10931(new_n11307, new_n11308);
nand_1 g10932(n12489, n11478, new_n11309);
not_1  g10933(new_n11309, new_n11310);
nand_1 g10934(n7159, n4805, new_n11311_1);
not_1  g10935(new_n11311_1, new_n11312);
nand_1 g10936(new_n11312, new_n11310, new_n11313);
nand_1 g10937(new_n11311_1, new_n11309, new_n11314);
nand_1 g10938(new_n11314, new_n11313, new_n11315);
nand_1 g10939(new_n11315, new_n11308, new_n11316);
xnor_1 g10940(new_n11315, new_n11307, new_n11317);
nand_1 g10941(n10990, n3992, new_n11318);
nand_1 g10942(n7236, n5760, new_n11319);
xnor_1 g10943(new_n11319, new_n11318, new_n11320);
nand_1 g10944(new_n11320, new_n11317, new_n11321);
nand_1 g10945(new_n11321, new_n11316, new_n11322);
nand_1 g10946(n10990, n8384, new_n11323);
nand_1 g10947(n7236, n1478, new_n11324);
nor_1  g10948(new_n11324, new_n11323, new_n11325);
not_1  g10949(new_n11306, new_n11326_1);
nor_1  g10950(new_n1466, new_n1835_1, new_n11327);
not_1  g10951(new_n11327, new_n11328);
nor_1  g10952(new_n11328, new_n11326_1, new_n11329);
nand_1 g10953(new_n11324, new_n11323, new_n11330);
nor_1  g10954(new_n11330, new_n11329, new_n11331);
nor_1  g10955(new_n11331, new_n11325, new_n11332);
nand_1 g10956(new_n11330, new_n11329, new_n11333);
nand_1 g10957(new_n11333, new_n11332, new_n11334);
nand_1 g10958(new_n11334, new_n11322, new_n11335);
not_1  g10959(new_n11334, new_n11336);
xnor_1 g10960(new_n11336, new_n11322, new_n11337);
nor_1  g10961(new_n1931, new_n1451, new_n11338);
nand_1 g10962(new_n11338, new_n11305, new_n11339);
not_1  g10963(new_n11339, new_n11340);
nor_1  g10964(new_n1539, new_n1923, new_n11341);
not_1  g10965(new_n11341, new_n11342);
nor_1  g10966(new_n8843, new_n1925, new_n11343);
not_1  g10967(new_n11343, new_n11344);
nand_1 g10968(new_n11344, new_n11342, new_n11345);
not_1  g10969(new_n11345, new_n11346);
nand_1 g10970(new_n11343, new_n11341, new_n11347);
not_1  g10971(new_n11347, new_n11348);
nor_1  g10972(new_n11348, new_n11346, new_n11349);
nor_1  g10973(new_n11349, new_n11340, new_n11350);
nor_1  g10974(new_n11346, new_n11339, new_n11351);
nor_1  g10975(new_n11351, new_n11350, new_n11352);
not_1  g10976(new_n11352, new_n11353);
nand_1 g10977(new_n11353, new_n11337, new_n11354);
nand_1 g10978(new_n11354, new_n11335, new_n11355);
nor_1  g10979(new_n1532, new_n1925, new_n11356);
nand_1 g10980(new_n11345, new_n11338, new_n11357);
nand_1 g10981(new_n11357, new_n11347, new_n11358);
nand_1 g10982(new_n11358, new_n11356, new_n11359);
not_1  g10983(new_n11359, new_n11360);
nor_1  g10984(new_n11358, new_n11356, new_n11361);
nor_1  g10985(new_n11361, new_n11360, new_n11362);
nor_1  g10986(new_n1451, new_n1923, new_n11363);
nand_1 g10987(n12489, n137, new_n11364);
nand_1 g10988(n12777, n11478, new_n11365);
xnor_1 g10989(new_n11365, new_n11364, new_n11366);
xnor_1 g10990(new_n11366, new_n11363, new_n11367);
xnor_1 g10991(new_n11367, new_n11362, new_n11368);
nor_1  g10992(new_n11349, new_n11313, new_n11369);
xnor_1 g10993(new_n11369, new_n11368, new_n11370);
not_1  g10994(new_n11370, new_n11371);
nor_1  g10995(new_n8748, new_n1833, new_n11372);
not_1  g10996(new_n11330, new_n11373);
nor_1  g10997(new_n11327, new_n11325, new_n11374);
nor_1  g10998(new_n11374, new_n11373, new_n11375);
nand_1 g10999(new_n11375, new_n11372, new_n11376);
not_1  g11000(new_n11376, new_n11377);
nor_1  g11001(new_n11375, new_n11372, new_n11378);
nor_1  g11002(new_n11378, new_n11377, new_n11379);
nor_1  g11003(new_n1837, new_n1466, new_n11380);
nand_1 g11004(n10990, n6358, new_n11381);
nand_1 g11005(n3992, n1478, new_n11382);
xnor_1 g11006(new_n11382, new_n11381, new_n11383);
xnor_1 g11007(new_n11383, new_n11380, new_n11384);
xnor_1 g11008(new_n11384, new_n11379, new_n11385);
nor_1  g11009(new_n11332, new_n11328, new_n11386);
xnor_1 g11010(new_n11386, new_n11385, new_n11387);
not_1  g11011(new_n11387, new_n11388);
nand_1 g11012(new_n11388, new_n11371, new_n11389);
nand_1 g11013(new_n11387, new_n11370, new_n11390);
nand_1 g11014(new_n11390, new_n11389, new_n11391);
xnor_1 g11015(new_n11391, new_n11355, new_n11392);
nor_1  g11016(new_n11392, new_n11304, new_n11393);
not_1  g11017(new_n11393, new_n11394);
not_1  g11018(new_n11304, new_n11395);
xnor_1 g11019(new_n11392, new_n11395, new_n11396);
xnor_1 g11020(new_n11353, new_n11337, new_n11397);
nor_1  g11021(new_n1402, new_n1350, new_n11398);
not_1  g11022(new_n11398, new_n11399);
nand_1 g11023(new_n11399, new_n11214, new_n11400);
not_1  g11024(new_n11400, new_n11401);
nor_1  g11025(new_n11401, new_n11229, new_n11402);
nor_1  g11026(new_n11400, new_n11228, new_n11403);
nor_1  g11027(new_n11403, new_n11402, new_n11404);
nand_1 g11028(new_n11404, new_n11397, new_n11405);
not_1  g11029(new_n11405, new_n11406);
nor_1  g11030(new_n11404, new_n11397, new_n11407_1);
nor_1  g11031(new_n11407_1, new_n11406, new_n11408);
xnor_1 g11032(new_n11320, new_n11317, new_n11409);
xnor_1 g11033(new_n11231, new_n11230, new_n11410);
not_1  g11034(new_n11410, new_n11411);
nand_1 g11035(new_n11411, new_n11409, new_n11412);
nand_1 g11036(new_n11306, new_n11305, new_n11413);
and_1  g11037(new_n11413, new_n11308, new_n11414);
and_1  g11038(new_n11414, new_n11398, new_n11415);
xnor_1 g11039(new_n11410, new_n11409, new_n11416);
nand_1 g11040(new_n11416, new_n11415, new_n11417);
nand_1 g11041(new_n11417, new_n11412, new_n11418);
nand_1 g11042(new_n11418, new_n11408, new_n11419);
nand_1 g11043(new_n11419, new_n11405, new_n11420);
nand_1 g11044(new_n11420, new_n11396, new_n11421);
nand_1 g11045(new_n11421, new_n11394, new_n11422);
not_1  g11046(new_n11422, new_n11423_1);
nand_1 g11047(new_n11423_1, new_n11303, new_n11424);
xnor_1 g11048(new_n11422, new_n11303, new_n11425);
not_1  g11049(new_n11368, new_n11426);
nand_1 g11050(new_n11369, new_n11426, new_n11427);
nor_1  g11051(new_n1451, new_n1959, new_n11428);
nand_1 g11052(n12777, n5283, new_n11429);
nand_1 g11053(n12489, n6294, new_n11430);
xnor_1 g11054(new_n11430, new_n11429, new_n11431);
nor_1  g11055(new_n11431, new_n11428, new_n11432);
not_1  g11056(new_n11432, new_n11433);
nand_1 g11057(new_n11431, new_n11428, new_n11434);
nand_1 g11058(new_n11434, new_n11433, new_n11435);
nor_1  g11059(new_n1931, new_n1532, new_n11436);
nand_1 g11060(new_n11365, new_n11364, new_n11437);
not_1  g11061(new_n11437, new_n11438);
nor_1  g11062(new_n11366, new_n11363, new_n11439);
nor_1  g11063(new_n11439, new_n11438, new_n11440);
nand_1 g11064(new_n11440, new_n11436, new_n11441);
not_1  g11065(new_n11441, new_n11442);
nor_1  g11066(new_n11440, new_n11436, new_n11443);
nor_1  g11067(new_n11443, new_n11442, new_n11444);
xnor_1 g11068(new_n11444, new_n11435, new_n11445);
not_1  g11069(new_n11445, new_n11446);
nor_1  g11070(new_n8888, new_n1925, new_n11447);
nand_1 g11071(new_n11367, new_n11362, new_n11448);
nand_1 g11072(new_n11448, new_n11359, new_n11449);
xnor_1 g11073(new_n11449, new_n11447, new_n11450);
xnor_1 g11074(new_n11450, new_n11446, new_n11451);
xnor_1 g11075(new_n11451, new_n11427, new_n11452);
not_1  g11076(new_n11452, new_n11453);
not_1  g11077(new_n11386, new_n11454);
nor_1  g11078(new_n11454, new_n11385, new_n11455);
not_1  g11079(new_n11455, new_n11456);
nor_1  g11080(new_n1866, new_n1466, new_n11457);
nand_1 g11081(n8384, n1478, new_n11458);
nand_1 g11082(n10990, n5198, new_n11459);
nand_1 g11083(new_n11459, new_n11458, new_n11460);
not_1  g11084(new_n11460, new_n11461);
nor_1  g11085(new_n11459, new_n11458, new_n11462);
nor_1  g11086(new_n11462, new_n11461, new_n11463);
xnor_1 g11087(new_n11463, new_n11457, new_n11464);
nor_1  g11088(new_n8748, new_n1835_1, new_n11465);
not_1  g11089(new_n11465, new_n11466);
nand_1 g11090(new_n11382, new_n11381, new_n11467);
not_1  g11091(new_n11467, new_n11468);
nor_1  g11092(new_n11383, new_n11380, new_n11469);
nor_1  g11093(new_n11469, new_n11468, new_n11470);
xnor_1 g11094(new_n11470, new_n11466, new_n11471);
xnor_1 g11095(new_n11471, new_n11464, new_n11472);
not_1  g11096(new_n11472, new_n11473);
nor_1  g11097(new_n8768, new_n1833, new_n11474);
nand_1 g11098(new_n11384, new_n11379, new_n11475);
nand_1 g11099(new_n11475, new_n11376, new_n11476);
xnor_1 g11100(new_n11476, new_n11474, new_n11477);
xnor_1 g11101(new_n11477, new_n11473, new_n11478_1);
nor_1  g11102(new_n11478_1, new_n11456, new_n11479);
not_1  g11103(new_n11479, new_n11480);
nand_1 g11104(new_n11478_1, new_n11456, new_n11481);
nand_1 g11105(new_n11481, new_n11480, new_n11482);
xnor_1 g11106(new_n11482, new_n11453, new_n11483);
not_1  g11107(new_n11391, new_n11484);
nand_1 g11108(new_n11484, new_n11355, new_n11485);
nand_1 g11109(new_n11485, new_n11389, new_n11486);
xnor_1 g11110(new_n11486, new_n11483, new_n11487);
nand_1 g11111(new_n11487, new_n11425, new_n11488);
nand_1 g11112(new_n11488, new_n11424, new_n11489);
nand_1 g11113(new_n11489, new_n11302, new_n11490);
nor_1  g11114(new_n1833, new_n8804, new_n11491);
not_1  g11115(new_n11491, new_n11492);
nand_1 g11116(new_n11470, new_n11465, new_n11493);
not_1  g11117(new_n11464, new_n11494);
nand_1 g11118(new_n11471, new_n11494, new_n11495);
nand_1 g11119(new_n11495, new_n11493, new_n11496);
nor_1  g11120(new_n8768, new_n1835_1, new_n11497);
not_1  g11121(new_n11497, new_n11498);
nor_1  g11122(new_n8748, new_n1837, new_n11499);
not_1  g11123(new_n11499, new_n11500);
nor_1  g11124(new_n11500, new_n11498, new_n11501);
not_1  g11125(new_n11501, new_n11502);
nand_1 g11126(new_n11500, new_n11498, new_n11503);
nand_1 g11127(new_n11503, new_n11502, new_n11504);
xnor_1 g11128(new_n11504, new_n11496, new_n11505);
nor_1  g11129(new_n1866, new_n8469, new_n11506);
not_1  g11130(new_n11506, new_n11507);
nand_1 g11131(n5760, n5198, new_n11508);
nand_1 g11132(n10990, n1471, new_n11509);
xnor_1 g11133(new_n11509, new_n11508, new_n11510);
nor_1  g11134(new_n11510, new_n11507, new_n11511);
not_1  g11135(new_n11511, new_n11512);
nand_1 g11136(new_n11510, new_n11507, new_n11513);
nand_1 g11137(new_n11513, new_n11512, new_n11514);
not_1  g11138(new_n11463, new_n11515);
nor_1  g11139(new_n11515, new_n11457, new_n11516);
nor_1  g11140(new_n11516, new_n11461, new_n11517);
xnor_1 g11141(new_n11517, new_n11514, new_n11518);
xnor_1 g11142(new_n11518, new_n11505, new_n11519);
nor_1  g11143(new_n11476, new_n11474, new_n11520);
nor_1  g11144(new_n11477, new_n11472, new_n11521);
nor_1  g11145(new_n11521, new_n11520, new_n11522);
xnor_1 g11146(new_n11522, new_n11519, new_n11523);
xnor_1 g11147(new_n11523, new_n11492, new_n11524);
xnor_1 g11148(new_n11524, new_n11480, new_n11525);
not_1  g11149(new_n11525, new_n11526);
not_1  g11150(new_n11451, new_n11527);
nor_1  g11151(new_n11527, new_n11427, new_n11528);
nor_1  g11152(new_n1925, new_n8942, new_n11529);
not_1  g11153(new_n11529, new_n11530);
nand_1 g11154(new_n11444, new_n11435, new_n11531);
nand_1 g11155(new_n11531, new_n11441, new_n11532);
nor_1  g11156(new_n8888, new_n1931, new_n11533);
not_1  g11157(new_n11533, new_n11534);
nor_1  g11158(new_n1532, new_n1923, new_n11535);
not_1  g11159(new_n11535, new_n11536_1);
nand_1 g11160(new_n11536_1, new_n11534, new_n11537);
nor_1  g11161(new_n11536_1, new_n11534, new_n11538);
not_1  g11162(new_n11538, new_n11539);
nand_1 g11163(new_n11539, new_n11537, new_n11540);
xnor_1 g11164(new_n11540, new_n11532, new_n11541);
nor_1  g11165(new_n8843, new_n1959, new_n11542);
not_1  g11166(new_n11542, new_n11543);
nand_1 g11167(n7159, n6294, new_n11544);
nand_1 g11168(n12489, n6797, new_n11545);
xnor_1 g11169(new_n11545, new_n11544, new_n11546);
xnor_1 g11170(new_n11546, new_n11543, new_n11547);
nand_1 g11171(new_n11430, new_n11429, new_n11548);
nand_1 g11172(new_n11433, new_n11548, new_n11549);
xnor_1 g11173(new_n11549, new_n11547, new_n11550);
not_1  g11174(new_n11550, new_n11551);
xnor_1 g11175(new_n11551, new_n11541, new_n11552);
nor_1  g11176(new_n11449, new_n11447, new_n11553);
nor_1  g11177(new_n11450, new_n11446, new_n11554);
nor_1  g11178(new_n11554, new_n11553, new_n11555);
xnor_1 g11179(new_n11555, new_n11552, new_n11556);
xnor_1 g11180(new_n11556, new_n11530, new_n11557);
xnor_1 g11181(new_n11557, new_n11528, new_n11558);
nor_1  g11182(new_n11482, new_n11453, new_n11559);
nor_1  g11183(new_n11486, new_n11483, new_n11560);
nor_1  g11184(new_n11560, new_n11559, new_n11561);
nand_1 g11185(new_n11561, new_n11558, new_n11562);
not_1  g11186(new_n11562, new_n11563);
nor_1  g11187(new_n11561, new_n11558, new_n11564);
nor_1  g11188(new_n11564, new_n11563, new_n11565);
nand_1 g11189(new_n11565, new_n11526, new_n11566);
not_1  g11190(new_n11566, new_n11567);
nor_1  g11191(new_n11565, new_n11526, new_n11568);
nor_1  g11192(new_n11568, new_n11567, new_n11569);
xnor_1 g11193(new_n11489, new_n11301, new_n11570);
nand_1 g11194(new_n11570, new_n11569, new_n11571);
nand_1 g11195(new_n11571, new_n11490, new_n11572);
not_1  g11196(new_n11296_1, new_n11573);
nand_1 g11197(new_n11298, new_n11573, new_n11574);
not_1  g11198(new_n11294, new_n11575);
nand_1 g11199(new_n11575, new_n11279, new_n11576);
nand_1 g11200(new_n11294, new_n11280, new_n11577);
nand_1 g11201(new_n11577, new_n11576, new_n11578);
nand_1 g11202(new_n11578, new_n11283, new_n11579);
not_1  g11203(new_n11267, new_n11580);
nand_1 g11204(new_n11580, new_n11261, new_n11581);
nand_1 g11205(new_n11272, new_n11268, new_n11582);
nand_1 g11206(new_n11582, new_n11581, new_n11583);
nor_1  g11207(new_n1735, new_n8602, new_n11584);
nand_1 g11208(n2464, n2433, new_n11585);
nand_1 g11209(n7730, n6877, new_n11586);
xnor_1 g11210(new_n11586, new_n11585, new_n11587);
xor_1  g11211(new_n11587, new_n11584, new_n11588);
xnor_1 g11212(new_n11588, new_n11583, new_n11589);
nand_1 g11213(n11311, n8819, new_n11590);
xnor_1 g11214(new_n11590, new_n11265, new_n11591);
nor_1  g11215(new_n1435, new_n2119, new_n11592);
nand_1 g11216(n6429, n4187, new_n11593);
nand_1 g11217(n12753, n12709, new_n11594);
xnor_1 g11218(new_n11594, new_n11593, new_n11595);
xor_1  g11219(new_n11595, new_n11592, new_n11596);
xnor_1 g11220(new_n11596, new_n11591, new_n11597);
xnor_1 g11221(new_n11597, new_n11589, new_n11598);
xnor_1 g11222(new_n11598, new_n11579, new_n11599);
xnor_1 g11223(new_n11599, new_n11574, new_n11600);
not_1  g11224(new_n11600, new_n11601);
nand_1 g11225(new_n11299, new_n11260, new_n11602);
not_1  g11226(new_n11260, new_n11603);
xnor_1 g11227(new_n11299, new_n11603, new_n11604);
nand_1 g11228(new_n11604, new_n11259, new_n11605);
nand_1 g11229(new_n11605, new_n11602, new_n11606);
xnor_1 g11230(new_n11606, new_n11601, new_n11607);
not_1  g11231(new_n11555, new_n11608);
nor_1  g11232(new_n11608, new_n11552, new_n11609);
not_1  g11233(new_n11609, new_n11610);
nor_1  g11234(new_n1931, new_n8942, new_n11611);
nand_1 g11235(n11967, n5283, new_n11612);
not_1  g11236(new_n11612, new_n11613);
nand_1 g11237(n4805, n1353, new_n11614);
xnor_1 g11238(new_n11614, new_n11613, new_n11615);
xnor_1 g11239(new_n11615, new_n11611, new_n11616);
nor_1  g11240(new_n11546, new_n11543, new_n11617);
nor_1  g11241(new_n11549, new_n11547, new_n11618);
nor_1  g11242(new_n11618, new_n11617, new_n11619);
not_1  g11243(new_n11619, new_n11620);
xnor_1 g11244(new_n11620, new_n11616, new_n11621);
nor_1  g11245(new_n11545, new_n11544, new_n11622);
nor_1  g11246(new_n1532, new_n1959, new_n11623);
xor_1  g11247(new_n11623, new_n11622, new_n11624);
nor_1  g11248(new_n1451, new_n2205, new_n11625);
nor_1  g11249(new_n8843, new_n3966, new_n11626);
not_1  g11250(new_n11626, new_n11627);
nor_1  g11251(new_n1539, new_n2363, new_n11628);
not_1  g11252(new_n11628, new_n11629);
nand_1 g11253(new_n11629, new_n11627, new_n11630);
nand_1 g11254(new_n11628, new_n11626, new_n11631);
nand_1 g11255(new_n11631, new_n11630, new_n11632);
xor_1  g11256(new_n11632, new_n11625, new_n11633);
xnor_1 g11257(new_n11633, new_n11624, new_n11634);
xnor_1 g11258(new_n11634, new_n11621, new_n11635);
not_1  g11259(new_n11540, new_n11636);
nand_1 g11260(new_n11636, new_n11532, new_n11637);
nand_1 g11261(new_n11551, new_n11541, new_n11638);
xnor_1 g11262(new_n11638, new_n11539, new_n11639);
nand_1 g11263(new_n11639, new_n11637, new_n11640);
xnor_1 g11264(new_n11640, new_n11635, new_n11641);
xnor_1 g11265(new_n11641, new_n11610, new_n11642);
nand_1 g11266(new_n11556, new_n11529, new_n11643);
nand_1 g11267(new_n11557, new_n11528, new_n11644);
nand_1 g11268(new_n11644, new_n11643, new_n11645);
xnor_1 g11269(new_n11645, new_n11642, new_n11646);
not_1  g11270(new_n11522, new_n11647);
nor_1  g11271(new_n11647, new_n11519, new_n11648);
not_1  g11272(new_n11514, new_n11649);
nand_1 g11273(new_n11517, new_n11649, new_n11650);
nand_1 g11274(new_n11650, new_n11512, new_n11651);
nor_1  g11275(new_n8804, new_n1835_1, new_n11652);
nand_1 g11276(n12947, n8384, new_n11653);
nand_1 g11277(n11999, n7236, new_n11654);
xnor_1 g11278(new_n11654, new_n11653, new_n11655);
xor_1  g11279(new_n11655, new_n11652, new_n11656);
xnor_1 g11280(new_n11656, new_n11651, new_n11657);
nor_1  g11281(new_n11509, new_n11508, new_n11658);
nor_1  g11282(new_n8748, new_n1866, new_n11659);
xor_1  g11283(new_n11659, new_n11658, new_n11660);
nor_1  g11284(new_n1466, new_n2154, new_n11661);
nand_1 g11285(n5198, n1478, new_n11662_1);
nand_1 g11286(n10990, n7646, new_n11663);
xnor_1 g11287(new_n11663, new_n11662_1, new_n11664);
xor_1  g11288(new_n11664, new_n11661, new_n11665);
xnor_1 g11289(new_n11665, new_n11660, new_n11666);
xnor_1 g11290(new_n11666, new_n11657, new_n11667);
not_1  g11291(new_n11504, new_n11668);
nand_1 g11292(new_n11668, new_n11496, new_n11669);
nand_1 g11293(new_n11518, new_n11505, new_n11670);
xnor_1 g11294(new_n11670, new_n11502, new_n11671);
nand_1 g11295(new_n11671, new_n11669, new_n11672);
xnor_1 g11296(new_n11672, new_n11667, new_n11673);
xnor_1 g11297(new_n11673, new_n11648, new_n11674);
nand_1 g11298(new_n11523, new_n11491, new_n11675);
nand_1 g11299(new_n11524, new_n11479, new_n11676);
nand_1 g11300(new_n11676, new_n11675, new_n11677);
xnor_1 g11301(new_n11677, new_n11674, new_n11678);
xnor_1 g11302(new_n11678, new_n11646, new_n11679);
nand_1 g11303(new_n11566, new_n11562, new_n11680);
xnor_1 g11304(new_n11680, new_n11679, new_n11681);
xnor_1 g11305(new_n11681, new_n11607, new_n11682);
xnor_1 g11306(new_n11682, new_n11572, new_n11683);
nand_1 g11307(new_n11683, new_n11204, new_n11684);
xnor_1 g11308(new_n11683, new_n11203, new_n11685);
xnor_1 g11309(new_n11199, new_n11196, new_n11686);
not_1  g11310(new_n11686, new_n11687);
xnor_1 g11311(new_n11195, new_n11194, new_n11688);
not_1  g11312(new_n11487, new_n11689);
xnor_1 g11313(new_n11689, new_n11425, new_n11690);
nand_1 g11314(new_n11690, new_n11688, new_n11691);
not_1  g11315(new_n11688, new_n11692);
xnor_1 g11316(new_n11690, new_n11692, new_n11693);
xor_1  g11317(new_n11193, new_n11188, new_n11694);
xnor_1 g11318(new_n11420, new_n11396, new_n11695);
not_1  g11319(new_n11695, new_n11696);
nor_1  g11320(new_n11696, new_n11694, new_n11697);
not_1  g11321(new_n11697, new_n11698);
xnor_1 g11322(new_n11418, new_n11408, new_n11699);
nand_1 g11323(new_n11143, new_n11141, new_n11700);
nor_1  g11324(new_n11700, new_n11138, new_n11701);
and_1  g11325(new_n11700, new_n11189, new_n11702);
nor_1  g11326(new_n11702, new_n11701, new_n11703);
nand_1 g11327(new_n11703, new_n11699, new_n11704);
not_1  g11328(new_n11704, new_n11705);
nor_1  g11329(new_n11703, new_n11699, new_n11706);
nor_1  g11330(new_n11706, new_n11705, new_n11707_1);
nor_1  g11331(new_n11414, new_n11398, new_n11708);
nor_1  g11332(new_n11708, new_n11415, new_n11709);
nand_1 g11333(new_n11709, new_n11140, new_n11710);
not_1  g11334(new_n11190, new_n11711);
xnor_1 g11335(new_n11191, new_n11711, new_n11712);
not_1  g11336(new_n11712, new_n11713);
nand_1 g11337(new_n11713, new_n11710, new_n11714);
not_1  g11338(new_n11714, new_n11715);
xnor_1 g11339(new_n11416, new_n11415, new_n11716);
not_1  g11340(new_n11716, new_n11717);
nor_1  g11341(new_n11713, new_n11710, new_n11718);
nor_1  g11342(new_n11718, new_n11715, new_n11719);
not_1  g11343(new_n11719, new_n11720);
nor_1  g11344(new_n11720, new_n11717, new_n11721);
nor_1  g11345(new_n11721, new_n11715, new_n11722);
not_1  g11346(new_n11722, new_n11723);
nand_1 g11347(new_n11723, new_n11707_1, new_n11724);
nand_1 g11348(new_n11724, new_n11704, new_n11725);
xnor_1 g11349(new_n11695, new_n11694, new_n11726);
nand_1 g11350(new_n11726, new_n11725, new_n11727);
nand_1 g11351(new_n11727, new_n11698, new_n11728_1);
nand_1 g11352(new_n11728_1, new_n11693, new_n11729);
nand_1 g11353(new_n11729, new_n11691, new_n11730);
nand_1 g11354(new_n11730, new_n11687, new_n11731);
not_1  g11355(new_n11569, new_n11732);
xnor_1 g11356(new_n11570, new_n11732, new_n11733);
xnor_1 g11357(new_n11730, new_n11686, new_n11734);
nand_1 g11358(new_n11734, new_n11733, new_n11735);
nand_1 g11359(new_n11735, new_n11731, new_n11736);
nand_1 g11360(new_n11736, new_n11685, new_n11737);
nand_1 g11361(new_n11737, new_n11684, new_n11738);
not_1  g11362(new_n11607, new_n11739);
not_1  g11363(new_n11681, new_n11740);
nor_1  g11364(new_n11740, new_n11739, new_n11741);
nor_1  g11365(new_n11681, new_n11607, new_n11742);
nor_1  g11366(new_n11742, new_n11572, new_n11743);
nor_1  g11367(new_n11743, new_n11741, new_n11744);
nand_1 g11368(new_n11181, new_n11155, new_n11745);
nand_1 g11369(new_n11201, new_n11182, new_n11746);
nand_1 g11370(new_n11746, new_n11745, new_n11747);
nor_1  g11371(new_n11638, new_n11539, new_n11748);
not_1  g11372(new_n11640, new_n11749);
nor_1  g11373(new_n11749, new_n11635, new_n11750);
nor_1  g11374(new_n11750, new_n11748, new_n11751);
nand_1 g11375(new_n11654, new_n11653, new_n11752);
not_1  g11376(new_n11752, new_n11753);
nor_1  g11377(new_n11655, new_n11652, new_n11754);
nor_1  g11378(new_n11754, new_n11753, new_n11755_1);
nand_1 g11379(n4805, n4436, new_n11756);
nand_1 g11380(n8384, n6441, new_n11757_1);
nand_1 g11381(n11791, n5198, new_n11758);
xnor_1 g11382(new_n11758, new_n11757_1, new_n11759);
xor_1  g11383(new_n11759, new_n11756, new_n11760);
xnor_1 g11384(new_n11760, new_n11755_1, new_n11761);
nand_1 g11385(n7159, n3146, new_n11762);
nand_1 g11386(n11967, n137, new_n11763);
xnor_1 g11387(new_n11763, new_n11762, new_n11764);
nand_1 g11388(n6294, n6254, new_n11765);
nand_1 g11389(n12947, n6358, new_n11766);
xnor_1 g11390(new_n11766, new_n11765, new_n11767);
nand_1 g11391(n11407, n6826, new_n11768);
nand_1 g11392(n7862, n6604, new_n11769);
xnor_1 g11393(new_n11769, new_n11768, new_n11770);
xnor_1 g11394(new_n11770, new_n11767, new_n11771);
xnor_1 g11395(new_n11771, new_n11764, new_n11772);
xnor_1 g11396(new_n11772, new_n11761, new_n11773);
nor_1  g11397(new_n11208, new_n2119, new_n11774);
nand_1 g11398(new_n11623, new_n11622, new_n11775);
not_1  g11399(new_n11633, new_n11776);
nand_1 g11400(new_n11776, new_n11624, new_n11777);
nand_1 g11401(new_n11777, new_n11775, new_n11778);
xnor_1 g11402(new_n11778, new_n11774, new_n11779);
xnor_1 g11403(new_n11779, new_n11773, new_n11780_1);
nand_1 g11404(new_n11619, new_n11616, new_n11781);
not_1  g11405(new_n11634, new_n11782);
nand_1 g11406(new_n11782, new_n11621, new_n11783);
nand_1 g11407(new_n11783, new_n11781, new_n11784);
not_1  g11408(new_n11651, new_n11785);
nand_1 g11409(new_n11656, new_n11785, new_n11786);
not_1  g11410(new_n11666, new_n11787);
nand_1 g11411(new_n11787, new_n11657, new_n11788);
nand_1 g11412(new_n11788, new_n11786, new_n11789);
nor_1  g11413(new_n1931, new_n8911, new_n11790);
not_1  g11414(new_n11615, new_n11791_1);
nor_1  g11415(new_n11791_1, new_n11611, new_n11792);
nor_1  g11416(new_n11792, new_n11612, new_n11793);
nand_1 g11417(new_n11793, new_n11790, new_n11794);
not_1  g11418(new_n11793, new_n11795);
nand_1 g11419(new_n11790, new_n11530, new_n11796);
nand_1 g11420(new_n11796, new_n11795, new_n11797);
nand_1 g11421(new_n11797, new_n11794, new_n11798);
nand_1 g11422(new_n11630, new_n11625, new_n11799);
nand_1 g11423(new_n11799, new_n11631, new_n11800);
xnor_1 g11424(new_n11800, new_n11798, new_n11801);
xnor_1 g11425(new_n11801, new_n11789, new_n11802);
xnor_1 g11426(new_n11802, new_n11784, new_n11803);
xnor_1 g11427(new_n11803, new_n11780_1, new_n11804);
nand_1 g11428(new_n11180, new_n11162, new_n11805);
nand_1 g11429(new_n11805, new_n11159, new_n11806);
nor_1  g11430(new_n8843, new_n2205, new_n11807);
xnor_1 g11431(new_n11807, new_n11806, new_n11808);
xnor_1 g11432(new_n11808, new_n11804, new_n11809);
xnor_1 g11433(new_n11809, new_n11751, new_n11810);
xnor_1 g11434(new_n11810, new_n11747, new_n11811);
xnor_1 g11435(new_n11811, new_n11744, new_n11812);
not_1  g11436(new_n11574, new_n11813);
nand_1 g11437(new_n11599, new_n11813, new_n11814);
nand_1 g11438(new_n11606, new_n11600, new_n11815);
nand_1 g11439(new_n11815, new_n11814, new_n11816);
nand_1 g11440(new_n11641, new_n11609, new_n11817);
nand_1 g11441(new_n11645, new_n11642, new_n11818);
nand_1 g11442(new_n11818, new_n11817, new_n11819);
xnor_1 g11443(new_n11819, new_n11816, new_n11820);
nand_1 g11444(new_n11673, new_n11648, new_n11821_1);
not_1  g11445(new_n11674, new_n11822);
nand_1 g11446(new_n11677, new_n11822, new_n11823);
nand_1 g11447(new_n11823, new_n11821_1, new_n11824);
not_1  g11448(new_n11588, new_n11825);
nand_1 g11449(new_n11825, new_n11583, new_n11826);
nand_1 g11450(new_n11597, new_n11589, new_n11827);
nand_1 g11451(new_n11827, new_n11826, new_n11828);
nand_1 g11452(new_n11586, new_n11585, new_n11829);
not_1  g11453(new_n11829, new_n11830);
nor_1  g11454(new_n11587, new_n11584, new_n11831);
nor_1  g11455(new_n11831, new_n11830, new_n11832);
nand_1 g11456(n5283, n447, new_n11833);
nand_1 g11457(n11999, n3992, new_n11834);
xnor_1 g11458(new_n11834, new_n11833, new_n11835);
xnor_1 g11459(new_n11835, new_n11832, new_n11836);
xnor_1 g11460(new_n11836, new_n11828, new_n11837);
nand_1 g11461(n7646, n5760, new_n11838);
nand_1 g11462(n10990, n4722, new_n11839);
xnor_1 g11463(new_n11839, new_n11838, new_n11840);
xnor_1 g11464(new_n11840, new_n11837, new_n11841);
xnor_1 g11465(new_n11841, new_n11824, new_n11842);
xnor_1 g11466(new_n11842, new_n11820, new_n11843);
not_1  g11467(new_n11646, new_n11844);
nand_1 g11468(new_n11678, new_n11844, new_n11845);
not_1  g11469(new_n11680, new_n11846);
nand_1 g11470(new_n11846, new_n11679, new_n11847);
nand_1 g11471(new_n11847, new_n11845, new_n11848);
not_1  g11472(new_n11598, new_n11849);
nand_1 g11473(new_n11849, new_n11579, new_n11850);
nand_1 g11474(new_n11850, new_n11576, new_n11851);
nand_1 g11475(new_n11178, new_n11172, new_n11852);
nand_1 g11476(new_n11179, new_n11170, new_n11853);
nand_1 g11477(new_n11853, new_n11852, new_n11854);
nand_1 g11478(new_n11594, new_n11593, new_n11855);
not_1  g11479(new_n11855, new_n11856);
nor_1  g11480(new_n11595, new_n11592, new_n11857);
nor_1  g11481(new_n11857, new_n11856, new_n11858);
nor_1  g11482(new_n8561, new_n1600, new_n11859);
nand_1 g11483(n9725, n1333, new_n11860);
nand_1 g11484(n12709, n10174, new_n11861);
xnor_1 g11485(new_n11861, new_n11860, new_n11862);
xnor_1 g11486(new_n11862, new_n11859, new_n11863);
xnor_1 g11487(new_n11863, new_n11858, new_n11864);
nor_1  g11488(new_n11590, new_n11266, new_n11865);
not_1  g11489(new_n11591, new_n11866);
nor_1  g11490(new_n11596, new_n11866, new_n11867);
nor_1  g11491(new_n11867, new_n11865, new_n11868);
nand_1 g11492(new_n11663, new_n11662_1, new_n11869);
not_1  g11493(new_n11869, new_n11870);
nor_1  g11494(new_n11664, new_n11661, new_n11871);
nor_1  g11495(new_n11871, new_n11870, new_n11872);
nand_1 g11496(n6877, n1198, new_n11873);
nor_1  g11497(new_n2450, new_n1435, new_n11874);
xnor_1 g11498(new_n11874, new_n11873, new_n11875);
xnor_1 g11499(new_n11875, new_n11872, new_n11876_1);
xnor_1 g11500(new_n11876_1, new_n11868, new_n11877_1);
xnor_1 g11501(new_n11877_1, new_n11864, new_n11878);
xnor_1 g11502(new_n11878, new_n11854, new_n11879);
nor_1  g11503(new_n1539, new_n7664, new_n11880);
nand_1 g11504(new_n11176, new_n11175, new_n11881);
not_1  g11505(new_n11881, new_n11882);
nor_1  g11506(new_n11177, new_n11174, new_n11883);
nor_1  g11507(new_n11883, new_n11882, new_n11884);
nand_1 g11508(n11757, n5320, new_n11885);
nand_1 g11509(n9080, n5212, new_n11886);
xnor_1 g11510(new_n11886, new_n11885, new_n11887);
nand_1 g11511(n11877, n11821, new_n11888);
nand_1 g11512(n5240, n4370, new_n11889);
xnor_1 g11513(new_n11889, new_n11888, new_n11890);
xnor_1 g11514(new_n11890, new_n11887, new_n11891);
xnor_1 g11515(new_n11891, new_n11884, new_n11892_1);
nand_1 g11516(n9400, n7730, new_n11893);
nor_1  g11517(new_n1747, new_n8622, new_n11894);
xnor_1 g11518(new_n11894, new_n11893, new_n11895);
xnor_1 g11519(new_n11895, new_n11892_1, new_n11896);
nand_1 g11520(new_n11167, new_n11166, new_n11897);
not_1  g11521(new_n11897, new_n11898);
not_1  g11522(new_n11165, new_n11899);
nor_1  g11523(new_n11168, new_n11899, new_n11900);
nor_1  g11524(new_n11900, new_n11898, new_n11901);
nand_1 g11525(new_n11163, new_n11080, new_n11902);
nand_1 g11526(new_n11169, new_n11164, new_n11903);
nand_1 g11527(new_n11903, new_n11902, new_n11904);
xnor_1 g11528(new_n11904, new_n11901, new_n11905);
xnor_1 g11529(new_n11905, new_n11896, new_n11906);
xnor_1 g11530(new_n11906, new_n11880, new_n11907);
xnor_1 g11531(new_n11907, new_n11879, new_n11908);
xnor_1 g11532(new_n11908, new_n11851, new_n11909);
or_1   g11533(new_n11670, new_n11502, new_n11910);
not_1  g11534(new_n11667, new_n11911);
nand_1 g11535(new_n11672, new_n11911, new_n11912);
nand_1 g11536(new_n11912, new_n11910, new_n11913);
nand_1 g11537(n8819, n4187, new_n11914);
nand_1 g11538(n1478, n1471, new_n11915);
xnor_1 g11539(new_n11915, new_n11914, new_n11916);
nand_1 g11540(n8717, n2464, new_n11917_1);
nand_1 g11541(n10022, n7236, new_n11918);
xnor_1 g11542(new_n11918, new_n11917_1, new_n11919_1);
xnor_1 g11543(new_n11919_1, new_n11916, new_n11920);
nand_1 g11544(new_n11659, new_n11658, new_n11921);
not_1  g11545(new_n11665, new_n11922_1);
nand_1 g11546(new_n11922_1, new_n11660, new_n11923);
nand_1 g11547(new_n11923, new_n11921, new_n11924);
xnor_1 g11548(new_n11924, new_n11920, new_n11925);
xnor_1 g11549(new_n11925, new_n11913, new_n11926);
xnor_1 g11550(new_n11926, new_n11909, new_n11927);
xnor_1 g11551(new_n11927, new_n11848, new_n11928);
xnor_1 g11552(new_n11928, new_n11843, new_n11929);
xnor_1 g11553(new_n11929, new_n11812, new_n11930);
xnor_1 g11554(new_n11930, new_n11738, n4378);
xnor_1 g11555(new_n4167, new_n4050, n4397);
xnor_1 g11556(new_n4501, new_n4270, n4553);
xnor_1 g11557(new_n977, new_n972, n4686);
xnor_1 g11558(new_n9907, new_n9887, n4689);
not_1  g11559(new_n5302, new_n11936);
xnor_1 g11560(new_n11936, new_n5301, n4733);
xnor_1 g11561(new_n2268, new_n2260, n4757);
xnor_1 g11562(new_n5297, new_n5296, n4971);
xnor_1 g11563(new_n7030, new_n7028, n5030);
xnor_1 g11564(new_n3147, new_n3115, n5034);
xnor_1 g11565(new_n3142, new_n3128, n5094);
nand_1 g11566(new_n10939, new_n10935, new_n11943);
nand_1 g11567(new_n10950, new_n11943, new_n11944);
nor_1  g11568(new_n8515, new_n1377, new_n11945);
not_1  g11569(new_n11945, new_n11946);
nor_1  g11570(new_n1365, new_n1367, new_n11947);
not_1  g11571(new_n11947, new_n11948);
nand_1 g11572(new_n11948, new_n11946, new_n11949);
nor_1  g11573(new_n11948, new_n11946, new_n11950);
not_1  g11574(new_n11950, new_n11951);
nand_1 g11575(new_n11951, new_n11949, new_n11952);
xnor_1 g11576(new_n11952, new_n11944, new_n11953);
nor_1  g11577(new_n1371, new_n4283, new_n11954);
nand_1 g11578(new_n10944, new_n10943, new_n11955);
not_1  g11579(new_n11955, new_n11956);
nor_1  g11580(new_n10947, new_n11956, new_n11957);
nand_1 g11581(new_n11957, new_n11954, new_n11958);
not_1  g11582(new_n11958, new_n11959);
nor_1  g11583(new_n11957, new_n11954, new_n11960);
nor_1  g11584(new_n11960, new_n11959, new_n11961);
nand_1 g11585(n9920, n5212, new_n11962);
nand_1 g11586(n11407, n3627, new_n11963);
xor_1  g11587(new_n11963, new_n11962, new_n11964);
xnor_1 g11588(new_n11964, new_n11961, new_n11965);
not_1  g11589(new_n11965, new_n11966);
nand_1 g11590(new_n11966, new_n11953, new_n11967_1);
not_1  g11591(new_n11967_1, new_n11968);
nor_1  g11592(new_n11966, new_n11953, new_n11969);
nor_1  g11593(new_n11969, new_n11968, new_n11970);
nand_1 g11594(new_n10933, new_n10932, new_n11971);
not_1  g11595(new_n11971, new_n11972);
nor_1  g11596(new_n10953, new_n10934, new_n11973);
nor_1  g11597(new_n11973, new_n11972, new_n11974);
not_1  g11598(new_n11974, new_n11975);
nand_1 g11599(new_n11975, new_n11970, new_n11976);
nand_1 g11600(new_n11964, new_n11961, new_n11977);
nand_1 g11601(new_n11977, new_n11958, new_n11978);
nor_1  g11602(new_n8561, new_n1377, new_n11979);
nor_1  g11603(new_n8515, new_n1367, new_n11980);
not_1  g11604(new_n11980, new_n11981);
nor_1  g11605(new_n9075, new_n378, new_n11982);
not_1  g11606(new_n11982, new_n11983);
nand_1 g11607(new_n11983, new_n11981, new_n11984);
nand_1 g11608(new_n11982, new_n11980, new_n11985);
nand_1 g11609(new_n11985, new_n11984, new_n11986);
xor_1  g11610(new_n11986, new_n11979, new_n11987);
xnor_1 g11611(new_n11987, new_n11978, new_n11988);
nor_1  g11612(new_n11963, new_n11962, new_n11989);
nor_1  g11613(new_n4283, new_n1365, new_n11990);
xor_1  g11614(new_n11990, new_n11989, new_n11991);
nor_1  g11615(new_n1378, new_n6617, new_n11992);
not_1  g11616(n9920, new_n11993);
nor_1  g11617(new_n1371, new_n11993, new_n11994);
not_1  g11618(new_n11994, new_n11995);
nand_1 g11619(n11407, n4516, new_n11996);
nand_1 g11620(new_n11996, new_n11995, new_n11997);
not_1  g11621(new_n11996, new_n11998);
nand_1 g11622(new_n11998, new_n11994, new_n11999_1);
nand_1 g11623(new_n11999_1, new_n11997, new_n12000_1);
xnor_1 g11624(new_n12000_1, new_n11992, new_n12001);
not_1  g11625(new_n12001, new_n12002);
xnor_1 g11626(new_n12002, new_n11991, new_n12003);
xnor_1 g11627(new_n12003, new_n11988, new_n12004);
not_1  g11628(new_n11952, new_n12005_1);
nand_1 g11629(new_n12005_1, new_n11944, new_n12006);
nand_1 g11630(new_n11968, new_n11950, new_n12007);
nand_1 g11631(new_n11967_1, new_n11951, new_n12008);
nand_1 g11632(new_n12008, new_n12007, new_n12009);
nand_1 g11633(new_n12009, new_n12006, new_n12010);
xnor_1 g11634(new_n12010, new_n12004, new_n12011);
xnor_1 g11635(new_n12011, new_n11976, new_n12012);
nor_1  g11636(new_n8561, new_n378, new_n12013);
not_1  g11637(new_n11976, new_n12014_1);
nor_1  g11638(new_n11975, new_n11970, new_n12015);
nor_1  g11639(new_n12015, new_n12014_1, new_n12016);
nand_1 g11640(new_n12016, new_n12013, new_n12017);
not_1  g11641(new_n10955, new_n12018);
nor_1  g11642(new_n12018, new_n10931, new_n12019);
not_1  g11643(new_n12013, new_n12020_1);
xnor_1 g11644(new_n12016, new_n12020_1, new_n12021);
nand_1 g11645(new_n12021, new_n12019, new_n12022);
nand_1 g11646(new_n12022, new_n12017, new_n12023);
xor_1  g11647(new_n12023, new_n12012, new_n12024);
nor_1  g11648(new_n8602, new_n382, new_n12025_1);
nor_1  g11649(new_n11208, new_n4529, new_n12026);
not_1  g11650(new_n12026, new_n12027);
nand_1 g11651(n11728, n1094, new_n12028);
nand_1 g11652(n12709, n10678, new_n12029);
xnor_1 g11653(new_n12029, new_n12028, new_n12030);
nor_1  g11654(new_n12030, new_n12027, new_n12031);
not_1  g11655(new_n12031, new_n12032);
nand_1 g11656(new_n12030, new_n12027, new_n12033);
nand_1 g11657(new_n12033, new_n12032, new_n12034);
not_1  g11658(new_n10965_1, new_n12035);
not_1  g11659(new_n10968, new_n12036);
nor_1  g11660(new_n12036, new_n10963, new_n12037);
nor_1  g11661(new_n12037, new_n12035, new_n12038);
xnor_1 g11662(new_n12038, new_n12034, new_n12039);
nand_1 g11663(n10928, n2433, new_n12040);
nand_1 g11664(n8819, n6986, new_n12041);
nand_1 g11665(new_n12041, new_n12040, new_n12042);
nor_1  g11666(new_n12041, new_n12040, new_n12043);
not_1  g11667(new_n12043, new_n12044_1);
nand_1 g11668(new_n12044_1, new_n12042, new_n12045);
xnor_1 g11669(new_n12045, new_n12039, new_n12046);
nand_1 g11670(new_n10961, new_n10958, new_n12047);
not_1  g11671(new_n12047, new_n12048);
not_1  g11672(new_n10970, new_n12049);
nor_1  g11673(new_n12049, new_n10962, new_n12050);
nor_1  g11674(new_n12050, new_n12048, new_n12051);
not_1  g11675(new_n12051, new_n12052);
xnor_1 g11676(new_n12052, new_n12046, new_n12053);
not_1  g11677(new_n12053, new_n12054);
nand_1 g11678(new_n10979, new_n10972, new_n12055);
nand_1 g11679(new_n12055, new_n12054, new_n12056);
not_1  g11680(new_n12056, new_n12057);
nor_1  g11681(new_n12055, new_n12054, new_n12058);
nor_1  g11682(new_n12058, new_n12057, new_n12059);
nand_1 g11683(new_n12059, new_n12025_1, new_n12060);
and_1  g11684(new_n10981, new_n1529, new_n12061);
not_1  g11685(new_n12025_1, new_n12062);
xnor_1 g11686(new_n12059, new_n12062, new_n12063);
nand_1 g11687(new_n12063, new_n12061, new_n12064);
nand_1 g11688(new_n12064, new_n12060, new_n12065);
not_1  g11689(new_n12034, new_n12066);
nand_1 g11690(new_n12038, new_n12066, new_n12067);
nand_1 g11691(new_n12067, new_n12032, new_n12068);
nor_1  g11692(new_n1434, new_n8602, new_n12069_1);
nand_1 g11693(n6986, n2433, new_n12070);
nand_1 g11694(n8336, n7730, new_n12071);
xnor_1 g11695(new_n12071, new_n12070, new_n12072);
xor_1  g11696(new_n12072, new_n12069_1, new_n12073);
xnor_1 g11697(new_n12073, new_n12068, new_n12074);
nor_1  g11698(new_n12029, new_n12028, new_n12075);
nor_1  g11699(new_n1506, new_n4529, new_n12076_1);
xor_1  g11700(new_n12076_1, new_n12075, new_n12077);
nor_1  g11701(new_n1435, new_n6725, new_n12078);
nand_1 g11702(n6429, n1094, new_n12079);
nand_1 g11703(n12709, n7320, new_n12080);
xnor_1 g11704(new_n12080, new_n12079, new_n12081);
xor_1  g11705(new_n12081, new_n12078, new_n12082);
xnor_1 g11706(new_n12082, new_n12077, new_n12083);
xnor_1 g11707(new_n12083, new_n12074, new_n12084);
not_1  g11708(new_n12045, new_n12085);
nand_1 g11709(new_n12085, new_n12039, new_n12086);
nand_1 g11710(new_n12052, new_n12046, new_n12087);
not_1  g11711(new_n12087, new_n12088);
nand_1 g11712(new_n12088, new_n12043, new_n12089);
nand_1 g11713(new_n12087, new_n12044_1, new_n12090);
nand_1 g11714(new_n12090, new_n12089, new_n12091);
nand_1 g11715(new_n12091, new_n12086, new_n12092);
xnor_1 g11716(new_n12092, new_n12084, new_n12093);
xnor_1 g11717(new_n12093, new_n12056, new_n12094);
xnor_1 g11718(new_n12094, new_n12065, new_n12095);
not_1  g11719(new_n12095, new_n12096);
xnor_1 g11720(new_n12063, new_n12061, new_n12097);
not_1  g11721(new_n10982, new_n12098);
nand_1 g11722(new_n10984, new_n12098, new_n12099);
nand_1 g11723(new_n11061, new_n12099, new_n12100);
not_1  g11724(new_n12100, new_n12101);
nand_1 g11725(new_n12101, new_n12097, new_n12102);
not_1  g11726(new_n11053, new_n12103);
nand_1 g11727(new_n12103, new_n11023_1, new_n12104);
nor_1  g11728(new_n385, new_n8804, new_n12105);
nand_1 g11729(new_n11030, new_n11025, new_n12106);
nand_1 g11730(new_n11041, new_n12106, new_n12107);
nor_1  g11731(new_n8768, new_n1467, new_n12108);
not_1  g11732(new_n12108, new_n12109);
nor_1  g11733(new_n8748, new_n1562, new_n12110);
not_1  g11734(new_n12110, new_n12111_1);
nand_1 g11735(new_n12111_1, new_n12109, new_n12112);
nor_1  g11736(new_n12111_1, new_n12109, new_n12113);
not_1  g11737(new_n12113, new_n12114);
nand_1 g11738(new_n12114, new_n12112, new_n12115);
xnor_1 g11739(new_n12115, new_n12107, new_n12116);
nor_1  g11740(new_n8469, new_n4542, new_n12117);
not_1  g11741(new_n12117, new_n12118);
nand_1 g11742(n10990, n5319, new_n12119);
nand_1 g11743(n5767, n5760, new_n12120);
xnor_1 g11744(new_n12120, new_n12119, new_n12121);
nor_1  g11745(new_n12121, new_n12118, new_n12122);
not_1  g11746(new_n12122, new_n12123);
nand_1 g11747(new_n12121, new_n12118, new_n12124);
nand_1 g11748(new_n12124, new_n12123, new_n12125);
not_1  g11749(new_n11037, new_n12126);
not_1  g11750(new_n11038, new_n12127);
nor_1  g11751(new_n12127, new_n11032, new_n12128);
nor_1  g11752(new_n12128, new_n12126, new_n12129);
xnor_1 g11753(new_n12129, new_n12125, new_n12130);
xnor_1 g11754(new_n12130, new_n12116, new_n12131);
not_1  g11755(new_n12131, new_n12132);
nand_1 g11756(new_n11052, new_n11048, new_n12133);
nand_1 g11757(new_n12133, new_n11045, new_n12134);
nand_1 g11758(new_n12134, new_n12132, new_n12135);
not_1  g11759(new_n12135, new_n12136);
nor_1  g11760(new_n12134, new_n12132, new_n12137);
nor_1  g11761(new_n12137, new_n12136, new_n12138);
nand_1 g11762(new_n12138, new_n12105, new_n12139);
not_1  g11763(new_n12139, new_n12140);
nor_1  g11764(new_n12138, new_n12105, new_n12141);
nor_1  g11765(new_n12141, new_n12140, new_n12142);
not_1  g11766(new_n12142, new_n12143);
nor_1  g11767(new_n12143, new_n12104, new_n12144);
not_1  g11768(new_n12104, new_n12145_1);
nor_1  g11769(new_n12142, new_n12145_1, new_n12146);
nor_1  g11770(new_n12146, new_n12144, new_n12147);
nand_1 g11771(new_n11019, new_n1552, new_n12148);
nor_1  g11772(new_n1533, new_n8942, new_n12149);
not_1  g11773(new_n12149, new_n12150);
nand_1 g11774(n12777, n7160, new_n12151);
nand_1 g11775(n7159, n4828, new_n12152);
nand_1 g11776(n12489, n2515, new_n12153);
xnor_1 g11777(new_n12153, new_n12152, new_n12154);
nor_1  g11778(new_n12154, new_n12151, new_n12155);
not_1  g11779(new_n12155, new_n12156);
nand_1 g11780(new_n12154, new_n12151, new_n12157);
nand_1 g11781(new_n12157, new_n12156, new_n12158);
not_1  g11782(new_n11002, new_n12159);
nor_1  g11783(new_n11003, new_n10997, new_n12160);
nor_1  g11784(new_n12160, new_n12159, new_n12161);
xnor_1 g11785(new_n12161, new_n12158, new_n12162);
nor_1  g11786(new_n1452, new_n8888, new_n12163);
not_1  g11787(new_n12163, new_n12164);
nor_1  g11788(new_n4386, new_n1532, new_n12165);
not_1  g11789(new_n12165, new_n12166);
nand_1 g11790(new_n12166, new_n12164, new_n12167);
nor_1  g11791(new_n12166, new_n12164, new_n12168);
not_1  g11792(new_n12168, new_n12169);
nand_1 g11793(new_n12169, new_n12167, new_n12170);
xnor_1 g11794(new_n12170, new_n12162, new_n12171);
nand_1 g11795(new_n11007, new_n10993, new_n12172);
xnor_1 g11796(new_n12172, new_n12171, new_n12173);
nand_1 g11797(new_n11010, new_n10986, new_n12174);
nand_1 g11798(new_n11016, new_n12174, new_n12175);
xnor_1 g11799(new_n12175, new_n12173, new_n12176);
xnor_1 g11800(new_n12176, new_n12150, new_n12177);
nor_1  g11801(new_n12177, new_n12148, new_n12178);
nand_1 g11802(new_n12177, new_n12148, new_n12179);
not_1  g11803(new_n12179, new_n12180);
nor_1  g11804(new_n12180, new_n12178, new_n12181);
not_1  g11805(new_n11058, new_n12182);
nand_1 g11806(new_n12182, new_n11054, new_n12183);
nand_1 g11807(new_n11059, new_n11020, new_n12184);
nand_1 g11808(new_n12184, new_n12183, new_n12185);
xnor_1 g11809(new_n12185, new_n12181, new_n12186);
xnor_1 g11810(new_n12186, new_n12147, new_n12187);
xnor_1 g11811(new_n12100, new_n12097, new_n12188);
nand_1 g11812(new_n12188, new_n12187, new_n12189);
nand_1 g11813(new_n12189, new_n12102, new_n12190);
xnor_1 g11814(new_n12190, new_n12096, new_n12191);
not_1  g11815(new_n12125, new_n12192);
nand_1 g11816(new_n12129, new_n12192, new_n12193);
nand_1 g11817(new_n12193, new_n12123, new_n12194);
nor_1  g11818(new_n1467, new_n8804, new_n12195);
nand_1 g11819(n12947, n5314, new_n12196);
nand_1 g11820(n11999, n11222, new_n12197);
xnor_1 g11821(new_n12197, new_n12196, new_n12198);
xor_1  g11822(new_n12198, new_n12195, new_n12199);
xnor_1 g11823(new_n12199, new_n12194, new_n12200);
nor_1  g11824(new_n12120, new_n12119, new_n12201);
nor_1  g11825(new_n8748, new_n4542, new_n12202);
xor_1  g11826(new_n12202, new_n12201, new_n12203);
nor_1  g11827(new_n1466, new_n6935, new_n12204);
nand_1 g11828(n5767, n1478, new_n12205);
nand_1 g11829(n10990, n9457, new_n12206);
xnor_1 g11830(new_n12206, new_n12205, new_n12207);
xnor_1 g11831(new_n12207, new_n12204, new_n12208);
not_1  g11832(new_n12208, new_n12209);
xnor_1 g11833(new_n12209, new_n12203, new_n12210);
xnor_1 g11834(new_n12210, new_n12200, new_n12211);
not_1  g11835(new_n12115, new_n12212);
nand_1 g11836(new_n12212, new_n12107, new_n12213);
nand_1 g11837(new_n12130, new_n12116, new_n12214);
xnor_1 g11838(new_n12214, new_n12114, new_n12215);
nand_1 g11839(new_n12215, new_n12213, new_n12216);
xnor_1 g11840(new_n12216, new_n12211, new_n12217);
xnor_1 g11841(new_n12217, new_n12135, new_n12218);
nor_1  g11842(new_n12144, new_n12140, new_n12219);
xnor_1 g11843(new_n12219, new_n12218, new_n12220);
not_1  g11844(new_n12173, new_n12221_1);
nand_1 g11845(new_n12175, new_n12221_1, new_n12222);
not_1  g11846(new_n12158, new_n12223);
nand_1 g11847(new_n12161, new_n12223, new_n12224);
nand_1 g11848(new_n12224, new_n12156, new_n12225);
nor_1  g11849(new_n1452, new_n8942, new_n12226);
nor_1  g11850(new_n8888, new_n4386, new_n12227);
not_1  g11851(new_n12227, new_n12228);
nor_1  g11852(new_n1533, new_n8911, new_n12229);
not_1  g11853(new_n12229, new_n12230);
nand_1 g11854(new_n12230, new_n12228, new_n12231);
nand_1 g11855(new_n12229, new_n12227, new_n12232);
nand_1 g11856(new_n12232, new_n12231, new_n12233);
xnor_1 g11857(new_n12233, new_n12226, new_n12234);
nand_1 g11858(new_n12234, new_n12225, new_n12235);
not_1  g11859(new_n12225, new_n12236);
not_1  g11860(new_n12234, new_n12237);
nand_1 g11861(new_n12237, new_n12236, new_n12238);
nand_1 g11862(new_n12238, new_n12235, new_n12239);
not_1  g11863(new_n12239, new_n12240);
nor_1  g11864(new_n12153, new_n12152, new_n12241);
nor_1  g11865(new_n1538, new_n1532, new_n12242);
xor_1  g11866(new_n12242, new_n12241, new_n12243);
nand_1 g11867(n7159, n2515, new_n12244);
nand_1 g11868(n12777, n4828, new_n12245);
nand_1 g11869(n12489, n1199, new_n12246);
xnor_1 g11870(new_n12246, new_n12245, new_n12247_1);
xnor_1 g11871(new_n12247_1, new_n12244, new_n12248);
xnor_1 g11872(new_n12248, new_n12243, new_n12249);
not_1  g11873(new_n12249, new_n12250);
nand_1 g11874(new_n12250, new_n12240, new_n12251);
nand_1 g11875(new_n12249, new_n12239, new_n12252);
nand_1 g11876(new_n12252, new_n12251, new_n12253);
not_1  g11877(new_n12253, new_n12254);
not_1  g11878(new_n12170, new_n12255);
nand_1 g11879(new_n12255, new_n12162, new_n12256);
nand_1 g11880(new_n12172, new_n12171, new_n12257);
not_1  g11881(new_n12257, new_n12258);
nand_1 g11882(new_n12258, new_n12168, new_n12259);
nand_1 g11883(new_n12257, new_n12169, new_n12260);
nand_1 g11884(new_n12260, new_n12259, new_n12261);
nand_1 g11885(new_n12261, new_n12256, new_n12262);
xnor_1 g11886(new_n12262, new_n12254, new_n12263);
xnor_1 g11887(new_n12263, new_n12222, new_n12264);
nor_1  g11888(new_n12176, new_n12149, new_n12265);
not_1  g11889(new_n12265, new_n12266);
nand_1 g11890(new_n12179, new_n12266, new_n12267);
xnor_1 g11891(new_n12267, new_n12264, new_n12268);
xnor_1 g11892(new_n12268, new_n12220, new_n12269);
not_1  g11893(new_n12181, new_n12270);
nand_1 g11894(new_n12185, new_n12270, new_n12271);
nand_1 g11895(new_n12186, new_n12147, new_n12272);
nand_1 g11896(new_n12272, new_n12271, new_n12273);
xnor_1 g11897(new_n12273, new_n12269, new_n12274);
xnor_1 g11898(new_n12274, new_n12191, new_n12275);
xnor_1 g11899(new_n12275, new_n12024, new_n12276);
xnor_1 g11900(new_n12021, new_n12019, new_n12277);
nand_1 g11901(new_n11073, new_n11068, new_n12278);
nand_1 g11902(new_n12278, new_n11066, new_n12279);
not_1  g11903(new_n12279, new_n12280);
nand_1 g11904(new_n12280, new_n12277, new_n12281);
xnor_1 g11905(new_n12279, new_n12277, new_n12282);
not_1  g11906(new_n12189, new_n12283);
nor_1  g11907(new_n12188, new_n12187, new_n12284);
nor_1  g11908(new_n12284, new_n12283, new_n12285);
nand_1 g11909(new_n12285, new_n12282, new_n12286);
nand_1 g11910(new_n12286, new_n12281, new_n12287);
xnor_1 g11911(new_n12287, new_n12276, n5132);
xnor_1 g11912(new_n11709, new_n11141, n5191);
not_1  g11913(new_n4042, new_n12290);
nor_1  g11914(new_n12290, new_n3906, new_n12291);
nor_1  g11915(new_n12291, new_n3905, new_n12292);
nor_1  g11916(new_n4038, new_n3950, new_n12293);
not_1  g11917(new_n4041, new_n12294);
nor_1  g11918(new_n12294, new_n4039, new_n12295);
nor_1  g11919(new_n12295, new_n12293, new_n12296);
nand_1 g11920(new_n3454, new_n3457, new_n12297);
nand_1 g11921(new_n3473, new_n3455, new_n12298);
nand_1 g11922(new_n12298, new_n12297, new_n12299_1);
nand_1 g11923(new_n3453, new_n3446, new_n12300);
nand_1 g11924(new_n12300, new_n3450, new_n12301);
nor_1  g11925(new_n1931, new_n3952, new_n12302);
nand_1 g11926(new_n3928, new_n3927, new_n12303);
not_1  g11927(new_n3934, new_n12304);
nand_1 g11928(new_n12304, new_n3929, new_n12305);
nand_1 g11929(new_n12305, new_n12303, new_n12306);
nand_1 g11930(n8433, n4722, new_n12307);
nand_1 g11931(n8065, n2464, new_n12308);
nand_1 g11932(n7646, n405, new_n12309);
xnor_1 g11933(new_n12309, new_n12308, new_n12310);
xor_1  g11934(new_n12310, new_n12307, new_n12311);
xnor_1 g11935(new_n12311, new_n12306, new_n12312);
xnor_1 g11936(new_n12312, new_n12302, new_n12313);
xnor_1 g11937(new_n12313, new_n12301, new_n12314);
not_1  g11938(new_n4000, new_n12315);
nand_1 g11939(new_n12315, new_n3997, new_n12316);
not_1  g11940(new_n4018, new_n12317);
nand_1 g11941(new_n12317, new_n4001, new_n12318);
nand_1 g11942(new_n12318, new_n12316, new_n12319);
nand_1 g11943(new_n3963, new_n3962, new_n12320);
nand_1 g11944(new_n3975, new_n3964, new_n12321);
nand_1 g11945(new_n12321, new_n12320, new_n12322);
nand_1 g11946(new_n4003, new_n4002, new_n12323);
nand_1 g11947(new_n4016, new_n4004, new_n12324);
nand_1 g11948(new_n12324, new_n12323, new_n12325);
xnor_1 g11949(new_n12325, new_n12322, new_n12326);
nand_1 g11950(n8384, n6359, new_n12327);
nand_1 g11951(n7546, n4805, new_n12328);
xnor_1 g11952(new_n12328, new_n12327, new_n12329);
nand_1 g11953(n12925, n4938, new_n12330);
nand_1 g11954(n11536, n7862, new_n12331);
xnor_1 g11955(new_n12331, new_n12330, new_n12332);
nand_1 g11956(new_n4013, new_n4005_1, new_n12333);
nand_1 g11957(new_n12333, new_n4014, new_n12334);
xnor_1 g11958(new_n12334, new_n12332, new_n12335);
xnor_1 g11959(new_n12335, new_n12329, new_n12336);
xnor_1 g11960(new_n12336, new_n12326, new_n12337);
xnor_1 g11961(new_n12337, new_n12319, new_n12338);
not_1  g11962(new_n3960, new_n12339);
nand_1 g11963(new_n12339, new_n3957, new_n12340);
nand_1 g11964(new_n3976, new_n3961, new_n12341);
nand_1 g11965(new_n12341, new_n12340, new_n12342);
nand_1 g11966(new_n3995, new_n3994, new_n12343);
not_1  g11967(new_n12343, new_n12344);
nor_1  g11968(new_n3996, new_n3993, new_n12345);
nor_1  g11969(new_n12345, new_n12344, new_n12346);
nand_1 g11970(n9956, n6826, new_n12347);
nand_1 g11971(n6797, n4826, new_n12348);
xnor_1 g11972(new_n12348, new_n12347, new_n12349);
nand_1 g11973(n7610, n6294, new_n12350);
nand_1 g11974(n6611, n6358, new_n12351);
xnor_1 g11975(new_n12351, new_n12350, new_n12352);
xnor_1 g11976(new_n12352, new_n12349, new_n12353);
xnor_1 g11977(new_n12353, new_n12346, new_n12354);
nand_1 g11978(n7733, n3146, new_n12355);
nand_1 g11979(new_n3955, new_n3954, new_n12356);
not_1  g11980(new_n12356, new_n12357);
nor_1  g11981(new_n3956, new_n3953, new_n12358);
nor_1  g11982(new_n12358, new_n12357, new_n12359);
xnor_1 g11983(new_n12359, new_n12355, new_n12360);
xnor_1 g11984(new_n12360, new_n12354, new_n12361);
nand_1 g11985(n5198, n217, new_n12362);
nand_1 g11986(n5283, n503, new_n12363);
xnor_1 g11987(new_n12363, new_n12362, new_n12364);
nand_1 g11988(n4970, n137, new_n12365);
nand_1 g11989(n11296, n3992, new_n12366);
xnor_1 g11990(new_n12366, new_n12365, new_n12367);
xnor_1 g11991(new_n12367, new_n12364, new_n12368);
nand_1 g11992(new_n3972, new_n3965, new_n12369);
nand_1 g11993(new_n12369, new_n3973, new_n12370);
nand_1 g11994(n11311, n10439, new_n12371);
nor_1  g11995(new_n2725, new_n2119, new_n12372);
xnor_1 g11996(new_n12372, new_n12371, new_n12373);
xnor_1 g11997(new_n12373, new_n12370, new_n12374);
xnor_1 g11998(new_n12374, new_n12368, new_n12375);
xnor_1 g11999(new_n12375, new_n12361, new_n12376);
xnor_1 g12000(new_n12376, new_n12342, new_n12377);
xnor_1 g12001(new_n12377, new_n12338, new_n12378);
not_1  g12002(new_n3936, new_n12379);
nand_1 g12003(new_n3944, new_n12379, new_n12380);
nand_1 g12004(new_n12380, new_n3941, new_n12381);
not_1  g12005(new_n3978, new_n12382);
nand_1 g12006(new_n3984, new_n12382, new_n12383);
nand_1 g12007(new_n12383, new_n3981, new_n12384);
xnor_1 g12008(new_n12384, new_n12381, new_n12385);
xnor_1 g12009(new_n12385, new_n12378, new_n12386);
xnor_1 g12010(new_n12386, new_n12314, new_n12387);
xnor_1 g12011(new_n12387, new_n12299_1, new_n12388);
nand_1 g12012(new_n3945, new_n3571, new_n12389);
not_1  g12013(new_n3949, new_n12390);
nand_1 g12014(new_n12390, new_n3946, new_n12391_1);
nand_1 g12015(new_n12391_1, new_n12389, new_n12392);
not_1  g12016(new_n3935, new_n12393);
nand_1 g12017(new_n12393, new_n3926, new_n12394);
nand_1 g12018(new_n12394, new_n3924, new_n12395);
nor_1  g12019(new_n3772, new_n2154, new_n12396);
nor_1  g12020(new_n3287_1, new_n1735, new_n12397);
nor_1  g12021(new_n3915, new_n3910, new_n12398);
nand_1 g12022(new_n12398, new_n12397, new_n12399);
not_1  g12023(new_n12398, new_n12400);
nand_1 g12024(new_n12397, new_n3538, new_n12401);
nand_1 g12025(new_n12401, new_n12400, new_n12402);
nand_1 g12026(new_n12402, new_n12399, new_n12403);
nor_1  g12027(new_n1592, new_n2481, new_n12404);
nand_1 g12028(n9637, n3172, new_n12405);
nand_1 g12029(n5240, n3842, new_n12406);
xnor_1 g12030(new_n12406, new_n12405, new_n12407);
xnor_1 g12031(new_n12407, new_n12404, new_n12408);
nor_1  g12032(new_n3428, new_n3424, new_n12409);
nor_1  g12033(new_n12409, new_n3429, new_n12410);
xnor_1 g12034(new_n12410, new_n12408, new_n12411);
xnor_1 g12035(new_n12411, new_n12403, new_n12412);
xnor_1 g12036(new_n12412, new_n12396, new_n12413);
nand_1 g12037(n7236, n1357, new_n12414);
nand_1 g12038(new_n3435, new_n3434, new_n12415);
nand_1 g12039(new_n3441, new_n3436, new_n12416);
nand_1 g12040(new_n12416, new_n12415, new_n12417);
xnor_1 g12041(new_n12417, new_n12414, new_n12418);
xnor_1 g12042(new_n12418, new_n12413, new_n12419);
xnor_1 g12043(new_n12419, new_n12395, new_n12420);
nand_1 g12044(n1835, n1333, new_n12421);
nand_1 g12045(n11917, n11821, new_n12422);
xnor_1 g12046(new_n12422, new_n12421, new_n12423);
nand_1 g12047(n12753, n3602, new_n12424);
nand_1 g12048(n8595, n4187, new_n12425);
xnor_1 g12049(new_n12425, new_n12424, new_n12426);
nand_1 g12050(n6877, n4190, new_n12427);
nand_1 g12051(n10174, n3719, new_n12428);
xnor_1 g12052(new_n12428, new_n12427, new_n12429);
xnor_1 g12053(new_n12429, new_n12426, new_n12430);
xnor_1 g12054(new_n12430, new_n12423, new_n12431);
nand_1 g12055(new_n3932_1, new_n3931, new_n12432);
not_1  g12056(new_n12432, new_n12433);
nor_1  g12057(new_n3933, new_n3930, new_n12434);
nor_1  g12058(new_n12434, new_n12433, new_n12435);
nand_1 g12059(n9080, n4921, new_n12436);
xnor_1 g12060(new_n12436, new_n12435, new_n12437);
xnor_1 g12061(new_n12437, new_n12431, new_n12438);
nand_1 g12062(new_n3431, new_n3423, new_n12439);
nand_1 g12063(new_n3443, new_n12439, new_n12440);
xnor_1 g12064(new_n12440, new_n12438, new_n12441);
xnor_1 g12065(new_n12441, new_n12420, new_n12442);
nor_1  g12066(new_n4023, new_n3792, new_n12443);
not_1  g12067(new_n4025, new_n12444_1);
nor_1  g12068(new_n12444_1, new_n4019, new_n12445);
nor_1  g12069(new_n12445, new_n12443, new_n12446);
xnor_1 g12070(new_n12446, new_n12442, new_n12447);
xnor_1 g12071(new_n12447, new_n12392, new_n12448);
not_1  g12072(new_n3951, new_n12449);
nand_1 g12073(new_n3985, new_n12449, new_n12450);
nand_1 g12074(new_n3991, new_n3986_1, new_n12451);
nand_1 g12075(new_n12451, new_n12450, new_n12452);
xnor_1 g12076(new_n12452, new_n12448, new_n12453);
xnor_1 g12077(new_n12453, new_n12388, new_n12454);
not_1  g12078(new_n4032, new_n12455);
nor_1  g12079(new_n12455, new_n3992_1, new_n12456);
not_1  g12080(new_n4033, new_n12457);
nor_1  g12081(new_n4037, new_n12457, new_n12458);
nor_1  g12082(new_n12458, new_n12456, new_n12459);
and_1  g12083(new_n4026, new_n3805, new_n12460);
not_1  g12084(new_n4027, new_n12461);
nor_1  g12085(new_n4031, new_n12461, new_n12462);
nor_1  g12086(new_n12462, new_n12460, new_n12463);
nand_1 g12087(new_n3439, new_n3438, new_n12464);
not_1  g12088(new_n12464, new_n12465);
nor_1  g12089(new_n3440, new_n3437, new_n12466);
nor_1  g12090(new_n12466, new_n12465, new_n12467);
xnor_1 g12091(new_n12467, new_n12463, new_n12468);
xnor_1 g12092(new_n12468, new_n12459, new_n12469);
xnor_1 g12093(new_n12469, new_n12454, new_n12470);
xnor_1 g12094(new_n12470, new_n12296, new_n12471);
xnor_1 g12095(new_n12471, new_n12292, n5257);
xnor_1 g12096(new_n11723, new_n11707_1, n5411);
xnor_1 g12097(new_n3891, new_n3880, n5435);
xnor_1 g12098(new_n6507, new_n10281, n5641);
xnor_1 g12099(new_n9052, new_n9040, n5670);
xnor_1 g12100(new_n5299, new_n5264, n5693);
xnor_1 g12101(new_n1502, new_n1491, n5934);
xnor_1 g12102(new_n11726, new_n11725, n6089);
not_1  g12103(new_n8233, new_n12480);
and_1  g12104(new_n8234, new_n12480, new_n12481);
not_1  g12105(new_n12481, new_n12482);
not_1  g12106(new_n8213, new_n12483);
nand_1 g12107(new_n8217, new_n12483, new_n12484);
nand_1 g12108(new_n12484, new_n8211, new_n12485);
nor_1  g12109(new_n1377, new_n5550, new_n12486);
nor_1  g12110(new_n5516, new_n1367, new_n12487);
not_1  g12111(new_n12487, new_n12488);
nand_1 g12112(n6687, n3865, new_n12489_1);
nand_1 g12113(new_n12489_1, new_n12488, new_n12490);
not_1  g12114(new_n12489_1, new_n12491);
nand_1 g12115(new_n12491, new_n12487, new_n12492);
and_1  g12116(new_n12492, new_n12490, new_n12493);
xnor_1 g12117(new_n12493, new_n12486, new_n12494);
xnor_1 g12118(new_n12494, new_n12485, new_n12495);
nand_1 g12119(n6770, n4634, new_n12496);
xnor_1 g12120(new_n12496, new_n8207, new_n12497);
not_1  g12121(new_n12497, new_n12498);
nor_1  g12122(new_n6617, new_n1130, new_n12499);
nand_1 g12123(n10223, n9920, new_n12500);
nand_1 g12124(n7265, n4516, new_n12501);
xnor_1 g12125(new_n12501, new_n12500, new_n12502);
and_1  g12126(new_n12502, new_n12499, new_n12503);
nor_1  g12127(new_n12502, new_n12499, new_n12504);
nor_1  g12128(new_n12504, new_n12503, new_n12505);
xnor_1 g12129(new_n12505, new_n12498, new_n12506);
xnor_1 g12130(new_n12506, new_n12495, new_n12507);
not_1  g12131(new_n8226, new_n12508);
nand_1 g12132(new_n12508, new_n8218, new_n12509);
nand_1 g12133(new_n8232, new_n8227, new_n12510);
not_1  g12134(new_n12510, new_n12511_1);
nand_1 g12135(new_n12511_1, new_n8224, new_n12512);
nand_1 g12136(new_n12510, new_n8225, new_n12513);
nand_1 g12137(new_n12513, new_n12512, new_n12514);
nand_1 g12138(new_n12514, new_n12509, new_n12515);
xor_1  g12139(new_n12515, new_n12507, new_n12516);
xnor_1 g12140(new_n12516, new_n12482, new_n12517);
nor_1  g12141(new_n8235, new_n8202_1, new_n12518);
nor_1  g12142(new_n8236_1, new_n6022, new_n12519);
nor_1  g12143(new_n12519, new_n12518, new_n12520);
not_1  g12144(new_n12520, new_n12521);
xnor_1 g12145(new_n12521, new_n12517, new_n12522);
not_1  g12146(new_n12522, new_n12523);
nand_1 g12147(new_n8288, new_n8284, new_n12524);
nand_1 g12148(new_n8368, new_n12524, new_n12525);
not_1  g12149(new_n12525, new_n12526);
nand_1 g12150(new_n8281, new_n8244, new_n12527);
nand_1 g12151(new_n8282, new_n8243, new_n12528);
nand_1 g12152(new_n12528, new_n12527, new_n12529);
not_1  g12153(new_n8246, new_n12530);
nor_1  g12154(new_n8252, new_n12530, new_n12531);
not_1  g12155(new_n12531, new_n12532);
nand_1 g12156(new_n8257, new_n8253, new_n12533);
nand_1 g12157(new_n12533, new_n12532, new_n12534);
nand_1 g12158(n12221, n10928, new_n12535);
nand_1 g12159(n12145, n6986, new_n12536);
nand_1 g12160(n10217, n8336, new_n12537);
nand_1 g12161(new_n12537, new_n12536, new_n12538);
not_1  g12162(new_n12538, new_n12539);
nor_1  g12163(new_n12537, new_n12536, new_n12540);
nor_1  g12164(new_n12540, new_n12539, new_n12541);
xor_1  g12165(new_n12541, new_n12535, new_n12542);
xnor_1 g12166(new_n12542, new_n12534, new_n12543);
nand_1 g12167(n2522, n2226, new_n12544);
xnor_1 g12168(new_n12544, new_n8250, new_n12545);
nor_1  g12169(new_n6725, new_n1192, new_n12546);
not_1  g12170(new_n12546, new_n12547);
nand_1 g12171(n9189, n1094, new_n12548);
nand_1 g12172(n7946, n7320, new_n12549);
xnor_1 g12173(new_n12549, new_n12548, new_n12550);
xnor_1 g12174(new_n12550, new_n12547, new_n12551);
xor_1  g12175(new_n12551, new_n12545, new_n12552);
xnor_1 g12176(new_n12552, new_n12543, new_n12553);
not_1  g12177(new_n12553, new_n12554);
not_1  g12178(new_n8258, new_n12555);
nand_1 g12179(new_n8267, new_n12555, new_n12556);
nand_1 g12180(new_n8273, new_n8268, new_n12557);
not_1  g12181(new_n12557, new_n12558);
nand_1 g12182(new_n12558, new_n8264, new_n12559);
nand_1 g12183(new_n12557, new_n8265, new_n12560);
nand_1 g12184(new_n12560, new_n12559, new_n12561);
nand_1 g12185(new_n12561, new_n12556, new_n12562);
xnor_1 g12186(new_n12562, new_n12554, new_n12563);
xnor_1 g12187(new_n12563, new_n8278, new_n12564);
xnor_1 g12188(new_n12564, new_n12529, new_n12565);
not_1  g12189(new_n8323, new_n12566);
nand_1 g12190(new_n12566, new_n8319, new_n12567);
nor_1  g12191(new_n8302, new_n8301, new_n12568);
nor_1  g12192(new_n1538, new_n1310, new_n12569);
not_1  g12193(new_n12569, new_n12570);
xnor_1 g12194(new_n12570, new_n12568, new_n12571);
nor_1  g12195(new_n6823, new_n1235, new_n12572);
not_1  g12196(new_n12572, new_n12573);
nand_1 g12197(n2558, n1199, new_n12574);
nand_1 g12198(n5579, n4828, new_n12575);
nand_1 g12199(new_n12575, new_n12574, new_n12576);
not_1  g12200(new_n12574, new_n12577);
not_1  g12201(new_n12575, new_n12578);
nand_1 g12202(new_n12578, new_n12577, new_n12579);
nand_1 g12203(new_n12579, new_n12576, new_n12580);
xnor_1 g12204(new_n12580, new_n12573, new_n12581);
xnor_1 g12205(new_n12581, new_n12571, new_n12582);
not_1  g12206(new_n8299, new_n12583);
not_1  g12207(new_n8303_1, new_n12584);
nand_1 g12208(new_n12584, new_n8300, new_n12585);
nand_1 g12209(new_n12585, new_n12583, new_n12586);
nor_1  g12210(new_n1452, new_n5727, new_n12587);
nand_1 g12211(n7891, n6016, new_n12588);
nand_1 g12212(n12069, n2347, new_n12589);
xnor_1 g12213(new_n12589, new_n12588, new_n12590);
xor_1  g12214(new_n12590, new_n12587, new_n12591_1);
xnor_1 g12215(new_n12591_1, new_n12586, new_n12592);
xnor_1 g12216(new_n12592, new_n12582, new_n12593);
not_1  g12217(new_n8312, new_n12594);
nand_1 g12218(new_n12594, new_n8304, new_n12595);
nand_1 g12219(new_n8317, new_n8310, new_n12596);
nand_1 g12220(new_n8316, new_n8311, new_n12597);
nand_1 g12221(new_n12597, new_n12596, new_n12598);
nand_1 g12222(new_n12598, new_n12595, new_n12599);
xnor_1 g12223(new_n12599, new_n12593, new_n12600);
xnor_1 g12224(new_n12600, new_n12567, new_n12601);
nand_1 g12225(new_n8324, new_n8291, new_n12602);
not_1  g12226(new_n8290, new_n12603);
nand_1 g12227(new_n8325, new_n12603, new_n12604);
nand_1 g12228(new_n12604, new_n12602, new_n12605);
xnor_1 g12229(new_n12605, new_n12601, new_n12606);
nand_1 g12230(new_n8353, new_n8352, new_n12607);
not_1  g12231(new_n8328, new_n12608);
nor_1  g12232(new_n8331, new_n12608, new_n12609);
not_1  g12233(new_n12609, new_n12610);
nand_1 g12234(new_n8336_1, new_n12610, new_n12611);
nor_1  g12235(new_n1467, new_n5924, new_n12612);
nand_1 g12236(n7270, n5314, new_n12613);
nand_1 g12237(n11222, n2507, new_n12614);
xnor_1 g12238(new_n12614, new_n12613, new_n12615);
and_1  g12239(new_n12615, new_n12612, new_n12616);
nor_1  g12240(new_n12615, new_n12612, new_n12617);
nor_1  g12241(new_n12617, new_n12616, new_n12618);
xnor_1 g12242(new_n12618, new_n12611, new_n12619);
nor_1  g12243(new_n8330, new_n8329, new_n12620);
nor_1  g12244(new_n4542, new_n1325, new_n12621);
xnor_1 g12245(new_n12621, new_n12620, new_n12622);
not_1  g12246(new_n12622, new_n12623);
nor_1  g12247(new_n1215, new_n6935, new_n12624);
nand_1 g12248(n5767, n3342, new_n12625);
nand_1 g12249(n9763, n9457, new_n12626);
xnor_1 g12250(new_n12626, new_n12625, new_n12627);
xnor_1 g12251(new_n12627, new_n12624, new_n12628);
xnor_1 g12252(new_n12628, new_n12623, new_n12629);
xnor_1 g12253(new_n12629, new_n12619, new_n12630);
not_1  g12254(new_n12630, new_n12631);
not_1  g12255(new_n8345, new_n12632);
nand_1 g12256(new_n12632, new_n8339, new_n12633);
nand_1 g12257(new_n8350, new_n8346, new_n12634);
not_1  g12258(new_n12634, new_n12635);
nand_1 g12259(new_n12635, new_n8343, new_n12636);
nand_1 g12260(new_n12634, new_n8344, new_n12637);
nand_1 g12261(new_n12637, new_n12636, new_n12638);
nand_1 g12262(new_n12638, new_n12633, new_n12639);
xnor_1 g12263(new_n12639, new_n12631, new_n12640);
xnor_1 g12264(new_n12640, new_n12607, new_n12641);
not_1  g12265(new_n8327, new_n12642);
nand_1 g12266(new_n8354, new_n12642, new_n12643);
nand_1 g12267(new_n8355, new_n6240, new_n12644);
nand_1 g12268(new_n12644, new_n12643, new_n12645);
xnor_1 g12269(new_n12645, new_n12641, new_n12646);
xnor_1 g12270(new_n12646, new_n12606, new_n12647);
not_1  g12271(new_n8356, new_n12648_1);
nand_1 g12272(new_n12648_1, new_n8326, new_n12649);
nand_1 g12273(new_n8362, new_n12649, new_n12650);
xnor_1 g12274(new_n12650, new_n12647, new_n12651);
xnor_1 g12275(new_n12651, new_n12565, new_n12652);
xnor_1 g12276(new_n12652, new_n12526, new_n12653);
nand_1 g12277(new_n12653, new_n12523, new_n12654);
nor_1  g12278(new_n8241, new_n8237, new_n12655);
nor_1  g12279(new_n8371, new_n12655, new_n12656);
xnor_1 g12280(new_n12653, new_n12522, new_n12657);
nand_1 g12281(new_n12657, new_n12656, new_n12658);
nand_1 g12282(new_n12658, new_n12654, new_n12659);
not_1  g12283(new_n12565, new_n12660);
not_1  g12284(new_n12651, new_n12661);
nor_1  g12285(new_n12661, new_n12660, new_n12662);
nor_1  g12286(new_n12652, new_n12525, new_n12663);
nor_1  g12287(new_n12663, new_n12662, new_n12664);
not_1  g12288(new_n12646, new_n12665);
nand_1 g12289(new_n12665, new_n12606, new_n12666);
not_1  g12290(new_n12650, new_n12667);
nand_1 g12291(new_n12667, new_n12647, new_n12668);
nand_1 g12292(new_n12668, new_n12666, new_n12669);
nand_1 g12293(new_n12562, new_n12553, new_n12670);
nand_1 g12294(new_n12670, new_n12559, new_n12671);
not_1  g12295(new_n12485, new_n12672);
nand_1 g12296(new_n12494, new_n12672, new_n12673);
nand_1 g12297(new_n12506, new_n12495, new_n12674);
nand_1 g12298(new_n12674, new_n12673, new_n12675);
nor_1  g12299(new_n1278, new_n8138_1, new_n12676);
nand_1 g12300(new_n12614, new_n12613, new_n12677);
not_1  g12301(new_n12677, new_n12678);
nor_1  g12302(new_n12617, new_n12678, new_n12679);
xnor_1 g12303(new_n12679, new_n12676, new_n12680);
xnor_1 g12304(new_n12680, new_n12675, new_n12681);
xnor_1 g12305(new_n12681, new_n12671, new_n12682);
not_1  g12306(new_n12534, new_n12683);
nand_1 g12307(new_n12542, new_n12683, new_n12684);
nand_1 g12308(new_n12552, new_n12543, new_n12685);
nand_1 g12309(new_n12685, new_n12684, new_n12686);
nor_1  g12310(new_n6725, new_n1199_1, new_n12687);
xnor_1 g12311(new_n12687, new_n12686, new_n12688);
nand_1 g12312(new_n12549, new_n12548, new_n12689);
not_1  g12313(new_n12689, new_n12690);
nor_1  g12314(new_n12550, new_n12546, new_n12691);
nor_1  g12315(new_n12691, new_n12690, new_n12692);
nor_1  g12316(new_n1196, new_n9946, new_n12693);
nand_1 g12317(n10223, n3627, new_n12694);
nand_1 g12318(n3865, n2564, new_n12695);
xnor_1 g12319(new_n12695, new_n12694, new_n12696);
xnor_1 g12320(new_n12696, new_n12693, new_n12697);
xnor_1 g12321(new_n12697, new_n12692, new_n12698);
nand_1 g12322(n12221, n6986, new_n12699);
nand_1 g12323(n8336, n7823, new_n12700);
xnor_1 g12324(new_n12700, new_n12699, new_n12701);
xnor_1 g12325(new_n12701, new_n12698, new_n12702);
nand_1 g12326(new_n12501, new_n12500, new_n12703);
not_1  g12327(new_n12703, new_n12704_1);
nor_1  g12328(new_n12504, new_n12704_1, new_n12705_1);
nand_1 g12329(new_n12544, new_n8251, new_n12706_1);
nand_1 g12330(new_n12551, new_n12545, new_n12707);
nand_1 g12331(new_n12707, new_n12706_1, new_n12708);
xnor_1 g12332(new_n12708, new_n12705_1, new_n12709_1);
nand_1 g12333(new_n12589, new_n12588, new_n12710);
not_1  g12334(new_n12710, new_n12711);
nor_1  g12335(new_n12590, new_n12587, new_n12712);
nor_1  g12336(new_n12712, new_n12711, new_n12713);
and_1  g12337(n6687, n2512, new_n12714);
nand_1 g12338(new_n12576, new_n12572, new_n12715);
nand_1 g12339(new_n12715, new_n12579, new_n12716);
xnor_1 g12340(new_n12716, new_n12714, new_n12717);
xnor_1 g12341(new_n12717, new_n12713, new_n12718);
xnor_1 g12342(new_n12718, new_n12709_1, new_n12719);
xnor_1 g12343(new_n12719, new_n12702, new_n12720_1);
nand_1 g12344(n11153, n2507, new_n12721);
nand_1 g12345(n7270, n996, new_n12722);
xnor_1 g12346(new_n12722, new_n12721, new_n12723);
nand_1 g12347(n7160, n6016, new_n12724);
nand_1 g12348(n5767, n806, new_n12725);
xnor_1 g12349(new_n12725, new_n12724, new_n12726);
xnor_1 g12350(new_n12726, new_n12723, new_n12727);
nand_1 g12351(n4828, n521, new_n12728);
nand_1 g12352(n5579, n2515, new_n12729);
xnor_1 g12353(new_n12729, new_n12728, new_n12730);
nand_1 g12354(n12069, n1576, new_n12731);
nand_1 g12355(n5314, n5153, new_n12732);
xnor_1 g12356(new_n12732, new_n12731, new_n12733);
xnor_1 g12357(new_n12733, new_n12730, new_n12734);
xnor_1 g12358(new_n12734, new_n12727, new_n12735);
nand_1 g12359(new_n12490, new_n12486, new_n12736);
nand_1 g12360(new_n12736, new_n12492, new_n12737);
nand_1 g12361(n4516, n2879, new_n12738);
nand_1 g12362(n4189, n2253, new_n12739);
nand_1 g12363(n9920, n4634, new_n12740);
xnor_1 g12364(new_n12740, new_n12739, new_n12741);
xnor_1 g12365(new_n12741, new_n12738, new_n12742);
xnor_1 g12366(new_n12742, new_n12737, new_n12743);
xnor_1 g12367(new_n12743, new_n12735, new_n12744);
nand_1 g12368(new_n12496, new_n8208, new_n12745);
nand_1 g12369(new_n12505, new_n12497, new_n12746);
nand_1 g12370(new_n12746, new_n12745, new_n12747);
nand_1 g12371(new_n12621, new_n12620, new_n12748);
nand_1 g12372(new_n12628, new_n12623, new_n12749);
nand_1 g12373(new_n12749, new_n12748, new_n12750);
xnor_1 g12374(new_n12750, new_n12747, new_n12751);
xnor_1 g12375(new_n12751, new_n12744, new_n12752);
xnor_1 g12376(new_n12752, new_n12720_1, new_n12753_1);
xnor_1 g12377(new_n12753_1, new_n12688, new_n12754);
xnor_1 g12378(new_n12754, new_n12682, new_n12755);
nand_1 g12379(new_n12639, new_n12630, new_n12756);
nand_1 g12380(new_n12756, new_n12636, new_n12757);
nand_1 g12381(n12145, n2226, new_n12758);
nor_1  g12382(new_n12539, new_n12535, new_n12759);
nor_1  g12383(new_n12759, new_n12540, new_n12760);
nand_1 g12384(n9195, n6770, new_n12761);
nand_1 g12385(n11222, n6431, new_n12762);
xnor_1 g12386(new_n12762, new_n12761, new_n12763);
nand_1 g12387(n10928, n10217, new_n12764);
nand_1 g12388(n7320, n2024, new_n12765);
xnor_1 g12389(new_n12765, new_n12764, new_n12766);
xnor_1 g12390(new_n12766, new_n12763, new_n12767);
nand_1 g12391(n5319, n3342, new_n12768);
nand_1 g12392(n9457, n9111, new_n12769);
nand_1 g12393(n9763, n4817, new_n12770);
xnor_1 g12394(new_n12770, new_n12769, new_n12771);
xnor_1 g12395(new_n12771, new_n12768, new_n12772);
xnor_1 g12396(new_n12772, new_n12767, new_n12773);
xnor_1 g12397(new_n12773, new_n12760, new_n12774);
xnor_1 g12398(new_n12774, new_n12758, new_n12775);
xnor_1 g12399(new_n12775, new_n12757, new_n12776);
xnor_1 g12400(new_n12776, new_n12755, new_n12777_1);
nand_1 g12401(new_n12563, new_n8279, new_n12778);
nand_1 g12402(new_n12564, new_n12529, new_n12779);
nand_1 g12403(new_n12779, new_n12778, new_n12780);
not_1  g12404(new_n12593, new_n12781);
nand_1 g12405(new_n12599, new_n12781, new_n12782);
nand_1 g12406(new_n12782, new_n12596, new_n12783);
nand_1 g12407(new_n12515, new_n12507, new_n12784);
nand_1 g12408(new_n12784, new_n12512, new_n12785);
not_1  g12409(new_n12611, new_n12786);
nand_1 g12410(new_n12618, new_n12786, new_n12787);
nand_1 g12411(new_n12629, new_n12619, new_n12788);
nand_1 g12412(new_n12788, new_n12787, new_n12789);
nand_1 g12413(new_n12569, new_n12568, new_n12790);
not_1  g12414(new_n12581, new_n12791);
nand_1 g12415(new_n12791, new_n12571, new_n12792);
nand_1 g12416(new_n12792, new_n12790, new_n12793);
nand_1 g12417(n7891, n5798, new_n12794);
xnor_1 g12418(new_n12794, new_n12793, new_n12795);
nand_1 g12419(n12391, n2347, new_n12796);
nand_1 g12420(n7265, n2087, new_n12797);
xnor_1 g12421(new_n12797, new_n12796, new_n12798);
xnor_1 g12422(new_n12798, new_n12795, new_n12799);
xnor_1 g12423(new_n12799, new_n12789, new_n12800);
nand_1 g12424(n2498, n1199, new_n12801);
nand_1 g12425(n6578, n2558, new_n12802);
xnor_1 g12426(new_n12802, new_n12801, new_n12803);
xnor_1 g12427(new_n12803, new_n12800, new_n12804);
xnor_1 g12428(new_n12804, new_n12785, new_n12805);
xnor_1 g12429(new_n12805, new_n12783, new_n12806);
xnor_1 g12430(new_n12806, new_n12780, new_n12807_1);
xnor_1 g12431(new_n12807_1, new_n12777_1, new_n12808);
not_1  g12432(new_n12640, new_n12809);
nor_1  g12433(new_n12809, new_n12607, new_n12810);
not_1  g12434(new_n12641, new_n12811);
nor_1  g12435(new_n12645, new_n12811, new_n12812);
nor_1  g12436(new_n12812, new_n12810, new_n12813);
nand_1 g12437(new_n12626, new_n12625, new_n12814);
not_1  g12438(new_n12814, new_n12815);
nor_1  g12439(new_n12627, new_n12624, new_n12816);
nor_1  g12440(new_n12816, new_n12815, new_n12817);
not_1  g12441(new_n12586, new_n12818);
nand_1 g12442(new_n12591_1, new_n12818, new_n12819);
not_1  g12443(new_n12582, new_n12820);
nand_1 g12444(new_n12592, new_n12820, new_n12821);
nand_1 g12445(new_n12821, new_n12819, new_n12822);
xnor_1 g12446(new_n12822, new_n12817, new_n12823);
xnor_1 g12447(new_n12823, new_n12813, new_n12824);
xnor_1 g12448(new_n12824, new_n12808, new_n12825);
xnor_1 g12449(new_n12825, new_n12669, new_n12826_1);
nand_1 g12450(new_n12516, new_n12481, new_n12827);
nand_1 g12451(new_n12520, new_n12517, new_n12828);
nand_1 g12452(new_n12828, new_n12827, new_n12829);
not_1  g12453(new_n12567, new_n12830);
nand_1 g12454(new_n12600, new_n12830, new_n12831);
nand_1 g12455(new_n12605, new_n12601, new_n12832);
nand_1 g12456(new_n12832, new_n12831, new_n12833);
xnor_1 g12457(new_n12833, new_n12829, new_n12834);
xnor_1 g12458(new_n12834, new_n12826_1, new_n12835);
xnor_1 g12459(new_n12835, new_n12664, new_n12836);
xnor_1 g12460(new_n12836, new_n12659, n6192);
xor_1  g12461(new_n996_1, new_n964, n6273);
not_1  g12462(new_n8003, new_n12839);
nand_1 g12463(new_n8002, new_n8001, new_n12840);
nand_1 g12464(new_n12840, new_n12839, n6445);
xnor_1 g12465(new_n9910, new_n9909, n6645);
xnor_1 g12466(new_n8410, new_n8409, n6689);
xor_1  g12467(new_n1492, new_n1396, n6742);
not_1  g12468(new_n2239, new_n12845);
xnor_1 g12469(new_n2278_1, new_n12845, n6809);
xnor_1 g12470(new_n7247, new_n7245, n6822);
xnor_1 g12471(new_n11719, new_n11716, n6860);
xnor_1 g12472(new_n9905, new_n9898, n7193);
not_1  g12473(new_n8004, new_n12850);
xnor_1 g12474(new_n8006, new_n12850, n7568);
xnor_1 g12475(new_n1500, new_n1499, n7676);
not_1  g12476(new_n550, new_n12853);
nand_1 g12477(new_n1001, new_n12853, new_n12854);
nand_1 g12478(new_n1119, new_n1002, new_n12855);
nand_1 g12479(new_n12855, new_n12854, new_n12856);
nor_1  g12480(new_n1112, new_n1034, new_n12857);
nor_1  g12481(new_n1118, new_n1113, new_n12858);
nor_1  g12482(new_n12858, new_n12857, new_n12859);
not_1  g12483(new_n1071, new_n12860);
nor_1  g12484(new_n1107, new_n12860, new_n12861);
not_1  g12485(new_n1108, new_n12862);
nor_1  g12486(new_n1111, new_n12862, new_n12863);
nor_1  g12487(new_n12863, new_n12861, new_n12864);
nor_1  g12488(new_n2723, new_n557, new_n12865);
nand_1 g12489(new_n1098, new_n1073, new_n12866);
not_1  g12490(new_n1099, new_n12867);
nand_1 g12491(new_n1106, new_n12867, new_n12868);
nand_1 g12492(new_n12868, new_n12866, new_n12869);
nor_1  g12493(new_n1094_1, new_n941, new_n12870);
nor_1  g12494(new_n1096, new_n1091, new_n12871);
nor_1  g12495(new_n12871, new_n12870, new_n12872);
nand_1 g12496(new_n519, new_n506, new_n12873);
nor_1  g12497(new_n509, new_n403, new_n12874);
not_1  g12498(new_n510, new_n12875);
nor_1  g12499(new_n516, new_n12875, new_n12876);
nor_1  g12500(new_n12876, new_n12874, new_n12877);
nor_1  g12501(new_n8505, new_n420, new_n12878);
nand_1 g12502(new_n499, new_n493, new_n12879);
nand_1 g12503(new_n12879, new_n500, new_n12880);
xnor_1 g12504(new_n12880, new_n12878, new_n12881);
nand_1 g12505(n3986, n1980, new_n12882);
nand_1 g12506(n10848, n5857, new_n12883);
xnor_1 g12507(new_n12883, new_n12882, new_n12884);
nand_1 g12508(n11257, n2509, new_n12885);
nand_1 g12509(n4005, n1097, new_n12886);
xnor_1 g12510(new_n12886, new_n12885, new_n12887);
xnor_1 g12511(new_n12887, new_n12884, new_n12888);
xnor_1 g12512(new_n12888, new_n12881, new_n12889);
xnor_1 g12513(new_n12889, new_n12877, new_n12890);
and_1  g12514(n8028, n45, new_n12891);
nand_1 g12515(new_n1008, new_n1007, new_n12892);
not_1  g12516(new_n12892, new_n12893);
nor_1  g12517(new_n1009, new_n1006, new_n12894);
nor_1  g12518(new_n12894, new_n12893, new_n12895);
xnor_1 g12519(new_n12895, new_n12891, new_n12896);
nor_1  g12520(new_n1017, new_n1016, new_n12897);
nand_1 g12521(new_n1017, new_n1016, new_n12898);
not_1  g12522(new_n12898, new_n12899);
nor_1  g12523(new_n12899, new_n1015, new_n12900);
nor_1  g12524(new_n12900, new_n12897, new_n12901);
xnor_1 g12525(new_n12901, new_n12896, new_n12902);
nand_1 g12526(n4312, n2585, new_n12903);
nand_1 g12527(new_n514, new_n513, new_n12904);
not_1  g12528(new_n12904, new_n12905);
nor_1  g12529(new_n515, new_n512, new_n12906);
nor_1  g12530(new_n12906, new_n12905, new_n12907);
nand_1 g12531(n10644, n7354, new_n12908);
nand_1 g12532(n12706, n5964, new_n12909);
nand_1 g12533(n12720, n12025, new_n12910);
xnor_1 g12534(new_n12910, new_n12909, new_n12911);
xnor_1 g12535(new_n12911, new_n12908, new_n12912);
xnor_1 g12536(new_n12912, new_n12907, new_n12913);
xnor_1 g12537(new_n12913, new_n12903, new_n12914);
xnor_1 g12538(new_n12914, new_n12902, new_n12915);
xnor_1 g12539(new_n12915, new_n12890, new_n12916);
xnor_1 g12540(new_n12916, new_n12873, new_n12917);
nand_1 g12541(n7436, n4141, new_n12918);
nand_1 g12542(new_n1013, new_n1012, new_n12919);
not_1  g12543(new_n1019, new_n12920);
nand_1 g12544(new_n12920, new_n1014, new_n12921);
nand_1 g12545(new_n12921, new_n12919, new_n12922);
xnor_1 g12546(new_n12922, new_n12918, new_n12923);
xnor_1 g12547(new_n12923, new_n12917, new_n12924);
xnor_1 g12548(new_n12924, new_n12872, new_n12925_1);
xnor_1 g12549(new_n12925_1, new_n12869, new_n12926);
xnor_1 g12550(new_n12926, new_n12865, new_n12927);
xnor_1 g12551(new_n12927, new_n12864, new_n12928);
nor_1  g12552(new_n3327, new_n377, new_n12929);
nand_1 g12553(new_n1041, new_n1040, new_n12930);
not_1  g12554(new_n12930, new_n12931);
nor_1  g12555(new_n1042, new_n1039, new_n12932);
nor_1  g12556(new_n12932, new_n12931, new_n12933);
xnor_1 g12557(new_n12933, new_n12929, new_n12934);
nand_1 g12558(new_n1051, new_n1050, new_n12935);
not_1  g12559(new_n12935, new_n12936);
nor_1  g12560(new_n1052, new_n1049, new_n12937);
nor_1  g12561(new_n12937, new_n12936, new_n12938);
nor_1  g12562(new_n2190, new_n712, new_n12939);
nand_1 g12563(n11892, n5814, new_n12940);
nand_1 g12564(n3616, n1512, new_n12941);
xnor_1 g12565(new_n12941, new_n12940, new_n12942);
xnor_1 g12566(new_n12942, new_n12939, new_n12943);
xnor_1 g12567(new_n12943, new_n12938, new_n12944);
xnor_1 g12568(new_n12944, new_n12934, new_n12945);
nand_1 g12569(n12299, n4928, new_n12946);
nand_1 g12570(new_n1087, new_n1086, new_n12947_1);
not_1  g12571(new_n12947_1, new_n12948);
nor_1  g12572(new_n1088, new_n1085, new_n12949);
nor_1  g12573(new_n12949, new_n12948, new_n12950);
xnor_1 g12574(new_n12950, new_n12946, new_n12951);
nand_1 g12575(n5069, n2530, new_n12952);
nand_1 g12576(n10545, n2802, new_n12953);
xnor_1 g12577(new_n12953, new_n12952, new_n12954);
xnor_1 g12578(new_n12954, new_n12951, new_n12955);
xnor_1 g12579(new_n12955, new_n12945, new_n12956);
nand_1 g12580(new_n1043, new_n1037, new_n12957);
nand_1 g12581(new_n1058, new_n1044, new_n12958);
nand_1 g12582(new_n12958, new_n12957, new_n12959);
nor_1  g12583(new_n1082, new_n923, new_n12960);
not_1  g12584(new_n1083, new_n12961);
nor_1  g12585(new_n1089, new_n12961, new_n12962);
nor_1  g12586(new_n12962, new_n12960, new_n12963);
nand_1 g12587(new_n1046, new_n1045, new_n12964);
nand_1 g12588(new_n1057, new_n12964, new_n12965);
nand_1 g12589(n7690, n533, new_n12966);
xnor_1 g12590(new_n12966, new_n12965, new_n12967);
xnor_1 g12591(new_n12967, new_n12963, new_n12968);
xnor_1 g12592(new_n12968, new_n12959, new_n12969);
xnor_1 g12593(new_n12969, new_n12956, new_n12970);
nand_1 g12594(n12704, n2393, new_n12971);
nor_1  g12595(new_n753_1, new_n802, new_n12972);
xnor_1 g12596(new_n12972, new_n12971, new_n12973);
nand_1 g12597(n12648, n6806, new_n12974);
nand_1 g12598(n4499, n1564, new_n12975);
xnor_1 g12599(new_n12975, new_n12974, new_n12976);
xnor_1 g12600(new_n12976, new_n12973, new_n12977);
nand_1 g12601(new_n1078, new_n1077, new_n12978);
not_1  g12602(new_n12978, new_n12979);
nor_1  g12603(new_n1079, new_n1076, new_n12980);
nor_1  g12604(new_n12980, new_n12979, new_n12981);
nand_1 g12605(n5694, n5331, new_n12982);
nand_1 g12606(n7388, n4903, new_n12983);
xnor_1 g12607(new_n12983, new_n12982, new_n12984);
xnor_1 g12608(new_n12984, new_n12981, new_n12985);
xnor_1 g12609(new_n12985, new_n12977, new_n12986);
nand_1 g12610(n8276, n5105, new_n12987);
nand_1 g12611(n5305, n615, new_n12988);
xnor_1 g12612(new_n12988, new_n12987, new_n12989);
xnor_1 g12613(new_n12989, new_n12986, new_n12990);
xnor_1 g12614(new_n12990, new_n12970, new_n12991);
not_1  g12615(new_n1022, new_n12992);
nand_1 g12616(new_n1028, new_n12992, new_n12993);
nand_1 g12617(new_n12993, new_n1025, new_n12994);
not_1  g12618(new_n1060, new_n12995);
nand_1 g12619(new_n1066, new_n12995, new_n12996);
nand_1 g12620(new_n12996, new_n1063, new_n12997);
xnor_1 g12621(new_n12997, new_n12994, new_n12998);
xnor_1 g12622(new_n12998, new_n12991, new_n12999);
nand_1 g12623(n8759, n783, new_n13000);
nand_1 g12624(n10510, n7500, new_n13001);
xnor_1 g12625(new_n13001, new_n13000, new_n13002);
nand_1 g12626(new_n528, new_n521_1, new_n13003);
nand_1 g12627(new_n13003, new_n525, new_n13004);
not_1  g12628(new_n1075, new_n13005);
nand_1 g12629(new_n1080, new_n13005, new_n13006);
not_1  g12630(new_n1090, new_n13007);
nand_1 g12631(new_n13007, new_n1081, new_n13008);
nand_1 g12632(new_n13008, new_n13006, new_n13009);
xnor_1 g12633(new_n13009, new_n13004, new_n13010);
xnor_1 g12634(new_n13010, new_n13002, new_n13011);
xnor_1 g12635(new_n13011, new_n12999, new_n13012);
not_1  g12636(new_n1035, new_n13013);
nand_1 g12637(new_n1067_1, new_n13013, new_n13014);
nand_1 g12638(new_n1070, new_n1068, new_n13015);
nand_1 g12639(new_n13015, new_n13014, new_n13016);
nand_1 g12640(n7965, n1906, new_n13017);
xnor_1 g12641(new_n13017, new_n13016, new_n13018);
xnor_1 g12642(new_n13018, new_n13012, new_n13019);
nand_1 g12643(new_n529, new_n487, new_n13020);
nand_1 g12644(new_n549, new_n530, new_n13021);
nand_1 g12645(new_n13021, new_n13020, new_n13022);
nand_1 g12646(new_n1029, new_n655, new_n13023);
nand_1 g12647(new_n1033, new_n1030, new_n13024);
nand_1 g12648(new_n13024, new_n13023, new_n13025);
nand_1 g12649(new_n1010, new_n1005, new_n13026);
not_1  g12650(new_n1011, new_n13027);
nand_1 g12651(new_n1021, new_n13027, new_n13028);
nand_1 g12652(new_n13028, new_n13026, new_n13029);
nand_1 g12653(n8236, n6776, new_n13030);
xor_1  g12654(new_n13030, new_n13029, new_n13031);
xnor_1 g12655(new_n13031, new_n13025, new_n13032);
xnor_1 g12656(new_n13032, new_n13022, new_n13033);
xnor_1 g12657(new_n13033, new_n13019, new_n13034);
xnor_1 g12658(new_n13034, new_n12928, new_n13035);
xnor_1 g12659(new_n13035, new_n12859, new_n13036);
xnor_1 g12660(new_n13036, new_n12856, n7966);
xnor_1 g12661(new_n12657, new_n12656, n7981);
not_1  g12662(new_n12024, new_n13039);
nand_1 g12663(new_n12275, new_n13039, new_n13040);
nand_1 g12664(new_n12287, new_n12276, new_n13041);
nand_1 g12665(new_n13041, new_n13040, new_n13042);
not_1  g12666(new_n12190, new_n13043);
nand_1 g12667(new_n13043, new_n12096, new_n13044);
nand_1 g12668(new_n12274, new_n12191, new_n13045);
nand_1 g12669(new_n13045, new_n13044, new_n13046);
nand_1 g12670(new_n12268, new_n12220, new_n13047);
not_1  g12671(new_n12218, new_n13048);
xnor_1 g12672(new_n12219, new_n13048, new_n13049);
xnor_1 g12673(new_n12268, new_n13049, new_n13050);
nand_1 g12674(new_n12273, new_n13050, new_n13051);
nand_1 g12675(new_n13051, new_n13047, new_n13052);
not_1  g12676(new_n12222, new_n13053);
nand_1 g12677(new_n12263, new_n13053, new_n13054);
not_1  g12678(new_n12267, new_n13055);
nand_1 g12679(new_n13055, new_n12264, new_n13056);
nand_1 g12680(new_n13056, new_n13054, new_n13057);
not_1  g12681(new_n12004, new_n13058);
nand_1 g12682(new_n12010, new_n13058, new_n13059);
nand_1 g12683(new_n13059, new_n12007, new_n13060);
nor_1  g12684(new_n12246, new_n12245, new_n13061);
nand_1 g12685(new_n12246, new_n12245, new_n13062);
not_1  g12686(new_n13062, new_n13063);
nor_1  g12687(new_n13063, new_n12244, new_n13064);
nor_1  g12688(new_n13064, new_n13061, new_n13065);
nand_1 g12689(n8717, n6986, new_n13066);
nand_1 g12690(n11222, n10022, new_n13067);
nand_1 g12691(n12391, n1353, new_n13068);
xnor_1 g12692(new_n13068, new_n13067, new_n13069);
xnor_1 g12693(new_n13069, new_n13066, new_n13070);
xnor_1 g12694(new_n13070, new_n13065, new_n13071);
xnor_1 g12695(new_n13071, new_n13060, new_n13072);
xnor_1 g12696(new_n13072, new_n13057, new_n13073);
xnor_1 g12697(new_n13073, new_n13052, new_n13074);
nand_1 g12698(new_n12262, new_n12253, new_n13075);
nand_1 g12699(new_n13075, new_n12259, new_n13076);
nand_1 g12700(new_n12251, new_n12238, new_n13077);
nand_1 g12701(n12069, n4436, new_n13078);
nand_1 g12702(n11999, n11153, new_n13079);
xnor_1 g12703(new_n13079, new_n13078, new_n13080);
nand_1 g12704(n7159, n1199, new_n13081);
nand_1 g12705(n11967, n7160, new_n13082);
xnor_1 g12706(new_n13082, new_n13081, new_n13083);
xnor_1 g12707(new_n13083, new_n13080, new_n13084);
nand_1 g12708(new_n12231, new_n12226, new_n13085);
nand_1 g12709(new_n13085, new_n12232, new_n13086);
nand_1 g12710(n6254, n4828, new_n13087);
nor_1  g12711(new_n1368, new_n10073, new_n13088);
xnor_1 g12712(new_n13088, new_n13087, new_n13089);
xnor_1 g12713(new_n13089, new_n13086, new_n13090);
xnor_1 g12714(new_n13090, new_n13084, new_n13091);
xnor_1 g12715(new_n13091, new_n13077, new_n13092);
xnor_1 g12716(new_n13092, new_n13076, new_n13093);
not_1  g12717(new_n12194, new_n13094);
nand_1 g12718(new_n12199, new_n13094, new_n13095);
not_1  g12719(new_n12210, new_n13096);
nand_1 g12720(new_n13096, new_n12200, new_n13097);
nand_1 g12721(new_n13097, new_n13095, new_n13098);
nand_1 g12722(n12489, n6578, new_n13099);
nand_1 g12723(n12947, n996, new_n13100);
nand_1 g12724(n9457, n5760, new_n13101);
xnor_1 g12725(new_n13101, new_n13100, new_n13102);
xnor_1 g12726(new_n13102, new_n13099, new_n13103);
xnor_1 g12727(new_n13103, new_n13098, new_n13104);
nand_1 g12728(new_n12242, new_n12241, new_n13105);
not_1  g12729(new_n12248, new_n13106);
nand_1 g12730(new_n13106, new_n12243, new_n13107);
nand_1 g12731(new_n13107, new_n13105, new_n13108);
nand_1 g12732(n7891, n447, new_n13109);
xnor_1 g12733(new_n13109, new_n13108, new_n13110);
nor_1  g12734(new_n8843, new_n6823, new_n13111);
nand_1 g12735(new_n12206, new_n12205, new_n13112);
not_1  g12736(new_n13112, new_n13113);
nor_1  g12737(new_n12207, new_n12204, new_n13114);
nor_1  g12738(new_n13114, new_n13113, new_n13115);
nand_1 g12739(new_n12197, new_n12196, new_n13116);
not_1  g12740(new_n13116, new_n13117);
nor_1  g12741(new_n12198, new_n12195, new_n13118);
nor_1  g12742(new_n13118, new_n13117, new_n13119);
xnor_1 g12743(new_n13119, new_n13115, new_n13120);
xnor_1 g12744(new_n13120, new_n13111, new_n13121);
xnor_1 g12745(new_n13121, new_n13110, new_n13122);
nand_1 g12746(n6441, n5314, new_n13123);
nand_1 g12747(n11791, n5767, new_n13124);
xnor_1 g12748(new_n13124, new_n13123, new_n13125);
nand_1 g12749(new_n12202, new_n12201, new_n13126);
nand_1 g12750(new_n12208, new_n12203, new_n13127);
nand_1 g12751(new_n13127, new_n13126, new_n13128);
and_1  g12752(n6687, n6604, new_n13129);
xnor_1 g12753(new_n13129, new_n13128, new_n13130);
xnor_1 g12754(new_n13130, new_n13125, new_n13131);
xnor_1 g12755(new_n13131, new_n13122, new_n13132);
xnor_1 g12756(new_n13132, new_n13104, new_n13133);
xnor_1 g12757(new_n13133, new_n13093, new_n13134);
not_1  g12758(new_n12084, new_n13135);
nand_1 g12759(new_n12092, new_n13135, new_n13136);
nand_1 g12760(new_n13136, new_n12089, new_n13137);
not_1  g12761(new_n12068, new_n13138);
nand_1 g12762(new_n12073, new_n13138, new_n13139);
not_1  g12763(new_n12083, new_n13140);
nand_1 g12764(new_n13140, new_n12074, new_n13141);
nand_1 g12765(new_n13141, new_n13139, new_n13142);
nor_1  g12766(new_n6725, new_n11208, new_n13143);
xnor_1 g12767(new_n13143, new_n13142, new_n13144);
nand_1 g12768(new_n12076_1, new_n12075, new_n13145);
not_1  g12769(new_n12082, new_n13146);
nand_1 g12770(new_n13146, new_n12077, new_n13147);
nand_1 g12771(new_n13147, new_n13145, new_n13148);
nor_1  g12772(new_n8622, new_n4529, new_n13149);
nand_1 g12773(n8819, n1094, new_n13150);
nand_1 g12774(n10928, n7730, new_n13151);
xnor_1 g12775(new_n13151, new_n13150, new_n13152);
xnor_1 g12776(new_n13152, new_n13149, new_n13153);
xnor_1 g12777(new_n13153, new_n13148, new_n13154);
xnor_1 g12778(new_n13154, new_n13144, new_n13155);
xnor_1 g12779(new_n13155, new_n13137, new_n13156);
xnor_1 g12780(new_n13156, new_n13134, new_n13157);
nor_1  g12781(new_n12214, new_n12114, new_n13158);
not_1  g12782(new_n12216, new_n13159);
nor_1  g12783(new_n13159, new_n12211, new_n13160);
nor_1  g12784(new_n13160, new_n13158, new_n13161);
nand_1 g12785(new_n12011, new_n12014_1, new_n13162);
nand_1 g12786(new_n12023, new_n12012, new_n13163);
nand_1 g12787(new_n13163, new_n13162, new_n13164);
xnor_1 g12788(new_n13164, new_n13161, new_n13165);
xnor_1 g12789(new_n13165, new_n13157, new_n13166);
and_1  g12790(new_n12217, new_n12136, new_n13167);
nor_1  g12791(new_n12219, new_n13048, new_n13168);
nor_1  g12792(new_n13168, new_n13167, new_n13169);
nand_1 g12793(new_n12093, new_n12057, new_n13170);
nand_1 g12794(new_n12094, new_n12065, new_n13171);
nand_1 g12795(new_n13171, new_n13170, new_n13172);
not_1  g12796(new_n11978, new_n13173);
nand_1 g12797(new_n11987, new_n13173, new_n13174);
not_1  g12798(new_n12003, new_n13175);
nand_1 g12799(new_n13175, new_n11988, new_n13176);
nand_1 g12800(new_n13176, new_n13174, new_n13177);
nand_1 g12801(new_n11984, new_n11979, new_n13178);
nand_1 g12802(new_n13178, new_n11985, new_n13179);
nand_1 g12803(n12709, n7523, new_n13180);
nor_1  g12804(new_n8561, new_n1367, new_n13181);
xnor_1 g12805(new_n13181, new_n13180, new_n13182);
xnor_1 g12806(new_n13182, new_n13179, new_n13183);
nand_1 g12807(n9725, n2564, new_n13184);
nand_1 g12808(n9920, n4370, new_n13185);
xnor_1 g12809(new_n13185, new_n13184, new_n13186);
nand_1 g12810(n5212, n4516, new_n13187);
nand_1 g12811(n6770, n5320, new_n13188);
nand_1 g12812(n5319, n1478, new_n13189);
xnor_1 g12813(new_n13189, new_n13188, new_n13190);
xnor_1 g12814(new_n13190, new_n13187, new_n13191);
xnor_1 g12815(new_n13191, new_n13186, new_n13192);
nand_1 g12816(n11728, n7320, new_n13193);
nand_1 g12817(new_n12080, new_n12079, new_n13194);
not_1  g12818(new_n13194, new_n13195);
nor_1  g12819(new_n12081, new_n12078, new_n13196);
nor_1  g12820(new_n13196, new_n13195, new_n13197);
xnor_1 g12821(new_n13197, new_n13193, new_n13198);
xnor_1 g12822(new_n13198, new_n13192, new_n13199);
xnor_1 g12823(new_n13199, new_n13183, new_n13200);
nand_1 g12824(new_n11997, new_n11992, new_n13201);
nand_1 g12825(new_n13201, new_n11999_1, new_n13202);
nand_1 g12826(n10990, n4817, new_n13203);
nand_1 g12827(n11877, n3627, new_n13204);
nand_1 g12828(n8336, n1198, new_n13205);
xnor_1 g12829(new_n13205, new_n13204, new_n13206);
xnor_1 g12830(new_n13206, new_n13203, new_n13207);
xnor_1 g12831(new_n13207, new_n13202, new_n13208);
nand_1 g12832(new_n11990, new_n11989, new_n13209);
nand_1 g12833(new_n12001, new_n11991, new_n13210);
nand_1 g12834(new_n13210, new_n13209, new_n13211);
nand_1 g12835(new_n12071, new_n12070, new_n13212);
not_1  g12836(new_n13212, new_n13213);
nor_1  g12837(new_n12072, new_n12069_1, new_n13214);
nor_1  g12838(new_n13214, new_n13213, new_n13215);
xnor_1 g12839(new_n13215, new_n13211, new_n13216);
xnor_1 g12840(new_n13216, new_n13208, new_n13217);
xnor_1 g12841(new_n13217, new_n13200, new_n13218);
xnor_1 g12842(new_n13218, new_n13177, new_n13219);
xnor_1 g12843(new_n13219, new_n13172, new_n13220);
xnor_1 g12844(new_n13220, new_n13169, new_n13221);
xnor_1 g12845(new_n13221, new_n13166, new_n13222);
xnor_1 g12846(new_n13222, new_n13074, new_n13223);
xnor_1 g12847(new_n13223, new_n13046, new_n13224);
xnor_1 g12848(new_n13224, new_n13042, n8100);
xnor_1 g12849(new_n9903, new_n9902, n8138);
xnor_1 g12850(new_n6268, new_n6267, n8202);
xor_1  g12851(new_n3881, new_n3870, n8303);
xnor_1 g12852(new_n3140, new_n3137, n8398);
xnor_1 g12853(new_n4508, new_n4507, n9137);
xnor_1 g12854(new_n7375, new_n7373, n9387);
xnor_1 g12855(new_n11734, new_n11733, n9571);
xor_1  g12856(new_n999, new_n998, n9578);
xor_1  g12857(new_n1274, new_n1272, n9706);
xnor_1 g12858(new_n4510, new_n4499_1, n9756);
nor_1  g12859(new_n7034, new_n7012, new_n13236);
nor_1  g12860(new_n13236, new_n7010, new_n13237);
nor_1  g12861(new_n4908, new_n4386, new_n13238);
or_1   g12862(new_n6736, new_n6680, new_n13239);
not_1  g12863(new_n6733, new_n13240);
nand_1 g12864(new_n6738, new_n13240, new_n13241);
nand_1 g12865(new_n13241, new_n13239, new_n13242);
xnor_1 g12866(new_n13242, new_n13238, new_n13243);
not_1  g12867(new_n6753, new_n13244);
nand_1 g12868(new_n6987, new_n13244, new_n13245);
nand_1 g12869(new_n7008, new_n6988, new_n13246);
nand_1 g12870(new_n13246, new_n13245, new_n13247);
and_1  g12871(n8336, n2278, new_n13248);
nand_1 g12872(new_n6636, new_n6639, new_n13249);
nand_1 g12873(new_n6651, new_n6637, new_n13250);
nand_1 g12874(new_n13250, new_n13249, new_n13251);
xnor_1 g12875(new_n13251, new_n13248, new_n13252);
nor_1  g12876(new_n6843, new_n6810, new_n13253);
nor_1  g12877(new_n6859, new_n6844, new_n13254);
nor_1  g12878(new_n13254, new_n13253, new_n13255);
not_1  g12879(new_n6579, new_n13256);
nor_1  g12880(new_n6615, new_n13256, new_n13257);
not_1  g12881(new_n6616, new_n13258);
nor_1  g12882(new_n6627, new_n13258, new_n13259);
nor_1  g12883(new_n13259, new_n13257, new_n13260);
not_1  g12884(new_n6713, new_n13261);
nand_1 g12885(new_n6720, new_n13261, new_n13262);
not_1  g12886(new_n6732, new_n13263);
nand_1 g12887(new_n13263, new_n6721, new_n13264);
nand_1 g12888(new_n13264, new_n13262, new_n13265);
nand_1 g12889(n11662, n6770, new_n13266);
nand_1 g12890(n10451, n2226, new_n13267);
nand_1 g12891(n5319, n3754, new_n13268);
xnor_1 g12892(new_n13268, new_n13267, new_n13269);
xnor_1 g12893(new_n13269, new_n13266, new_n13270);
nand_1 g12894(new_n6729, new_n6728, new_n13271);
not_1  g12895(new_n13271, new_n13272);
nor_1  g12896(new_n6730, new_n6726, new_n13273);
nor_1  g12897(new_n13273, new_n13272, new_n13274);
xnor_1 g12898(new_n13274, new_n13270, new_n13275);
nand_1 g12899(new_n6622, new_n6618, new_n13276);
nand_1 g12900(new_n13276, new_n6625, new_n13277);
nand_1 g12901(n10278, n6986, new_n13278);
nand_1 g12902(n10678, n3022, new_n13279);
xnor_1 g12903(new_n13279, new_n13278, new_n13280);
xnor_1 g12904(new_n13280, new_n13277, new_n13281);
xnor_1 g12905(new_n13281, new_n13275, new_n13282);
nand_1 g12906(new_n6722, new_n6659, new_n13283);
not_1  g12907(new_n6731, new_n13284);
nand_1 g12908(new_n13284, new_n6724, new_n13285);
nand_1 g12909(new_n13285, new_n13283, new_n13286);
nand_1 g12910(new_n6716, new_n6715, new_n13287);
not_1  g12911(new_n13287, new_n13288);
nor_1  g12912(new_n6719, new_n13288, new_n13289);
xnor_1 g12913(new_n13289, new_n13286, new_n13290);
xnor_1 g12914(new_n13290, new_n13282, new_n13291);
xnor_1 g12915(new_n13291, new_n13265, new_n13292);
xnor_1 g12916(new_n13292, new_n13260, new_n13293);
nand_1 g12917(new_n6609, new_n6608, new_n13294);
not_1  g12918(new_n13294, new_n13295);
nor_1  g12919(new_n6612, new_n13295, new_n13296);
nand_1 g12920(n8665, n2515, new_n13297);
nand_1 g12921(n10898, n9457, new_n13298);
nand_1 g12922(n12511, n11222, new_n13299);
xnor_1 g12923(new_n13299, new_n13298, new_n13300);
xnor_1 g12924(new_n13300, new_n13297, new_n13301);
xnor_1 g12925(new_n13301, new_n13296, new_n13302);
xnor_1 g12926(new_n13302, new_n13293, new_n13303);
nand_1 g12927(n12391, n4094, new_n13304);
not_1  g12928(new_n6606, new_n13305);
nand_1 g12929(new_n6613, new_n13305, new_n13306);
not_1  g12930(new_n6628, new_n13307);
nand_1 g12931(new_n13307, new_n6614, new_n13308);
nand_1 g12932(new_n13308, new_n13306, new_n13309);
nand_1 g12933(n4516, n3932, new_n13310);
nand_1 g12934(n7523, n6703, new_n13311);
xnor_1 g12935(new_n13311, new_n13310, new_n13312);
nand_1 g12936(n11423, n10928, new_n13313);
nand_1 g12937(n12591, n3627, new_n13314);
xnor_1 g12938(new_n13314, new_n13313, new_n13315);
xnor_1 g12939(new_n13315, new_n13312, new_n13316);
xnor_1 g12940(new_n13316, new_n13309, new_n13317);
nand_1 g12941(n11876, n4817, new_n13318);
nand_1 g12942(new_n6831, new_n6824, new_n13319);
nand_1 g12943(new_n13319, new_n6832, new_n13320);
nand_1 g12944(n10327, n4189, new_n13321);
nor_1  g12945(new_n11993, new_n4044, new_n13322);
xnor_1 g12946(new_n13322, new_n13321, new_n13323);
xnor_1 g12947(new_n13323, new_n13320, new_n13324);
xnor_1 g12948(new_n13324, new_n13318, new_n13325);
xnor_1 g12949(new_n13325, new_n13317, new_n13326);
xnor_1 g12950(new_n13326, new_n13304, new_n13327);
xnor_1 g12951(new_n13327, new_n13303, new_n13328);
xnor_1 g12952(new_n13328, new_n13255, new_n13329);
xnor_1 g12953(new_n13329, new_n13252, new_n13330);
not_1  g12954(new_n6629, new_n13331);
nand_1 g12955(new_n6635, new_n13331, new_n13332);
nand_1 g12956(new_n13332, new_n6632, new_n13333);
nor_1  g12957(new_n6840, new_n6782, new_n13334);
not_1  g12958(new_n6836, new_n13335);
not_1  g12959(new_n6842, new_n13336);
nor_1  g12960(new_n13336, new_n13335, new_n13337);
nor_1  g12961(new_n13337, new_n13334, new_n13338);
xnor_1 g12962(new_n13338, new_n13333, new_n13339);
nand_1 g12963(new_n6949, new_n6921, new_n13340);
nand_1 g12964(new_n13340, new_n6918, new_n13341);
nor_1  g12965(new_n4232, new_n8138_1, new_n13342);
xnor_1 g12966(new_n13342, new_n13341, new_n13343);
not_1  g12967(new_n6929, new_n13344);
nor_1  g12968(new_n13344, new_n6924, new_n13345);
nor_1  g12969(new_n6947, new_n13345, new_n13346);
nand_1 g12970(new_n6820, new_n6819, new_n13347);
nand_1 g12971(new_n6834, new_n6822_1, new_n13348);
nand_1 g12972(new_n13348, new_n13347, new_n13349);
nand_1 g12973(new_n6927, new_n6926, new_n13350);
not_1  g12974(new_n13350, new_n13351);
nor_1  g12975(new_n6928, new_n6925, new_n13352);
nor_1  g12976(new_n13352, new_n13351, new_n13353);
nand_1 g12977(new_n6938, new_n6937, new_n13354);
not_1  g12978(new_n13354, new_n13355);
nor_1  g12979(new_n6939, new_n6936, new_n13356);
nor_1  g12980(new_n13356, new_n13355, new_n13357);
xnor_1 g12981(new_n13357, new_n13353, new_n13358);
nand_1 g12982(n12069, n10685, new_n13359);
nor_1  g12983(new_n8087, new_n4195, new_n13360);
xnor_1 g12984(new_n13360, new_n13359, new_n13361);
nand_1 g12985(n5767, n2749, new_n13362);
nand_1 g12986(n996, n159, new_n13363);
nand_1 g12987(n5314, n1510, new_n13364);
xnor_1 g12988(new_n13364, new_n13363, new_n13365);
xnor_1 g12989(new_n13365, new_n13362, new_n13366);
xnor_1 g12990(new_n13366, new_n13361, new_n13367);
xnor_1 g12991(new_n13367, new_n13358, new_n13368);
nand_1 g12992(new_n6933, new_n6932, new_n13369);
nand_1 g12993(new_n6944, new_n13369, new_n13370);
nor_1  g12994(new_n1538, new_n4951, new_n13371);
nand_1 g12995(n9583, n2564, new_n13372);
nand_1 g12996(n9640, n7320, new_n13373);
xnor_1 g12997(new_n13373, new_n13372, new_n13374);
xnor_1 g12998(new_n13374, new_n13371, new_n13375);
nand_1 g12999(n1199, n1067, new_n13376);
nand_1 g13000(n12247, n11153, new_n13377);
xnor_1 g13001(new_n13377, new_n13376, new_n13378);
xnor_1 g13002(new_n13378, new_n13375, new_n13379);
xnor_1 g13003(new_n13379, new_n13370, new_n13380);
xnor_1 g13004(new_n13380, new_n13368, new_n13381);
xnor_1 g13005(new_n13381, new_n13349, new_n13382);
not_1  g13006(new_n6811, new_n13383);
nand_1 g13007(new_n6817, new_n13383, new_n13384);
nand_1 g13008(new_n6835, new_n6818, new_n13385);
nand_1 g13009(new_n13385, new_n13384, new_n13386);
nand_1 g13010(new_n6814, new_n6813, new_n13387);
not_1  g13011(new_n13387, new_n13388);
nor_1  g13012(new_n6815, new_n6812, new_n13389);
nor_1  g13013(new_n13389, new_n13388, new_n13390);
nand_1 g13014(n6687, n753, new_n13391);
nand_1 g13015(n2087, n1798, new_n13392);
xnor_1 g13016(new_n13392, new_n13391, new_n13393);
xnor_1 g13017(new_n13393, new_n13390, new_n13394);
xnor_1 g13018(new_n13394, new_n13386, new_n13395);
xnor_1 g13019(new_n13395, new_n13382, new_n13396);
xnor_1 g13020(new_n13396, new_n13346, new_n13397);
xnor_1 g13021(new_n13397, new_n13343, new_n13398);
xnor_1 g13022(new_n13398, new_n13339, new_n13399);
nand_1 g13023(new_n6951, new_n6954, new_n13400);
nand_1 g13024(new_n6965, new_n6952, new_n13401);
nand_1 g13025(new_n13401, new_n13400, new_n13402);
nor_1  g13026(new_n6740, new_n6712, new_n13403);
nor_1  g13027(new_n6752, new_n6741, new_n13404);
nor_1  g13028(new_n13404, new_n13403, new_n13405);
xnor_1 g13029(new_n13405, new_n13402, new_n13406);
xnor_1 g13030(new_n13406, new_n13399, new_n13407);
xnor_1 g13031(new_n13407, new_n13330, new_n13408);
nand_1 g13032(n11922, n4828, new_n13409);
not_1  g13033(new_n6985, new_n13410);
nand_1 g13034(new_n13410, new_n6966, new_n13411);
nand_1 g13035(new_n6986_1, new_n6860_1, new_n13412);
nand_1 g13036(new_n13412, new_n13411, new_n13413);
xnor_1 g13037(new_n13413, new_n13409, new_n13414);
xnor_1 g13038(new_n13414, new_n13408, new_n13415);
xnor_1 g13039(new_n13415, new_n13247, new_n13416);
xnor_1 g13040(new_n13416, new_n13243, new_n13417);
xnor_1 g13041(new_n13417, new_n13237, n9767);
xnor_1 g13042(new_n2266, new_n2265, n9820);
xnor_1 g13043(new_n9918, new_n9917, n9938);
xnor_1 g13044(new_n993, new_n992_1, n10476);
xnor_1 g13045(new_n990, new_n976, n10589);
xnor_1 g13046(new_n1270, new_n1267, n10695);
not_1  g13047(new_n3901, new_n13424);
nand_1 g13048(new_n3857, new_n3856, new_n13425);
xnor_1 g13049(new_n13425, new_n13424, n10789);
xor_1  g13050(new_n3130, new_n3122, n10851);
xnor_1 g13051(new_n5294, new_n5281, n10913);
xnor_1 g13052(new_n7496, new_n7380, n10949);
xnor_1 g13053(new_n11736, new_n11685, n11216);
xnor_1 g13054(new_n5282, new_n5274, n11326);
nand_1 g13055(new_n5835, new_n5589, new_n13432);
nand_1 g13056(new_n5966, new_n5836, new_n13433);
nand_1 g13057(new_n13433, new_n13432, new_n13434);
not_1  g13058(new_n5872, new_n13435);
nand_1 g13059(new_n5876, new_n13435, new_n13436);
nand_1 g13060(new_n5965, new_n5877, new_n13437);
nand_1 g13061(new_n13437, new_n13436, new_n13438);
not_1  g13062(new_n5870, new_n13439);
nand_1 g13063(new_n13439, new_n5841, new_n13440);
nand_1 g13064(new_n5871, new_n5839, new_n13441);
nand_1 g13065(new_n13441, new_n13440, new_n13442);
nand_1 g13066(new_n5869, new_n5861, new_n13443);
nand_1 g13067(new_n13443, new_n5866, new_n13444);
nand_1 g13068(n9763, n45, new_n13445);
nand_1 g13069(n8759, n7823, new_n13446);
xor_1  g13070(new_n13446, new_n13445, new_n13447);
xnor_1 g13071(new_n13447, new_n13444, new_n13448);
nand_1 g13072(new_n5562, new_n5561, new_n13449);
not_1  g13073(new_n13449, new_n13450);
nor_1  g13074(new_n5563, new_n5560, new_n13451);
nor_1  g13075(new_n13451, new_n13450, new_n13452);
nor_1  g13076(new_n2723, new_n1199_1, new_n13453);
xnor_1 g13077(new_n13453, new_n13452, new_n13454);
nand_1 g13078(n12705, n4634, new_n13455);
nand_1 g13079(n12145, n7436, new_n13456);
xnor_1 g13080(new_n13456, new_n13455, new_n13457);
nand_1 g13081(n9195, n4312, new_n13458);
nand_1 g13082(n10217, n6776, new_n13459);
xnor_1 g13083(new_n13459, new_n13458, new_n13460);
xnor_1 g13084(new_n13460, new_n13457, new_n13461);
xnor_1 g13085(new_n13461, new_n13454, new_n13462);
nand_1 g13086(new_n5851, new_n5850, new_n13463);
not_1  g13087(new_n5858, new_n13464);
nand_1 g13088(new_n13464, new_n5852, new_n13465);
nand_1 g13089(new_n13465, new_n13463, new_n13466);
nand_1 g13090(new_n5846, new_n5845, new_n13467);
not_1  g13091(new_n13467, new_n13468);
nor_1  g13092(new_n5847, new_n5844, new_n13469);
nor_1  g13093(new_n13469, new_n13468, new_n13470);
xnor_1 g13094(new_n13470, new_n13466, new_n13471);
xnor_1 g13095(new_n13471, new_n13462, new_n13472);
nor_1  g13096(new_n5856, new_n5855, new_n13473);
nand_1 g13097(new_n5856, new_n5855, new_n13474);
and_1  g13098(new_n13474, new_n5853, new_n13475);
nor_1  g13099(new_n13475, new_n13473, new_n13476);
xnor_1 g13100(new_n13476, new_n13472, new_n13477);
nor_1  g13101(new_n1084, new_n1219, new_n13478);
nand_1 g13102(n8276, n2522, new_n13479);
nand_1 g13103(n12299, n12221, new_n13480);
xnor_1 g13104(new_n13480, new_n13479, new_n13481);
xnor_1 g13105(new_n13481, new_n13478, new_n13482);
xnor_1 g13106(new_n13482, new_n13477, new_n13483);
not_1  g13107(new_n5843, new_n13484);
nand_1 g13108(new_n5848, new_n13484, new_n13485);
not_1  g13109(new_n5859, new_n13486);
nand_1 g13110(new_n13486, new_n5849, new_n13487);
nand_1 g13111(new_n13487, new_n13485, new_n13488);
nand_1 g13112(new_n5952, new_n5944, new_n13489);
nand_1 g13113(new_n13489, new_n5949, new_n13490);
xnor_1 g13114(new_n13490, new_n13488, new_n13491);
xnor_1 g13115(new_n13491, new_n13483, new_n13492);
xnor_1 g13116(new_n13492, new_n13448, new_n13493);
xnor_1 g13117(new_n13493, new_n13442, new_n13494);
nor_1  g13118(new_n511, new_n1139, new_n13495);
nand_1 g13119(new_n5558, new_n5557, new_n13496);
not_1  g13120(new_n5564, new_n13497);
nand_1 g13121(new_n13497, new_n5559, new_n13498);
nand_1 g13122(new_n13498, new_n13496, new_n13499);
xnor_1 g13123(new_n13499, new_n13495, new_n13500);
xnor_1 g13124(new_n13500, new_n13494, new_n13501);
or_1   g13125(new_n5929, new_n5923, new_n13502);
nand_1 g13126(new_n5942, new_n13502, new_n13503);
nand_1 g13127(n7690, n5579, new_n13504);
nand_1 g13128(n7388, n2507, new_n13505);
xnor_1 g13129(new_n13505, new_n13504, new_n13506);
nand_1 g13130(n7270, n2393, new_n13507);
nand_1 g13131(n5331, n1576, new_n13508);
xnor_1 g13132(new_n13508, new_n13507, new_n13509);
xnor_1 g13133(new_n13509, new_n13506, new_n13510);
nand_1 g13134(n3616, n2498, new_n13511);
nand_1 g13135(n12648, n6016, new_n13512);
xnor_1 g13136(new_n13512, new_n13511, new_n13513);
xnor_1 g13137(new_n13513, new_n13510, new_n13514);
nor_1  g13138(new_n5727, new_n740, new_n13515);
nand_1 g13139(n10644, n7946, new_n13516);
xnor_1 g13140(new_n13516, new_n13515, new_n13517);
nand_1 g13141(new_n5927, new_n5926, new_n13518);
not_1  g13142(new_n13518, new_n13519);
nor_1  g13143(new_n5928, new_n5925, new_n13520);
nor_1  g13144(new_n13520, new_n13519, new_n13521);
nand_1 g13145(new_n5553, new_n5552, new_n13522);
not_1  g13146(new_n13522, new_n13523);
nor_1  g13147(new_n5554, new_n5551, new_n13524);
nor_1  g13148(new_n13524, new_n13523, new_n13525);
xnor_1 g13149(new_n13525, new_n13521, new_n13526);
xnor_1 g13150(new_n13526, new_n13517, new_n13527);
xnor_1 g13151(new_n13527, new_n13514, new_n13528);
xnor_1 g13152(new_n13528, new_n13503, new_n13529);
not_1  g13153(new_n5905, new_n13530);
nand_1 g13154(new_n5913, new_n13530, new_n13531);
nand_1 g13155(new_n13531, new_n5910, new_n13532);
nand_1 g13156(new_n5937, new_n5936, new_n13533);
not_1  g13157(new_n13533, new_n13534);
nor_1  g13158(new_n5938, new_n5935, new_n13535);
nor_1  g13159(new_n13535, new_n13534, new_n13536);
nand_1 g13160(new_n5933, new_n5932, new_n13537);
not_1  g13161(new_n5939, new_n13538);
nand_1 g13162(new_n13538, new_n5934_1, new_n13539);
nand_1 g13163(new_n13539, new_n13537, new_n13540);
nand_1 g13164(n7965, n6431, new_n13541);
nor_1  g13165(new_n1215, new_n3280, new_n13542);
xnor_1 g13166(new_n13542, new_n13541, new_n13543);
nand_1 g13167(n11892, n5153, new_n13544);
nand_1 g13168(n5860, n806, new_n13545);
xnor_1 g13169(new_n13545, new_n13544, new_n13546);
nand_1 g13170(n10545, n521, new_n13547);
nand_1 g13171(n10547, n7265, new_n13548);
xnor_1 g13172(new_n13548, new_n13547, new_n13549);
xnor_1 g13173(new_n13549, new_n13546, new_n13550);
xnor_1 g13174(new_n13550, new_n13543, new_n13551);
xnor_1 g13175(new_n13551, new_n13540, new_n13552);
xnor_1 g13176(new_n13552, new_n13536, new_n13553);
xnor_1 g13177(new_n13553, new_n13532, new_n13554);
nand_1 g13178(new_n5555, new_n5548, new_n13555);
not_1  g13179(new_n5565, new_n13556);
nand_1 g13180(new_n13556, new_n5556, new_n13557);
nand_1 g13181(new_n13557, new_n13555, new_n13558);
nor_1  g13182(new_n5897, new_n5736, new_n13559);
not_1  g13183(new_n5898, new_n13560);
nor_1  g13184(new_n5903, new_n13560, new_n13561);
nor_1  g13185(new_n13561, new_n13559, new_n13562);
xnor_1 g13186(new_n13562, new_n13558, new_n13563);
xnor_1 g13187(new_n13563, new_n13554, new_n13564);
xnor_1 g13188(new_n13564, new_n13529, new_n13565);
nand_1 g13189(new_n5914, new_n5767_1, new_n13566);
nand_1 g13190(new_n5919, new_n5915, new_n13567);
nand_1 g13191(new_n13567, new_n13566, new_n13568);
not_1  g13192(new_n5566, new_n13569);
nand_1 g13193(new_n5574, new_n13569, new_n13570);
nand_1 g13194(new_n13570, new_n5571, new_n13571);
not_1  g13195(new_n5904, new_n13572);
nand_1 g13196(new_n13572, new_n5896, new_n13573);
nand_1 g13197(new_n13573, new_n5894, new_n13574);
nand_1 g13198(new_n5901, new_n5900, new_n13575);
not_1  g13199(new_n13575, new_n13576);
nor_1  g13200(new_n5902, new_n5899, new_n13577);
nor_1  g13201(new_n13577, new_n13576, new_n13578);
nand_1 g13202(n4499, n2558, new_n13579);
nand_1 g13203(n5305, n2512, new_n13580);
xnor_1 g13204(new_n13580, new_n13579, new_n13581);
xnor_1 g13205(new_n13581, new_n13578, new_n13582);
nor_1  g13206(new_n5885, new_n5879, new_n13583);
nor_1  g13207(new_n712, new_n5880, new_n13584);
nand_1 g13208(new_n13584, new_n13583, new_n13585);
not_1  g13209(new_n13583, new_n13586);
nand_1 g13210(new_n13584, new_n5729, new_n13587);
nand_1 g13211(new_n13587, new_n13586, new_n13588);
nand_1 g13212(new_n13588, new_n13585, new_n13589);
nand_1 g13213(n2253, n1097, new_n13590);
nand_1 g13214(n5964, n3865, new_n13591);
xnor_1 g13215(new_n13591, new_n13590, new_n13592);
xnor_1 g13216(new_n13592, new_n13589, new_n13593);
xnor_1 g13217(new_n13593, new_n13582, new_n13594);
xnor_1 g13218(new_n13594, new_n13574, new_n13595);
nand_1 g13219(n10510, n2024, new_n13596);
nand_1 g13220(n11257, n2879, new_n13597);
xnor_1 g13221(new_n13597, new_n13596, new_n13598);
xnor_1 g13222(new_n13598, new_n13595, new_n13599);
xnor_1 g13223(new_n13599, new_n13571, new_n13600);
xnor_1 g13224(new_n13600, new_n13568, new_n13601);
xnor_1 g13225(new_n13601, new_n13565, new_n13602);
xnor_1 g13226(new_n13602, new_n13501, new_n13603);
not_1  g13227(new_n5959, new_n13604);
nand_1 g13228(new_n13604, new_n5920, new_n13605);
nand_1 g13229(new_n5964_1, new_n5960, new_n13606);
nand_1 g13230(new_n13606, new_n13605, new_n13607);
nand_1 g13231(new_n5575, new_n5578, new_n13608);
nand_1 g13232(new_n5588, new_n5576, new_n13609);
nand_1 g13233(new_n13609, new_n13608, new_n13610);
nor_1  g13234(new_n5953, new_n5807, new_n13611);
not_1  g13235(new_n5954, new_n13612);
nor_1  g13236(new_n5958, new_n13612, new_n13613);
nor_1  g13237(new_n13613, new_n13611, new_n13614);
xnor_1 g13238(new_n13614, new_n13610, new_n13615);
xnor_1 g13239(new_n13615, new_n13607, new_n13616);
xnor_1 g13240(new_n13616, new_n13603, new_n13617);
xnor_1 g13241(new_n13617, new_n13438, new_n13618);
xnor_1 g13242(new_n13618, new_n13434, n11707);
xnor_1 g13243(new_n6491, new_n6489, n11755);
xor_1  g13244(new_n3894, new_n3893, n11780);
xnor_1 g13245(new_n10292, new_n10291, n11919);
xnor_1 g13246(new_n10294, new_n10279, n12005);
xnor_1 g13247(new_n10739, new_n10736, n12014);
not_1  g13248(new_n9056, new_n13625);
xnor_1 g13249(new_n13625, new_n9028, n12020);
xnor_1 g13250(new_n11728_1, new_n11693, n12076);
xnor_1 g13251(new_n12285, new_n12282, n12111);
xnor_1 g13252(new_n10741, new_n10729, n12444);
xnor_1 g13253(new_n5833, new_n5822, n12807);
endmodule


