// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Thu Jun 27 13:50:34 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533_1, new_n2534,
    new_n2535_1, new_n2536, new_n2537_1, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2546, new_n2547_1,
    new_n2548, new_n2549, new_n2550, new_n2552, new_n2553_1, new_n2554,
    new_n2555_1, new_n2557, new_n2558, new_n2559, new_n2560_1, new_n2561_1,
    new_n2562, new_n2563, new_n2564, new_n2565, new_n2566, new_n2567,
    new_n2568, new_n2569, new_n2570_1, new_n2571, new_n2572, new_n2573_1,
    new_n2574, new_n2575, new_n2576, new_n2577, new_n2578_1, new_n2579,
    new_n2580, new_n2581, new_n2582_1, new_n2583, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602_1, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619_1, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826_1, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886_1,
    new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945, new_n2946,
    new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971_1, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978_1, new_n2979_1, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985_1, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1,
    new_n3019, new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067_1, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3075, new_n3076_1, new_n3077, new_n3078, new_n3079,
    new_n3080, new_n3081, new_n3082, new_n3083, new_n3084, new_n3085,
    new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090, new_n3091,
    new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097,
    new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3162, new_n3163,
    new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235_1,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253_1,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260_1, new_n3261, new_n3262, new_n3263_1, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279_1, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289_1,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301_1,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306_1, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319,
    new_n3320_1, new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332_1, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505, new_n3506_1,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528_1, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541_1, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555_1, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561_1, new_n3562, new_n3563_1, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570_1, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582_1, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617_1, new_n3618_1, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642_1, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649_1, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665_1, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679_1, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710_1,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3724, new_n3725_1, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733_1, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740_1, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755_1, new_n3756, new_n3757, new_n3758_1, new_n3759,
    new_n3760_1, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781_1, new_n3782, new_n3783,
    new_n3784, new_n3785_1, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794_1, new_n3795_1,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828_1, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850_1, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869_1, new_n3870, new_n3871_1, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891_1,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909_1,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918_1, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925_1, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934_1, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945_1, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952_1,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959_1, new_n3960, new_n3961, new_n3962_1, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971_1, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983_1, new_n3984_1, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000_1,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010_1, new_n4011, new_n4012,
    new_n4013, new_n4014_1, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071_1, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085_1, new_n4086, new_n4087, new_n4088_1, new_n4089_1, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100_1, new_n4101, new_n4102,
    new_n4103_1, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119_1, new_n4120, new_n4121,
    new_n4122, new_n4123_1, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134_1, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146_1, new_n4147, new_n4148, new_n4149, new_n4150_1, new_n4151_1,
    new_n4152_1, new_n4153_1, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4165_1, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172_1, new_n4173_1, new_n4174, new_n4175, new_n4176_1,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186_1, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204_1, new_n4205_1, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215_1, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221_1, new_n4222, new_n4223, new_n4224_1,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231_1, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256_1, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266_1,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272_1,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4301, new_n4302, new_n4303,
    new_n4304, new_n4305, new_n4306_1, new_n4307, new_n4308, new_n4309,
    new_n4310, new_n4311, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319_1, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325_1, new_n4326_1, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340_1, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374_1, new_n4375,
    new_n4376_1, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401_1, new_n4402, new_n4403, new_n4404, new_n4405,
    new_n4406, new_n4407, new_n4408, new_n4409_1, new_n4410, new_n4411,
    new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4417,
    new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423,
    new_n4424_1, new_n4425, new_n4426_1, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4431, new_n4432_1, new_n4433, new_n4434, new_n4435,
    new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441_1,
    new_n4442, new_n4443, new_n4444, new_n4445, new_n4446, new_n4447,
    new_n4448, new_n4449, new_n4450, new_n4451_1, new_n4452, new_n4453,
    new_n4454, new_n4455, new_n4456, new_n4457, new_n4458, new_n4459,
    new_n4460, new_n4461, new_n4462, new_n4463, new_n4464, new_n4465,
    new_n4466, new_n4467, new_n4468, new_n4469, new_n4470, new_n4471,
    new_n4472, new_n4473, new_n4474, new_n4475, new_n4476_1, new_n4477,
    new_n4478_1, new_n4479, new_n4480, new_n4481, new_n4482, new_n4483,
    new_n4484, new_n4485, new_n4486, new_n4487, new_n4488, new_n4489,
    new_n4490, new_n4491, new_n4492, new_n4493, new_n4494, new_n4495,
    new_n4496, new_n4497, new_n4498, new_n4499, new_n4500, new_n4501,
    new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507,
    new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513,
    new_n4514_1, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519,
    new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525,
    new_n4526, new_n4527, new_n4528, new_n4529_1, new_n4530, new_n4531,
    new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537,
    new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543,
    new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549,
    new_n4550, new_n4551, new_n4552_1, new_n4553, new_n4554, new_n4555,
    new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561,
    new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567,
    new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573,
    new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588_1, new_n4589, new_n4590_1, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595_1, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624_1, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646_1,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652,
    new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658,
    new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665_1, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670,
    new_n4671, new_n4672, new_n4673, new_n4674_1, new_n4675, new_n4676,
    new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682,
    new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4689, new_n4690, new_n4691, new_n4692, new_n4693_1, new_n4694,
    new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731_1, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745_1, new_n4746, new_n4747_1, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760,
    new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766_1,
    new_n4767, new_n4769, new_n4770_1, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777_1, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785_1,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804_1, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810_1, new_n4811, new_n4812_1, new_n4813, new_n4814_1, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850_1, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858_1, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891_1, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913_1, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921, new_n4922, new_n4923,
    new_n4924, new_n4925_1, new_n4926, new_n4927, new_n4928, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938, new_n4939_1, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947_1,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952_1, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957_1, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964_1, new_n4965,
    new_n4966_1, new_n4967_1, new_n4968, new_n4969, new_n4970, new_n4971,
    new_n4972_1, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011_1, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020_1, new_n5021, new_n5022, new_n5023, new_n5024_1, new_n5025_1,
    new_n5026_1, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031_1,
    new_n5032, new_n5033, new_n5034, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046_1, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060_1, new_n5061, new_n5062_1,
    new_n5063, new_n5064_1, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077_1, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082_1, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098_1,
    new_n5099, new_n5100, new_n5101_1, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5107, new_n5108, new_n5109, new_n5110, new_n5111,
    new_n5112, new_n5113, new_n5114, new_n5115_1, new_n5116, new_n5117,
    new_n5118, new_n5119, new_n5120_1, new_n5121, new_n5122, new_n5123,
    new_n5124, new_n5125, new_n5126, new_n5127, new_n5128_1, new_n5129,
    new_n5130, new_n5131_1, new_n5132, new_n5133, new_n5134, new_n5135,
    new_n5136, new_n5137, new_n5138, new_n5139, new_n5140_1, new_n5141,
    new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147,
    new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153,
    new_n5154, new_n5155, new_n5156, new_n5157, new_n5158_1, new_n5159,
    new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168_1, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184_1, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211_1, new_n5212, new_n5213_1,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5218, new_n5219,
    new_n5220, new_n5221, new_n5222, new_n5223, new_n5224, new_n5225,
    new_n5226_1, new_n5227, new_n5228_1, new_n5229, new_n5230, new_n5231,
    new_n5232, new_n5233, new_n5234, new_n5235, new_n5236, new_n5237,
    new_n5238, new_n5239, new_n5240, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255_1, new_n5256_1,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265_1, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273_1, new_n5274_1,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300_1, new_n5301, new_n5302_1, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325_1, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330_1, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337_1, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351_1, new_n5352,
    new_n5353_1, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376_1,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386_1, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399_1, new_n5400_1,
    new_n5401, new_n5402, new_n5403_1, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430_1,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438_1, new_n5439_1, new_n5440, new_n5441, new_n5442,
    new_n5443_1, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451_1, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472_1,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5480, new_n5481, new_n5482, new_n5483, new_n5484, new_n5485_1,
    new_n5486, new_n5487, new_n5488, new_n5489, new_n5490, new_n5491,
    new_n5492, new_n5493, new_n5494, new_n5495, new_n5496, new_n5497,
    new_n5498, new_n5499, new_n5500, new_n5501, new_n5502, new_n5503,
    new_n5504, new_n5505, new_n5506, new_n5507, new_n5508, new_n5509,
    new_n5510, new_n5511, new_n5512, new_n5513, new_n5514, new_n5515,
    new_n5516, new_n5517_1, new_n5518, new_n5519, new_n5520, new_n5521_1,
    new_n5522, new_n5523, new_n5524_1, new_n5525, new_n5526, new_n5527,
    new_n5528, new_n5529, new_n5530, new_n5531, new_n5532_1, new_n5533,
    new_n5534, new_n5535, new_n5536, new_n5537, new_n5538, new_n5539,
    new_n5540, new_n5541, new_n5542, new_n5543, new_n5544, new_n5545,
    new_n5546, new_n5547, new_n5548, new_n5549, new_n5550, new_n5551,
    new_n5552, new_n5553, new_n5554, new_n5555, new_n5556, new_n5557,
    new_n5558, new_n5559, new_n5560, new_n5561, new_n5562, new_n5563,
    new_n5564_1, new_n5565, new_n5566, new_n5567, new_n5568, new_n5569,
    new_n5570, new_n5571, new_n5572, new_n5573, new_n5574, new_n5575,
    new_n5576, new_n5577, new_n5578, new_n5579_1, new_n5580, new_n5581,
    new_n5582, new_n5583, new_n5584, new_n5585, new_n5586, new_n5587,
    new_n5588, new_n5589, new_n5590, new_n5591, new_n5592, new_n5593_1,
    new_n5594, new_n5595, new_n5596, new_n5597, new_n5598, new_n5599,
    new_n5600, new_n5601, new_n5602, new_n5603_1, new_n5604, new_n5605_1,
    new_n5606, new_n5607, new_n5608, new_n5609_1, new_n5610, new_n5611,
    new_n5612, new_n5613, new_n5614, new_n5615, new_n5616, new_n5617,
    new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623,
    new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629,
    new_n5630, new_n5631, new_n5632, new_n5633, new_n5634_1, new_n5635,
    new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641,
    new_n5642, new_n5643_1, new_n5644, new_n5645, new_n5646, new_n5647,
    new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680_1, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687_1, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696_1, new_n5697, new_n5698, new_n5699, new_n5700_1, new_n5701,
    new_n5702, new_n5703, new_n5704_1, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732_1, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742_1, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752_1, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765_1, new_n5766, new_n5767,
    new_n5768, new_n5769, new_n5770, new_n5771, new_n5772, new_n5773,
    new_n5774, new_n5775, new_n5776_1, new_n5777, new_n5778, new_n5779,
    new_n5780, new_n5781, new_n5782_1, new_n5783, new_n5784, new_n5785,
    new_n5786, new_n5787, new_n5788, new_n5789, new_n5790, new_n5791,
    new_n5792, new_n5793, new_n5794, new_n5795, new_n5796, new_n5797,
    new_n5798, new_n5799, new_n5800, new_n5801, new_n5802, new_n5803,
    new_n5804, new_n5805, new_n5806, new_n5807, new_n5808, new_n5809,
    new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815,
    new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821,
    new_n5822_1, new_n5823, new_n5824, new_n5825, new_n5826, new_n5827,
    new_n5829, new_n5830, new_n5831, new_n5832, new_n5833_1, new_n5834_1,
    new_n5835, new_n5836, new_n5837, new_n5838, new_n5839, new_n5840_1,
    new_n5841_1, new_n5842_1, new_n5843, new_n5844, new_n5845, new_n5846,
    new_n5847, new_n5848, new_n5849, new_n5851, new_n5852, new_n5853,
    new_n5856, new_n5857, new_n5858, new_n5859, new_n5860, new_n5861,
    new_n5862, new_n5863, new_n5864, new_n5865, new_n5866, new_n5867,
    new_n5868, new_n5869, new_n5870, new_n5871, new_n5872, new_n5873,
    new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879,
    new_n5880, new_n5882_1, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903_1, new_n5904_1,
    new_n5905, new_n5906, new_n5910, new_n5911_1, new_n5912, new_n5913,
    new_n5914, new_n5915, new_n5916, new_n5917, new_n5918, new_n5919,
    new_n5920, new_n5921, new_n5922, new_n5923, new_n5924, new_n5925,
    new_n5926, new_n5927, new_n5928, new_n5929, new_n5930, new_n5931,
    new_n5932, new_n5933, new_n5934, new_n5935, new_n5936_1, new_n5937,
    new_n5938, new_n5939, new_n5940, new_n5941, new_n5942, new_n5943_1,
    new_n5944, new_n5945, new_n5946, new_n5947, new_n5948, new_n5949,
    new_n5950, new_n5951, new_n5952, new_n5953, new_n5954, new_n5955,
    new_n5956, new_n5957, new_n5958, new_n5959, new_n5960, new_n5961,
    new_n5962, new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967,
    new_n5968, new_n5969, new_n5970, new_n5971, new_n5972, new_n5973,
    new_n5974, new_n5975, new_n5976, new_n5977, new_n5978, new_n5979,
    new_n5980_1, new_n5981, new_n5982, new_n5983, new_n5984, new_n5985,
    new_n5986, new_n5987, new_n5988, new_n5989, new_n5990, new_n5991,
    new_n5992, new_n5993, new_n5994, new_n5995, new_n5996, new_n5997,
    new_n5998, new_n5999, new_n6000, new_n6001, new_n6002, new_n6003,
    new_n6004, new_n6005, new_n6006, new_n6007, new_n6008, new_n6009,
    new_n6010, new_n6011, new_n6012_1, new_n6013, new_n6014, new_n6015,
    new_n6016, new_n6017, new_n6018, new_n6019, new_n6020, new_n6021,
    new_n6022_1, new_n6023, new_n6024, new_n6025, new_n6026, new_n6027,
    new_n6028, new_n6029, new_n6030, new_n6031_1, new_n6032, new_n6033,
    new_n6034, new_n6035, new_n6036, new_n6037, new_n6038, new_n6039,
    new_n6040, new_n6041, new_n6042, new_n6043, new_n6044_1, new_n6045,
    new_n6046_1, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051,
    new_n6052, new_n6053, new_n6054, new_n6055, new_n6056, new_n6057,
    new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063,
    new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069,
    new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075,
    new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081,
    new_n6082, new_n6083, new_n6084_1, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104_1, new_n6105_1,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153,
    new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159,
    new_n6160_1, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165,
    new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171_1,
    new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183_1,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189_1,
    new_n6190, new_n6191, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204_1, new_n6205, new_n6206, new_n6207, new_n6208,
    new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214,
    new_n6215, new_n6216, new_n6217, new_n6218_1, new_n6219, new_n6220,
    new_n6221, new_n6222, new_n6223_1, new_n6224, new_n6225, new_n6226,
    new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232,
    new_n6233_1, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238,
    new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6244,
    new_n6245_1, new_n6246, new_n6247, new_n6248_1, new_n6249, new_n6250,
    new_n6251, new_n6252, new_n6253, new_n6254, new_n6255, new_n6256_1,
    new_n6257, new_n6258, new_n6259, new_n6260, new_n6261, new_n6262,
    new_n6263, new_n6264, new_n6265, new_n6266, new_n6267, new_n6268,
    new_n6269, new_n6270, new_n6271_1, new_n6272, new_n6273, new_n6274,
    new_n6275, new_n6276_1, new_n6277, new_n6278, new_n6279, new_n6280,
    new_n6281, new_n6282, new_n6283, new_n6284, new_n6285, new_n6286,
    new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292,
    new_n6293, new_n6294, new_n6295, new_n6296, new_n6297, new_n6298,
    new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304,
    new_n6305, new_n6306, new_n6307, new_n6308_1, new_n6309, new_n6310,
    new_n6311_1, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316,
    new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322,
    new_n6323_1, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328,
    new_n6329, new_n6330_1, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339_1, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354_1, new_n6355, new_n6356_1, new_n6357, new_n6358,
    new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369_1, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375_1, new_n6376,
    new_n6377, new_n6378, new_n6379_1, new_n6380, new_n6381_1, new_n6382,
    new_n6383_1, new_n6384, new_n6385_1, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397_1, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407_1, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427_1, new_n6428, new_n6429, new_n6430,
    new_n6431_1, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437_1, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442,
    new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6457_1, new_n6458, new_n6459, new_n6460, new_n6461,
    new_n6462, new_n6463, new_n6464, new_n6465_1, new_n6466, new_n6467,
    new_n6468, new_n6469, new_n6470_1, new_n6471, new_n6472, new_n6473,
    new_n6474, new_n6475, new_n6476_1, new_n6477, new_n6478, new_n6479,
    new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485_1,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502_1, new_n6503,
    new_n6504, new_n6505, new_n6506_1, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513_1, new_n6514_1, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542_1, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556_1, new_n6557,
    new_n6558_1, new_n6559, new_n6560_1, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567_1, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576_1, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587_1,
    new_n6588, new_n6589, new_n6590_1, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596_1, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611_1,
    new_n6612_1, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6629, new_n6630_1,
    new_n6631_1, new_n6632, new_n6634_1, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6650, new_n6651, new_n6652_1, new_n6653, new_n6654, new_n6655_1,
    new_n6656, new_n6657, new_n6658, new_n6659_1, new_n6660, new_n6661,
    new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667,
    new_n6668, new_n6669_1, new_n6670, new_n6671_1, new_n6672, new_n6673_1,
    new_n6674_1, new_n6675, new_n6676, new_n6677, new_n6678, new_n6679,
    new_n6680, new_n6681, new_n6682, new_n6683, new_n6684_1, new_n6685,
    new_n6686, new_n6687, new_n6688, new_n6689, new_n6690, new_n6691_1,
    new_n6692, new_n6693, new_n6694, new_n6695, new_n6696, new_n6697,
    new_n6698, new_n6699, new_n6700, new_n6701, new_n6702, new_n6703,
    new_n6704, new_n6705, new_n6706_1, new_n6707_1, new_n6708, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729_1, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736_1, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6743, new_n6744, new_n6745, new_n6746,
    new_n6747, new_n6748, new_n6749, new_n6750, new_n6751, new_n6752,
    new_n6753, new_n6754, new_n6755, new_n6756, new_n6757, new_n6758,
    new_n6759, new_n6760, new_n6761, new_n6762, new_n6763, new_n6764,
    new_n6765, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770,
    new_n6771, new_n6772, new_n6773_1, new_n6775_1, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785_1, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790_1, new_n6791_1, new_n6792, new_n6793, new_n6794_1, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802_1, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814_1, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835_1, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853_1, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861_1,
    new_n6862_1, new_n6863_1, new_n6864, new_n6865, new_n6866, new_n6867_1,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965_1, new_n6966, new_n6967_1, new_n6968, new_n6969,
    new_n6970, new_n6971_1, new_n6972, new_n6973, new_n6974, new_n6975_1,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983_1, new_n6984, new_n6985_1, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6995, new_n6996, new_n6997, new_n6998_1, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026_1, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032_1, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038_1, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057_1, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072,
    new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078,
    new_n7079_1, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084,
    new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090,
    new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096,
    new_n7097, new_n7098, new_n7099_1, new_n7100, new_n7101, new_n7102,
    new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108,
    new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114,
    new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120,
    new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139_1, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149_1, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190_1, new_n7191, new_n7192,
    new_n7193, new_n7194, new_n7195, new_n7196, new_n7197, new_n7198,
    new_n7199, new_n7200, new_n7201, new_n7202, new_n7203, new_n7204,
    new_n7205, new_n7206, new_n7207, new_n7208, new_n7209, new_n7210,
    new_n7211, new_n7212, new_n7213, new_n7214, new_n7215, new_n7216,
    new_n7217, new_n7218, new_n7219, new_n7220, new_n7221, new_n7222,
    new_n7223, new_n7224, new_n7225, new_n7226, new_n7227, new_n7228,
    new_n7229_1, new_n7230_1, new_n7231, new_n7232, new_n7233_1, new_n7234,
    new_n7235, new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240,
    new_n7241, new_n7242, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7250, new_n7251, new_n7252, new_n7253_1, new_n7254,
    new_n7255, new_n7256_1, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268_1, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277_1, new_n7278,
    new_n7279, new_n7280_1, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298_1, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305_1, new_n7306, new_n7307, new_n7308_1,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313_1, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330_1, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335_1, new_n7336, new_n7337, new_n7338,
    new_n7339_1, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346_1, new_n7347, new_n7348, new_n7349_1, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363_1, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377_1, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390_1, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403_1, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408_1, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421_1, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428_1,
    new_n7429, new_n7430, new_n7431, new_n7432_1, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437_1, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460_1, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475_1, new_n7476,
    new_n7477_1, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7513,
    new_n7514_1, new_n7515, new_n7516, new_n7517, new_n7518, new_n7519,
    new_n7520, new_n7521, new_n7522, new_n7523, new_n7524_1, new_n7525,
    new_n7526, new_n7527, new_n7528, new_n7529, new_n7530, new_n7531,
    new_n7532, new_n7533, new_n7534, new_n7535, new_n7536, new_n7537,
    new_n7538, new_n7539, new_n7540, new_n7541, new_n7542, new_n7543,
    new_n7544, new_n7545, new_n7546, new_n7547, new_n7548, new_n7549,
    new_n7550, new_n7551, new_n7552, new_n7553, new_n7554, new_n7555,
    new_n7556, new_n7557, new_n7558_1, new_n7559, new_n7560, new_n7561,
    new_n7562, new_n7563, new_n7564, new_n7565, new_n7566_1, new_n7567,
    new_n7568, new_n7569_1, new_n7570, new_n7571, new_n7572_1, new_n7573,
    new_n7574, new_n7575_1, new_n7576, new_n7577, new_n7578, new_n7579,
    new_n7580, new_n7581, new_n7582, new_n7583, new_n7584, new_n7585_1,
    new_n7586, new_n7587, new_n7588_1, new_n7589, new_n7590, new_n7591,
    new_n7592, new_n7593_1, new_n7594, new_n7595, new_n7596, new_n7597,
    new_n7598_1, new_n7599, new_n7600, new_n7601, new_n7602, new_n7603,
    new_n7604, new_n7605, new_n7606, new_n7607_1, new_n7608, new_n7609,
    new_n7610_1, new_n7611, new_n7612, new_n7613, new_n7614, new_n7615,
    new_n7616_1, new_n7617, new_n7618, new_n7619, new_n7620, new_n7621,
    new_n7622, new_n7623, new_n7624, new_n7625, new_n7626, new_n7627,
    new_n7628, new_n7629, new_n7630_1, new_n7631, new_n7632, new_n7633,
    new_n7634, new_n7635, new_n7636, new_n7637, new_n7638, new_n7639,
    new_n7640, new_n7641, new_n7642, new_n7643_1, new_n7644, new_n7645,
    new_n7646, new_n7647_1, new_n7648, new_n7649, new_n7650, new_n7651,
    new_n7652, new_n7653, new_n7654, new_n7655, new_n7656, new_n7657_1,
    new_n7658, new_n7659, new_n7660, new_n7661, new_n7662, new_n7663,
    new_n7664, new_n7665, new_n7666, new_n7667, new_n7668, new_n7669,
    new_n7670_1, new_n7671, new_n7672, new_n7673, new_n7674_1, new_n7675,
    new_n7676, new_n7677, new_n7678_1, new_n7679_1, new_n7680, new_n7681,
    new_n7682, new_n7683, new_n7684, new_n7685, new_n7686_1, new_n7687,
    new_n7688, new_n7689, new_n7690, new_n7691, new_n7692_1, new_n7693_1,
    new_n7694, new_n7695, new_n7696, new_n7697, new_n7698_1, new_n7699,
    new_n7700, new_n7701, new_n7702, new_n7703, new_n7704, new_n7705,
    new_n7706, new_n7707, new_n7708_1, new_n7709, new_n7710, new_n7711,
    new_n7712, new_n7713, new_n7714, new_n7715, new_n7716, new_n7717,
    new_n7718, new_n7719, new_n7720, new_n7721_1, new_n7722, new_n7723,
    new_n7724, new_n7725, new_n7726, new_n7728, new_n7729, new_n7730,
    new_n7731_1, new_n7732, new_n7733, new_n7734, new_n7735, new_n7736,
    new_n7737, new_n7738, new_n7739, new_n7740, new_n7741, new_n7742,
    new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748,
    new_n7749, new_n7750, new_n7751_1, new_n7752, new_n7753, new_n7754,
    new_n7755, new_n7756, new_n7757, new_n7758, new_n7759_1, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769_1, new_n7770, new_n7771, new_n7772,
    new_n7773_1, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780_1, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788_1, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794_1, new_n7795, new_n7796,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811_1, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820,
    new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826,
    new_n7827, new_n7828, new_n7829, new_n7830_1, new_n7831, new_n7832,
    new_n7833, new_n7834_1, new_n7835, new_n7836, new_n7837, new_n7838,
    new_n7839, new_n7840, new_n7841_1, new_n7842, new_n7843, new_n7844,
    new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850,
    new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856,
    new_n7857, new_n7858, new_n7859, new_n7860, new_n7861, new_n7862,
    new_n7863, new_n7864, new_n7865, new_n7866, new_n7867, new_n7868,
    new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874,
    new_n7875, new_n7876_1, new_n7877, new_n7878, new_n7879, new_n7880,
    new_n7881, new_n7882, new_n7883, new_n7884_1, new_n7885, new_n7886,
    new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892,
    new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898,
    new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917_1, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937_1, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943_1, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949_1, new_n7950_1, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959_1, new_n7960, new_n7961, new_n7962, new_n7963_1, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968_1, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992_1, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999_1, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006_1,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027_1, new_n8028, new_n8029, new_n8030,
    new_n8031_1, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042_1,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8050, new_n8051, new_n8052_1, new_n8053, new_n8054, new_n8055,
    new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061,
    new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067_1,
    new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073,
    new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079,
    new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085,
    new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091,
    new_n8092, new_n8093, new_n8094, new_n8095_1, new_n8096, new_n8097,
    new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8103_1,
    new_n8104, new_n8105, new_n8106, new_n8107, new_n8108, new_n8109_1,
    new_n8110, new_n8111, new_n8112, new_n8113, new_n8114, new_n8115,
    new_n8116, new_n8117, new_n8118, new_n8119, new_n8120, new_n8121,
    new_n8122, new_n8123, new_n8124, new_n8125, new_n8126, new_n8127_1,
    new_n8128, new_n8129, new_n8130_1, new_n8131, new_n8132, new_n8133,
    new_n8134, new_n8135_1, new_n8136, new_n8137, new_n8138, new_n8139_1,
    new_n8140, new_n8141, new_n8142, new_n8143, new_n8144, new_n8145,
    new_n8146, new_n8147, new_n8148_1, new_n8149_1, new_n8150, new_n8151,
    new_n8152, new_n8153, new_n8154, new_n8155, new_n8156, new_n8157,
    new_n8158, new_n8159_1, new_n8160, new_n8161, new_n8162, new_n8163,
    new_n8164, new_n8165, new_n8166, new_n8167, new_n8168, new_n8169,
    new_n8170, new_n8171, new_n8172, new_n8173, new_n8174, new_n8175,
    new_n8176, new_n8177, new_n8178, new_n8179_1, new_n8180, new_n8181,
    new_n8182, new_n8183, new_n8184, new_n8185, new_n8186, new_n8187,
    new_n8188, new_n8189, new_n8190, new_n8191, new_n8192, new_n8193,
    new_n8194_1, new_n8195, new_n8196, new_n8197, new_n8198, new_n8199,
    new_n8200, new_n8201, new_n8202, new_n8203, new_n8204, new_n8205,
    new_n8206, new_n8207, new_n8208, new_n8209, new_n8210, new_n8211,
    new_n8212, new_n8213, new_n8214, new_n8215_1, new_n8216, new_n8217,
    new_n8218, new_n8219, new_n8220, new_n8221, new_n8222, new_n8223,
    new_n8224, new_n8225, new_n8226, new_n8227, new_n8228, new_n8229,
    new_n8230, new_n8231, new_n8232, new_n8233, new_n8234, new_n8235,
    new_n8236, new_n8237, new_n8238, new_n8239, new_n8240, new_n8241,
    new_n8242, new_n8243, new_n8244_1, new_n8245, new_n8246, new_n8247,
    new_n8248, new_n8249, new_n8250, new_n8251, new_n8252, new_n8253,
    new_n8254, new_n8255_1, new_n8256_1, new_n8257, new_n8258, new_n8259_1,
    new_n8260, new_n8261, new_n8262, new_n8263, new_n8264, new_n8265,
    new_n8266, new_n8267_1, new_n8268, new_n8269, new_n8270, new_n8271,
    new_n8272, new_n8273, new_n8274, new_n8275, new_n8276_1, new_n8277,
    new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283,
    new_n8284, new_n8285_1, new_n8286, new_n8287, new_n8288_1, new_n8289,
    new_n8290, new_n8291, new_n8292, new_n8293, new_n8294, new_n8295,
    new_n8296, new_n8297, new_n8298, new_n8299, new_n8300, new_n8301,
    new_n8302, new_n8303, new_n8304, new_n8305_1, new_n8306_1, new_n8307,
    new_n8308, new_n8309_1, new_n8310, new_n8311, new_n8312, new_n8313,
    new_n8314, new_n8315, new_n8316, new_n8317, new_n8318, new_n8319,
    new_n8320_1, new_n8321_1, new_n8322, new_n8323, new_n8324_1, new_n8325,
    new_n8326, new_n8327, new_n8328, new_n8329, new_n8330, new_n8331,
    new_n8332, new_n8333, new_n8334, new_n8335, new_n8336, new_n8337,
    new_n8338, new_n8339_1, new_n8340, new_n8341, new_n8342, new_n8343,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363_1,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376_1, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381_1,
    new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398, new_n8399_1,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405_1,
    new_n8406, new_n8407, new_n8408_1, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417_1,
    new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423,
    new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432_1, new_n8433, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439_1, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453_1,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476, new_n8477,
    new_n8478, new_n8479, new_n8480_1, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489_1,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505_1, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510_1, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519_1,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526_1, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535_1, new_n8536, new_n8537,
    new_n8538, new_n8540, new_n8541, new_n8542, new_n8543, new_n8544,
    new_n8545, new_n8546, new_n8547, new_n8548, new_n8549, new_n8550_1,
    new_n8551, new_n8552, new_n8553, new_n8554, new_n8555, new_n8556,
    new_n8557, new_n8558, new_n8559, new_n8560, new_n8561, new_n8562,
    new_n8563_1, new_n8564, new_n8565, new_n8566, new_n8567, new_n8568,
    new_n8569, new_n8570, new_n8571, new_n8572, new_n8573, new_n8574,
    new_n8575, new_n8576, new_n8577, new_n8579, new_n8580, new_n8581_1,
    new_n8582, new_n8583, new_n8584, new_n8585, new_n8586, new_n8587,
    new_n8588, new_n8589, new_n8590, new_n8591, new_n8592, new_n8593,
    new_n8594_1, new_n8595, new_n8596, new_n8597, new_n8598, new_n8599,
    new_n8600, new_n8601, new_n8602, new_n8603, new_n8604, new_n8605,
    new_n8606, new_n8607, new_n8608_1, new_n8609, new_n8610, new_n8611,
    new_n8612, new_n8613, new_n8614_1, new_n8615, new_n8616, new_n8617,
    new_n8618, new_n8619, new_n8620_1, new_n8621, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637_1, new_n8638_1, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656_1, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662_1, new_n8663, new_n8664, new_n8665, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678_1,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687_1, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694_1, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716_1, new_n8717, new_n8718, new_n8719, new_n8720,
    new_n8721_1, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8730, new_n8731, new_n8732, new_n8733,
    new_n8734, new_n8735, new_n8736, new_n8737, new_n8738, new_n8739,
    new_n8740, new_n8741, new_n8742, new_n8743, new_n8744_1, new_n8745_1,
    new_n8746, new_n8747, new_n8748, new_n8749, new_n8750, new_n8751,
    new_n8752, new_n8753, new_n8754, new_n8755, new_n8756, new_n8757,
    new_n8758, new_n8759, new_n8760, new_n8761, new_n8762, new_n8763,
    new_n8764, new_n8765, new_n8766, new_n8767, new_n8768, new_n8769,
    new_n8770, new_n8771, new_n8772, new_n8773, new_n8774, new_n8775,
    new_n8776, new_n8777, new_n8778, new_n8779, new_n8780, new_n8781,
    new_n8782_1, new_n8783, new_n8784, new_n8785, new_n8786, new_n8787,
    new_n8788, new_n8789, new_n8790, new_n8791, new_n8792, new_n8793,
    new_n8794, new_n8795, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803_1, new_n8804, new_n8805, new_n8806_1,
    new_n8807, new_n8808, new_n8809_1, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819, new_n8820, new_n8821_1, new_n8822, new_n8823, new_n8824_1,
    new_n8825, new_n8826, new_n8827_1, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849_1, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856_1, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861_1, new_n8862_1, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869_1, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884_1,
    new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890,
    new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896,
    new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902,
    new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908,
    new_n8909_1, new_n8910, new_n8911_1, new_n8912, new_n8913, new_n8914,
    new_n8915, new_n8916, new_n8917, new_n8918, new_n8919, new_n8920_1,
    new_n8921, new_n8922, new_n8923, new_n8924, new_n8925, new_n8926,
    new_n8927, new_n8928, new_n8929, new_n8930, new_n8931, new_n8932,
    new_n8933, new_n8934, new_n8935, new_n8936, new_n8937, new_n8938,
    new_n8939, new_n8940, new_n8941, new_n8942, new_n8943_1, new_n8944,
    new_n8945, new_n8946, new_n8947, new_n8948, new_n8949, new_n8950,
    new_n8951, new_n8952, new_n8953, new_n8954, new_n8955, new_n8956,
    new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962,
    new_n8963, new_n8964_1, new_n8965, new_n8966, new_n8967, new_n8968,
    new_n8969, new_n8970, new_n8971_1, new_n8972, new_n8973, new_n8974,
    new_n8975, new_n8976, new_n8977, new_n8978, new_n8979, new_n8980,
    new_n8981, new_n8982_1, new_n8983, new_n8984, new_n8985, new_n8986,
    new_n8987, new_n8988, new_n8989, new_n8990, new_n8991, new_n8992,
    new_n8993_1, new_n8994, new_n8995, new_n8996, new_n8997, new_n8998,
    new_n8999, new_n9000, new_n9001, new_n9002, new_n9003_1, new_n9004,
    new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010,
    new_n9011, new_n9012_1, new_n9013, new_n9014, new_n9015, new_n9016,
    new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022,
    new_n9023, new_n9024, new_n9025, new_n9026, new_n9027, new_n9028,
    new_n9029, new_n9030, new_n9031, new_n9032_1, new_n9033, new_n9034,
    new_n9035, new_n9036, new_n9037, new_n9038, new_n9039, new_n9040,
    new_n9041, new_n9042_1, new_n9043, new_n9044, new_n9045, new_n9046_1,
    new_n9047_1, new_n9048, new_n9049, new_n9050, new_n9051, new_n9052,
    new_n9053, new_n9054, new_n9055, new_n9056, new_n9057, new_n9058,
    new_n9059, new_n9060, new_n9061, new_n9062, new_n9063, new_n9064,
    new_n9065, new_n9066, new_n9067, new_n9068, new_n9069, new_n9070,
    new_n9071, new_n9072, new_n9073, new_n9074, new_n9075, new_n9076,
    new_n9077, new_n9078, new_n9079, new_n9080, new_n9081, new_n9082,
    new_n9083, new_n9084, new_n9085, new_n9086, new_n9087, new_n9089,
    new_n9090_1, new_n9091, new_n9092, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104_1, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129_1, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146_1, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164_1, new_n9165, new_n9166_1, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172_1, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182_1, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191_1, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217_1, new_n9218, new_n9219, new_n9220_1, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246_1,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251_1, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259_1, new_n9260, new_n9261_1, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287_1, new_n9288,
    new_n9289, new_n9291, new_n9292, new_n9293, new_n9294, new_n9295,
    new_n9296, new_n9297, new_n9298, new_n9299, new_n9300, new_n9301,
    new_n9302, new_n9303, new_n9304, new_n9305, new_n9306, new_n9307,
    new_n9308_1, new_n9309, new_n9310, new_n9311, new_n9312, new_n9313,
    new_n9314, new_n9315, new_n9316, new_n9317, new_n9318_1, new_n9319,
    new_n9320, new_n9321, new_n9322, new_n9323_1, new_n9324, new_n9325,
    new_n9326, new_n9327, new_n9328, new_n9329, new_n9330, new_n9331,
    new_n9332, new_n9333, new_n9334, new_n9335, new_n9336, new_n9337,
    new_n9338, new_n9339, new_n9340, new_n9341, new_n9342, new_n9343,
    new_n9344_1, new_n9345, new_n9346, new_n9347, new_n9348, new_n9349,
    new_n9350, new_n9351, new_n9352, new_n9353, new_n9354, new_n9355,
    new_n9356, new_n9357, new_n9358, new_n9359, new_n9360, new_n9361,
    new_n9362, new_n9363, new_n9364_1, new_n9365, new_n9366, new_n9367,
    new_n9368, new_n9369, new_n9370, new_n9371_1, new_n9372_1, new_n9373,
    new_n9374, new_n9375, new_n9376, new_n9377, new_n9378, new_n9379,
    new_n9380_1, new_n9381, new_n9382_1, new_n9383, new_n9384, new_n9385,
    new_n9386, new_n9387, new_n9388, new_n9389, new_n9390, new_n9391,
    new_n9392, new_n9393, new_n9394, new_n9395, new_n9396_1, new_n9397,
    new_n9398, new_n9399_1, new_n9400, new_n9401, new_n9402, new_n9403_1,
    new_n9404, new_n9405, new_n9406, new_n9407, new_n9408, new_n9409,
    new_n9410, new_n9411, new_n9412, new_n9413, new_n9414, new_n9415,
    new_n9416, new_n9417, new_n9418, new_n9419_1, new_n9420, new_n9421,
    new_n9422, new_n9423_1, new_n9424, new_n9425, new_n9426, new_n9427,
    new_n9428, new_n9429, new_n9430_1, new_n9431, new_n9432, new_n9433,
    new_n9434, new_n9435_1, new_n9436, new_n9437, new_n9438, new_n9439,
    new_n9440, new_n9441, new_n9442, new_n9443, new_n9444, new_n9445_1,
    new_n9446, new_n9447, new_n9448, new_n9449, new_n9450, new_n9451_1,
    new_n9452, new_n9453, new_n9454, new_n9455, new_n9456, new_n9457,
    new_n9458_1, new_n9459_1, new_n9460_1, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493_1, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507_1, new_n9508_1, new_n9509,
    new_n9510, new_n9511, new_n9512_1, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552_1, new_n9553, new_n9554_1, new_n9555, new_n9556_1,
    new_n9557_1, new_n9558_1, new_n9559, new_n9560, new_n9561, new_n9562,
    new_n9563, new_n9564, new_n9565, new_n9566, new_n9567, new_n9568,
    new_n9569, new_n9570, new_n9571, new_n9572, new_n9573, new_n9574,
    new_n9575, new_n9576, new_n9577, new_n9578, new_n9579, new_n9580,
    new_n9581, new_n9582, new_n9583, new_n9584, new_n9585, new_n9586,
    new_n9587, new_n9588, new_n9589, new_n9590, new_n9591, new_n9592,
    new_n9593, new_n9594, new_n9595, new_n9596, new_n9597, new_n9598_1,
    new_n9599, new_n9600, new_n9601, new_n9602, new_n9603, new_n9604,
    new_n9605, new_n9606, new_n9607, new_n9608, new_n9609, new_n9610,
    new_n9611, new_n9612, new_n9613, new_n9614, new_n9615, new_n9616_1,
    new_n9617, new_n9618, new_n9619, new_n9620, new_n9621, new_n9622_1,
    new_n9623, new_n9624, new_n9625, new_n9626_1, new_n9627, new_n9628,
    new_n9629, new_n9630, new_n9631, new_n9633_1, new_n9634, new_n9635_1,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646_1, new_n9647,
    new_n9648_1, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655_1, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689_1,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695_1,
    new_n9696, new_n9697, new_n9698, new_n9699_1, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725, new_n9726_1, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739,
    new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753_1, new_n9754, new_n9755, new_n9756, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761_1, new_n9762, new_n9763_1,
    new_n9764, new_n9765, new_n9766, new_n9767_1, new_n9768, new_n9769,
    new_n9770, new_n9771_1, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778_1, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783_1, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799,
    new_n9800, new_n9801, new_n9802, new_n9803_1, new_n9804, new_n9805,
    new_n9806, new_n9807, new_n9808, new_n9809, new_n9811, new_n9812,
    new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818,
    new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832_1, new_n9833_1, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838_1, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848,
    new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867_1, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872_1,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890_1,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896,
    new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902,
    new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908,
    new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914,
    new_n9915, new_n9916, new_n9917_1, new_n9918, new_n9919_1, new_n9920,
    new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926_1,
    new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932,
    new_n9933, new_n9934_1, new_n9935, new_n9936, new_n9937, new_n9938_1,
    new_n9939, new_n9940, new_n9941, new_n9942_1, new_n9943, new_n9944,
    new_n9945, new_n9947, new_n9948, new_n9950, new_n9951, new_n9952,
    new_n9953, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967_1, new_n9968_1, new_n9969, new_n9970, new_n9971,
    new_n9973, new_n9974, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009_1, new_n10010_1, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017_1, new_n10018_1,
    new_n10019_1, new_n10020, new_n10021_1, new_n10022, new_n10023,
    new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10048, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053_1, new_n10054, new_n10055_1, new_n10056, new_n10057_1,
    new_n10058, new_n10059, new_n10060, new_n10061, new_n10062, new_n10063,
    new_n10064, new_n10065, new_n10066, new_n10067, new_n10068, new_n10069,
    new_n10070, new_n10071, new_n10072, new_n10073, new_n10074, new_n10075,
    new_n10076, new_n10077, new_n10078, new_n10079, new_n10080, new_n10081,
    new_n10082, new_n10083, new_n10084, new_n10085, new_n10086, new_n10087,
    new_n10088, new_n10089, new_n10090, new_n10091, new_n10092, new_n10093,
    new_n10094, new_n10095, new_n10096_1, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101_1, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111_1, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117_1, new_n10118, new_n10119,
    new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125_1, new_n10126, new_n10127, new_n10128, new_n10129,
    new_n10130, new_n10131, new_n10132, new_n10133, new_n10134, new_n10135,
    new_n10136, new_n10137, new_n10138, new_n10139, new_n10140, new_n10141,
    new_n10142, new_n10143, new_n10144, new_n10145, new_n10146, new_n10147,
    new_n10148, new_n10149, new_n10150, new_n10151, new_n10152, new_n10153,
    new_n10154, new_n10155, new_n10156, new_n10157, new_n10158_1,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165_1, new_n10166, new_n10167, new_n10168, new_n10169,
    new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201_1, new_n10202, new_n10203, new_n10204,
    new_n10205, new_n10206, new_n10207, new_n10208, new_n10209, new_n10210,
    new_n10211, new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217, new_n10218, new_n10219, new_n10220, new_n10221, new_n10222,
    new_n10223, new_n10224, new_n10225, new_n10226, new_n10227, new_n10228,
    new_n10229, new_n10230, new_n10231, new_n10232, new_n10233, new_n10234,
    new_n10235, new_n10236_1, new_n10237, new_n10238, new_n10239_1,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244_1,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249,
    new_n10250_1, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261_1, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275_1, new_n10276, new_n10277,
    new_n10278, new_n10279, new_n10280, new_n10281, new_n10282, new_n10283,
    new_n10284, new_n10285, new_n10286, new_n10287_1, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295_1, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10321_1, new_n10322,
    new_n10323, new_n10324, new_n10325, new_n10326_1, new_n10327_1,
    new_n10328, new_n10329, new_n10330_1, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340_1, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345_1, new_n10346, new_n10347, new_n10348,
    new_n10349, new_n10350, new_n10351, new_n10352, new_n10353, new_n10354,
    new_n10355, new_n10356_1, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372_1, new_n10373, new_n10374, new_n10375, new_n10376,
    new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385_1, new_n10386, new_n10387_1,
    new_n10388_1, new_n10389, new_n10390_1, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404_1, new_n10405_1, new_n10406, new_n10407, new_n10408,
    new_n10409_1, new_n10410, new_n10411_1, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420_1, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432_1, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484_1, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489_1, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505,
    new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514_1, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525_1, new_n10526, new_n10527,
    new_n10528, new_n10529, new_n10530, new_n10531, new_n10532, new_n10533,
    new_n10534, new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540_1, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561_1,
    new_n10562, new_n10563, new_n10564_1, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577_1,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588_1,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593_1,
    new_n10594, new_n10595_1, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611_1, new_n10612, new_n10613, new_n10614_1, new_n10615,
    new_n10616, new_n10617_1, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628_1, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647_1, new_n10648,
    new_n10649, new_n10650_1, new_n10651, new_n10652, new_n10653_1,
    new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671,
    new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683,
    new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689,
    new_n10690, new_n10691, new_n10692_1, new_n10693, new_n10694_1,
    new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700,
    new_n10701_1, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710_1,
    new_n10711, new_n10712_1, new_n10713, new_n10714, new_n10715,
    new_n10716, new_n10717, new_n10718, new_n10720, new_n10721, new_n10722,
    new_n10723, new_n10724, new_n10725, new_n10726, new_n10727, new_n10728,
    new_n10729, new_n10730, new_n10731, new_n10732, new_n10733, new_n10734,
    new_n10735, new_n10736, new_n10737, new_n10738, new_n10739_1,
    new_n10740, new_n10741, new_n10742, new_n10743, new_n10744, new_n10745,
    new_n10746, new_n10747, new_n10748, new_n10749, new_n10750, new_n10751,
    new_n10752, new_n10753, new_n10754, new_n10755, new_n10756_1,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763_1, new_n10764, new_n10765, new_n10766, new_n10767,
    new_n10768, new_n10769, new_n10770, new_n10771, new_n10772, new_n10773,
    new_n10774, new_n10775_1, new_n10776, new_n10777, new_n10778,
    new_n10779, new_n10780_1, new_n10781, new_n10782, new_n10783,
    new_n10784, new_n10785, new_n10786, new_n10787, new_n10788, new_n10789,
    new_n10790, new_n10791, new_n10792_1, new_n10793, new_n10794,
    new_n10795, new_n10796, new_n10797, new_n10798, new_n10799, new_n10800,
    new_n10801, new_n10802, new_n10803, new_n10804, new_n10805, new_n10806,
    new_n10807, new_n10808, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817_1, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834_1, new_n10835,
    new_n10836, new_n10837, new_n10838, new_n10839, new_n10840, new_n10841,
    new_n10842, new_n10843, new_n10844, new_n10845, new_n10846, new_n10847,
    new_n10848, new_n10849, new_n10850, new_n10851_1, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874_1, new_n10875,
    new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881,
    new_n10882, new_n10883, new_n10884, new_n10885, new_n10886, new_n10887,
    new_n10888, new_n10889, new_n10890, new_n10891, new_n10892, new_n10893,
    new_n10894, new_n10895, new_n10896, new_n10897, new_n10898, new_n10899,
    new_n10900, new_n10901, new_n10902, new_n10903, new_n10904, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923,
    new_n10924_1, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943_1, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961_1, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005_1, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011_1, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023_1, new_n11024, new_n11025_1,
    new_n11026, new_n11027, new_n11028, new_n11029, new_n11030, new_n11031,
    new_n11032, new_n11033, new_n11034, new_n11035, new_n11036, new_n11037,
    new_n11038, new_n11039, new_n11040, new_n11041, new_n11042, new_n11043,
    new_n11044_1, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056_1, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063_1, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11072, new_n11073, new_n11075, new_n11076, new_n11077,
    new_n11078_1, new_n11079, new_n11080_1, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094_1, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101_1, new_n11102, new_n11103_1,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109,
    new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115,
    new_n11116, new_n11117, new_n11118, new_n11119, new_n11120_1,
    new_n11121_1, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127_1, new_n11128, new_n11129, new_n11130,
    new_n11131, new_n11132_1, new_n11133, new_n11134_1, new_n11135,
    new_n11136, new_n11137, new_n11138_1, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11146,
    new_n11147, new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153, new_n11154, new_n11155, new_n11156, new_n11157, new_n11158,
    new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164,
    new_n11165, new_n11167, new_n11168, new_n11169, new_n11170, new_n11171,
    new_n11172, new_n11173, new_n11174, new_n11175, new_n11176, new_n11177,
    new_n11178, new_n11179, new_n11180, new_n11181, new_n11182_1,
    new_n11183, new_n11184_1, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192_1,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201_1, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216, new_n11217, new_n11218, new_n11219, new_n11220_1,
    new_n11221, new_n11222, new_n11223_1, new_n11224, new_n11225,
    new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231,
    new_n11232, new_n11233, new_n11234_1, new_n11235, new_n11236,
    new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242,
    new_n11243, new_n11244, new_n11245_1, new_n11246, new_n11247,
    new_n11248, new_n11249, new_n11250, new_n11251, new_n11252, new_n11253,
    new_n11254, new_n11255, new_n11256, new_n11257, new_n11258, new_n11259,
    new_n11260, new_n11261_1, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266_1, new_n11267, new_n11268, new_n11269,
    new_n11270, new_n11271, new_n11272, new_n11273_1, new_n11274,
    new_n11275_1, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290_1,
    new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301,
    new_n11302_1, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313_1, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325_1, new_n11326_1, new_n11327, new_n11328,
    new_n11329, new_n11330_1, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347_1, new_n11348_1, new_n11349, new_n11350,
    new_n11351, new_n11352_1, new_n11353, new_n11354, new_n11355,
    new_n11356_1, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375_1, new_n11376, new_n11377,
    new_n11378, new_n11379_1, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386_1, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391_1, new_n11392,
    new_n11393, new_n11394, new_n11395, new_n11396, new_n11397, new_n11399,
    new_n11400, new_n11401, new_n11402, new_n11403_1, new_n11404,
    new_n11405, new_n11406, new_n11407, new_n11408, new_n11409, new_n11410,
    new_n11411, new_n11412, new_n11413, new_n11414, new_n11415, new_n11416,
    new_n11417, new_n11418, new_n11419_1, new_n11420, new_n11421,
    new_n11422, new_n11423, new_n11424_1, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439_1, new_n11440, new_n11441, new_n11442, new_n11443,
    new_n11444, new_n11445, new_n11446, new_n11447, new_n11448, new_n11449,
    new_n11450, new_n11451, new_n11452, new_n11453, new_n11454, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11463,
    new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470_1, new_n11471, new_n11472_1, new_n11473_1, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479_1,
    new_n11480, new_n11481_1, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486_1, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496_1, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503_1, new_n11504, new_n11505,
    new_n11506_1, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515_1,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537, new_n11538_1,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548_1, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564_1, new_n11565, new_n11566_1,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579_1, new_n11580_1, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589,
    new_n11590, new_n11591_1, new_n11592, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607_1, new_n11608, new_n11609,
    new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615_1, new_n11616, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627, new_n11628, new_n11629, new_n11630_1,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647_1,
    new_n11648, new_n11649, new_n11650, new_n11651, new_n11652, new_n11653,
    new_n11654, new_n11655, new_n11656, new_n11657, new_n11658, new_n11659,
    new_n11660, new_n11661, new_n11662, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667_1, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674_1, new_n11675,
    new_n11676, new_n11677, new_n11678, new_n11679, new_n11680, new_n11681,
    new_n11682_1, new_n11683, new_n11684, new_n11685, new_n11686,
    new_n11687, new_n11688, new_n11689, new_n11690, new_n11691, new_n11692,
    new_n11693, new_n11694, new_n11695, new_n11696, new_n11697, new_n11698,
    new_n11699, new_n11700, new_n11701, new_n11702, new_n11703, new_n11704,
    new_n11705, new_n11706, new_n11707, new_n11708, new_n11709,
    new_n11710_1, new_n11711, new_n11712_1, new_n11713, new_n11714,
    new_n11715, new_n11716, new_n11717, new_n11718, new_n11719, new_n11720,
    new_n11721, new_n11722, new_n11723, new_n11724_1, new_n11725,
    new_n11726, new_n11727, new_n11728, new_n11729, new_n11730, new_n11731,
    new_n11732, new_n11733, new_n11734, new_n11735, new_n11736_1,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741_1,
    new_n11742, new_n11743, new_n11744, new_n11745, new_n11746, new_n11747,
    new_n11748, new_n11749_1, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11756, new_n11757, new_n11758, new_n11759,
    new_n11760, new_n11761, new_n11762, new_n11763, new_n11764, new_n11765,
    new_n11766, new_n11767, new_n11768, new_n11769, new_n11770_1,
    new_n11771_1, new_n11772, new_n11773, new_n11774, new_n11775_1,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780, new_n11781,
    new_n11782, new_n11783, new_n11784, new_n11785, new_n11786, new_n11787,
    new_n11788, new_n11789, new_n11790, new_n11791, new_n11792, new_n11793,
    new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799,
    new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805,
    new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811,
    new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818_1, new_n11819, new_n11820, new_n11821, new_n11822,
    new_n11823, new_n11824, new_n11825, new_n11826, new_n11827, new_n11828,
    new_n11829, new_n11830, new_n11831, new_n11832, new_n11833, new_n11834,
    new_n11835, new_n11836, new_n11837_1, new_n11838, new_n11839,
    new_n11840, new_n11841_1, new_n11842_1, new_n11843_1, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897,
    new_n11898_1, new_n11899, new_n11900, new_n11901, new_n11902,
    new_n11903, new_n11904, new_n11905_1, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926_1, new_n11927, new_n11928, new_n11929, new_n11930,
    new_n11931, new_n11932, new_n11933, new_n11934, new_n11935, new_n11936,
    new_n11937, new_n11938, new_n11939, new_n11940, new_n11941, new_n11942,
    new_n11943, new_n11944, new_n11945, new_n11946, new_n11947, new_n11948,
    new_n11949, new_n11950, new_n11951, new_n11952, new_n11953, new_n11954,
    new_n11955, new_n11956, new_n11957, new_n11958, new_n11962, new_n11963,
    new_n11964, new_n11965_1, new_n11966, new_n11967, new_n11968,
    new_n11969, new_n11970, new_n11971, new_n11972, new_n11976, new_n11977,
    new_n11978, new_n11979, new_n11980_1, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999,
    new_n12000_1, new_n12001, new_n12002, new_n12003_1, new_n12006,
    new_n12007, new_n12008, new_n12009, new_n12010, new_n12011_1,
    new_n12012, new_n12013, new_n12014, new_n12015, new_n12016, new_n12017,
    new_n12018, new_n12019, new_n12020, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044, new_n12045, new_n12046, new_n12047,
    new_n12048, new_n12049, new_n12050, new_n12051, new_n12052, new_n12053,
    new_n12054, new_n12055, new_n12056, new_n12057, new_n12058, new_n12059,
    new_n12060, new_n12061, new_n12062, new_n12063, new_n12064, new_n12065,
    new_n12066, new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072_1, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12108, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113_1, new_n12114, new_n12115, new_n12116, new_n12117,
    new_n12118, new_n12119, new_n12120, new_n12121_1, new_n12122,
    new_n12123, new_n12124, new_n12125, new_n12126, new_n12127, new_n12128,
    new_n12129, new_n12130, new_n12131_1, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145,
    new_n12146_1, new_n12147, new_n12148, new_n12149, new_n12150,
    new_n12151, new_n12152_1, new_n12153_1, new_n12154, new_n12155,
    new_n12156, new_n12157_1, new_n12158_1, new_n12159, new_n12160,
    new_n12161_1, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166, new_n12167, new_n12168, new_n12169, new_n12170, new_n12171,
    new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177,
    new_n12178, new_n12179_1, new_n12180, new_n12181, new_n12182,
    new_n12183, new_n12184, new_n12185, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192_1, new_n12193, new_n12194, new_n12195,
    new_n12196, new_n12197, new_n12198, new_n12199, new_n12200, new_n12201,
    new_n12202, new_n12203, new_n12204, new_n12205, new_n12206, new_n12207,
    new_n12208, new_n12209_1, new_n12210, new_n12211, new_n12212,
    new_n12213, new_n12214, new_n12215, new_n12216, new_n12217, new_n12218,
    new_n12219, new_n12220, new_n12221, new_n12222, new_n12223_1,
    new_n12224, new_n12225_1, new_n12226, new_n12227, new_n12228_1,
    new_n12229, new_n12230, new_n12231, new_n12232, new_n12233, new_n12234,
    new_n12235_1, new_n12236, new_n12237, new_n12238, new_n12239,
    new_n12240, new_n12241, new_n12242, new_n12243, new_n12244, new_n12245,
    new_n12246, new_n12247, new_n12248, new_n12249, new_n12250, new_n12251,
    new_n12252, new_n12253, new_n12254, new_n12255, new_n12256, new_n12257,
    new_n12258, new_n12259, new_n12260, new_n12261, new_n12262, new_n12263,
    new_n12264, new_n12265, new_n12266, new_n12267, new_n12268, new_n12269,
    new_n12270, new_n12271, new_n12272, new_n12273, new_n12274, new_n12275,
    new_n12276, new_n12277, new_n12278, new_n12279, new_n12280, new_n12281,
    new_n12282, new_n12283, new_n12284, new_n12285, new_n12286, new_n12287,
    new_n12288, new_n12289, new_n12290, new_n12291, new_n12292, new_n12293,
    new_n12294, new_n12295, new_n12296, new_n12297, new_n12298, new_n12299,
    new_n12300, new_n12301, new_n12302_1, new_n12303, new_n12304_1,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315_1,
    new_n12316, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324_1, new_n12325_1, new_n12326, new_n12327,
    new_n12328, new_n12329_1, new_n12330_1, new_n12331, new_n12332,
    new_n12333, new_n12334, new_n12335, new_n12336, new_n12337, new_n12338,
    new_n12339, new_n12340, new_n12341_1, new_n12342, new_n12343,
    new_n12344, new_n12345, new_n12346_1, new_n12347, new_n12348,
    new_n12349_1, new_n12350, new_n12351, new_n12352, new_n12353,
    new_n12354, new_n12355, new_n12356, new_n12357, new_n12358, new_n12359,
    new_n12360, new_n12361, new_n12362, new_n12363, new_n12364_1,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370,
    new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380_1, new_n12381,
    new_n12382, new_n12383_1, new_n12384_1, new_n12385, new_n12386,
    new_n12387, new_n12388, new_n12389, new_n12390, new_n12391, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397_1,
    new_n12398_1, new_n12399, new_n12400, new_n12401, new_n12402,
    new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408_1, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444, new_n12445, new_n12446_1, new_n12447, new_n12448,
    new_n12449_1, new_n12450, new_n12451, new_n12452, new_n12453,
    new_n12454, new_n12455, new_n12456, new_n12457, new_n12458, new_n12459,
    new_n12460, new_n12461_1, new_n12462_1, new_n12463, new_n12464,
    new_n12468, new_n12469_1, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490,
    new_n12491, new_n12492, new_n12493, new_n12494, new_n12495_1,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506,
    new_n12507_1, new_n12508, new_n12509, new_n12510, new_n12511,
    new_n12512, new_n12513, new_n12514, new_n12515_1, new_n12516_1,
    new_n12517, new_n12518, new_n12519, new_n12520, new_n12521, new_n12522,
    new_n12523, new_n12524, new_n12525, new_n12526, new_n12527, new_n12528,
    new_n12529, new_n12530, new_n12531, new_n12532, new_n12533, new_n12534,
    new_n12535, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540_1, new_n12541, new_n12542, new_n12543, new_n12546_1,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552_1, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562_1, new_n12563, new_n12564, new_n12565, new_n12566_1,
    new_n12567, new_n12568, new_n12569_1, new_n12570, new_n12571,
    new_n12572, new_n12573, new_n12574, new_n12575, new_n12576, new_n12577,
    new_n12578, new_n12579, new_n12580, new_n12581, new_n12582, new_n12583,
    new_n12584, new_n12585, new_n12586, new_n12587_1, new_n12588,
    new_n12589, new_n12590, new_n12591, new_n12592, new_n12593_1,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607_1, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620_1, new_n12621_1,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626_1,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649,
    new_n12650_1, new_n12651, new_n12652, new_n12653, new_n12654_1,
    new_n12655, new_n12656, new_n12657_1, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665_1, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670_1, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702_1, new_n12703,
    new_n12704, new_n12705, new_n12706, new_n12707_1, new_n12708,
    new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714,
    new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725_1,
    new_n12726, new_n12727_1, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12740_1, new_n12741,
    new_n12742_1, new_n12743, new_n12744, new_n12745, new_n12746_1,
    new_n12747, new_n12748, new_n12749, new_n12750, new_n12751, new_n12752,
    new_n12753, new_n12754, new_n12755, new_n12756_1, new_n12757,
    new_n12758, new_n12759, new_n12760, new_n12761, new_n12762, new_n12763,
    new_n12764, new_n12765, new_n12766, new_n12767, new_n12768, new_n12769,
    new_n12770, new_n12771, new_n12772, new_n12773, new_n12774, new_n12775,
    new_n12776, new_n12777, new_n12778, new_n12779, new_n12782,
    new_n12783_1, new_n12784, new_n12785, new_n12786, new_n12787,
    new_n12788, new_n12789, new_n12790, new_n12791, new_n12792, new_n12793,
    new_n12794, new_n12795, new_n12796, new_n12797, new_n12798, new_n12799,
    new_n12800, new_n12801_1, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811_1, new_n12812_1, new_n12813, new_n12814, new_n12815,
    new_n12816_1, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821_1, new_n12822, new_n12824, new_n12825, new_n12826,
    new_n12827, new_n12828, new_n12829, new_n12830, new_n12831, new_n12832,
    new_n12833, new_n12834, new_n12835, new_n12836, new_n12837, new_n12838,
    new_n12839, new_n12840, new_n12841, new_n12842, new_n12843_1,
    new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849,
    new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855,
    new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861_1, new_n12862, new_n12863, new_n12864_1, new_n12865_1,
    new_n12866, new_n12867, new_n12868, new_n12869, new_n12870_1,
    new_n12871_1, new_n12872, new_n12873_1, new_n12874, new_n12875_1,
    new_n12876, new_n12877, new_n12878, new_n12879, new_n12880, new_n12881,
    new_n12882, new_n12883, new_n12884, new_n12885, new_n12886, new_n12887,
    new_n12888, new_n12889, new_n12890, new_n12891, new_n12892_1,
    new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898,
    new_n12899, new_n12900_1, new_n12901, new_n12902, new_n12903,
    new_n12904_1, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917_1, new_n12918, new_n12919,
    new_n12920, new_n12921, new_n12922, new_n12923, new_n12924, new_n12925,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941_1, new_n12942_1,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956_1, new_n12957, new_n12958, new_n12959,
    new_n12960, new_n12961, new_n12962, new_n12963, new_n12964, new_n12965,
    new_n12966, new_n12967, new_n12968, new_n12969, new_n12970, new_n12971,
    new_n12972, new_n12973, new_n12974, new_n12975, new_n12976, new_n12977,
    new_n12978_1, new_n12979, new_n12980_1, new_n12981, new_n12982,
    new_n12983, new_n12984, new_n12985_1, new_n12986, new_n12987_1,
    new_n12988, new_n12989, new_n12990, new_n12991, new_n12992_1,
    new_n12993, new_n12994, new_n12995, new_n12996, new_n12997, new_n12998,
    new_n12999, new_n13000, new_n13001, new_n13002, new_n13003, new_n13004,
    new_n13005_1, new_n13006, new_n13007, new_n13008, new_n13009,
    new_n13010, new_n13011, new_n13012, new_n13013, new_n13014, new_n13015,
    new_n13016, new_n13017, new_n13018, new_n13019, new_n13020, new_n13021,
    new_n13022, new_n13023, new_n13024, new_n13025, new_n13026_1,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043_1,
    new_n13044_1, new_n13045, new_n13046, new_n13047, new_n13048_1,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053,
    new_n13054_1, new_n13055, new_n13056, new_n13057, new_n13058,
    new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064,
    new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13072, new_n13073, new_n13074_1, new_n13075,
    new_n13076, new_n13077, new_n13078, new_n13079, new_n13080, new_n13081,
    new_n13082_1, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096_1, new_n13097,
    new_n13098, new_n13099, new_n13100, new_n13101, new_n13102, new_n13103,
    new_n13104, new_n13105, new_n13106, new_n13107, new_n13108, new_n13109,
    new_n13110_1, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116_1, new_n13117, new_n13118, new_n13119,
    new_n13120, new_n13121, new_n13122_1, new_n13123, new_n13124,
    new_n13125, new_n13126, new_n13127, new_n13128, new_n13129, new_n13130,
    new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137_1, new_n13138, new_n13139, new_n13140, new_n13141_1,
    new_n13142, new_n13143, new_n13144_1, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13151, new_n13152, new_n13153, new_n13154,
    new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160,
    new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166,
    new_n13167, new_n13168_1, new_n13169, new_n13170, new_n13171,
    new_n13172, new_n13173, new_n13174, new_n13175, new_n13176, new_n13177,
    new_n13178, new_n13179, new_n13180, new_n13181, new_n13182, new_n13183,
    new_n13184, new_n13185, new_n13186, new_n13187, new_n13188, new_n13189,
    new_n13190_1, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198_1, new_n13199_1,
    new_n13200, new_n13201, new_n13202, new_n13203, new_n13204_1,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209_1,
    new_n13210, new_n13211, new_n13212, new_n13213, new_n13214, new_n13215,
    new_n13216, new_n13217, new_n13218, new_n13219, new_n13220, new_n13225,
    new_n13226, new_n13227, new_n13228, new_n13229, new_n13230, new_n13231,
    new_n13232, new_n13233, new_n13234, new_n13235, new_n13236, new_n13237,
    new_n13238, new_n13239, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252,
    new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258,
    new_n13259, new_n13260, new_n13261, new_n13262, new_n13263_1,
    new_n13264, new_n13265, new_n13269, new_n13270_1, new_n13271,
    new_n13272, new_n13273_1, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285_1, new_n13286, new_n13287,
    new_n13288, new_n13289, new_n13290, new_n13291, new_n13292, new_n13293,
    new_n13294, new_n13295, new_n13296, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312,
    new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318,
    new_n13319_1, new_n13320, new_n13321, new_n13322, new_n13323,
    new_n13324, new_n13325, new_n13326, new_n13327, new_n13328, new_n13329,
    new_n13330, new_n13334, new_n13335, new_n13336, new_n13337,
    new_n13338_1, new_n13339, new_n13340, new_n13341, new_n13342,
    new_n13343, new_n13344, new_n13345, new_n13346, new_n13347, new_n13348,
    new_n13349, new_n13350, new_n13351, new_n13352, new_n13353, new_n13354,
    new_n13355, new_n13356, new_n13357, new_n13358, new_n13359, new_n13360,
    new_n13361, new_n13362, new_n13363, new_n13364, new_n13365, new_n13366,
    new_n13367_1, new_n13368, new_n13369, new_n13370, new_n13371,
    new_n13372, new_n13373, new_n13374, new_n13375, new_n13376, new_n13379,
    new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385,
    new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391,
    new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397,
    new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407_1, new_n13408,
    new_n13409_1, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419_1, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424_1, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453_1, new_n13454, new_n13455, new_n13456_1, new_n13457_1,
    new_n13458, new_n13459, new_n13460_1, new_n13461, new_n13462,
    new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468,
    new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474,
    new_n13475, new_n13476, new_n13477_1, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13483, new_n13484_1,
    new_n13485, new_n13486_1, new_n13487_1, new_n13488, new_n13489,
    new_n13490_1, new_n13491, new_n13492, new_n13493, new_n13494_1,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13500_1,
    new_n13501_1, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506_1, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534,
    new_n13535, new_n13536, new_n13537, new_n13538, new_n13539, new_n13540,
    new_n13541, new_n13542, new_n13543, new_n13544, new_n13545, new_n13546,
    new_n13547, new_n13548_1, new_n13549_1, new_n13550, new_n13551_1,
    new_n13552, new_n13553, new_n13554, new_n13555, new_n13556, new_n13557,
    new_n13558, new_n13559, new_n13560, new_n13561, new_n13562, new_n13563,
    new_n13564, new_n13565, new_n13566, new_n13567, new_n13568, new_n13569,
    new_n13570, new_n13571, new_n13572, new_n13573, new_n13574, new_n13575,
    new_n13576, new_n13577, new_n13578, new_n13579, new_n13580, new_n13581,
    new_n13582, new_n13583, new_n13584, new_n13585, new_n13586, new_n13587,
    new_n13588, new_n13589, new_n13590, new_n13591, new_n13592, new_n13593,
    new_n13594, new_n13595, new_n13596, new_n13597, new_n13598, new_n13599,
    new_n13600, new_n13601, new_n13602_1, new_n13603, new_n13604,
    new_n13605, new_n13606, new_n13607, new_n13608, new_n13609, new_n13610,
    new_n13611, new_n13612, new_n13613, new_n13615, new_n13616, new_n13617,
    new_n13618, new_n13619, new_n13620, new_n13621, new_n13622, new_n13623,
    new_n13624, new_n13625, new_n13626_1, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634,
    new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640,
    new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646,
    new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652,
    new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658,
    new_n13659, new_n13660, new_n13661, new_n13662, new_n13665, new_n13666,
    new_n13667, new_n13668_1, new_n13669, new_n13670, new_n13671,
    new_n13672, new_n13673, new_n13675, new_n13676, new_n13677_1,
    new_n13678, new_n13679, new_n13680, new_n13681, new_n13682,
    new_n13683_1, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708_1, new_n13709, new_n13710_1,
    new_n13711, new_n13712, new_n13713, new_n13714_1, new_n13715,
    new_n13716, new_n13717, new_n13718, new_n13719_1, new_n13720,
    new_n13721, new_n13722_1, new_n13723, new_n13724, new_n13725,
    new_n13726, new_n13727, new_n13728, new_n13729, new_n13730, new_n13731,
    new_n13732, new_n13733, new_n13734, new_n13735, new_n13736, new_n13737,
    new_n13738, new_n13739, new_n13740, new_n13741, new_n13742, new_n13743,
    new_n13744, new_n13745, new_n13746, new_n13747, new_n13748, new_n13749,
    new_n13750, new_n13751, new_n13752, new_n13753, new_n13754_1,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764_1, new_n13765,
    new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771,
    new_n13772, new_n13773, new_n13774, new_n13775_1, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781_1,
    new_n13782, new_n13783_1, new_n13784, new_n13785, new_n13786,
    new_n13787, new_n13788, new_n13789, new_n13790, new_n13791, new_n13792,
    new_n13793, new_n13794, new_n13795, new_n13796, new_n13797,
    new_n13798_1, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835_1, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13842, new_n13843, new_n13844, new_n13845,
    new_n13846, new_n13847, new_n13848, new_n13849, new_n13850_1,
    new_n13851_1, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912_1, new_n13913, new_n13914_1,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922_1, new_n13923_1, new_n13924, new_n13925,
    new_n13926, new_n13927, new_n13928, new_n13929, new_n13931, new_n13932,
    new_n13933, new_n13934, new_n13935, new_n13936, new_n13937, new_n13940,
    new_n13941, new_n13942, new_n13943, new_n13944, new_n13945, new_n13946,
    new_n13947, new_n13948, new_n13949, new_n13950, new_n13951_1,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004_1,
    new_n14005, new_n14006, new_n14007, new_n14008, new_n14009, new_n14010,
    new_n14011, new_n14012, new_n14013, new_n14014, new_n14015, new_n14016,
    new_n14017, new_n14018, new_n14019, new_n14020, new_n14021, new_n14022,
    new_n14023, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036_1, new_n14037, new_n14038, new_n14039, new_n14040,
    new_n14041, new_n14042, new_n14043, new_n14044, new_n14045, new_n14046,
    new_n14047, new_n14048, new_n14049, new_n14050, new_n14051, new_n14052,
    new_n14053, new_n14054, new_n14055, new_n14056, new_n14057, new_n14058,
    new_n14059_1, new_n14060, new_n14061, new_n14062, new_n14063,
    new_n14064, new_n14065, new_n14066, new_n14067, new_n14068, new_n14069,
    new_n14070, new_n14071_1, new_n14072, new_n14073, new_n14074,
    new_n14075, new_n14076, new_n14077, new_n14078, new_n14079, new_n14080,
    new_n14081_1, new_n14082, new_n14083, new_n14084, new_n14085,
    new_n14086, new_n14087, new_n14088, new_n14089, new_n14090_1,
    new_n14091, new_n14092, new_n14093, new_n14094, new_n14095_1,
    new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101,
    new_n14102, new_n14103, new_n14104, new_n14105, new_n14106,
    new_n14107_1, new_n14108, new_n14109, new_n14110, new_n14111,
    new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117,
    new_n14118, new_n14119, new_n14120, new_n14121_1, new_n14122,
    new_n14123, new_n14124, new_n14125, new_n14126_1, new_n14127,
    new_n14128, new_n14129, new_n14130_1, new_n14131, new_n14132,
    new_n14133, new_n14134, new_n14135, new_n14136_1, new_n14137,
    new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143,
    new_n14144, new_n14145, new_n14146, new_n14147_1, new_n14148_1,
    new_n14149, new_n14152, new_n14153, new_n14154, new_n14155, new_n14156,
    new_n14157, new_n14158, new_n14159, new_n14160, new_n14161, new_n14162,
    new_n14163, new_n14164, new_n14165, new_n14166, new_n14167, new_n14168,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173,
    new_n14174_1, new_n14175, new_n14176, new_n14177, new_n14178,
    new_n14179, new_n14180, new_n14181, new_n14182, new_n14183, new_n14184,
    new_n14185, new_n14186, new_n14187, new_n14188, new_n14189,
    new_n14190_1, new_n14191, new_n14192, new_n14193, new_n14194,
    new_n14195, new_n14196, new_n14197, new_n14198, new_n14199, new_n14200,
    new_n14201, new_n14202, new_n14205, new_n14206, new_n14207, new_n14208,
    new_n14209, new_n14210, new_n14211_1, new_n14212, new_n14213,
    new_n14214, new_n14215, new_n14216, new_n14217, new_n14218, new_n14219,
    new_n14220, new_n14221, new_n14222_1, new_n14223, new_n14224,
    new_n14225, new_n14226, new_n14227, new_n14228, new_n14229,
    new_n14230_1, new_n14231, new_n14232, new_n14233, new_n14234,
    new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267_1, new_n14268, new_n14269,
    new_n14270, new_n14271_1, new_n14272, new_n14273, new_n14274,
    new_n14275_1, new_n14276, new_n14277_1, new_n14278, new_n14279,
    new_n14280, new_n14281, new_n14282, new_n14283, new_n14284, new_n14285,
    new_n14286, new_n14287, new_n14288, new_n14289, new_n14290, new_n14291,
    new_n14292, new_n14293, new_n14294_1, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310_1, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14320, new_n14321, new_n14322, new_n14323_1, new_n14324,
    new_n14325, new_n14326_1, new_n14327, new_n14328, new_n14329,
    new_n14330, new_n14331, new_n14332, new_n14333, new_n14334, new_n14335,
    new_n14336, new_n14337, new_n14338, new_n14339, new_n14340, new_n14341,
    new_n14342_1, new_n14343, new_n14344, new_n14345_1, new_n14346,
    new_n14347, new_n14348, new_n14349, new_n14350, new_n14351, new_n14352,
    new_n14353_1, new_n14355, new_n14356, new_n14357, new_n14358,
    new_n14359, new_n14360, new_n14361, new_n14362, new_n14363,
    new_n14364_1, new_n14365, new_n14366, new_n14367, new_n14368,
    new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374,
    new_n14375_1, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14384, new_n14385, new_n14386,
    new_n14387, new_n14388, new_n14389, new_n14390, new_n14391, new_n14392,
    new_n14393, new_n14394, new_n14395, new_n14396, new_n14397, new_n14398,
    new_n14399, new_n14400, new_n14401, new_n14402, new_n14403, new_n14404,
    new_n14405, new_n14406, new_n14407, new_n14408, new_n14409, new_n14410,
    new_n14411, new_n14412_1, new_n14413, new_n14414_1, new_n14415,
    new_n14416, new_n14417, new_n14418, new_n14419, new_n14420, new_n14421,
    new_n14422, new_n14423, new_n14424, new_n14425, new_n14426, new_n14427,
    new_n14428, new_n14429, new_n14430, new_n14431, new_n14432, new_n14433,
    new_n14434, new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440_1, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457_1, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464_1, new_n14465, new_n14466,
    new_n14467, new_n14468, new_n14469, new_n14470, new_n14471_1,
    new_n14472, new_n14473, new_n14474, new_n14475_1, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510_1, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540,
    new_n14541_1, new_n14542, new_n14543, new_n14544, new_n14545,
    new_n14546_1, new_n14547_1, new_n14548, new_n14549, new_n14550,
    new_n14551, new_n14552, new_n14553, new_n14554, new_n14555, new_n14556,
    new_n14557, new_n14558, new_n14559, new_n14560, new_n14561, new_n14562,
    new_n14563, new_n14564, new_n14565, new_n14566, new_n14567, new_n14568,
    new_n14569, new_n14570_1, new_n14571, new_n14572, new_n14573,
    new_n14574, new_n14575_1, new_n14576_1, new_n14577, new_n14578,
    new_n14579, new_n14580, new_n14581, new_n14582, new_n14583, new_n14584,
    new_n14585, new_n14586, new_n14587, new_n14588, new_n14589, new_n14590,
    new_n14591, new_n14592, new_n14593_1, new_n14594, new_n14595,
    new_n14596, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602,
    new_n14603_1, new_n14604, new_n14605, new_n14606, new_n14607,
    new_n14608, new_n14609, new_n14610, new_n14611, new_n14612, new_n14613,
    new_n14614, new_n14615, new_n14616, new_n14617, new_n14618, new_n14619,
    new_n14620, new_n14621, new_n14622, new_n14623, new_n14624, new_n14625,
    new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631,
    new_n14632, new_n14633_1, new_n14634, new_n14635, new_n14636_1,
    new_n14637, new_n14638, new_n14639, new_n14640, new_n14641, new_n14642,
    new_n14643, new_n14644, new_n14645, new_n14646, new_n14647, new_n14648,
    new_n14649, new_n14650, new_n14651, new_n14652, new_n14653, new_n14654,
    new_n14655, new_n14656, new_n14657, new_n14658, new_n14659, new_n14660,
    new_n14661, new_n14662, new_n14663, new_n14664, new_n14665, new_n14666,
    new_n14667, new_n14668, new_n14669, new_n14670, new_n14671, new_n14672,
    new_n14673, new_n14674, new_n14675, new_n14676, new_n14677, new_n14678,
    new_n14679, new_n14680_1, new_n14681, new_n14682, new_n14683,
    new_n14684_1, new_n14685, new_n14686, new_n14687, new_n14688,
    new_n14689, new_n14690, new_n14691, new_n14692_1, new_n14693,
    new_n14694, new_n14695, new_n14696, new_n14697, new_n14698, new_n14699,
    new_n14700, new_n14701_1, new_n14702_1, new_n14703, new_n14704_1,
    new_n14705, new_n14706, new_n14707, new_n14708, new_n14709, new_n14710,
    new_n14711, new_n14712, new_n14713, new_n14714, new_n14715, new_n14716,
    new_n14717, new_n14718, new_n14719, new_n14720, new_n14721, new_n14722,
    new_n14723, new_n14724, new_n14725, new_n14726, new_n14727, new_n14728,
    new_n14729, new_n14730, new_n14731, new_n14732, new_n14733,
    new_n14734_1, new_n14735, new_n14736, new_n14737, new_n14738,
    new_n14739, new_n14740, new_n14741, new_n14742, new_n14743, new_n14744,
    new_n14745, new_n14746_1, new_n14747, new_n14748, new_n14749,
    new_n14750, new_n14751, new_n14752, new_n14753, new_n14754, new_n14756,
    new_n14757, new_n14758, new_n14759, new_n14760, new_n14761, new_n14762,
    new_n14763_1, new_n14764, new_n14765, new_n14766, new_n14767,
    new_n14768, new_n14769, new_n14770, new_n14771, new_n14772_1,
    new_n14773, new_n14774, new_n14775, new_n14776, new_n14777, new_n14778,
    new_n14779, new_n14780, new_n14781, new_n14782, new_n14783, new_n14784,
    new_n14785, new_n14786, new_n14787, new_n14788, new_n14789,
    new_n14790_1, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800,
    new_n14801_1, new_n14802, new_n14803, new_n14804, new_n14805,
    new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819_1, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826_1, new_n14827_1,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839_1, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14848,
    new_n14849_1, new_n14850, new_n14851, new_n14852, new_n14853,
    new_n14854, new_n14855, new_n14856, new_n14857, new_n14858, new_n14859,
    new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865,
    new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871,
    new_n14872, new_n14873, new_n14874, new_n14875, new_n14876, new_n14877,
    new_n14878, new_n14879, new_n14880, new_n14881, new_n14882, new_n14883,
    new_n14884, new_n14885, new_n14886, new_n14887, new_n14888, new_n14889,
    new_n14890, new_n14891_1, new_n14892, new_n14893, new_n14894,
    new_n14895, new_n14896, new_n14897, new_n14898, new_n14900, new_n14901,
    new_n14902, new_n14903, new_n14904, new_n14905, new_n14906, new_n14907,
    new_n14908, new_n14909, new_n14910, new_n14911, new_n14912, new_n14913,
    new_n14914, new_n14915, new_n14916, new_n14917, new_n14918, new_n14919,
    new_n14920, new_n14921, new_n14922, new_n14923, new_n14924, new_n14925,
    new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931_1, new_n14932, new_n14933, new_n14934, new_n14935,
    new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941,
    new_n14942, new_n14943, new_n14944_1, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954_1, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977_1, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986,
    new_n14987, new_n14988, new_n14989_1, new_n14990, new_n14991,
    new_n14992, new_n14993, new_n14994, new_n14995, new_n14996, new_n14997,
    new_n14998, new_n14999, new_n15000, new_n15001, new_n15002_1,
    new_n15003, new_n15004_1, new_n15005, new_n15006, new_n15007,
    new_n15008, new_n15009, new_n15010, new_n15011_1, new_n15012,
    new_n15013, new_n15014, new_n15015, new_n15016, new_n15017,
    new_n15019_1, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031_1, new_n15032, new_n15033_1, new_n15034,
    new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040,
    new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046,
    new_n15047, new_n15048, new_n15049, new_n15050, new_n15051,
    new_n15052_1, new_n15053_1, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077_1, new_n15078, new_n15079,
    new_n15080, new_n15081, new_n15082_1, new_n15083, new_n15084,
    new_n15085, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092,
    new_n15093, new_n15094_1, new_n15095, new_n15096, new_n15097,
    new_n15098, new_n15099, new_n15100, new_n15101, new_n15102, new_n15103,
    new_n15104, new_n15105, new_n15106, new_n15107, new_n15108, new_n15109,
    new_n15110, new_n15111, new_n15112, new_n15113, new_n15114, new_n15115,
    new_n15116, new_n15117, new_n15118_1, new_n15119, new_n15120,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128_1, new_n15129, new_n15130, new_n15131,
    new_n15132, new_n15133, new_n15134, new_n15135, new_n15136, new_n15137,
    new_n15138, new_n15139_1, new_n15140, new_n15141, new_n15142,
    new_n15143, new_n15144, new_n15145_1, new_n15146_1, new_n15147,
    new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153,
    new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159,
    new_n15160, new_n15161, new_n15162, new_n15163, new_n15164,
    new_n15165_1, new_n15166, new_n15167_1, new_n15168, new_n15169,
    new_n15170, new_n15171, new_n15172, new_n15173, new_n15174, new_n15175,
    new_n15176_1, new_n15177, new_n15178, new_n15179, new_n15180_1,
    new_n15181, new_n15182_1, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205_1, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230_1, new_n15231,
    new_n15232, new_n15233, new_n15235, new_n15236, new_n15237, new_n15238,
    new_n15239, new_n15240, new_n15241_1, new_n15242, new_n15243,
    new_n15244, new_n15245, new_n15246, new_n15247, new_n15248, new_n15249,
    new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255_1, new_n15256, new_n15257, new_n15258_1, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271_1, new_n15272, new_n15273, new_n15274, new_n15275_1,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289_1, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300_1, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307_1, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327_1, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332_1, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342,
    new_n15343, new_n15344, new_n15345_1, new_n15346, new_n15347,
    new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353_1, new_n15359, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15367, new_n15368, new_n15369, new_n15370, new_n15371,
    new_n15372, new_n15373, new_n15374, new_n15375, new_n15376, new_n15377,
    new_n15378_1, new_n15379, new_n15380, new_n15381, new_n15382_1,
    new_n15383, new_n15384, new_n15385, new_n15386, new_n15387, new_n15388,
    new_n15389, new_n15390, new_n15391, new_n15392, new_n15393, new_n15394,
    new_n15395, new_n15398, new_n15399, new_n15400, new_n15401, new_n15402,
    new_n15403, new_n15404, new_n15405, new_n15406, new_n15407_1,
    new_n15408, new_n15409, new_n15410, new_n15411, new_n15412, new_n15413,
    new_n15414, new_n15415, new_n15416, new_n15417, new_n15418, new_n15419,
    new_n15420, new_n15421, new_n15422, new_n15423, new_n15424_1,
    new_n15425, new_n15426, new_n15427, new_n15428_1, new_n15429,
    new_n15430, new_n15431, new_n15432, new_n15433, new_n15434,
    new_n15435_1, new_n15436, new_n15437, new_n15438_1, new_n15439,
    new_n15440, new_n15441, new_n15442, new_n15443, new_n15444, new_n15445,
    new_n15446, new_n15447, new_n15448, new_n15449, new_n15450, new_n15451,
    new_n15452, new_n15453, new_n15454, new_n15455, new_n15456, new_n15457,
    new_n15458, new_n15459, new_n15460, new_n15461, new_n15462, new_n15463,
    new_n15464, new_n15465_1, new_n15466, new_n15467_1, new_n15468,
    new_n15469, new_n15470_1, new_n15471, new_n15472, new_n15478,
    new_n15479, new_n15480, new_n15481_1, new_n15482, new_n15483,
    new_n15484, new_n15485, new_n15486, new_n15487, new_n15488, new_n15489,
    new_n15490_1, new_n15491, new_n15492, new_n15493, new_n15494,
    new_n15495, new_n15496_1, new_n15497, new_n15498, new_n15499,
    new_n15500, new_n15501_1, new_n15502, new_n15503, new_n15504,
    new_n15505, new_n15506_1, new_n15507, new_n15508_1, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527,
    new_n15528, new_n15529, new_n15530, new_n15531, new_n15532, new_n15533,
    new_n15534, new_n15535, new_n15536, new_n15537, new_n15538,
    new_n15539_1, new_n15540, new_n15541, new_n15542, new_n15543,
    new_n15544, new_n15545, new_n15546_1, new_n15547, new_n15548,
    new_n15549, new_n15550, new_n15551, new_n15552, new_n15553, new_n15554,
    new_n15555_1, new_n15556, new_n15557, new_n15558_1, new_n15559_1,
    new_n15560, new_n15561, new_n15562, new_n15563, new_n15564, new_n15565,
    new_n15566, new_n15567, new_n15568, new_n15569, new_n15570_1,
    new_n15571, new_n15572, new_n15573_1, new_n15574, new_n15575,
    new_n15576, new_n15577, new_n15578, new_n15579, new_n15580, new_n15581,
    new_n15582, new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588_1, new_n15589, new_n15590_1, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598_1, new_n15599, new_n15600, new_n15601, new_n15602_1,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613, new_n15616,
    new_n15617, new_n15618, new_n15619, new_n15620, new_n15621, new_n15622,
    new_n15623, new_n15624, new_n15625, new_n15626, new_n15627, new_n15628,
    new_n15629, new_n15630, new_n15631, new_n15632, new_n15633, new_n15634,
    new_n15635, new_n15636_1, new_n15637, new_n15638, new_n15639,
    new_n15640, new_n15641, new_n15642, new_n15643, new_n15644, new_n15645,
    new_n15646, new_n15647, new_n15648, new_n15649, new_n15650, new_n15651,
    new_n15652_1, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661,
    new_n15662_1, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15680, new_n15681, new_n15682, new_n15683, new_n15684, new_n15685,
    new_n15686, new_n15687, new_n15688, new_n15689, new_n15690, new_n15691,
    new_n15692, new_n15693, new_n15694, new_n15695, new_n15696, new_n15697,
    new_n15698, new_n15699, new_n15700, new_n15701, new_n15702, new_n15703,
    new_n15704, new_n15705, new_n15706, new_n15707, new_n15708, new_n15709,
    new_n15710, new_n15713, new_n15714, new_n15715, new_n15716_1,
    new_n15717, new_n15718, new_n15719, new_n15720, new_n15721, new_n15722,
    new_n15723, new_n15724, new_n15725, new_n15726, new_n15727, new_n15728,
    new_n15729, new_n15730, new_n15731, new_n15732, new_n15733, new_n15734,
    new_n15735, new_n15736, new_n15737, new_n15738, new_n15739, new_n15740,
    new_n15741, new_n15742, new_n15743_1, new_n15744, new_n15745,
    new_n15746, new_n15747, new_n15748, new_n15749_1, new_n15750,
    new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756,
    new_n15758, new_n15759, new_n15760, new_n15761_1, new_n15762_1,
    new_n15763, new_n15764, new_n15765, new_n15766_1, new_n15767,
    new_n15768, new_n15769, new_n15770, new_n15771, new_n15772, new_n15773,
    new_n15774, new_n15775, new_n15776, new_n15777, new_n15778, new_n15779,
    new_n15780_1, new_n15781, new_n15782, new_n15783, new_n15784,
    new_n15785, new_n15786, new_n15787, new_n15788, new_n15789, new_n15790,
    new_n15791, new_n15792, new_n15793_1, new_n15794, new_n15795,
    new_n15796, new_n15797, new_n15799, new_n15800, new_n15801, new_n15802,
    new_n15803, new_n15804, new_n15805, new_n15806, new_n15807, new_n15808,
    new_n15809, new_n15810, new_n15811, new_n15812_1, new_n15813,
    new_n15814, new_n15815_1, new_n15816_1, new_n15817, new_n15818,
    new_n15819, new_n15820, new_n15821, new_n15822, new_n15823, new_n15824,
    new_n15825, new_n15826, new_n15827, new_n15828, new_n15829, new_n15830,
    new_n15831_1, new_n15832, new_n15833, new_n15834, new_n15835,
    new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841,
    new_n15842, new_n15843, new_n15844, new_n15845, new_n15846_1,
    new_n15847, new_n15848, new_n15849, new_n15850, new_n15851, new_n15852,
    new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859_1, new_n15860, new_n15861, new_n15862, new_n15863,
    new_n15864, new_n15865, new_n15866, new_n15867, new_n15868,
    new_n15869_1, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884_1,
    new_n15885_1, new_n15886, new_n15887, new_n15888, new_n15889_1,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917_1, new_n15918_1,
    new_n15919, new_n15920, new_n15921, new_n15922_1, new_n15923,
    new_n15924, new_n15925, new_n15926, new_n15927, new_n15928, new_n15929,
    new_n15930, new_n15931, new_n15932, new_n15933, new_n15934, new_n15935,
    new_n15936_1, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947_1, new_n15948, new_n15949, new_n15950, new_n15951,
    new_n15952, new_n15953, new_n15954, new_n15955, new_n15956_1,
    new_n15957, new_n15958_1, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967_1, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15974, new_n15975, new_n15976, new_n15977,
    new_n15978, new_n15979_1, new_n15980, new_n15981, new_n15982,
    new_n15983, new_n15984, new_n15985, new_n15986_1, new_n15987,
    new_n15988, new_n15989, new_n15990, new_n15991, new_n15992, new_n15993,
    new_n15994, new_n15995, new_n15996, new_n15997, new_n15998, new_n15999,
    new_n16000, new_n16001, new_n16002, new_n16004, new_n16008, new_n16009,
    new_n16010, new_n16011, new_n16012, new_n16013_1, new_n16014,
    new_n16015, new_n16016, new_n16017, new_n16018, new_n16019, new_n16020,
    new_n16021, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029_1, new_n16030, new_n16031, new_n16032, new_n16033,
    new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039,
    new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045,
    new_n16046, new_n16047, new_n16048, new_n16049, new_n16050, new_n16051,
    new_n16052, new_n16053, new_n16054, new_n16055, new_n16056, new_n16057,
    new_n16058, new_n16059, new_n16060_1, new_n16061, new_n16062_1,
    new_n16063, new_n16064, new_n16065, new_n16066, new_n16067,
    new_n16068_1, new_n16069, new_n16070, new_n16071, new_n16072,
    new_n16073, new_n16074, new_n16075, new_n16076, new_n16077, new_n16078,
    new_n16079, new_n16080_1, new_n16081, new_n16082, new_n16083,
    new_n16084, new_n16085, new_n16086, new_n16087, new_n16088, new_n16089,
    new_n16090, new_n16091, new_n16092, new_n16093, new_n16094, new_n16095,
    new_n16096, new_n16097, new_n16098_1, new_n16099, new_n16100,
    new_n16101, new_n16102, new_n16103, new_n16104, new_n16105, new_n16106,
    new_n16107, new_n16108, new_n16109, new_n16110_1, new_n16111,
    new_n16112, new_n16113, new_n16114, new_n16115, new_n16116, new_n16117,
    new_n16118, new_n16119, new_n16120, new_n16121, new_n16122, new_n16123,
    new_n16124, new_n16125, new_n16126, new_n16129, new_n16130, new_n16131,
    new_n16132, new_n16133, new_n16134, new_n16135, new_n16136, new_n16137,
    new_n16138, new_n16139, new_n16140, new_n16141, new_n16142_1,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16156, new_n16157, new_n16158_1, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167_1, new_n16168, new_n16169, new_n16170, new_n16171,
    new_n16172, new_n16173, new_n16174, new_n16175, new_n16176, new_n16177,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185_1, new_n16186, new_n16187, new_n16188, new_n16189,
    new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195,
    new_n16196_1, new_n16197, new_n16198, new_n16199, new_n16200,
    new_n16201, new_n16202, new_n16203, new_n16204, new_n16205,
    new_n16206_1, new_n16207, new_n16208, new_n16209, new_n16210,
    new_n16211, new_n16212, new_n16213, new_n16214, new_n16215_1,
    new_n16216, new_n16217_1, new_n16218_1, new_n16219_1, new_n16221,
    new_n16222, new_n16223_1, new_n16224, new_n16225, new_n16226,
    new_n16227, new_n16228, new_n16229, new_n16230_1, new_n16231,
    new_n16232, new_n16233, new_n16234, new_n16235, new_n16236, new_n16237,
    new_n16238, new_n16239, new_n16240, new_n16241, new_n16242,
    new_n16243_1, new_n16244, new_n16245, new_n16246, new_n16247_1,
    new_n16248, new_n16249, new_n16250, new_n16251, new_n16252, new_n16253,
    new_n16254, new_n16255, new_n16256, new_n16257, new_n16258, new_n16259,
    new_n16260, new_n16261, new_n16262, new_n16263, new_n16264, new_n16265,
    new_n16266, new_n16267, new_n16268, new_n16269, new_n16270, new_n16271,
    new_n16272, new_n16273, new_n16274, new_n16275_1, new_n16276,
    new_n16277, new_n16278, new_n16279_1, new_n16280, new_n16281,
    new_n16282, new_n16283, new_n16284, new_n16285, new_n16286, new_n16287,
    new_n16288, new_n16289, new_n16290, new_n16291, new_n16292, new_n16293,
    new_n16294, new_n16295, new_n16296, new_n16297, new_n16298, new_n16299,
    new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305,
    new_n16306, new_n16307, new_n16308, new_n16309, new_n16310, new_n16311,
    new_n16312, new_n16313, new_n16314, new_n16315, new_n16316, new_n16317,
    new_n16318, new_n16319, new_n16320, new_n16321, new_n16322_1,
    new_n16323, new_n16324, new_n16325, new_n16326, new_n16327_1,
    new_n16328, new_n16329, new_n16330, new_n16331, new_n16332, new_n16333,
    new_n16334, new_n16335, new_n16336, new_n16337, new_n16338, new_n16339,
    new_n16340, new_n16341, new_n16342, new_n16343, new_n16344, new_n16345,
    new_n16346, new_n16347, new_n16348, new_n16349, new_n16350_1,
    new_n16351, new_n16352, new_n16353, new_n16354, new_n16355, new_n16356,
    new_n16357, new_n16358, new_n16359, new_n16360, new_n16361, new_n16362,
    new_n16363, new_n16364, new_n16365, new_n16366, new_n16367_1,
    new_n16368, new_n16369, new_n16370, new_n16371, new_n16372, new_n16373,
    new_n16374, new_n16375, new_n16376_1, new_n16377, new_n16378,
    new_n16379_1, new_n16380, new_n16381, new_n16382, new_n16383,
    new_n16384, new_n16385, new_n16386, new_n16387, new_n16388, new_n16389,
    new_n16390, new_n16391, new_n16392, new_n16393, new_n16395,
    new_n16396_1, new_n16397, new_n16398_1, new_n16399, new_n16400,
    new_n16401, new_n16402, new_n16403, new_n16404, new_n16405,
    new_n16406_1, new_n16407_1, new_n16408, new_n16409, new_n16410,
    new_n16411, new_n16412, new_n16413, new_n16414, new_n16415, new_n16416,
    new_n16417, new_n16418, new_n16419_1, new_n16420, new_n16421,
    new_n16422, new_n16423, new_n16424_1, new_n16425, new_n16426,
    new_n16427, new_n16428_1, new_n16429, new_n16430, new_n16431,
    new_n16432, new_n16433_1, new_n16434, new_n16435, new_n16436,
    new_n16437, new_n16438, new_n16439_1, new_n16440_1, new_n16441,
    new_n16442, new_n16443, new_n16444, new_n16445_1, new_n16446,
    new_n16447, new_n16448, new_n16449, new_n16450, new_n16451, new_n16452,
    new_n16453, new_n16454, new_n16455, new_n16456, new_n16457, new_n16458,
    new_n16459, new_n16460_1, new_n16461, new_n16462, new_n16463,
    new_n16464, new_n16465, new_n16466, new_n16467, new_n16468, new_n16469,
    new_n16470, new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476_1, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481_1, new_n16482_1, new_n16483, new_n16484, new_n16485,
    new_n16486, new_n16487, new_n16488, new_n16489, new_n16490, new_n16491,
    new_n16494, new_n16495, new_n16496, new_n16497, new_n16498, new_n16499,
    new_n16500, new_n16501, new_n16502_1, new_n16503, new_n16504,
    new_n16505, new_n16506_1, new_n16507_1, new_n16508, new_n16509,
    new_n16510, new_n16511, new_n16512, new_n16513, new_n16514, new_n16515,
    new_n16516_1, new_n16517_1, new_n16518, new_n16519, new_n16520,
    new_n16521_1, new_n16522, new_n16523, new_n16524_1, new_n16525,
    new_n16526, new_n16527_1, new_n16528, new_n16529, new_n16530,
    new_n16531, new_n16532, new_n16533, new_n16534, new_n16535, new_n16536,
    new_n16537, new_n16538, new_n16539, new_n16540, new_n16541, new_n16542,
    new_n16543, new_n16544_1, new_n16545, new_n16546, new_n16547,
    new_n16548, new_n16549, new_n16550, new_n16551, new_n16552, new_n16553,
    new_n16554_1, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583_1, new_n16584_1, new_n16585, new_n16586, new_n16587,
    new_n16588, new_n16589_1, new_n16590, new_n16591, new_n16592,
    new_n16593, new_n16594, new_n16595, new_n16596_1, new_n16597,
    new_n16599, new_n16600, new_n16601, new_n16602, new_n16603, new_n16604,
    new_n16605, new_n16606, new_n16607, new_n16608_1, new_n16609,
    new_n16610, new_n16611, new_n16612, new_n16613, new_n16614, new_n16615,
    new_n16616, new_n16617_1, new_n16618, new_n16619, new_n16620,
    new_n16621, new_n16622, new_n16623, new_n16624, new_n16625, new_n16626,
    new_n16627, new_n16628, new_n16629, new_n16630_1, new_n16631,
    new_n16632, new_n16633, new_n16634, new_n16635, new_n16636, new_n16637,
    new_n16638, new_n16639, new_n16640_1, new_n16641, new_n16642,
    new_n16643, new_n16644, new_n16645, new_n16646, new_n16647, new_n16648,
    new_n16649, new_n16650, new_n16651, new_n16652, new_n16653, new_n16654,
    new_n16655, new_n16656_1, new_n16658, new_n16659, new_n16660,
    new_n16661, new_n16662, new_n16663, new_n16664, new_n16665, new_n16666,
    new_n16667, new_n16668, new_n16669, new_n16670, new_n16671, new_n16672,
    new_n16673, new_n16674_1, new_n16675, new_n16676, new_n16679,
    new_n16680, new_n16681, new_n16682_1, new_n16683, new_n16684_1,
    new_n16685, new_n16686, new_n16687, new_n16688_1, new_n16689,
    new_n16690, new_n16691, new_n16692, new_n16693, new_n16694, new_n16695,
    new_n16696, new_n16697, new_n16698, new_n16699, new_n16700, new_n16701,
    new_n16702, new_n16703, new_n16704, new_n16705, new_n16706, new_n16707,
    new_n16708, new_n16709, new_n16710, new_n16711, new_n16712, new_n16713,
    new_n16714, new_n16715, new_n16716, new_n16717, new_n16718, new_n16719,
    new_n16720, new_n16721, new_n16722_1, new_n16723, new_n16724,
    new_n16725, new_n16726, new_n16727, new_n16728, new_n16729, new_n16730,
    new_n16731, new_n16732, new_n16733_1, new_n16734, new_n16735,
    new_n16736, new_n16737, new_n16738, new_n16739, new_n16740, new_n16741,
    new_n16742, new_n16743_1, new_n16744, new_n16745, new_n16746,
    new_n16747, new_n16748, new_n16749, new_n16750, new_n16751, new_n16752,
    new_n16753, new_n16754, new_n16755, new_n16756, new_n16757, new_n16761,
    new_n16762, new_n16763, new_n16764, new_n16765, new_n16766, new_n16767,
    new_n16768, new_n16769, new_n16770, new_n16771, new_n16772, new_n16776,
    new_n16777, new_n16778, new_n16779, new_n16780, new_n16781, new_n16782,
    new_n16783, new_n16784, new_n16785, new_n16786, new_n16787, new_n16788,
    new_n16789, new_n16790, new_n16791, new_n16792, new_n16793, new_n16794,
    new_n16795, new_n16796, new_n16797, new_n16798_1, new_n16799,
    new_n16800, new_n16803, new_n16804, new_n16805, new_n16806, new_n16807,
    new_n16808, new_n16809, new_n16810, new_n16811, new_n16812_1,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817,
    new_n16818_1, new_n16819, new_n16820, new_n16821, new_n16822,
    new_n16823, new_n16824_1, new_n16825, new_n16826, new_n16827,
    new_n16828, new_n16829, new_n16830, new_n16831, new_n16832, new_n16833,
    new_n16834_1, new_n16835, new_n16836, new_n16837_1, new_n16838,
    new_n16839, new_n16840, new_n16841_1, new_n16842, new_n16843,
    new_n16844, new_n16845, new_n16846, new_n16847, new_n16848, new_n16849,
    new_n16850, new_n16851, new_n16852, new_n16853, new_n16854, new_n16855,
    new_n16856, new_n16857, new_n16858, new_n16859, new_n16860, new_n16861,
    new_n16862, new_n16863, new_n16864, new_n16865, new_n16866, new_n16867,
    new_n16868, new_n16869, new_n16870, new_n16871, new_n16872, new_n16873,
    new_n16874, new_n16875, new_n16876, new_n16877, new_n16878, new_n16879,
    new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885_1, new_n16886, new_n16887, new_n16888, new_n16889,
    new_n16890, new_n16891, new_n16892, new_n16893, new_n16894, new_n16895,
    new_n16896, new_n16897, new_n16898, new_n16899, new_n16900, new_n16901,
    new_n16902, new_n16903, new_n16904, new_n16905_1, new_n16906,
    new_n16907, new_n16908, new_n16909, new_n16910, new_n16911_1,
    new_n16912, new_n16913, new_n16914, new_n16915, new_n16916, new_n16917,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951_1, new_n16952, new_n16953, new_n16954_1, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968_1, new_n16969, new_n16970, new_n16971_1, new_n16972,
    new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978,
    new_n16979, new_n16980, new_n16981, new_n16982, new_n16983, new_n16984,
    new_n16985, new_n16986, new_n16987, new_n16988_1, new_n16989_1,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994_1,
    new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000,
    new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006_1, new_n17007, new_n17008, new_n17009, new_n17010,
    new_n17011, new_n17012, new_n17013, new_n17014, new_n17015, new_n17016,
    new_n17017, new_n17018, new_n17019, new_n17020, new_n17021, new_n17022,
    new_n17023, new_n17024, new_n17025, new_n17026, new_n17027, new_n17028,
    new_n17029, new_n17030, new_n17031, new_n17032, new_n17033, new_n17034,
    new_n17035_1, new_n17036, new_n17037_1, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045,
    new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051,
    new_n17052, new_n17053, new_n17055, new_n17056, new_n17057, new_n17058,
    new_n17059, new_n17060, new_n17061, new_n17062, new_n17063, new_n17064,
    new_n17065, new_n17067, new_n17068_1, new_n17069_1, new_n17070_1,
    new_n17071, new_n17072, new_n17073, new_n17074, new_n17075_1,
    new_n17076, new_n17077_1, new_n17078, new_n17079, new_n17080,
    new_n17081, new_n17082, new_n17083, new_n17084_1, new_n17085,
    new_n17086, new_n17087, new_n17088, new_n17089, new_n17090_1,
    new_n17091, new_n17092, new_n17093, new_n17094, new_n17095_1,
    new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101,
    new_n17102, new_n17103, new_n17104_1, new_n17105, new_n17106_1,
    new_n17107, new_n17108, new_n17109, new_n17111, new_n17112, new_n17113,
    new_n17114, new_n17115, new_n17116, new_n17117, new_n17118,
    new_n17119_1, new_n17120, new_n17121, new_n17122, new_n17123,
    new_n17124, new_n17125, new_n17126, new_n17127, new_n17128, new_n17129,
    new_n17130_1, new_n17131, new_n17132, new_n17133, new_n17134,
    new_n17135, new_n17136, new_n17137, new_n17138_1, new_n17139,
    new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17147, new_n17148, new_n17149, new_n17150, new_n17152,
    new_n17153, new_n17154, new_n17155, new_n17156, new_n17157, new_n17158,
    new_n17159, new_n17160, new_n17161, new_n17162, new_n17163_1,
    new_n17164, new_n17165, new_n17166, new_n17167, new_n17168_1,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174,
    new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180,
    new_n17181, new_n17184, new_n17185, new_n17186, new_n17187, new_n17188,
    new_n17189, new_n17190, new_n17191, new_n17192, new_n17193, new_n17194,
    new_n17195, new_n17196, new_n17197, new_n17198, new_n17199, new_n17200,
    new_n17201, new_n17202_1, new_n17203, new_n17204, new_n17205,
    new_n17206, new_n17207, new_n17209, new_n17210, new_n17211, new_n17212,
    new_n17213, new_n17214, new_n17215, new_n17216, new_n17217, new_n17218,
    new_n17219_1, new_n17220, new_n17221, new_n17222, new_n17223,
    new_n17224, new_n17225, new_n17226, new_n17227, new_n17228, new_n17229,
    new_n17230, new_n17231, new_n17232_1, new_n17233, new_n17234,
    new_n17235, new_n17236_1, new_n17237, new_n17238, new_n17239,
    new_n17240, new_n17241, new_n17242, new_n17243_1, new_n17244,
    new_n17245, new_n17246, new_n17247, new_n17248, new_n17249,
    new_n17250_1, new_n17251_1, new_n17252, new_n17253, new_n17254,
    new_n17255, new_n17256, new_n17257, new_n17258, new_n17259, new_n17260,
    new_n17261, new_n17262, new_n17263_1, new_n17264, new_n17265,
    new_n17266, new_n17267, new_n17268, new_n17269, new_n17270, new_n17271,
    new_n17272, new_n17273, new_n17274, new_n17275, new_n17276, new_n17278,
    new_n17279, new_n17280, new_n17281, new_n17282, new_n17283, new_n17284,
    new_n17285_1, new_n17286, new_n17287, new_n17288, new_n17289,
    new_n17290, new_n17291, new_n17292, new_n17293, new_n17294, new_n17295,
    new_n17296, new_n17297, new_n17298, new_n17299, new_n17300, new_n17301,
    new_n17302_1, new_n17303, new_n17304, new_n17305, new_n17306,
    new_n17307, new_n17308, new_n17309, new_n17310, new_n17311, new_n17312,
    new_n17313, new_n17314, new_n17315, new_n17316, new_n17317, new_n17318,
    new_n17319, new_n17320_1, new_n17321, new_n17322, new_n17323,
    new_n17324, new_n17325, new_n17326, new_n17327, new_n17328, new_n17329,
    new_n17330, new_n17331, new_n17332, new_n17333, new_n17334, new_n17335,
    new_n17336, new_n17337_1, new_n17338, new_n17339, new_n17340,
    new_n17341, new_n17342, new_n17343, new_n17344_1, new_n17345,
    new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351_1, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359_1, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387_1, new_n17388, new_n17389,
    new_n17390, new_n17391_1, new_n17392_1, new_n17393, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421_1, new_n17422, new_n17423,
    new_n17424, new_n17425, new_n17426, new_n17427, new_n17428, new_n17429,
    new_n17430, new_n17431, new_n17432_1, new_n17433, new_n17434,
    new_n17435, new_n17436_1, new_n17437, new_n17438, new_n17439,
    new_n17440_1, new_n17441, new_n17442, new_n17443, new_n17444,
    new_n17445, new_n17446, new_n17448, new_n17449, new_n17450_1,
    new_n17451, new_n17452, new_n17453, new_n17454, new_n17455, new_n17456,
    new_n17457, new_n17458_1, new_n17459, new_n17460, new_n17461_1,
    new_n17464, new_n17465, new_n17466_1, new_n17467, new_n17468,
    new_n17469, new_n17470, new_n17471, new_n17472, new_n17473, new_n17474,
    new_n17475, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17486, new_n17487, new_n17488, new_n17489, new_n17490,
    new_n17491, new_n17492, new_n17493_1, new_n17494, new_n17501,
    new_n17502, new_n17503, new_n17504, new_n17505, new_n17506, new_n17507,
    new_n17508, new_n17509, new_n17510, new_n17511, new_n17512, new_n17513,
    new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519,
    new_n17520, new_n17521, new_n17522, new_n17523, new_n17524_1,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529_1,
    new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535,
    new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541,
    new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547,
    new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553,
    new_n17554, new_n17555, new_n17556, new_n17557_1, new_n17558,
    new_n17559, new_n17560, new_n17561, new_n17562, new_n17563, new_n17564,
    new_n17565, new_n17566, new_n17567, new_n17568, new_n17569, new_n17570,
    new_n17571, new_n17572, new_n17573, new_n17574, new_n17575, new_n17576,
    new_n17577, new_n17578, new_n17579, new_n17580, new_n17581, new_n17582,
    new_n17583_1, new_n17584, new_n17585, new_n17586, new_n17587,
    new_n17588, new_n17589, new_n17590, new_n17591, new_n17592_1,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17599,
    new_n17600, new_n17601, new_n17602, new_n17603, new_n17604, new_n17605,
    new_n17606, new_n17607, new_n17608, new_n17609, new_n17610, new_n17611,
    new_n17612, new_n17613, new_n17614, new_n17615, new_n17616, new_n17617,
    new_n17618, new_n17619, new_n17620, new_n17621, new_n17622, new_n17623,
    new_n17624, new_n17625, new_n17626, new_n17627, new_n17628, new_n17629,
    new_n17630, new_n17631, new_n17632, new_n17633, new_n17634, new_n17635,
    new_n17636, new_n17637, new_n17638_1, new_n17639, new_n17640,
    new_n17641, new_n17642, new_n17643, new_n17644, new_n17646, new_n17647,
    new_n17648, new_n17649, new_n17650, new_n17651, new_n17652, new_n17653,
    new_n17654, new_n17655, new_n17656, new_n17657, new_n17658, new_n17659,
    new_n17660, new_n17661, new_n17662, new_n17663, new_n17664_1,
    new_n17665, new_n17666, new_n17667, new_n17668, new_n17669, new_n17670,
    new_n17671, new_n17672, new_n17673, new_n17674, new_n17675, new_n17676,
    new_n17677, new_n17678, new_n17679, new_n17680, new_n17681, new_n17682,
    new_n17683, new_n17684, new_n17685, new_n17686, new_n17687_1,
    new_n17688, new_n17689, new_n17690, new_n17691, new_n17692, new_n17693,
    new_n17694, new_n17695, new_n17696, new_n17697, new_n17698, new_n17699,
    new_n17700, new_n17701, new_n17702, new_n17703, new_n17704, new_n17705,
    new_n17706, new_n17707, new_n17708, new_n17709, new_n17710, new_n17711,
    new_n17712, new_n17713, new_n17714, new_n17715, new_n17716, new_n17717,
    new_n17718, new_n17719, new_n17720, new_n17721_1, new_n17722,
    new_n17723, new_n17724, new_n17725, new_n17726, new_n17727, new_n17728,
    new_n17729, new_n17730, new_n17731, new_n17732, new_n17733, new_n17734,
    new_n17735_1, new_n17736, new_n17737, new_n17738_1, new_n17739,
    new_n17740, new_n17741, new_n17742, new_n17743, new_n17744, new_n17745,
    new_n17746_1, new_n17747, new_n17748, new_n17749_1, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17782, new_n17783, new_n17784_1, new_n17785,
    new_n17786, new_n17787, new_n17788, new_n17789, new_n17790, new_n17791,
    new_n17792, new_n17793, new_n17794, new_n17795, new_n17796, new_n17797,
    new_n17798, new_n17799, new_n17800, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17807, new_n17808, new_n17809, new_n17810,
    new_n17811, new_n17812, new_n17813, new_n17814, new_n17815, new_n17816,
    new_n17817, new_n17818, new_n17819, new_n17820_1, new_n17821,
    new_n17822, new_n17823, new_n17824, new_n17825, new_n17826, new_n17827,
    new_n17828, new_n17829, new_n17830, new_n17831, new_n17832, new_n17833,
    new_n17834, new_n17835, new_n17836, new_n17837, new_n17838, new_n17839,
    new_n17840, new_n17841, new_n17842, new_n17843, new_n17844, new_n17845,
    new_n17846, new_n17847, new_n17848, new_n17849, new_n17852, new_n17853,
    new_n17854, new_n17855_1, new_n17856, new_n17857, new_n17858,
    new_n17859, new_n17860, new_n17861, new_n17862, new_n17863, new_n17864,
    new_n17865, new_n17866, new_n17867, new_n17868, new_n17871, new_n17872,
    new_n17873, new_n17874, new_n17875, new_n17876, new_n17877_1,
    new_n17878, new_n17879, new_n17883, new_n17884, new_n17885, new_n17886,
    new_n17887, new_n17888, new_n17889_1, new_n17890, new_n17891,
    new_n17892, new_n17893, new_n17894, new_n17895, new_n17896, new_n17897,
    new_n17898, new_n17899, new_n17900, new_n17901, new_n17902, new_n17903,
    new_n17904, new_n17905, new_n17906, new_n17907, new_n17908, new_n17909,
    new_n17910, new_n17911_1, new_n17912_1, new_n17913, new_n17914,
    new_n17915, new_n17916, new_n17917, new_n17918, new_n17919, new_n17920,
    new_n17921, new_n17922, new_n17923, new_n17924, new_n17925, new_n17926,
    new_n17929, new_n17930, new_n17931_1, new_n17932, new_n17933,
    new_n17934, new_n17935, new_n17936, new_n17937, new_n17938, new_n17939,
    new_n17940, new_n17941, new_n17942, new_n17943, new_n17944, new_n17945,
    new_n17946, new_n17947, new_n17948_1, new_n17949, new_n17950,
    new_n17951, new_n17952, new_n17953, new_n17954_1, new_n17955,
    new_n17956_1, new_n17957, new_n17958, new_n17959_1, new_n17960,
    new_n17961, new_n17962, new_n17963_1, new_n17964, new_n17965,
    new_n17966, new_n17967, new_n17968_1, new_n17969, new_n17970,
    new_n17971, new_n17972, new_n17973, new_n17974, new_n17975,
    new_n17976_1, new_n17977, new_n17978, new_n17979, new_n17980,
    new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986,
    new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992,
    new_n17993, new_n17994, new_n17995, new_n17996, new_n17997,
    new_n17998_1, new_n17999, new_n18000, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18016, new_n18017, new_n18018, new_n18019, new_n18020, new_n18021,
    new_n18022, new_n18023, new_n18024, new_n18025_1, new_n18026,
    new_n18027, new_n18028, new_n18029, new_n18030, new_n18031, new_n18032,
    new_n18033, new_n18034, new_n18035_1, new_n18036, new_n18037,
    new_n18038, new_n18039, new_n18040, new_n18041, new_n18042,
    new_n18043_1, new_n18044, new_n18045_1, new_n18046, new_n18047,
    new_n18048, new_n18049, new_n18050, new_n18051, new_n18052, new_n18053,
    new_n18055, new_n18056, new_n18057, new_n18058, new_n18059_1,
    new_n18060, new_n18061_1, new_n18062, new_n18063, new_n18064,
    new_n18065, new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071_1, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18078, new_n18079, new_n18080, new_n18081,
    new_n18082, new_n18083, new_n18084, new_n18085, new_n18086, new_n18087,
    new_n18088, new_n18089, new_n18090, new_n18091, new_n18092, new_n18093,
    new_n18094, new_n18095, new_n18096, new_n18097, new_n18098, new_n18099,
    new_n18100, new_n18101, new_n18102, new_n18103, new_n18104,
    new_n18105_1, new_n18106, new_n18107, new_n18108, new_n18109,
    new_n18110, new_n18111, new_n18112, new_n18113, new_n18114, new_n18115,
    new_n18116, new_n18117, new_n18118, new_n18119, new_n18120, new_n18121,
    new_n18122, new_n18123, new_n18124, new_n18125, new_n18126, new_n18132,
    new_n18133, new_n18134, new_n18135, new_n18136, new_n18137, new_n18138,
    new_n18139, new_n18140, new_n18141, new_n18142, new_n18143_1,
    new_n18144, new_n18145_1, new_n18146, new_n18147, new_n18148,
    new_n18149, new_n18150, new_n18151_1, new_n18152_1, new_n18153,
    new_n18154, new_n18155, new_n18156, new_n18157_1, new_n18158,
    new_n18159, new_n18160, new_n18161, new_n18162, new_n18163, new_n18164,
    new_n18165, new_n18166, new_n18167, new_n18168, new_n18169, new_n18170,
    new_n18171_1, new_n18172, new_n18173, new_n18174, new_n18175,
    new_n18176, new_n18177, new_n18178, new_n18179, new_n18180, new_n18181,
    new_n18182, new_n18183, new_n18184, new_n18185, new_n18186, new_n18187,
    new_n18188, new_n18189, new_n18190, new_n18191, new_n18192,
    new_n18193_1, new_n18194, new_n18195, new_n18196, new_n18197,
    new_n18198, new_n18201, new_n18202, new_n18203, new_n18204, new_n18205,
    new_n18206, new_n18207, new_n18208, new_n18209, new_n18210, new_n18211,
    new_n18212, new_n18213, new_n18214, new_n18215, new_n18216, new_n18217,
    new_n18218, new_n18219, new_n18220, new_n18221, new_n18222, new_n18223,
    new_n18224, new_n18225, new_n18226, new_n18227_1, new_n18228,
    new_n18229, new_n18230, new_n18233, new_n18234, new_n18235, new_n18236,
    new_n18237, new_n18238_1, new_n18239, new_n18240, new_n18241_1,
    new_n18242, new_n18243, new_n18244, new_n18245, new_n18246, new_n18247,
    new_n18248, new_n18249, new_n18250, new_n18251, new_n18252, new_n18253,
    new_n18254_1, new_n18256, new_n18261, new_n18262, new_n18263,
    new_n18264, new_n18265, new_n18266, new_n18267, new_n18268, new_n18269,
    new_n18270, new_n18271, new_n18272, new_n18273, new_n18274_1,
    new_n18275, new_n18276, new_n18277, new_n18278, new_n18279, new_n18280,
    new_n18281, new_n18282, new_n18283, new_n18284, new_n18285, new_n18286,
    new_n18287, new_n18288_1, new_n18289, new_n18290_1, new_n18291,
    new_n18292, new_n18293, new_n18294, new_n18295_1, new_n18296,
    new_n18297, new_n18298, new_n18299, new_n18300, new_n18301_1,
    new_n18302, new_n18303, new_n18304_1, new_n18305, new_n18306,
    new_n18307, new_n18308, new_n18309, new_n18310_1, new_n18311_1,
    new_n18312, new_n18313, new_n18314, new_n18315, new_n18316, new_n18317,
    new_n18318, new_n18319, new_n18320, new_n18321, new_n18322,
    new_n18323_1, new_n18324, new_n18325, new_n18326, new_n18327,
    new_n18328, new_n18329, new_n18330, new_n18331, new_n18332_1,
    new_n18333, new_n18334, new_n18335, new_n18336, new_n18337, new_n18338,
    new_n18339, new_n18340, new_n18341, new_n18342, new_n18343_1,
    new_n18344, new_n18345_1, new_n18346, new_n18347, new_n18348,
    new_n18349, new_n18350_1, new_n18351, new_n18352, new_n18353,
    new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359,
    new_n18360, new_n18361, new_n18362_1, new_n18363, new_n18364,
    new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370,
    new_n18371, new_n18372, new_n18376, new_n18377_1, new_n18378,
    new_n18379, new_n18380, new_n18381, new_n18382, new_n18383, new_n18384,
    new_n18385, new_n18386, new_n18387, new_n18388, new_n18389, new_n18390,
    new_n18391, new_n18392, new_n18393, new_n18394, new_n18395, new_n18396,
    new_n18397, new_n18398, new_n18399, new_n18400, new_n18401, new_n18402,
    new_n18409_1, new_n18410, new_n18411, new_n18412, new_n18413,
    new_n18414_1, new_n18415, new_n18416, new_n18417, new_n18418_1,
    new_n18419, new_n18420, new_n18421, new_n18422, new_n18423, new_n18424,
    new_n18425, new_n18426, new_n18427, new_n18428, new_n18429, new_n18430,
    new_n18431, new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437_1, new_n18438, new_n18439_1, new_n18440, new_n18441,
    new_n18442, new_n18443, new_n18444_1, new_n18445_1, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451,
    new_n18452_1, new_n18453, new_n18454, new_n18455, new_n18456,
    new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462,
    new_n18463, new_n18464, new_n18465, new_n18466, new_n18467_1,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482_1, new_n18483_1, new_n18484,
    new_n18485, new_n18488, new_n18489, new_n18490, new_n18491, new_n18492,
    new_n18493, new_n18494, new_n18495, new_n18496_1, new_n18497,
    new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503,
    new_n18504, new_n18505, new_n18506, new_n18507, new_n18508,
    new_n18509_1, new_n18510, new_n18511, new_n18512, new_n18513_1,
    new_n18514, new_n18515_1, new_n18516, new_n18517, new_n18518,
    new_n18519, new_n18520, new_n18521, new_n18522, new_n18523, new_n18524,
    new_n18525, new_n18526, new_n18527, new_n18528, new_n18529, new_n18530,
    new_n18531, new_n18532, new_n18533, new_n18534, new_n18535, new_n18536,
    new_n18537_1, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18555, new_n18556, new_n18557, new_n18558_1,
    new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564,
    new_n18565, new_n18566, new_n18567, new_n18569, new_n18570, new_n18571,
    new_n18572_1, new_n18573, new_n18574_1, new_n18575, new_n18576_1,
    new_n18577, new_n18578_1, new_n18579, new_n18580, new_n18581,
    new_n18582_1, new_n18583_1, new_n18584_1, new_n18585, new_n18586,
    new_n18587, new_n18588, new_n18589, new_n18590, new_n18591, new_n18592,
    new_n18593, new_n18594, new_n18595, new_n18596, new_n18597, new_n18598,
    new_n18599, new_n18600, new_n18601, new_n18602, new_n18603, new_n18604,
    new_n18605, new_n18606, new_n18607, new_n18608, new_n18609,
    new_n18610_1, new_n18611, new_n18612, new_n18613, new_n18614,
    new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620,
    new_n18621, new_n18622, new_n18623, new_n18625, new_n18626, new_n18627,
    new_n18628, new_n18629, new_n18630, new_n18631, new_n18632, new_n18633,
    new_n18634, new_n18635_1, new_n18636, new_n18637, new_n18638,
    new_n18639, new_n18640, new_n18641, new_n18642, new_n18643, new_n18644,
    new_n18645, new_n18646, new_n18647, new_n18648, new_n18649_1,
    new_n18650, new_n18651, new_n18652, new_n18653_1, new_n18654,
    new_n18655, new_n18656, new_n18657, new_n18658, new_n18659, new_n18660,
    new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666,
    new_n18667, new_n18668, new_n18669, new_n18674, new_n18675, new_n18676,
    new_n18677, new_n18678, new_n18679_1, new_n18680, new_n18681,
    new_n18682, new_n18683, new_n18684, new_n18685, new_n18686, new_n18687,
    new_n18692, new_n18693_1, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707,
    new_n18708_1, new_n18709, new_n18710, new_n18711, new_n18712,
    new_n18713, new_n18714, new_n18715, new_n18716, new_n18717, new_n18718,
    new_n18719, new_n18720, new_n18721_1, new_n18722, new_n18723,
    new_n18724, new_n18725_1, new_n18726, new_n18727, new_n18728,
    new_n18729, new_n18730, new_n18731, new_n18732, new_n18733, new_n18734,
    new_n18735, new_n18736, new_n18737_1, new_n18738, new_n18739,
    new_n18740, new_n18741, new_n18742, new_n18744, new_n18745_1,
    new_n18746, new_n18747, new_n18748, new_n18750, new_n18751_1,
    new_n18752, new_n18753, new_n18754, new_n18755, new_n18756, new_n18757,
    new_n18758, new_n18759, new_n18760, new_n18761, new_n18762, new_n18766,
    new_n18767, new_n18768, new_n18769, new_n18770, new_n18771, new_n18772,
    new_n18773, new_n18774, new_n18775, new_n18776, new_n18777, new_n18778,
    new_n18779, new_n18780_1, new_n18781, new_n18782_1, new_n18783,
    new_n18784, new_n18785, new_n18786, new_n18787, new_n18788, new_n18789,
    new_n18791, new_n18792, new_n18793, new_n18794, new_n18795, new_n18796,
    new_n18797, new_n18798, new_n18799, new_n18800, new_n18801,
    new_n18802_1, new_n18803, new_n18804, new_n18805, new_n18806,
    new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812,
    new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818,
    new_n18819, new_n18820, new_n18821, new_n18822, new_n18823, new_n18824,
    new_n18825, new_n18826, new_n18827, new_n18828, new_n18829,
    new_n18830_1, new_n18831_1, new_n18832, new_n18833, new_n18834,
    new_n18835, new_n18836, new_n18837, new_n18838, new_n18839, new_n18840,
    new_n18841, new_n18842, new_n18843_1, new_n18844, new_n18845,
    new_n18846, new_n18847, new_n18848, new_n18849, new_n18850, new_n18851,
    new_n18852, new_n18853, new_n18854, new_n18855, new_n18856, new_n18857,
    new_n18858_1, new_n18859_1, new_n18860, new_n18861, new_n18862,
    new_n18864_1, new_n18865_1, new_n18866, new_n18867, new_n18868,
    new_n18869, new_n18870, new_n18871, new_n18872, new_n18873, new_n18874,
    new_n18876, new_n18877, new_n18878, new_n18879, new_n18880_1,
    new_n18881, new_n18882, new_n18883, new_n18884, new_n18885,
    new_n18886_1, new_n18887_1, new_n18888, new_n18889, new_n18890,
    new_n18891, new_n18892, new_n18893, new_n18894, new_n18895, new_n18896,
    new_n18897, new_n18898, new_n18899, new_n18900, new_n18901_1,
    new_n18902, new_n18903, new_n18904, new_n18905, new_n18906,
    new_n18907_1, new_n18908, new_n18909, new_n18910, new_n18911,
    new_n18912, new_n18913, new_n18914, new_n18915, new_n18916, new_n18917,
    new_n18918, new_n18919_1, new_n18920, new_n18921, new_n18922,
    new_n18923, new_n18924, new_n18925, new_n18926_1, new_n18927,
    new_n18928, new_n18929, new_n18930, new_n18931, new_n18932, new_n18933,
    new_n18934, new_n18935, new_n18936, new_n18937, new_n18938, new_n18939,
    new_n18940_1, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945_1, new_n18946, new_n18947, new_n18948, new_n18949,
    new_n18950, new_n18951, new_n18952, new_n18953, new_n18954, new_n18955,
    new_n18956, new_n18957, new_n18958, new_n18959, new_n18960, new_n18961,
    new_n18962_1, new_n18963, new_n18964, new_n18965, new_n18966,
    new_n18967, new_n18968, new_n18969, new_n18970_1, new_n18971,
    new_n18972, new_n18973, new_n18974, new_n18975, new_n18976,
    new_n18977_1, new_n18978, new_n18979, new_n18980, new_n18981,
    new_n18982_1, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999_1, new_n19000, new_n19001, new_n19002, new_n19003,
    new_n19004, new_n19005_1, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033_1, new_n19034, new_n19035, new_n19036, new_n19037,
    new_n19038, new_n19039, new_n19040, new_n19041, new_n19042_1,
    new_n19043, new_n19044_1, new_n19045, new_n19046, new_n19047,
    new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053,
    new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065,
    new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071,
    new_n19072, new_n19073, new_n19074, new_n19075, new_n19076, new_n19077,
    new_n19078, new_n19079, new_n19080, new_n19081_1, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19090,
    new_n19091, new_n19092, new_n19093, new_n19094, new_n19095, new_n19096,
    new_n19097, new_n19098, new_n19099, new_n19100, new_n19101, new_n19102,
    new_n19103, new_n19104, new_n19105, new_n19106, new_n19107_1,
    new_n19108, new_n19109, new_n19110, new_n19111, new_n19112, new_n19113,
    new_n19114, new_n19115, new_n19116_1, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123,
    new_n19125_1, new_n19126, new_n19127, new_n19128, new_n19129,
    new_n19130, new_n19131, new_n19132, new_n19133, new_n19134, new_n19135,
    new_n19136, new_n19137, new_n19138, new_n19139, new_n19140,
    new_n19141_1, new_n19142, new_n19143, new_n19144_1, new_n19145,
    new_n19148, new_n19149, new_n19150, new_n19151, new_n19152, new_n19153,
    new_n19158, new_n19159, new_n19160, new_n19161, new_n19162,
    new_n19163_1, new_n19164_1, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174_1, new_n19175, new_n19176_1, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190,
    new_n19191, new_n19192, new_n19193, new_n19194, new_n19195,
    new_n19196_1, new_n19197, new_n19198, new_n19199, new_n19200,
    new_n19201, new_n19202_1, new_n19203, new_n19204, new_n19205,
    new_n19206, new_n19207, new_n19208, new_n19209, new_n19210, new_n19211,
    new_n19212, new_n19213, new_n19214, new_n19215, new_n19216, new_n19217,
    new_n19218, new_n19219, new_n19220_1, new_n19221_1, new_n19222,
    new_n19223_1, new_n19224_1, new_n19225, new_n19226, new_n19227,
    new_n19228_1, new_n19229, new_n19230, new_n19231, new_n19232,
    new_n19233_1, new_n19234_1, new_n19235, new_n19236, new_n19237,
    new_n19238, new_n19239, new_n19240, new_n19241, new_n19242, new_n19243,
    new_n19244_1, new_n19245, new_n19246, new_n19247, new_n19248,
    new_n19249, new_n19250, new_n19251, new_n19252, new_n19253, new_n19254,
    new_n19255, new_n19256, new_n19257, new_n19258, new_n19259, new_n19260,
    new_n19261, new_n19262, new_n19263, new_n19264, new_n19265, new_n19268,
    new_n19269, new_n19270_1, new_n19271, new_n19272, new_n19273,
    new_n19274, new_n19275, new_n19276, new_n19277, new_n19278, new_n19279,
    new_n19280, new_n19281, new_n19282_1, new_n19283, new_n19284,
    new_n19285, new_n19286, new_n19287, new_n19288, new_n19289, new_n19290,
    new_n19291, new_n19292, new_n19293, new_n19295, new_n19296, new_n19297,
    new_n19298, new_n19299, new_n19300, new_n19301, new_n19302, new_n19303,
    new_n19304, new_n19305, new_n19306, new_n19307, new_n19308, new_n19309,
    new_n19310, new_n19311, new_n19312, new_n19313, new_n19314_1,
    new_n19315_1, new_n19316, new_n19317, new_n19318, new_n19319,
    new_n19320, new_n19321, new_n19322, new_n19323_1, new_n19324,
    new_n19325, new_n19326, new_n19327_1, new_n19328, new_n19329,
    new_n19330, new_n19331, new_n19332, new_n19333_1, new_n19334,
    new_n19335, new_n19336, new_n19337, new_n19338, new_n19339, new_n19340,
    new_n19341, new_n19342, new_n19343, new_n19344, new_n19347,
    new_n19348_1, new_n19349, new_n19350, new_n19351, new_n19352,
    new_n19353, new_n19354_1, new_n19355, new_n19356, new_n19357_1,
    new_n19358, new_n19359, new_n19360, new_n19361_1, new_n19362,
    new_n19363, new_n19364, new_n19365, new_n19366, new_n19367_1,
    new_n19368, new_n19369, new_n19370, new_n19371, new_n19372, new_n19373,
    new_n19374, new_n19375, new_n19376, new_n19377, new_n19378, new_n19379,
    new_n19380, new_n19381, new_n19382, new_n19383, new_n19384,
    new_n19385_1, new_n19387, new_n19388, new_n19389_1, new_n19390,
    new_n19391, new_n19392, new_n19393, new_n19394, new_n19395, new_n19396,
    new_n19397, new_n19398, new_n19399, new_n19400, new_n19401_1,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414_1, new_n19415, new_n19416, new_n19417, new_n19418,
    new_n19419, new_n19420, new_n19421, new_n19422, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19442, new_n19443, new_n19444, new_n19445, new_n19446,
    new_n19447, new_n19448, new_n19453, new_n19454_1, new_n19455,
    new_n19456, new_n19457, new_n19458_1, new_n19459, new_n19460,
    new_n19461, new_n19462, new_n19463, new_n19464, new_n19465, new_n19466,
    new_n19467_1, new_n19468, new_n19469, new_n19470, new_n19471,
    new_n19472_1, new_n19473, new_n19474, new_n19475, new_n19476,
    new_n19477_1, new_n19478, new_n19479, new_n19480, new_n19481,
    new_n19482, new_n19483, new_n19484, new_n19485, new_n19486, new_n19487,
    new_n19488, new_n19489, new_n19490, new_n19491, new_n19492, new_n19493,
    new_n19494_1, new_n19495, new_n19496_1, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510,
    new_n19511, new_n19512, new_n19513, new_n19514_1, new_n19515_1,
    new_n19516, new_n19517, new_n19518, new_n19519, new_n19520, new_n19521,
    new_n19522, new_n19523_1, new_n19524, new_n19525, new_n19526,
    new_n19527, new_n19528, new_n19529, new_n19530, new_n19531_1,
    new_n19532, new_n19533, new_n19534, new_n19535, new_n19536, new_n19542,
    new_n19543, new_n19544, new_n19545, new_n19546, new_n19547, new_n19548,
    new_n19549, new_n19550, new_n19551, new_n19552, new_n19553, new_n19554,
    new_n19555, new_n19556, new_n19557, new_n19558, new_n19559, new_n19560,
    new_n19561, new_n19563, new_n19564, new_n19565, new_n19566, new_n19567,
    new_n19568, new_n19569, new_n19570_1, new_n19571, new_n19572,
    new_n19573, new_n19574, new_n19575_1, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641_1, new_n19642, new_n19643,
    new_n19648_1, new_n19649, new_n19650, new_n19651, new_n19652_1,
    new_n19653, new_n19654, new_n19655, new_n19656, new_n19657, new_n19658,
    new_n19659, new_n19660, new_n19661, new_n19662, new_n19663,
    new_n19664_1, new_n19665, new_n19666, new_n19667, new_n19668,
    new_n19669, new_n19670, new_n19671, new_n19672, new_n19673, new_n19674,
    new_n19675, new_n19676, new_n19677, new_n19678, new_n19679,
    new_n19680_1, new_n19681, new_n19682, new_n19683, new_n19684,
    new_n19685, new_n19686, new_n19687, new_n19688, new_n19689, new_n19690,
    new_n19691, new_n19692, new_n19693, new_n19694, new_n19695, new_n19696,
    new_n19697, new_n19698, new_n19699, new_n19700, new_n19701_1,
    new_n19702, new_n19703, new_n19704, new_n19705, new_n19706, new_n19707,
    new_n19708, new_n19709, new_n19710, new_n19711, new_n19712, new_n19713,
    new_n19714, new_n19715, new_n19716, new_n19717, new_n19718, new_n19721,
    new_n19722, new_n19723, new_n19724, new_n19725, new_n19726, new_n19727,
    new_n19728, new_n19729, new_n19730, new_n19731, new_n19732, new_n19733,
    new_n19734, new_n19735, new_n19736_1, new_n19737, new_n19738,
    new_n19739, new_n19740, new_n19741, new_n19742, new_n19743, new_n19744,
    new_n19745, new_n19746, new_n19747, new_n19748, new_n19749_1,
    new_n19750, new_n19751, new_n19752, new_n19753, new_n19754, new_n19755,
    new_n19756_1, new_n19757, new_n19758, new_n19759, new_n19760,
    new_n19761, new_n19762, new_n19763, new_n19764, new_n19765, new_n19766,
    new_n19767_1, new_n19768, new_n19769, new_n19770_1, new_n19771,
    new_n19772, new_n19773, new_n19774, new_n19775, new_n19776, new_n19777,
    new_n19778, new_n19779, new_n19780_1, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789_1, new_n19790, new_n19791, new_n19792_1, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798_1,
    new_n19801, new_n19802, new_n19803_1, new_n19804, new_n19805,
    new_n19806, new_n19807, new_n19808, new_n19809, new_n19810, new_n19811,
    new_n19812, new_n19813, new_n19814, new_n19815, new_n19816, new_n19817,
    new_n19818, new_n19820, new_n19821, new_n19822, new_n19823, new_n19824,
    new_n19825, new_n19826, new_n19827, new_n19828, new_n19829, new_n19830,
    new_n19831, new_n19832, new_n19833, new_n19834, new_n19835, new_n19836,
    new_n19837, new_n19838, new_n19839, new_n19840, new_n19841, new_n19842,
    new_n19844, new_n19845, new_n19846, new_n19847, new_n19848, new_n19849,
    new_n19850, new_n19851, new_n19852, new_n19853, new_n19854, new_n19855,
    new_n19856, new_n19857, new_n19858, new_n19859, new_n19860, new_n19861,
    new_n19862, new_n19863, new_n19864, new_n19865, new_n19866, new_n19867,
    new_n19868, new_n19869, new_n19870, new_n19871, new_n19872,
    new_n19873_1, new_n19874, new_n19875, new_n19876, new_n19877,
    new_n19878, new_n19879, new_n19880, new_n19881, new_n19882, new_n19883,
    new_n19884, new_n19885, new_n19889, new_n19890, new_n19891, new_n19892,
    new_n19893, new_n19894, new_n19895, new_n19896, new_n19897, new_n19898,
    new_n19899, new_n19900, new_n19901, new_n19902, new_n19903, new_n19904,
    new_n19905_1, new_n19906, new_n19907, new_n19908, new_n19909_1,
    new_n19910, new_n19911_1, new_n19912, new_n19913, new_n19914,
    new_n19915, new_n19916_1, new_n19917, new_n19918, new_n19919,
    new_n19920, new_n19921, new_n19922_1, new_n19923_1, new_n19924,
    new_n19925, new_n19926, new_n19927, new_n19928, new_n19929,
    new_n19930_1, new_n19931, new_n19932, new_n19933, new_n19934,
    new_n19935, new_n19936, new_n19937, new_n19938, new_n19939, new_n19940,
    new_n19942, new_n19943, new_n19944, new_n19945, new_n19946, new_n19947,
    new_n19948, new_n19949, new_n19950, new_n19951, new_n19952, new_n19953,
    new_n19954, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959,
    new_n19960, new_n19961, new_n19962, new_n19963, new_n19964, new_n19965,
    new_n19966, new_n19967, new_n19968_1, new_n19970, new_n19971,
    new_n19972, new_n19973, new_n19974, new_n19975, new_n19976, new_n19977,
    new_n19978, new_n19979, new_n19980, new_n19981, new_n19982, new_n19983,
    new_n19984, new_n19985, new_n19986, new_n19991, new_n19992, new_n19993,
    new_n19994, new_n19995, new_n19996, new_n19997, new_n19998, new_n19999,
    new_n20000, new_n20003, new_n20004_1, new_n20005, new_n20006,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013_1, new_n20014, new_n20015, new_n20016, new_n20017_1,
    new_n20018, new_n20019, new_n20020, new_n20021, new_n20022, new_n20023,
    new_n20024, new_n20025, new_n20026, new_n20027, new_n20028, new_n20029,
    new_n20030, new_n20031, new_n20032, new_n20033_1, new_n20034,
    new_n20035, new_n20036_1, new_n20037, new_n20038, new_n20039,
    new_n20040_1, new_n20041, new_n20042, new_n20043, new_n20044,
    new_n20045, new_n20046, new_n20047, new_n20048, new_n20049, new_n20050,
    new_n20051, new_n20052, new_n20053, new_n20054, new_n20055, new_n20056,
    new_n20057, new_n20058, new_n20059, new_n20060, new_n20061_1,
    new_n20062, new_n20063, new_n20064, new_n20065, new_n20066, new_n20067,
    new_n20068, new_n20073, new_n20074, new_n20075, new_n20076,
    new_n20077_1, new_n20078, new_n20079, new_n20080, new_n20081,
    new_n20082, new_n20083, new_n20084, new_n20085, new_n20086_1,
    new_n20087, new_n20088, new_n20089, new_n20090, new_n20091, new_n20092,
    new_n20093, new_n20094, new_n20095, new_n20096_1, new_n20097,
    new_n20098, new_n20099, new_n20103_1, new_n20104, new_n20105,
    new_n20106, new_n20107, new_n20108, new_n20109, new_n20110, new_n20111,
    new_n20112, new_n20113, new_n20114, new_n20115, new_n20116, new_n20117,
    new_n20118, new_n20119, new_n20120, new_n20121, new_n20122, new_n20123,
    new_n20124, new_n20125, new_n20126_1, new_n20127, new_n20128,
    new_n20129, new_n20130, new_n20131, new_n20132, new_n20133, new_n20134,
    new_n20135, new_n20136, new_n20137, new_n20138_1, new_n20139,
    new_n20140, new_n20141, new_n20142, new_n20143, new_n20144, new_n20145,
    new_n20146, new_n20147, new_n20148, new_n20149_1, new_n20150,
    new_n20151_1, new_n20152, new_n20153, new_n20154, new_n20155,
    new_n20156, new_n20157, new_n20158, new_n20159, new_n20160, new_n20161,
    new_n20162, new_n20163, new_n20164, new_n20165, new_n20166, new_n20167,
    new_n20168, new_n20169_1, new_n20170, new_n20171, new_n20172,
    new_n20173, new_n20174, new_n20175, new_n20176, new_n20177, new_n20178,
    new_n20179_1, new_n20180, new_n20181, new_n20182, new_n20183,
    new_n20184, new_n20185, new_n20186, new_n20187_1, new_n20188,
    new_n20189, new_n20190, new_n20191, new_n20192, new_n20193, new_n20194,
    new_n20195, new_n20196, new_n20197, new_n20198, new_n20199, new_n20200,
    new_n20201, new_n20202, new_n20203, new_n20204, new_n20212,
    new_n20213_1, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229,
    new_n20230, new_n20231, new_n20232, new_n20233, new_n20234,
    new_n20235_1, new_n20236, new_n20237, new_n20238, new_n20239,
    new_n20240, new_n20241, new_n20242, new_n20243, new_n20244, new_n20245,
    new_n20246, new_n20247, new_n20248, new_n20249, new_n20250_1,
    new_n20251, new_n20252, new_n20256, new_n20257, new_n20258,
    new_n20259_1, new_n20260, new_n20261, new_n20262, new_n20263,
    new_n20264, new_n20265, new_n20266, new_n20267, new_n20268, new_n20269,
    new_n20270, new_n20271, new_n20272, new_n20273, new_n20274, new_n20275,
    new_n20276, new_n20277, new_n20278, new_n20279_1, new_n20280,
    new_n20281, new_n20282, new_n20283, new_n20284, new_n20285, new_n20286,
    new_n20287_1, new_n20288, new_n20289, new_n20290, new_n20291,
    new_n20292, new_n20293, new_n20294, new_n20295, new_n20296, new_n20297,
    new_n20298, new_n20299, new_n20300, new_n20301_1, new_n20302,
    new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308,
    new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314,
    new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320,
    new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326,
    new_n20327, new_n20328, new_n20329, new_n20330_1, new_n20331,
    new_n20332, new_n20333_1, new_n20334, new_n20335, new_n20336,
    new_n20337, new_n20338, new_n20339, new_n20340, new_n20341, new_n20342,
    new_n20343, new_n20344, new_n20346, new_n20347, new_n20348,
    new_n20349_1, new_n20350, new_n20351, new_n20352, new_n20353,
    new_n20354, new_n20355_1, new_n20356, new_n20360, new_n20361,
    new_n20362, new_n20363, new_n20364, new_n20365, new_n20366_1,
    new_n20367, new_n20368, new_n20369, new_n20370, new_n20371, new_n20372,
    new_n20373, new_n20374, new_n20375, new_n20376, new_n20377, new_n20378,
    new_n20379, new_n20380, new_n20381, new_n20382, new_n20383, new_n20384,
    new_n20385_1, new_n20386, new_n20388_1, new_n20389, new_n20390,
    new_n20391, new_n20392, new_n20393, new_n20394, new_n20395, new_n20396,
    new_n20397, new_n20398, new_n20399, new_n20400, new_n20401,
    new_n20402_1, new_n20403_1, new_n20404, new_n20405, new_n20406,
    new_n20407, new_n20408, new_n20409_1, new_n20410, new_n20411_1,
    new_n20412, new_n20413, new_n20414, new_n20415, new_n20416, new_n20417,
    new_n20418, new_n20419, new_n20420, new_n20421, new_n20422, new_n20423,
    new_n20424_1, new_n20425, new_n20426, new_n20427, new_n20428,
    new_n20429_1, new_n20430, new_n20431, new_n20432, new_n20433,
    new_n20434, new_n20435, new_n20436_1, new_n20437, new_n20438,
    new_n20439, new_n20440, new_n20441_1, new_n20442, new_n20443,
    new_n20444, new_n20445_1, new_n20446, new_n20447, new_n20448,
    new_n20449, new_n20450_1, new_n20451, new_n20452, new_n20453,
    new_n20454, new_n20455_1, new_n20456, new_n20457, new_n20458,
    new_n20459, new_n20460, new_n20462, new_n20465, new_n20466, new_n20467,
    new_n20468, new_n20469, new_n20470_1, new_n20471, new_n20472,
    new_n20473, new_n20474, new_n20475, new_n20476, new_n20477,
    new_n20478_1, new_n20479, new_n20480, new_n20481, new_n20482,
    new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489_1, new_n20490_1, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495_1, new_n20496, new_n20497, new_n20498,
    new_n20499, new_n20500, new_n20501, new_n20502, new_n20503, new_n20504,
    new_n20505, new_n20506, new_n20507, new_n20508, new_n20509, new_n20510,
    new_n20511, new_n20512, new_n20513, new_n20514, new_n20515_1,
    new_n20516, new_n20517, new_n20518, new_n20519, new_n20520, new_n20521,
    new_n20522, new_n20523, new_n20524, new_n20525, new_n20526, new_n20527,
    new_n20528, new_n20529, new_n20530, new_n20531, new_n20532,
    new_n20533_1, new_n20534, new_n20535, new_n20536, new_n20537,
    new_n20538, new_n20539, new_n20540, new_n20541, new_n20542, new_n20543,
    new_n20544, new_n20545, new_n20546, new_n20547, new_n20548, new_n20549,
    new_n20550, new_n20551, new_n20552, new_n20553, new_n20554, new_n20555,
    new_n20556, new_n20557, new_n20558, new_n20559, new_n20560, new_n20561,
    new_n20562, new_n20563, new_n20564, new_n20565, new_n20566, new_n20567,
    new_n20568, new_n20569, new_n20570, new_n20573, new_n20574, new_n20575,
    new_n20576, new_n20577, new_n20578, new_n20579, new_n20580, new_n20581,
    new_n20582_1, new_n20583, new_n20584, new_n20585, new_n20586,
    new_n20587, new_n20588, new_n20589, new_n20590_1, new_n20591,
    new_n20592, new_n20593, new_n20594, new_n20595, new_n20596, new_n20597,
    new_n20598, new_n20599, new_n20600, new_n20601, new_n20602_1,
    new_n20603, new_n20604_1, new_n20605, new_n20606, new_n20607,
    new_n20608, new_n20609_1, new_n20610, new_n20611, new_n20612,
    new_n20613, new_n20614, new_n20615, new_n20616, new_n20617, new_n20618,
    new_n20619, new_n20620, new_n20621, new_n20622, new_n20623_1,
    new_n20624, new_n20625, new_n20626, new_n20627, new_n20628,
    new_n20629_1, new_n20630, new_n20631, new_n20632, new_n20633,
    new_n20634, new_n20635, new_n20636, new_n20637, new_n20638, new_n20639,
    new_n20640, new_n20647, new_n20648, new_n20649, new_n20653, new_n20654,
    new_n20655, new_n20656, new_n20657, new_n20658_1, new_n20659,
    new_n20660, new_n20661_1, new_n20662, new_n20663, new_n20664,
    new_n20665, new_n20666, new_n20667, new_n20668, new_n20669, new_n20670,
    new_n20671, new_n20672, new_n20673_1, new_n20674, new_n20675,
    new_n20676, new_n20677, new_n20678_1, new_n20679, new_n20680_1,
    new_n20681, new_n20682, new_n20683, new_n20684, new_n20685_1,
    new_n20686, new_n20687, new_n20688, new_n20689, new_n20690,
    new_n20691_1, new_n20692, new_n20693, new_n20694, new_n20695,
    new_n20696_1, new_n20697, new_n20698, new_n20699, new_n20700_1,
    new_n20701, new_n20702, new_n20703, new_n20704_1, new_n20705_1,
    new_n20706, new_n20707, new_n20708, new_n20709_1, new_n20710,
    new_n20711, new_n20712, new_n20713_1, new_n20714, new_n20715,
    new_n20716, new_n20717, new_n20718, new_n20719, new_n20720, new_n20721,
    new_n20722_1, new_n20723_1, new_n20724, new_n20725, new_n20726,
    new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732,
    new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738,
    new_n20739, new_n20740, new_n20741, new_n20742, new_n20743, new_n20744,
    new_n20745, new_n20746, new_n20747, new_n20748_1, new_n20749,
    new_n20750, new_n20751, new_n20752, new_n20753, new_n20754, new_n20755,
    new_n20756, new_n20757, new_n20758, new_n20759, new_n20760,
    new_n20761_1, new_n20762, new_n20763, new_n20764, new_n20765,
    new_n20766, new_n20767, new_n20768, new_n20769, new_n20770, new_n20771,
    new_n20772, new_n20773, new_n20774_1, new_n20775, new_n20776,
    new_n20777, new_n20778, new_n20779, new_n20780, new_n20781, new_n20782,
    new_n20783, new_n20784, new_n20785, new_n20786, new_n20787,
    new_n20788_1, new_n20789, new_n20790, new_n20791, new_n20792,
    new_n20795_1, new_n20796, new_n20797, new_n20798, new_n20799,
    new_n20800, new_n20801, new_n20802, new_n20803_1, new_n20804,
    new_n20805, new_n20806, new_n20807, new_n20808, new_n20809, new_n20810,
    new_n20811, new_n20812, new_n20813, new_n20814, new_n20815, new_n20816,
    new_n20817, new_n20818, new_n20819, new_n20820, new_n20821, new_n20822,
    new_n20823, new_n20824, new_n20825, new_n20826_1, new_n20827,
    new_n20828, new_n20829, new_n20830, new_n20831, new_n20832, new_n20833,
    new_n20834, new_n20835, new_n20836, new_n20837, new_n20838, new_n20839,
    new_n20840, new_n20841, new_n20842, new_n20843, new_n20844, new_n20845,
    new_n20846, new_n20847, new_n20848, new_n20849, new_n20850, new_n20851,
    new_n20852, new_n20853, new_n20854, new_n20855, new_n20856, new_n20857,
    new_n20858, new_n20859, new_n20860, new_n20861, new_n20862, new_n20863,
    new_n20864, new_n20865, new_n20866, new_n20867, new_n20868,
    new_n20869_1, new_n20870, new_n20871, new_n20872, new_n20873,
    new_n20874, new_n20875, new_n20876, new_n20877, new_n20878,
    new_n20879_1, new_n20880, new_n20881, new_n20882, new_n20883,
    new_n20884, new_n20889, new_n20890, new_n20891, new_n20892, new_n20893,
    new_n20894, new_n20895, new_n20896, new_n20897, new_n20898, new_n20899,
    new_n20900, new_n20901, new_n20902, new_n20903, new_n20904, new_n20905,
    new_n20906, new_n20907, new_n20908, new_n20909, new_n20910, new_n20911,
    new_n20912, new_n20913, new_n20914, new_n20915_1, new_n20916,
    new_n20917, new_n20918, new_n20919, new_n20920, new_n20921, new_n20922,
    new_n20923_1, new_n20924, new_n20925, new_n20926, new_n20927,
    new_n20928, new_n20929_1, new_n20930, new_n20931, new_n20932,
    new_n20933, new_n20934, new_n20935_1, new_n20936_1, new_n20937,
    new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943,
    new_n20944, new_n20945, new_n20946_1, new_n20947, new_n20948,
    new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20954,
    new_n20955, new_n20956, new_n20957, new_n20958, new_n20959, new_n20960,
    new_n20961, new_n20962, new_n20963, new_n20964, new_n20965, new_n20966,
    new_n20967, new_n20968, new_n20969, new_n20970, new_n20971, new_n20972,
    new_n20973, new_n20974, new_n20975, new_n20976, new_n20977, new_n20978,
    new_n20979, new_n20980, new_n20981, new_n20982, new_n20983, new_n20984,
    new_n20985, new_n20986_1, new_n20987, new_n20988, new_n20989,
    new_n20990, new_n20992, new_n20993, new_n20994, new_n20995, new_n20996,
    new_n20997, new_n20998, new_n20999, new_n21000, new_n21002, new_n21003,
    new_n21004, new_n21005, new_n21006, new_n21007, new_n21008_1,
    new_n21009, new_n21010, new_n21011, new_n21012, new_n21013, new_n21014,
    new_n21015, new_n21016, new_n21017_1, new_n21018, new_n21019,
    new_n21020, new_n21021, new_n21022, new_n21023, new_n21024, new_n21025,
    new_n21026, new_n21027, new_n21028, new_n21035, new_n21036, new_n21037,
    new_n21038, new_n21039, new_n21040, new_n21041, new_n21042, new_n21043,
    new_n21044, new_n21045, new_n21046_1, new_n21047, new_n21048,
    new_n21049, new_n21050, new_n21051, new_n21052, new_n21053, new_n21054,
    new_n21066, new_n21067, new_n21068, new_n21069, new_n21070, new_n21071,
    new_n21072, new_n21073, new_n21074, new_n21075, new_n21076, new_n21077,
    new_n21078_1, new_n21079, new_n21080, new_n21081, new_n21082,
    new_n21083, new_n21084, new_n21085, new_n21086, new_n21087, new_n21088,
    new_n21089, new_n21090, new_n21091, new_n21092, new_n21093_1,
    new_n21094_1, new_n21095_1, new_n21096, new_n21097, new_n21098,
    new_n21099, new_n21100, new_n21101, new_n21102, new_n21103, new_n21104,
    new_n21105, new_n21107, new_n21108, new_n21109, new_n21110, new_n21111,
    new_n21112, new_n21113, new_n21114, new_n21115, new_n21116, new_n21117,
    new_n21118, new_n21119, new_n21120, new_n21121, new_n21122,
    new_n21123_1, new_n21124, new_n21125, new_n21126, new_n21127,
    new_n21128, new_n21129, new_n21130, new_n21131, new_n21132, new_n21133,
    new_n21134_1, new_n21136, new_n21137, new_n21138_1, new_n21139,
    new_n21140, new_n21141, new_n21142, new_n21143, new_n21144, new_n21145,
    new_n21146, new_n21147, new_n21148, new_n21149, new_n21150, new_n21151,
    new_n21152, new_n21153, new_n21154_1, new_n21155, new_n21156,
    new_n21157_1, new_n21158, new_n21159, new_n21160, new_n21161,
    new_n21162, new_n21163, new_n21164, new_n21165, new_n21166, new_n21167,
    new_n21168_1, new_n21169, new_n21170, new_n21171, new_n21172,
    new_n21173_1, new_n21174, new_n21175, new_n21176_1, new_n21177,
    new_n21178, new_n21179, new_n21180, new_n21181, new_n21182_1,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193_1,
    new_n21194, new_n21195, new_n21196, new_n21197, new_n21198, new_n21199,
    new_n21200, new_n21201, new_n21202, new_n21203_1, new_n21204,
    new_n21205, new_n21206, new_n21207, new_n21208, new_n21209, new_n21210,
    new_n21211, new_n21212, new_n21213, new_n21214, new_n21215, new_n21216,
    new_n21217, new_n21218, new_n21219, new_n21220, new_n21221,
    new_n21222_1, new_n21223, new_n21224, new_n21225_1, new_n21226_1,
    new_n21227, new_n21228, new_n21229, new_n21230, new_n21231, new_n21232,
    new_n21233, new_n21234, new_n21235, new_n21236, new_n21237,
    new_n21238_1, new_n21239, new_n21240, new_n21241, new_n21242,
    new_n21243, new_n21244, new_n21245, new_n21246, new_n21247, new_n21248,
    new_n21249, new_n21250, new_n21251, new_n21252, new_n21253,
    new_n21254_1, new_n21255, new_n21256, new_n21257, new_n21258,
    new_n21259, new_n21260, new_n21261, new_n21262, new_n21263, new_n21264,
    new_n21265, new_n21266, new_n21267, new_n21268, new_n21269, new_n21270,
    new_n21271, new_n21272, new_n21273, new_n21274, new_n21275,
    new_n21276_1, new_n21277, new_n21278, new_n21279, new_n21280,
    new_n21281, new_n21282, new_n21283, new_n21284, new_n21285, new_n21286,
    new_n21287_1, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298_1, new_n21299, new_n21300, new_n21301, new_n21302_1,
    new_n21303, new_n21304, new_n21305, new_n21306, new_n21307, new_n21308,
    new_n21309, new_n21310, new_n21311, new_n21312, new_n21313, new_n21314,
    new_n21315, new_n21316, new_n21321, new_n21322, new_n21323, new_n21324,
    new_n21325, new_n21326, new_n21327, new_n21328, new_n21329, new_n21330,
    new_n21331, new_n21332, new_n21333, new_n21334, new_n21335, new_n21336,
    new_n21337, new_n21338, new_n21339, new_n21340, new_n21341, new_n21342,
    new_n21345, new_n21346, new_n21347, new_n21348, new_n21349_1,
    new_n21350, new_n21351, new_n21352, new_n21353, new_n21354, new_n21355,
    new_n21356, new_n21357, new_n21358, new_n21359, new_n21360, new_n21361,
    new_n21362, new_n21363, new_n21364, new_n21365_1, new_n21366,
    new_n21367_1, new_n21368, new_n21369, new_n21372, new_n21373,
    new_n21374, new_n21375, new_n21376, new_n21377, new_n21378, new_n21379,
    new_n21380, new_n21381, new_n21386, new_n21387, new_n21391, new_n21392,
    new_n21393, new_n21394, new_n21395, new_n21396_1, new_n21397,
    new_n21398_1, new_n21399_1, new_n21400, new_n21401, new_n21402,
    new_n21403, new_n21404_1, new_n21405, new_n21406, new_n21407,
    new_n21408, new_n21409, new_n21413, new_n21414, new_n21415, new_n21416,
    new_n21417, new_n21418, new_n21419, new_n21420, new_n21421, new_n21422,
    new_n21424, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429,
    new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435,
    new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441,
    new_n21442, new_n21443, new_n21445, new_n21446_1, new_n21447,
    new_n21448, new_n21449, new_n21450, new_n21451, new_n21452, new_n21453,
    new_n21454, new_n21455, new_n21456, new_n21457, new_n21458, new_n21459,
    new_n21460, new_n21461, new_n21462, new_n21463, new_n21464, new_n21465,
    new_n21466, new_n21467, new_n21468, new_n21469, new_n21470,
    new_n21471_1, new_n21472_1, new_n21473, new_n21474, new_n21475,
    new_n21476, new_n21477, new_n21478, new_n21479, new_n21480, new_n21481,
    new_n21482, new_n21483, new_n21484, new_n21485, new_n21486, new_n21487,
    new_n21488, new_n21490, new_n21491, new_n21492, new_n21493, new_n21494,
    new_n21495, new_n21496, new_n21497, new_n21498, new_n21499, new_n21500,
    new_n21501, new_n21502, new_n21503, new_n21504, new_n21505, new_n21506,
    new_n21507, new_n21508, new_n21509, new_n21510, new_n21511, new_n21512,
    new_n21513, new_n21514, new_n21515, new_n21516, new_n21517, new_n21518,
    new_n21519, new_n21520, new_n21521, new_n21522, new_n21523, new_n21524,
    new_n21525_1, new_n21526, new_n21527, new_n21528, new_n21529,
    new_n21530, new_n21531, new_n21532, new_n21533, new_n21534, new_n21535,
    new_n21536, new_n21537, new_n21538_1, new_n21539, new_n21540,
    new_n21541, new_n21542, new_n21543, new_n21544, new_n21545, new_n21546,
    new_n21547, new_n21548, new_n21549_1, new_n21550, new_n21551,
    new_n21552, new_n21553, new_n21554, new_n21555, new_n21556, new_n21557,
    new_n21558, new_n21559, new_n21560, new_n21561, new_n21562, new_n21563,
    new_n21564, new_n21565, new_n21566, new_n21571, new_n21572, new_n21573,
    new_n21574, new_n21575, new_n21576, new_n21577, new_n21578, new_n21579,
    new_n21580, new_n21581, new_n21582, new_n21583, new_n21584, new_n21585,
    new_n21586, new_n21587, new_n21588, new_n21589, new_n21590, new_n21591,
    new_n21592, new_n21593, new_n21594, new_n21595, new_n21596, new_n21597,
    new_n21598, new_n21599_1, new_n21600, new_n21601, new_n21602,
    new_n21603, new_n21604, new_n21605, new_n21606, new_n21607, new_n21608,
    new_n21609, new_n21610, new_n21611, new_n21612, new_n21613, new_n21614,
    new_n21615_1, new_n21616, new_n21617, new_n21618, new_n21619,
    new_n21620, new_n21621, new_n21622, new_n21623, new_n21624, new_n21625,
    new_n21626, new_n21627, new_n21628_1, new_n21629, new_n21630,
    new_n21631, new_n21632, new_n21633, new_n21634, new_n21635, new_n21636,
    new_n21637_1, new_n21638, new_n21639, new_n21640, new_n21641,
    new_n21642, new_n21643, new_n21644, new_n21645_1, new_n21646,
    new_n21647, new_n21648, new_n21649_1, new_n21650, new_n21651,
    new_n21652, new_n21653, new_n21654_1, new_n21655, new_n21656,
    new_n21657, new_n21658, new_n21659, new_n21660, new_n21661, new_n21662,
    new_n21663, new_n21664, new_n21665_1, new_n21666, new_n21667,
    new_n21668, new_n21669, new_n21670, new_n21671, new_n21672, new_n21673,
    new_n21674_1, new_n21675, new_n21676, new_n21677, new_n21678,
    new_n21679, new_n21680_1, new_n21681, new_n21682, new_n21683,
    new_n21684, new_n21685_1, new_n21686, new_n21687_1, new_n21688,
    new_n21689, new_n21690, new_n21691, new_n21692, new_n21694, new_n21695,
    new_n21696, new_n21701, new_n21704, new_n21705, new_n21706, new_n21707,
    new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713,
    new_n21714, new_n21715, new_n21716, new_n21717_1, new_n21718,
    new_n21719_1, new_n21720, new_n21721, new_n21722, new_n21723,
    new_n21724, new_n21725, new_n21726, new_n21727, new_n21728, new_n21729,
    new_n21730, new_n21731, new_n21732, new_n21733, new_n21734,
    new_n21735_1, new_n21736, new_n21737, new_n21738, new_n21739,
    new_n21740, new_n21741, new_n21743, new_n21744, new_n21745, new_n21746,
    new_n21747, new_n21748, new_n21749_1, new_n21750_1, new_n21751,
    new_n21752, new_n21753_1, new_n21754, new_n21755, new_n21756,
    new_n21757, new_n21758, new_n21759, new_n21760, new_n21761, new_n21762,
    new_n21763, new_n21764, new_n21765_1, new_n21766, new_n21767,
    new_n21768, new_n21769, new_n21770, new_n21771, new_n21772, new_n21773,
    new_n21774, new_n21775, new_n21776, new_n21777, new_n21786, new_n21787,
    new_n21788, new_n21789, new_n21790, new_n21791, new_n21792, new_n21793,
    new_n21794, new_n21795, new_n21796, new_n21797, new_n21798, new_n21799,
    new_n21803, new_n21804, new_n21805, new_n21806, new_n21807, new_n21808,
    new_n21809, new_n21810, new_n21811, new_n21812, new_n21813, new_n21814,
    new_n21815, new_n21816, new_n21817, new_n21818, new_n21819,
    new_n21820_1, new_n21821, new_n21822, new_n21823, new_n21824,
    new_n21825, new_n21826, new_n21827, new_n21828, new_n21829, new_n21830,
    new_n21831, new_n21832_1, new_n21833, new_n21834, new_n21835,
    new_n21836, new_n21837, new_n21838, new_n21839_1, new_n21840,
    new_n21843, new_n21844, new_n21845, new_n21846, new_n21847, new_n21848,
    new_n21849, new_n21850, new_n21851, new_n21852, new_n21853, new_n21854,
    new_n21855, new_n21856, new_n21857, new_n21858, new_n21859, new_n21860,
    new_n21861, new_n21862, new_n21863, new_n21864, new_n21865, new_n21866,
    new_n21867, new_n21868, new_n21869, new_n21870, new_n21871, new_n21872,
    new_n21873, new_n21874_1, new_n21875, new_n21876, new_n21877,
    new_n21878, new_n21879, new_n21880, new_n21881, new_n21882, new_n21883,
    new_n21884, new_n21885, new_n21886, new_n21887, new_n21888, new_n21889,
    new_n21890, new_n21891, new_n21892, new_n21893, new_n21894, new_n21895,
    new_n21896, new_n21897, new_n21898_1, new_n21899, new_n21900,
    new_n21901, new_n21902, new_n21903, new_n21904, new_n21905_1,
    new_n21906, new_n21907, new_n21908, new_n21909, new_n21910, new_n21911,
    new_n21912, new_n21914, new_n21915_1, new_n21916, new_n21917,
    new_n21918, new_n21919, new_n21920, new_n21921, new_n21922, new_n21923,
    new_n21924, new_n21925, new_n21926, new_n21927, new_n21928, new_n21929,
    new_n21930, new_n21931, new_n21932, new_n21933, new_n21934_1,
    new_n21935, new_n21936, new_n21937, new_n21938, new_n21939, new_n21940,
    new_n21941, new_n21942, new_n21943_1, new_n21944, new_n21945,
    new_n21947, new_n21948, new_n21950, new_n21951, new_n21952, new_n21953,
    new_n21954, new_n21955, new_n21956, new_n21957_1, new_n21958,
    new_n21959, new_n21960_1, new_n21961, new_n21962, new_n21963,
    new_n21964, new_n21965, new_n21966, new_n21967, new_n21968, new_n21969,
    new_n21970, new_n21971, new_n21972, new_n21973, new_n21974, new_n21975,
    new_n21976_1, new_n21977, new_n21978, new_n21979, new_n21980,
    new_n21981_1, new_n21982, new_n21983, new_n21984, new_n21985,
    new_n21986_1, new_n21987, new_n21988, new_n21989, new_n21990,
    new_n21991, new_n21992, new_n21995, new_n21996, new_n21999, new_n22000,
    new_n22001, new_n22002, new_n22003, new_n22004, new_n22005, new_n22006,
    new_n22007, new_n22008, new_n22009, new_n22010, new_n22011, new_n22012,
    new_n22013, new_n22014, new_n22015, new_n22016_1, new_n22017,
    new_n22018, new_n22019, new_n22020, new_n22021, new_n22022, new_n22023,
    new_n22024, new_n22025, new_n22026, new_n22027_1, new_n22028,
    new_n22029, new_n22030, new_n22031, new_n22032, new_n22033, new_n22034,
    new_n22035, new_n22036, new_n22037, new_n22038, new_n22039, new_n22042,
    new_n22043_1, new_n22044, new_n22045, new_n22046, new_n22047,
    new_n22048, new_n22049, new_n22050_1, new_n22051, new_n22052,
    new_n22053, new_n22054, new_n22055, new_n22056, new_n22057, new_n22058,
    new_n22059, new_n22060, new_n22061, new_n22062, new_n22063_1,
    new_n22064, new_n22065, new_n22066, new_n22074, new_n22075,
    new_n22076_1, new_n22077, new_n22078, new_n22079, new_n22080,
    new_n22081, new_n22082, new_n22083, new_n22084, new_n22085, new_n22086,
    new_n22087, new_n22088, new_n22089, new_n22090_1, new_n22091,
    new_n22092, new_n22093, new_n22094, new_n22095, new_n22096, new_n22097,
    new_n22098, new_n22099, new_n22100, new_n22101, new_n22102, new_n22103,
    new_n22104, new_n22105, new_n22106, new_n22107_1, new_n22108,
    new_n22109, new_n22110, new_n22111, new_n22112, new_n22113_1,
    new_n22114, new_n22115, new_n22116, new_n22117, new_n22118, new_n22119,
    new_n22120, new_n22121, new_n22122, new_n22123, new_n22124_1,
    new_n22125, new_n22126_1, new_n22127, new_n22128, new_n22129,
    new_n22130_1, new_n22131, new_n22132, new_n22133, new_n22134,
    new_n22135, new_n22136, new_n22137, new_n22147, new_n22148, new_n22149,
    new_n22150_1, new_n22151, new_n22152, new_n22153, new_n22154,
    new_n22155, new_n22156, new_n22157_1, new_n22173_1, new_n22175,
    new_n22176, new_n22177, new_n22178, new_n22179, new_n22180, new_n22181,
    new_n22182, new_n22183, new_n22184, new_n22185, new_n22186, new_n22187,
    new_n22188, new_n22189, new_n22190, new_n22191, new_n22192, new_n22193,
    new_n22194, new_n22195, new_n22196, new_n22197, new_n22199, new_n22200,
    new_n22201_1, new_n22202, new_n22203, new_n22204, new_n22205,
    new_n22206, new_n22207, new_n22208, new_n22209, new_n22210, new_n22211,
    new_n22212, new_n22213_1, new_n22214, new_n22215, new_n22216,
    new_n22218, new_n22219, new_n22220, new_n22221, new_n22222, new_n22223,
    new_n22224, new_n22225, new_n22226, new_n22227, new_n22228, new_n22229,
    new_n22230, new_n22231, new_n22232, new_n22233, new_n22234, new_n22235,
    new_n22240, new_n22241, new_n22242, new_n22243, new_n22244, new_n22245,
    new_n22246, new_n22247, new_n22248, new_n22249, new_n22250, new_n22251,
    new_n22252, new_n22253_1, new_n22254, new_n22255, new_n22256,
    new_n22257, new_n22258, new_n22259, new_n22260, new_n22269,
    new_n22270_1, new_n22271, new_n22272, new_n22273, new_n22274_1,
    new_n22275, new_n22276, new_n22277, new_n22283_1, new_n22284,
    new_n22285, new_n22286, new_n22287, new_n22288, new_n22289,
    new_n22290_1, new_n22291, new_n22296, new_n22302, new_n22303,
    new_n22304, new_n22305, new_n22306, new_n22307, new_n22308,
    new_n22309_1, new_n22310, new_n22311_1, new_n22312, new_n22313,
    new_n22314, new_n22315, new_n22316, new_n22317_1, new_n22318,
    new_n22319, new_n22320, new_n22325, new_n22326, new_n22327, new_n22328,
    new_n22329, new_n22330, new_n22331, new_n22332_1, new_n22339,
    new_n22340, new_n22341_1, new_n22342, new_n22343, new_n22344,
    new_n22345, new_n22346, new_n22347, new_n22348, new_n22349, new_n22350,
    new_n22351, new_n22352, new_n22353_1, new_n22354, new_n22355,
    new_n22356, new_n22357, new_n22358_1, new_n22359_1, new_n22360,
    new_n22361, new_n22362, new_n22363, new_n22364, new_n22365, new_n22366,
    new_n22367, new_n22368, new_n22369, new_n22370, new_n22371, new_n22372,
    new_n22373, new_n22374, new_n22375, new_n22376, new_n22377, new_n22378,
    new_n22379_1, new_n22380, new_n22381, new_n22382, new_n22383,
    new_n22384, new_n22385, new_n22386, new_n22389, new_n22390, new_n22391,
    new_n22392, new_n22393, new_n22394, new_n22395, new_n22396, new_n22397,
    new_n22398, new_n22399, new_n22401, new_n22402, new_n22403, new_n22404,
    new_n22405, new_n22406, new_n22407, new_n22408, new_n22409, new_n22410,
    new_n22411, new_n22412, new_n22413, new_n22414, new_n22415, new_n22416,
    new_n22417, new_n22427, new_n22428, new_n22429, new_n22430, new_n22431,
    new_n22432, new_n22433_1, new_n22434, new_n22435, new_n22436,
    new_n22437, new_n22438, new_n22439, new_n22440, new_n22441,
    new_n22442_1, new_n22443, new_n22444_1, new_n22445, new_n22446,
    new_n22447, new_n22448, new_n22449, new_n22450, new_n22451, new_n22452,
    new_n22453, new_n22454, new_n22455, new_n22456, new_n22462, new_n22463,
    new_n22464, new_n22465, new_n22475, new_n22476, new_n22477, new_n22478,
    new_n22479, new_n22480, new_n22481, new_n22482, new_n22483,
    new_n22484_1, new_n22485, new_n22486, new_n22487, new_n22488,
    new_n22489_1, new_n22490, new_n22491, new_n22492_1, new_n22493,
    new_n22494_1, new_n22495, new_n22496, new_n22497, new_n22498,
    new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504,
    new_n22505, new_n22506, new_n22507, new_n22508, new_n22509, new_n22510,
    new_n22511, new_n22512, new_n22513, new_n22514, new_n22515, new_n22516,
    new_n22517, new_n22518, new_n22519, new_n22520, new_n22521, new_n22522,
    new_n22523, new_n22524, new_n22525, new_n22526, new_n22527, new_n22528,
    new_n22529, new_n22530, new_n22531, new_n22532, new_n22533_1,
    new_n22534, new_n22535, new_n22536, new_n22537, new_n22538, new_n22539,
    new_n22540, new_n22541, new_n22542, new_n22543, new_n22544, new_n22545,
    new_n22546, new_n22547, new_n22548, new_n22549, new_n22550, new_n22551,
    new_n22552, new_n22553, new_n22554_1, new_n22555, new_n22556,
    new_n22558, new_n22559, new_n22560, new_n22561, new_n22562, new_n22563,
    new_n22564, new_n22565, new_n22566, new_n22567, new_n22568, new_n22569,
    new_n22570, new_n22571, new_n22572, new_n22573, new_n22574, new_n22575,
    new_n22576, new_n22577, new_n22578, new_n22579, new_n22580, new_n22581,
    new_n22582, new_n22583, new_n22584_1, new_n22585, new_n22586,
    new_n22587, new_n22588_1, new_n22589_1, new_n22590, new_n22591_1,
    new_n22592, new_n22593, new_n22594, new_n22595, new_n22596,
    new_n22597_1, new_n22598, new_n22599, new_n22600, new_n22601,
    new_n22602, new_n22603, new_n22604, new_n22605, new_n22606, new_n22607,
    new_n22608, new_n22609, new_n22610, new_n22611, new_n22612, new_n22613,
    new_n22614, new_n22615, new_n22616, new_n22617, new_n22618,
    new_n22619_1, new_n22620_1, new_n22621, new_n22622, new_n22623_1,
    new_n22624, new_n22625, new_n22626_1, new_n22627, new_n22628,
    new_n22631_1, new_n22632, new_n22633, new_n22634, new_n22635,
    new_n22636, new_n22637, new_n22638, new_n22639, new_n22640, new_n22641,
    new_n22642, new_n22643, new_n22644, new_n22650, new_n22651, new_n22652,
    new_n22653, new_n22654, new_n22655, new_n22656, new_n22657, new_n22658,
    new_n22659, new_n22660_1, new_n22661, new_n22662, new_n22663,
    new_n22664, new_n22665, new_n22666, new_n22667, new_n22668, new_n22669,
    new_n22670, new_n22671, new_n22672, new_n22673, new_n22674, new_n22675,
    new_n22676, new_n22677, new_n22678, new_n22679, new_n22680, new_n22681,
    new_n22682, new_n22683, new_n22684, new_n22685, new_n22686, new_n22687,
    new_n22688, new_n22689, new_n22690, new_n22691, new_n22692, new_n22693,
    new_n22694, new_n22695, new_n22696, new_n22697_1, new_n22698,
    new_n22699, new_n22700, new_n22701, new_n22702, new_n22703, new_n22704,
    new_n22705, new_n22706, new_n22707, new_n22708, new_n22709, new_n22710,
    new_n22711, new_n22712, new_n22713, new_n22714_1, new_n22715,
    new_n22716, new_n22717, new_n22718, new_n22719, new_n22720, new_n22721,
    new_n22722, new_n22724, new_n22725, new_n22726, new_n22727, new_n22728,
    new_n22729, new_n22730, new_n22731, new_n22732, new_n22733, new_n22736,
    new_n22737, new_n22738, new_n22739, new_n22740, new_n22741, new_n22742,
    new_n22743, new_n22744, new_n22745, new_n22751, new_n22752, new_n22753,
    new_n22754, new_n22755, new_n22756, new_n22757, new_n22758, new_n22759,
    new_n22760, new_n22761_1, new_n22762, new_n22763, new_n22764_1,
    new_n22765, new_n22766, new_n22767, new_n22768, new_n22769, new_n22770,
    new_n22771, new_n22772, new_n22773, new_n22774, new_n22775, new_n22776,
    new_n22777, new_n22778, new_n22779_1, new_n22780, new_n22781,
    new_n22782, new_n22783, new_n22784, new_n22785, new_n22786,
    new_n22787_1, new_n22788, new_n22789, new_n22790, new_n22791,
    new_n22792, new_n22793_1, new_n22794, new_n22795, new_n22796,
    new_n22797, new_n22798, new_n22799, new_n22800, new_n22801, new_n22802,
    new_n22803, new_n22804, new_n22805, new_n22806, new_n22807, new_n22808,
    new_n22809, new_n22810, new_n22811, new_n22812, new_n22813, new_n22814,
    new_n22815, new_n22816, new_n22817, new_n22818, new_n22819_1,
    new_n22820, new_n22821, new_n22822, new_n22823, new_n22824, new_n22832,
    new_n22833, new_n22834, new_n22835, new_n22836, new_n22837, new_n22842,
    new_n22845, new_n22847, new_n22848, new_n22849, new_n22850, new_n22851,
    new_n22852, new_n22853, new_n22854, new_n22855, new_n22856, new_n22857,
    new_n22858_1, new_n22859, new_n22860, new_n22861, new_n22862,
    new_n22863, new_n22864, new_n22865, new_n22866, new_n22867, new_n22868,
    new_n22869, new_n22870_1, new_n22871_1, new_n22872, new_n22873,
    new_n22874, new_n22875, new_n22876, new_n22877, new_n22878,
    new_n22879_1, new_n22880, new_n22881, new_n22882, new_n22883,
    new_n22884, new_n22885, new_n22886, new_n22887, new_n22888, new_n22889,
    new_n22890, new_n22891_1, new_n22892, new_n22893, new_n22894,
    new_n22895, new_n22896, new_n22897_1, new_n22898, new_n22899,
    new_n22900, new_n22901, new_n22902, new_n22903_1, new_n22906,
    new_n22907_1, new_n22908, new_n22909, new_n22917, new_n22918_1,
    new_n22919, new_n22920, new_n22921, new_n22922, new_n22923, new_n22924,
    new_n22925, new_n22926, new_n22930, new_n22938, new_n22939_1,
    new_n22940, new_n22941, new_n22942, new_n22943, new_n22944, new_n22945,
    new_n22946, new_n22947, new_n22948, new_n22949, new_n22950, new_n22951,
    new_n22952, new_n22953, new_n22954, new_n22955, new_n22956, new_n22958,
    new_n22959, new_n22960, new_n22961, new_n22962, new_n22963, new_n22964,
    new_n22965, new_n22966, new_n22967, new_n22968, new_n22969, new_n22970,
    new_n22971, new_n22972, new_n22973, new_n22974, new_n22980, new_n22981,
    new_n22982, new_n22983, new_n22984, new_n22985, new_n22986, new_n22987,
    new_n22988, new_n22989, new_n22990, new_n22991, new_n22992, new_n22993,
    new_n22994, new_n22995, new_n22996, new_n22997, new_n22998_1,
    new_n22999, new_n23000, new_n23001, new_n23002, new_n23003, new_n23004,
    new_n23005, new_n23006_1, new_n23007_1, new_n23008, new_n23009_1,
    new_n23012, new_n23013, new_n23014_1, new_n23015, new_n23016,
    new_n23017, new_n23018, new_n23019, new_n23020, new_n23021, new_n23022,
    new_n23023, new_n23024, new_n23025, new_n23026, new_n23027, new_n23028,
    new_n23029, new_n23030, new_n23031, new_n23032, new_n23033,
    new_n23035_1, new_n23036, new_n23037, new_n23038, new_n23039_1,
    new_n23040, new_n23041, new_n23042, new_n23043, new_n23044, new_n23045,
    new_n23046, new_n23047_1, new_n23051, new_n23053, new_n23054,
    new_n23059, new_n23060, new_n23061, new_n23062, new_n23063, new_n23064,
    new_n23065_1, new_n23066_1, new_n23067_1, new_n23068_1, new_n23069,
    new_n23070, new_n23071, new_n23072, new_n23073, new_n23074, new_n23075,
    new_n23076, new_n23077, new_n23078, new_n23079, new_n23080, new_n23081,
    new_n23082, new_n23083, new_n23084, new_n23085, new_n23086, new_n23087,
    new_n23088, new_n23089, new_n23090, new_n23091, new_n23092, new_n23093,
    new_n23094, new_n23095, new_n23096, new_n23097, new_n23098, new_n23099,
    new_n23100, new_n23101, new_n23102, new_n23103, new_n23104, new_n23105,
    new_n23106, new_n23107, new_n23108, new_n23109, new_n23110, new_n23111,
    new_n23113, new_n23114, new_n23115, new_n23116, new_n23117, new_n23118,
    new_n23119, new_n23120_1, new_n23121, new_n23122, new_n23123,
    new_n23124, new_n23125, new_n23126, new_n23127, new_n23128, new_n23129,
    new_n23130, new_n23131, new_n23132, new_n23133, new_n23134, new_n23135,
    new_n23136, new_n23137, new_n23138, new_n23139, new_n23140, new_n23141,
    new_n23142, new_n23143, new_n23144, new_n23145, new_n23146_1,
    new_n23147, new_n23148, new_n23149, new_n23150, new_n23151, new_n23152,
    new_n23153, new_n23154, new_n23155, new_n23156, new_n23157, new_n23158,
    new_n23159, new_n23160_1, new_n23161, new_n23162, new_n23163,
    new_n23164, new_n23165, new_n23166_1, new_n23167, new_n23168,
    new_n23169, new_n23170, new_n23171, new_n23177, new_n23186, new_n23187,
    new_n23188, new_n23189, new_n23195, new_n23202, new_n23203, new_n23204,
    new_n23205, new_n23206, new_n23207, new_n23208, new_n23209, new_n23210,
    new_n23211, new_n23212, new_n23213, new_n23214, new_n23215, new_n23216,
    new_n23217, new_n23218, new_n23219, new_n23220, new_n23221, new_n23222,
    new_n23223, new_n23224, new_n23225, new_n23226, new_n23227, new_n23228,
    new_n23229, new_n23230, new_n23231, new_n23232, new_n23233, new_n23234,
    new_n23235, new_n23236, new_n23237, new_n23238_1, new_n23239,
    new_n23240, new_n23243, new_n23244, new_n23245, new_n23246,
    new_n23247_1, new_n23248_1, new_n23249, new_n23250_1, new_n23251,
    new_n23252, new_n23253, new_n23254, new_n23261, new_n23262, new_n23263,
    new_n23264, new_n23265, new_n23266, new_n23267, new_n23268, new_n23269,
    new_n23270_1, new_n23271, new_n23272_1, new_n23273, new_n23274,
    new_n23275, new_n23276, new_n23277, new_n23278, new_n23279, new_n23280,
    new_n23281, new_n23282, new_n23283, new_n23284, new_n23285, new_n23286,
    new_n23287, new_n23288, new_n23289_1, new_n23290, new_n23291,
    new_n23292, new_n23293, new_n23294, new_n23295, new_n23296, new_n23297,
    new_n23298, new_n23299, new_n23300, new_n23301, new_n23302, new_n23303,
    new_n23304_1, new_n23305_1, new_n23306, new_n23307, new_n23308,
    new_n23309, new_n23310, new_n23311, new_n23312, new_n23313, new_n23314,
    new_n23315, new_n23316, new_n23317, new_n23318, new_n23319, new_n23320,
    new_n23321, new_n23322, new_n23323, new_n23324, new_n23325, new_n23326,
    new_n23327, new_n23328, new_n23329, new_n23330, new_n23331, new_n23332,
    new_n23333_1, new_n23334, new_n23335, new_n23336, new_n23337,
    new_n23338, new_n23339, new_n23340, new_n23341_1, new_n23342_1,
    new_n23343, new_n23344, new_n23345, new_n23346, new_n23347, new_n23348,
    new_n23349, new_n23350, new_n23351, new_n23352, new_n23353, new_n23354,
    new_n23355_1, new_n23356, new_n23357, new_n23358, new_n23359,
    new_n23360, new_n23361, new_n23362, new_n23363, new_n23364, new_n23365,
    new_n23366, new_n23367, new_n23368, new_n23369_1, new_n23370,
    new_n23371_1, new_n23372, new_n23373, new_n23374, new_n23375,
    new_n23376, new_n23377, new_n23378, new_n23379, new_n23380, new_n23381,
    new_n23382, new_n23383, new_n23384, new_n23385, new_n23386, new_n23387,
    new_n23388, new_n23389, new_n23390, new_n23391, new_n23392, new_n23393,
    new_n23394, new_n23395, new_n23399, new_n23402, new_n23403, new_n23404,
    new_n23405, new_n23406, new_n23407, new_n23408, new_n23409, new_n23410,
    new_n23411, new_n23412, new_n23413, new_n23414_1, new_n23415,
    new_n23416, new_n23417, new_n23418, new_n23419, new_n23420, new_n23421,
    new_n23422, new_n23427, new_n23428, new_n23429_1, new_n23430_1,
    new_n23431, new_n23432, new_n23433_1, new_n23434_1, new_n23435,
    new_n23436, new_n23437, new_n23438, new_n23439, new_n23440, new_n23441,
    new_n23442, new_n23443, new_n23444, new_n23445, new_n23446, new_n23447,
    new_n23448, new_n23449, new_n23450_1, new_n23451, new_n23452,
    new_n23453, new_n23455, new_n23456, new_n23457, new_n23458, new_n23459,
    new_n23460, new_n23461, new_n23465, new_n23466, new_n23467, new_n23468,
    new_n23478, new_n23479, new_n23480_1, new_n23481, new_n23482,
    new_n23483, new_n23484, new_n23485, new_n23486, new_n23487, new_n23488,
    new_n23489, new_n23490, new_n23491, new_n23492, new_n23493_1,
    new_n23494, new_n23495, new_n23496, new_n23497, new_n23498, new_n23499,
    new_n23500, new_n23501, new_n23502, new_n23503, new_n23504, new_n23505,
    new_n23526, new_n23527, new_n23528, new_n23529_1, new_n23530,
    new_n23531, new_n23532, new_n23533, new_n23534, new_n23535, new_n23536,
    new_n23537, new_n23538, new_n23539, new_n23540, new_n23541_1,
    new_n23542, new_n23543, new_n23544, new_n23545, new_n23546_1,
    new_n23547, new_n23548, new_n23549, new_n23550_1, new_n23551,
    new_n23552, new_n23553, new_n23554, new_n23555, new_n23556, new_n23557,
    new_n23558, new_n23559, new_n23560, new_n23561, new_n23562, new_n23563,
    new_n23564, new_n23565, new_n23573, new_n23574, new_n23575, new_n23576,
    new_n23577, new_n23578, new_n23579, new_n23580, new_n23581, new_n23582,
    new_n23583, new_n23584, new_n23585_1, new_n23586_1, new_n23587,
    new_n23588_1, new_n23589, new_n23590, new_n23591, new_n23595,
    new_n23596, new_n23599, new_n23600, new_n23601, new_n23602, new_n23603,
    new_n23604, new_n23605, new_n23606, new_n23609, new_n23610, new_n23611,
    new_n23612, new_n23613, new_n23614, new_n23615, new_n23616, new_n23617,
    new_n23618, new_n23619_1, new_n23620, new_n23621, new_n23622,
    new_n23623, new_n23624_1, new_n23625, new_n23626, new_n23627,
    new_n23630, new_n23631, new_n23632, new_n23633, new_n23634, new_n23635,
    new_n23636, new_n23637_1, new_n23638, new_n23639, new_n23640,
    new_n23641, new_n23642, new_n23643, new_n23644, new_n23645, new_n23646,
    new_n23647, new_n23648, new_n23649, new_n23650, new_n23651, new_n23652,
    new_n23653, new_n23654, new_n23655, new_n23656, new_n23657_1,
    new_n23658, new_n23659, new_n23660, new_n23661, new_n23662,
    new_n23663_1, new_n23664, new_n23665, new_n23666, new_n23667,
    new_n23668, new_n23669_1, new_n23670, new_n23671, new_n23672,
    new_n23673, new_n23674, new_n23695, new_n23699, new_n23700, new_n23701,
    new_n23702, new_n23703, new_n23704, new_n23705, new_n23706, new_n23707,
    new_n23708, new_n23709, new_n23710, new_n23711, new_n23712, new_n23715,
    new_n23716, new_n23717_1, new_n23718, new_n23719_1, new_n23720,
    new_n23721, new_n23722, new_n23723, new_n23724, new_n23725, new_n23726,
    new_n23727, new_n23728, new_n23729, new_n23730, new_n23731, new_n23732,
    new_n23733, new_n23734, new_n23738, new_n23739, new_n23740, new_n23741,
    new_n23742, new_n23743, new_n23744, new_n23748_1, new_n23753,
    new_n23754, new_n23755_1, new_n23756, new_n23757, new_n23758,
    new_n23759, new_n23760, new_n23761, new_n23763, new_n23764, new_n23765,
    new_n23766, new_n23767, new_n23768, new_n23769, new_n23770, new_n23771,
    new_n23772, new_n23773, new_n23774, new_n23775_1, new_n23776,
    new_n23777, new_n23778, new_n23779, new_n23780, new_n23781, new_n23802,
    new_n23805, new_n23806, new_n23807, new_n23808, new_n23809, new_n23810,
    new_n23811, new_n23812, new_n23813, new_n23814, new_n23815, new_n23816,
    new_n23817, new_n23818, new_n23819, new_n23820, new_n23821, new_n23822,
    new_n23823, new_n23824, new_n23825, new_n23826, new_n23827, new_n23832,
    new_n23833, new_n23834, new_n23835, new_n23847, new_n23850, new_n23865,
    new_n23866, new_n23867, new_n23868, new_n23869, new_n23870, new_n23884,
    new_n23885, new_n23886, new_n23887, new_n23888_1, new_n23889,
    new_n23890, new_n23891, new_n23895_1, new_n23896, new_n23897,
    new_n23898, new_n23899_1, new_n23900, new_n23901, new_n23902,
    new_n23903_1, new_n23908, new_n23909, new_n23910, new_n23911,
    new_n23912_1, new_n23913_1, new_n23914, new_n23915, new_n23916,
    new_n23919, new_n23920, new_n23921, new_n23936, new_n23937, new_n23938,
    new_n23941, new_n23942_1, new_n23943, new_n23944, new_n23952,
    new_n23953, new_n23962, new_n23972, new_n23973, new_n23974_1,
    new_n23975, new_n23976, new_n23977, new_n23978, new_n23979, new_n23980,
    new_n23981, new_n23990, new_n23991, new_n23992, new_n23993, new_n23994,
    new_n23995, new_n23996, new_n23997, new_n23998, new_n23999, new_n24000,
    new_n24001, new_n24002_1, new_n24003, new_n24004_1, new_n24006,
    new_n24007, new_n24008, new_n24009, new_n24020, new_n24021, new_n24023,
    new_n24024, new_n24025, new_n24026, new_n24027, new_n24028, new_n24029,
    new_n24030, new_n24031, new_n24032_1, new_n24033, new_n24034,
    new_n24035, new_n24036, new_n24054, new_n24055, new_n24056, new_n24057,
    new_n24058, new_n24059, new_n24060, new_n24061, new_n24062, new_n24063,
    new_n24064, new_n24065, new_n24066, new_n24067, new_n24068, new_n24071,
    new_n24072, new_n24073, new_n24078, new_n24079, new_n24080, new_n24081,
    new_n24082, new_n24083, new_n24084, new_n24085_1, new_n24088,
    new_n24089, new_n24090, new_n24091, new_n24092_1, new_n24093_1,
    new_n24094, new_n24097_1, new_n24098, new_n24099, new_n24100,
    new_n24101, new_n24103, new_n24104, new_n24105_1, new_n24106,
    new_n24107, new_n24108, new_n24109, new_n24110, new_n24111, new_n24112,
    new_n24113, new_n24114, new_n24115, new_n24116, new_n24117, new_n24118,
    new_n24119_1, new_n24120, new_n24121, new_n24122, new_n24123,
    new_n24124, new_n24125, new_n24126, new_n24127, new_n24131, new_n24132,
    new_n24133_1, new_n24134, new_n24135, new_n24136, new_n24137,
    new_n24138, new_n24152, new_n24153, new_n24164, new_n24171,
    new_n24172_1, new_n24173, new_n24174, new_n24175, new_n24176,
    new_n24184, new_n24203, new_n24225, new_n24226, new_n24240, new_n24241,
    new_n24242, new_n24243, new_n24244, new_n24245, new_n24246, new_n24247,
    new_n24254, new_n24262, new_n24263, new_n24264, new_n24265, new_n24266,
    new_n24267, new_n24268, new_n24269, new_n24270, new_n24271, new_n24272,
    new_n24273, new_n24279, new_n24280, new_n24281, new_n24282, new_n24283,
    new_n24284, new_n24285, new_n24286, new_n24289_1, new_n24290,
    new_n24291, new_n24292, new_n24298, new_n24299, new_n24300, new_n24301,
    new_n24303, new_n24304, new_n24305, new_n24306, new_n24307_1,
    new_n24308, new_n24309, new_n24310, new_n24311, new_n24312, new_n24313,
    new_n24314, new_n24315, new_n24316, new_n24317, new_n24318,
    new_n24319_1, new_n24331, new_n24359, new_n24360, new_n24361,
    new_n24362, new_n24373_1, new_n24379, new_n24380, new_n24381,
    new_n24382, new_n24383, new_n24398, new_n24405, new_n24406_1,
    new_n24407, new_n24408, new_n24409, new_n24410, new_n24411, new_n24412,
    new_n24413, new_n24414, new_n24429, new_n24430, new_n24431_1,
    new_n24432, new_n24433, new_n24434, new_n24435, new_n24440, new_n24446,
    new_n24447, new_n24448, new_n24449, new_n24450, new_n24451, new_n24452,
    new_n24453, new_n24454, new_n24455, new_n24456, new_n24457, new_n24470,
    new_n24471, new_n24472_1, new_n24476_1, new_n24481, new_n24482,
    new_n24483_1, new_n24490, new_n24491, new_n24492, new_n24493,
    new_n24494, new_n24495, new_n24496, new_n24497, new_n24503, new_n24504,
    new_n24512_1, new_n24513, new_n24514, new_n24515, new_n24516,
    new_n24517, new_n24520, new_n24523, new_n24524, new_n24525, new_n24526,
    new_n24539, new_n24540, new_n24541, new_n24542, new_n24544, new_n24555,
    new_n24556, new_n24557, new_n24558_1, new_n24561, new_n24569,
    new_n24570, new_n24571, new_n24572, new_n24573, new_n24574, new_n24575,
    new_n24576_1, new_n24578, new_n24583, new_n24584, new_n24585,
    new_n24586, new_n24588, new_n24589, new_n24590, new_n24591, new_n24596,
    new_n24597, new_n24598, new_n24599, new_n24600, new_n24601,
    new_n24602_1, new_n24603, new_n24604_1, new_n24605, new_n24606,
    new_n24607, new_n24608, new_n24609, new_n24610, new_n24611, new_n24612,
    new_n24613, new_n24614, new_n24615, new_n24616, new_n24617,
    new_n24618_1, new_n24619, new_n24620_1, new_n24621, new_n24622,
    new_n24627, new_n24628, new_n24629_1, new_n24630, new_n24634,
    new_n24644, new_n24645, new_n24646, new_n24647, new_n24648, new_n24667,
    new_n24668, new_n24669, new_n24670, new_n24671, new_n24672, new_n24674,
    new_n24675, new_n24676, new_n24677, new_n24678, new_n24679, new_n24690,
    new_n24702, new_n24703, new_n24707, new_n24708, new_n24709, new_n24710,
    new_n24712, new_n24713, new_n24715_1, new_n24725, new_n24726,
    new_n24727, new_n24728, new_n24729, new_n24730, new_n24731,
    new_n24732_1, new_n24741, new_n24752, new_n24761, new_n24770,
    new_n24771, new_n24781, new_n24782, new_n24783, new_n24784_1,
    new_n24790, new_n24791, new_n24792, new_n24795, new_n24796, new_n24797,
    new_n24798, new_n24815, new_n24820, new_n24840_1, new_n24850,
    new_n24851, new_n24852, new_n24866, new_n24867, new_n24882, new_n24898,
    new_n24903, new_n24906, new_n24907, new_n24908, new_n24914, new_n24915,
    new_n24916, new_n24920, new_n24921, new_n24922, new_n24923, new_n24925,
    new_n24938, new_n24941, new_n24942, new_n24943, new_n24944, new_n24947,
    new_n24950, new_n24951, new_n24952, new_n24953, new_n24954, new_n24968,
    new_n24969, new_n24972, new_n24984, new_n24986, new_n24987, new_n24988,
    new_n24989, new_n24992, new_n24993, new_n24994, new_n25004,
    new_n25006_1, new_n25011, new_n25012, new_n25013, new_n25014,
    new_n25020, new_n25021, new_n25031, new_n25045, new_n25054, new_n25055,
    new_n25056, new_n25059;
xnor_4 g00000(n10739, n9942, new_n2349);
not_10 g00001(n21753, new_n2350);
or_5   g00002(n25643, new_n2350, new_n2351);
xnor_4 g00003(n25643, n21753, new_n2352);
not_10 g00004(new_n2352, new_n2353);
not_10 g00005(n21832, new_n2354);
or_5   g00006(new_n2354, n9557, new_n2355_1);
xnor_4 g00007(n21832, n9557, new_n2356);
not_10 g00008(new_n2356, new_n2357);
not_10 g00009(n26913, new_n2358);
or_5   g00010(new_n2358, n3136, new_n2359);
xnor_4 g00011(n26913, n3136, new_n2360);
not_10 g00012(n6385, new_n2361_1);
or_5   g00013(n16223, new_n2361_1, new_n2362);
not_10 g00014(n16223, new_n2363_1);
or_5   g00015(new_n2363_1, n6385, new_n2364);
not_10 g00016(n19494, new_n2365);
and_5  g00017(n20138, new_n2365, new_n2366);
not_10 g00018(n20138, new_n2367);
and_5  g00019(new_n2367, n19494, new_n2368);
not_10 g00020(new_n2368, new_n2369);
not_10 g00021(n2387, new_n2370);
and_5  g00022(n9251, new_n2370, new_n2371);
and_5  g00023(new_n2371, new_n2369, new_n2372);
nor_5  g00024(new_n2372, new_n2366, new_n2373);
not_10 g00025(new_n2373, new_n2374_1);
nand_5 g00026(new_n2374_1, new_n2364, new_n2375);
and_5  g00027(new_n2375, new_n2362, new_n2376);
nand_5 g00028(new_n2376, new_n2360, new_n2377);
and_5  g00029(new_n2377, new_n2359, new_n2378);
or_5   g00030(new_n2378, new_n2357, new_n2379);
and_5  g00031(new_n2379, new_n2355_1, new_n2380);
or_5   g00032(new_n2380, new_n2353, new_n2381);
and_5  g00033(new_n2381, new_n2351, new_n2382);
xor_4  g00034(new_n2382, new_n2349, new_n2383);
xor_4  g00035(n13781, n5704, new_n2384);
and_5  g00036(n13781, n5704, new_n2385);
xnor_4 g00037(n18409, n11486, new_n2386);
xor_4  g00038(new_n2386, new_n2385, new_n2387_1);
not_10 g00039(new_n2387_1, new_n2388_1);
nor_5  g00040(new_n2388_1, new_n2384, new_n2389);
not_10 g00041(new_n2389, new_n2390);
xor_4  g00042(n16722, n13708, new_n2391);
not_10 g00043(new_n2391, new_n2392);
nor_5  g00044(n18409, n11486, new_n2393);
nor_5  g00045(new_n2386, new_n2385, new_n2394);
nor_5  g00046(new_n2394, new_n2393, new_n2395);
xor_4  g00047(new_n2395, new_n2392, new_n2396);
not_10 g00048(new_n2396, new_n2397);
nor_5  g00049(new_n2397, new_n2390, new_n2398);
xor_4  g00050(n19911, n3480, new_n2399);
not_10 g00051(new_n2399, new_n2400);
or_5   g00052(n16722, n13708, new_n2401);
or_5   g00053(new_n2395, new_n2392, new_n2402);
and_5  g00054(new_n2402, new_n2401, new_n2403);
xor_4  g00055(new_n2403, new_n2400, new_n2404);
and_5  g00056(new_n2404, new_n2398, new_n2405);
not_10 g00057(new_n2405, new_n2406);
xor_4  g00058(n3018, n2731, new_n2407);
not_10 g00059(new_n2407, new_n2408);
or_5   g00060(n19911, n3480, new_n2409_1);
or_5   g00061(new_n2403, new_n2400, new_n2410);
and_5  g00062(new_n2410, new_n2409_1, new_n2411);
xor_4  g00063(new_n2411, new_n2408, new_n2412);
not_10 g00064(new_n2412, new_n2413);
nor_5  g00065(new_n2413, new_n2406, new_n2414);
xor_4  g00066(n26660, n18907, new_n2415);
not_10 g00067(new_n2415, new_n2416_1);
or_5   g00068(n3018, n2731, new_n2417);
or_5   g00069(new_n2411, new_n2408, new_n2418);
and_5  g00070(new_n2418, new_n2417, new_n2419);
xor_4  g00071(new_n2419, new_n2416_1, new_n2420_1);
and_5  g00072(new_n2420_1, new_n2414, new_n2421_1);
xnor_4 g00073(n22332, n13783, new_n2422);
or_5   g00074(n26660, n18907, new_n2423);
or_5   g00075(new_n2419, new_n2416_1, new_n2424);
and_5  g00076(new_n2424, new_n2423, new_n2425);
xor_4  g00077(new_n2425, new_n2422, new_n2426);
xor_4  g00078(new_n2426, new_n2421_1, new_n2427);
not_10 g00079(new_n2427, new_n2428);
xnor_4 g00080(n13490, n7751, new_n2429);
or_5   g00081(n26823, n22660, new_n2430);
xnor_4 g00082(n26823, n22660, new_n2431);
or_5   g00083(n4812, n1777, new_n2432);
xnor_4 g00084(n4812, n1777, new_n2433);
or_5   g00085(n24278, n8745, new_n2434);
xnor_4 g00086(n24278, n8745, new_n2435);
or_5   g00087(n24618, n15636, new_n2436);
xor_4  g00088(n24618, n15636, new_n2437);
nand_5 g00089(n20077, n3952, new_n2438);
nor_5  g00090(n20077, n3952, new_n2439);
nand_5 g00091(n12315, n6794, new_n2440_1);
or_5   g00092(new_n2440_1, new_n2439, new_n2441);
and_5  g00093(new_n2441, new_n2438, new_n2442);
nand_5 g00094(new_n2442, new_n2437, new_n2443);
and_5  g00095(new_n2443, new_n2436, new_n2444_1);
or_5   g00096(new_n2444_1, new_n2435, new_n2445);
and_5  g00097(new_n2445, new_n2434, new_n2446);
or_5   g00098(new_n2446, new_n2433, new_n2447);
and_5  g00099(new_n2447, new_n2432, new_n2448);
or_5   g00100(new_n2448, new_n2431, new_n2449);
and_5  g00101(new_n2449, new_n2430, new_n2450);
xor_4  g00102(new_n2450, new_n2429, new_n2451);
xor_4  g00103(new_n2451, new_n2428, new_n2452);
not_10 g00104(new_n2420_1, new_n2453);
xor_4  g00105(new_n2453, new_n2414, new_n2454);
xor_4  g00106(new_n2448, new_n2431, new_n2455);
nand_5 g00107(new_n2455, new_n2454, new_n2456);
xor_4  g00108(new_n2413, new_n2406, new_n2457);
xnor_4 g00109(new_n2446, new_n2433, new_n2458);
nor_5  g00110(new_n2458, new_n2457, new_n2459);
not_10 g00111(new_n2459, new_n2460);
xor_4  g00112(new_n2446, new_n2433, new_n2461);
xnor_4 g00113(new_n2461, new_n2457, new_n2462);
not_10 g00114(new_n2462, new_n2463);
not_10 g00115(new_n2404, new_n2464);
xor_4  g00116(new_n2464, new_n2398, new_n2465);
xor_4  g00117(new_n2444_1, new_n2435, new_n2466);
nand_5 g00118(new_n2466, new_n2465, new_n2467);
xor_4  g00119(new_n2397, new_n2390, new_n2468);
xnor_4 g00120(new_n2442, new_n2437, new_n2469);
nor_5  g00121(new_n2469, new_n2468, new_n2470);
not_10 g00122(new_n2470, new_n2471);
xor_4  g00123(new_n2442, new_n2437, new_n2472);
xnor_4 g00124(new_n2472, new_n2468, new_n2473);
not_10 g00125(new_n2473, new_n2474);
xor_4  g00126(n12315, n6794, new_n2475);
and_5  g00127(new_n2475, new_n2384, new_n2476);
xor_4  g00128(n20077, n3952, new_n2477);
xnor_4 g00129(new_n2477, new_n2440_1, new_n2478);
or_5   g00130(new_n2478, new_n2476, new_n2479_1);
nor_5  g00131(n13781, n5704, new_n2480);
not_10 g00132(new_n2394, new_n2481);
nor_5  g00133(new_n2481, new_n2480, new_n2482);
nor_5  g00134(new_n2482, new_n2389, new_n2483);
not_10 g00135(new_n2483, new_n2484);
nand_5 g00136(new_n2477, new_n2476, new_n2485);
and_5  g00137(new_n2485, new_n2479_1, new_n2486);
nand_5 g00138(new_n2486, new_n2484, new_n2487);
and_5  g00139(new_n2487, new_n2479_1, new_n2488);
nor_5  g00140(new_n2488, new_n2474, new_n2489);
not_10 g00141(new_n2489, new_n2490);
and_5  g00142(new_n2490, new_n2471, new_n2491);
xnor_4 g00143(new_n2466, new_n2465, new_n2492);
or_5   g00144(new_n2492, new_n2491, new_n2493);
and_5  g00145(new_n2493, new_n2467, new_n2494);
nor_5  g00146(new_n2494, new_n2463, new_n2495);
not_10 g00147(new_n2495, new_n2496);
and_5  g00148(new_n2496, new_n2460, new_n2497);
xnor_4 g00149(new_n2455, new_n2454, new_n2498);
or_5   g00150(new_n2498, new_n2497, new_n2499);
and_5  g00151(new_n2499, new_n2456, new_n2500);
xnor_4 g00152(new_n2500, new_n2452, new_n2501);
xor_4  g00153(new_n2501, new_n2383, new_n2502);
xor_4  g00154(new_n2380, new_n2353, new_n2503);
xor_4  g00155(new_n2455, new_n2454, new_n2504);
xnor_4 g00156(new_n2504, new_n2497, new_n2505);
not_10 g00157(new_n2505, new_n2506);
or_5   g00158(new_n2506, new_n2503, new_n2507);
xor_4  g00159(new_n2506, new_n2503, new_n2508);
not_10 g00160(new_n2508, new_n2509);
xor_4  g00161(new_n2378, new_n2357, new_n2510);
xor_4  g00162(new_n2494, new_n2463, new_n2511);
not_10 g00163(new_n2511, new_n2512);
or_5   g00164(new_n2512, new_n2510, new_n2513_1);
xor_4  g00165(new_n2512, new_n2510, new_n2514);
xor_4  g00166(new_n2376, new_n2360, new_n2515_1);
xor_4  g00167(new_n2492, new_n2491, new_n2516);
not_10 g00168(new_n2516, new_n2517);
or_5   g00169(new_n2517, new_n2515_1, new_n2518);
xor_4  g00170(new_n2517, new_n2515_1, new_n2519);
xor_4  g00171(new_n2488, new_n2474, new_n2520);
xnor_4 g00172(n16223, n6385, new_n2521);
xor_4  g00173(new_n2521, new_n2374_1, new_n2522);
nand_5 g00174(new_n2522, new_n2520, new_n2523);
not_10 g00175(new_n2520, new_n2524);
xnor_4 g00176(new_n2522, new_n2524, new_n2525);
xnor_4 g00177(n9251, n2387, new_n2526);
xor_4  g00178(new_n2475, new_n2384, new_n2527);
not_10 g00179(new_n2527, new_n2528);
nor_5  g00180(new_n2528, new_n2526, new_n2529);
xnor_4 g00181(n20138, n19494, new_n2530);
xnor_4 g00182(new_n2530, new_n2371, new_n2531);
or_5   g00183(new_n2531, new_n2529, new_n2532);
xor_4  g00184(new_n2486, new_n2484, new_n2533_1);
xor_4  g00185(new_n2531, new_n2529, new_n2534);
nand_5 g00186(new_n2534, new_n2533_1, new_n2535_1);
nand_5 g00187(new_n2535_1, new_n2532, new_n2536);
nand_5 g00188(new_n2536, new_n2525, new_n2537_1);
nand_5 g00189(new_n2537_1, new_n2523, new_n2538);
nand_5 g00190(new_n2538, new_n2519, new_n2539);
nand_5 g00191(new_n2539, new_n2518, new_n2540);
nand_5 g00192(new_n2540, new_n2514, new_n2541);
and_5  g00193(new_n2541, new_n2513_1, new_n2542);
or_5   g00194(new_n2542, new_n2509, new_n2543);
and_5  g00195(new_n2543, new_n2507, new_n2544);
xor_4  g00196(new_n2544, new_n2502, n7);
xor_4  g00197(n3618, n1681, new_n2546);
xor_4  g00198(new_n2546, n4588, new_n2547_1);
not_10 g00199(n22201, new_n2548);
xnor_4 g00200(n22843, n583, new_n2549);
xor_4  g00201(new_n2549, new_n2548, new_n2550);
xor_4  g00202(new_n2550, new_n2547_1, n50);
xor_4  g00203(n19922, n6773, new_n2552);
xor_4  g00204(new_n2552, n21687, new_n2553_1);
xor_4  g00205(n21398, n14090, new_n2554);
xor_4  g00206(new_n2554, n25926, new_n2555_1);
xor_4  g00207(new_n2555_1, new_n2553_1, n55);
not_10 g00208(n25365, new_n2557);
xnor_4 g00209(n20040, n9396, new_n2558);
or_5   g00210(n19531, n1999, new_n2559);
xnor_4 g00211(n19531, n1999, new_n2560_1);
or_5   g00212(n25168, n18345, new_n2561_1);
xnor_4 g00213(n25168, n18345, new_n2562);
or_5   g00214(n13190, n9318, new_n2563);
xnor_4 g00215(n13190, n9318, new_n2564);
or_5   g00216(n19477, n3460, new_n2565);
xnor_4 g00217(n19477, n3460, new_n2566);
or_5   g00218(n11223, n5226, new_n2567);
xnor_4 g00219(n11223, n5226, new_n2568);
or_5   g00220(n17664, n5115, new_n2569);
xnor_4 g00221(n17664, n5115, new_n2570_1);
or_5   g00222(n26572, n23369, new_n2571);
xnor_4 g00223(n26572, n23369, new_n2572);
or_5   g00224(n11667, n1136, new_n2573_1);
nand_5 g00225(n21398, n19234, new_n2574);
xor_4  g00226(n11667, n1136, new_n2575);
nand_5 g00227(new_n2575, new_n2574, new_n2576);
and_5  g00228(new_n2576, new_n2573_1, new_n2577);
or_5   g00229(new_n2577, new_n2572, new_n2578_1);
and_5  g00230(new_n2578_1, new_n2571, new_n2579);
or_5   g00231(new_n2579, new_n2570_1, new_n2580);
and_5  g00232(new_n2580, new_n2569, new_n2581);
or_5   g00233(new_n2581, new_n2568, new_n2582_1);
and_5  g00234(new_n2582_1, new_n2567, new_n2583);
or_5   g00235(new_n2583, new_n2566, new_n2584);
and_5  g00236(new_n2584, new_n2565, new_n2585);
or_5   g00237(new_n2585, new_n2564, new_n2586);
and_5  g00238(new_n2586, new_n2563, new_n2587);
or_5   g00239(new_n2587, new_n2562, new_n2588);
and_5  g00240(new_n2588, new_n2561_1, new_n2589);
or_5   g00241(new_n2589, new_n2560_1, new_n2590);
and_5  g00242(new_n2590, new_n2559, new_n2591);
xor_4  g00243(new_n2591, new_n2558, new_n2592);
xor_4  g00244(new_n2592, new_n2557, new_n2593);
not_10 g00245(new_n2593, new_n2594);
not_10 g00246(n14704, new_n2595);
xor_4  g00247(new_n2589, new_n2560_1, new_n2596);
or_5   g00248(new_n2596, new_n2595, new_n2597);
xor_4  g00249(new_n2596, new_n2595, new_n2598);
not_10 g00250(new_n2598, new_n2599);
not_10 g00251(n19270, new_n2600);
xor_4  g00252(new_n2587, new_n2562, new_n2601);
or_5   g00253(new_n2601, new_n2600, new_n2602_1);
xor_4  g00254(new_n2601, new_n2600, new_n2603);
not_10 g00255(new_n2603, new_n2604);
not_10 g00256(n8687, new_n2605);
xor_4  g00257(new_n2585, new_n2564, new_n2606);
or_5   g00258(new_n2606, new_n2605, new_n2607);
not_10 g00259(n24768, new_n2608);
xor_4  g00260(new_n2583, new_n2566, new_n2609);
and_5  g00261(new_n2609, new_n2608, new_n2610);
xor_4  g00262(new_n2609, new_n2608, new_n2611);
not_10 g00263(new_n2611, new_n2612);
not_10 g00264(n26483, new_n2613);
xor_4  g00265(new_n2581, new_n2568, new_n2614);
nand_5 g00266(new_n2614, new_n2613, new_n2615);
xor_4  g00267(new_n2614, new_n2613, new_n2616);
not_10 g00268(n15979, new_n2617);
xor_4  g00269(new_n2579, new_n2570_1, new_n2618);
or_5   g00270(new_n2618, new_n2617, new_n2619_1);
xor_4  g00271(new_n2618, new_n2617, new_n2620);
not_10 g00272(new_n2620, new_n2621);
not_10 g00273(n8638, new_n2622);
xor_4  g00274(new_n2577, new_n2572, new_n2623);
or_5   g00275(new_n2623, new_n2622, new_n2624);
not_10 g00276(n16247, new_n2625);
xor_4  g00277(new_n2575, new_n2574, new_n2626);
nand_5 g00278(new_n2626, new_n2625, new_n2627);
xor_4  g00279(n21398, n19234, new_n2628);
nand_5 g00280(new_n2628, n23541, new_n2629);
xor_4  g00281(new_n2626, new_n2625, new_n2630);
nand_5 g00282(new_n2630, new_n2629, new_n2631);
and_5  g00283(new_n2631, new_n2627, new_n2632);
xor_4  g00284(new_n2623, new_n2622, new_n2633);
nand_5 g00285(new_n2633, new_n2632, new_n2634);
and_5  g00286(new_n2634, new_n2624, new_n2635);
or_5   g00287(new_n2635, new_n2621, new_n2636);
and_5  g00288(new_n2636, new_n2619_1, new_n2637);
nand_5 g00289(new_n2637, new_n2616, new_n2638);
and_5  g00290(new_n2638, new_n2615, new_n2639);
nor_5  g00291(new_n2639, new_n2612, new_n2640);
nor_5  g00292(new_n2640, new_n2610, new_n2641);
xor_4  g00293(new_n2606, new_n2605, new_n2642);
nand_5 g00294(new_n2642, new_n2641, new_n2643);
and_5  g00295(new_n2643, new_n2607, new_n2644);
or_5   g00296(new_n2644, new_n2604, new_n2645);
and_5  g00297(new_n2645, new_n2602_1, new_n2646_1);
or_5   g00298(new_n2646_1, new_n2599, new_n2647);
and_5  g00299(new_n2647, new_n2597, new_n2648);
xor_4  g00300(new_n2648, new_n2594, new_n2649);
not_10 g00301(n13951, new_n2650);
not_10 g00302(n22793, new_n2651);
not_10 g00303(n8439, new_n2652);
not_10 g00304(n25523, new_n2653);
not_10 g00305(n5579, new_n2654);
not_10 g00306(n23430, new_n2655);
not_10 g00307(n10411, new_n2656);
not_10 g00308(n16971, new_n2657);
nor_5  g00309(n18151, n11503, new_n2658);
and_5  g00310(new_n2658, new_n2657, new_n2659_1);
and_5  g00311(new_n2659_1, new_n2656, new_n2660);
and_5  g00312(new_n2660, new_n2655, new_n2661_1);
and_5  g00313(new_n2661_1, new_n2654, new_n2662);
and_5  g00314(new_n2662, new_n2653, new_n2663);
and_5  g00315(new_n2663, new_n2652, new_n2664);
and_5  g00316(new_n2664, new_n2651, new_n2665);
xor_4  g00317(new_n2665, new_n2650, new_n2666);
xor_4  g00318(n22270, n2944, new_n2667);
not_10 g00319(new_n2667, new_n2668);
or_5   g00320(n8806, n767, new_n2669);
xor_4  g00321(n8806, n767, new_n2670);
not_10 g00322(new_n2670, new_n2671);
or_5   g00323(n7330, n2479, new_n2672);
xor_4  g00324(n7330, n2479, new_n2673);
not_10 g00325(new_n2673, new_n2674);
or_5   g00326(n22492, n9372, new_n2675);
xor_4  g00327(n22492, n9372, new_n2676);
not_10 g00328(new_n2676, new_n2677);
or_5   g00329(n12821, n6596, new_n2678);
xor_4  g00330(n12821, n6596, new_n2679);
not_10 g00331(new_n2679, new_n2680_1);
or_5   g00332(n15289, n3468, new_n2681);
xor_4  g00333(n15289, n3468, new_n2682);
not_10 g00334(new_n2682, new_n2683);
or_5   g00335(n18558, n6556, new_n2684);
xor_4  g00336(n18558, n6556, new_n2685);
not_10 g00337(new_n2685, new_n2686);
or_5   g00338(n22871, n7149, new_n2687);
xor_4  g00339(n22871, n7149, new_n2688);
not_10 g00340(new_n2688, new_n2689);
or_5   g00341(n14275, n14148, new_n2690);
and_5  g00342(n25023, n1152, new_n2691);
xnor_4 g00343(n14275, n14148, new_n2692);
or_5   g00344(new_n2692, new_n2691, new_n2693_1);
and_5  g00345(new_n2693_1, new_n2690, new_n2694);
or_5   g00346(new_n2694, new_n2689, new_n2695);
and_5  g00347(new_n2695, new_n2687, new_n2696);
or_5   g00348(new_n2696, new_n2686, new_n2697);
and_5  g00349(new_n2697, new_n2684, new_n2698);
or_5   g00350(new_n2698, new_n2683, new_n2699);
and_5  g00351(new_n2699, new_n2681, new_n2700);
or_5   g00352(new_n2700, new_n2680_1, new_n2701);
and_5  g00353(new_n2701, new_n2678, new_n2702);
or_5   g00354(new_n2702, new_n2677, new_n2703_1);
and_5  g00355(new_n2703_1, new_n2675, new_n2704);
or_5   g00356(new_n2704, new_n2674, new_n2705);
and_5  g00357(new_n2705, new_n2672, new_n2706_1);
or_5   g00358(new_n2706_1, new_n2671, new_n2707);
and_5  g00359(new_n2707, new_n2669, new_n2708);
xor_4  g00360(new_n2708, new_n2668, new_n2709);
not_10 g00361(new_n2709, new_n2710);
xor_4  g00362(new_n2710, new_n2666, new_n2711_1);
xor_4  g00363(new_n2664, new_n2651, new_n2712);
xor_4  g00364(new_n2706_1, new_n2671, new_n2713);
nand_5 g00365(new_n2713, new_n2712, new_n2714);
not_10 g00366(new_n2713, new_n2715);
xnor_4 g00367(new_n2715, new_n2712, new_n2716);
xor_4  g00368(new_n2663, new_n2652, new_n2717);
xor_4  g00369(new_n2704, new_n2674, new_n2718);
or_5   g00370(new_n2718, new_n2717, new_n2719);
not_10 g00371(new_n2718, new_n2720);
xor_4  g00372(new_n2720, new_n2717, new_n2721);
xor_4  g00373(new_n2662, new_n2653, new_n2722);
xor_4  g00374(new_n2702, new_n2677, new_n2723);
or_5   g00375(new_n2723, new_n2722, new_n2724);
not_10 g00376(new_n2723, new_n2725);
xor_4  g00377(new_n2725, new_n2722, new_n2726);
xor_4  g00378(new_n2661_1, new_n2654, new_n2727);
xor_4  g00379(new_n2700, new_n2680_1, new_n2728);
or_5   g00380(new_n2728, new_n2727, new_n2729);
not_10 g00381(new_n2728, new_n2730);
xor_4  g00382(new_n2730, new_n2727, new_n2731_1);
xor_4  g00383(new_n2660, new_n2655, new_n2732);
xor_4  g00384(new_n2698, new_n2683, new_n2733);
or_5   g00385(new_n2733, new_n2732, new_n2734);
xor_4  g00386(new_n2659_1, new_n2656, new_n2735);
not_10 g00387(new_n2735, new_n2736);
xor_4  g00388(new_n2696, new_n2686, new_n2737);
not_10 g00389(new_n2737, new_n2738);
and_5  g00390(new_n2738, new_n2736, new_n2739);
xor_4  g00391(new_n2738, new_n2736, new_n2740);
xor_4  g00392(new_n2658, new_n2657, new_n2741);
not_10 g00393(new_n2741, new_n2742);
xor_4  g00394(new_n2694, new_n2689, new_n2743_1);
not_10 g00395(new_n2743_1, new_n2744);
nand_5 g00396(new_n2744, new_n2742, new_n2745);
xor_4  g00397(new_n2744, new_n2742, new_n2746);
xor_4  g00398(n18151, n11503, new_n2747);
xor_4  g00399(n14275, n14148, new_n2748);
xnor_4 g00400(new_n2748, new_n2691, new_n2749);
or_5   g00401(new_n2749, new_n2747, new_n2750);
not_10 g00402(n18151, new_n2751);
xor_4  g00403(n25023, n1152, new_n2752);
and_5  g00404(new_n2752, new_n2751, new_n2753);
not_10 g00405(new_n2749, new_n2754);
xnor_4 g00406(new_n2754, new_n2747, new_n2755);
nand_5 g00407(new_n2755, new_n2753, new_n2756);
nand_5 g00408(new_n2756, new_n2750, new_n2757);
nand_5 g00409(new_n2757, new_n2746, new_n2758);
nand_5 g00410(new_n2758, new_n2745, new_n2759);
and_5  g00411(new_n2759, new_n2740, new_n2760);
or_5   g00412(new_n2760, new_n2739, new_n2761_1);
not_10 g00413(new_n2733, new_n2762);
xnor_4 g00414(new_n2762, new_n2732, new_n2763);
nand_5 g00415(new_n2763, new_n2761_1, new_n2764);
and_5  g00416(new_n2764, new_n2734, new_n2765);
or_5   g00417(new_n2765, new_n2731_1, new_n2766);
and_5  g00418(new_n2766, new_n2729, new_n2767);
or_5   g00419(new_n2767, new_n2726, new_n2768);
and_5  g00420(new_n2768, new_n2724, new_n2769);
or_5   g00421(new_n2769, new_n2721, new_n2770);
and_5  g00422(new_n2770, new_n2719, new_n2771);
nand_5 g00423(new_n2771, new_n2716, new_n2772);
and_5  g00424(new_n2772, new_n2714, new_n2773);
xor_4  g00425(new_n2773, new_n2711_1, new_n2774_1);
xor_4  g00426(new_n2774_1, new_n2649, new_n2775);
xor_4  g00427(new_n2646_1, new_n2599, new_n2776);
xor_4  g00428(new_n2771, new_n2716, new_n2777);
and_5  g00429(new_n2777, new_n2776, new_n2778);
xor_4  g00430(new_n2777, new_n2776, new_n2779_1);
xor_4  g00431(new_n2644, new_n2604, new_n2780);
not_10 g00432(new_n2780, new_n2781);
xor_4  g00433(new_n2769, new_n2721, new_n2782);
nand_5 g00434(new_n2782, new_n2781, new_n2783_1);
xnor_4 g00435(new_n2782, new_n2780, new_n2784);
not_10 g00436(new_n2784, new_n2785);
xor_4  g00437(new_n2642, new_n2641, new_n2786);
not_10 g00438(new_n2786, new_n2787);
xor_4  g00439(new_n2767, new_n2726, new_n2788);
nand_5 g00440(new_n2788, new_n2787, new_n2789);
xor_4  g00441(new_n2788, new_n2787, new_n2790);
xor_4  g00442(new_n2639, new_n2612, new_n2791);
xor_4  g00443(new_n2765, new_n2731_1, new_n2792);
nor_5  g00444(new_n2792, new_n2791, new_n2793);
xor_4  g00445(new_n2792, new_n2791, new_n2794);
xor_4  g00446(new_n2637, new_n2616, new_n2795);
xor_4  g00447(new_n2763, new_n2761_1, new_n2796);
nand_5 g00448(new_n2796, new_n2795, new_n2797);
not_10 g00449(new_n2795, new_n2798);
xnor_4 g00450(new_n2796, new_n2798, new_n2799);
not_10 g00451(new_n2799, new_n2800);
xor_4  g00452(new_n2759, new_n2740, new_n2801);
xor_4  g00453(new_n2635, new_n2621, new_n2802);
not_10 g00454(new_n2802, new_n2803);
nand_5 g00455(new_n2803, new_n2801, new_n2804);
xnor_4 g00456(new_n2802, new_n2801, new_n2805);
xnor_4 g00457(new_n2757, new_n2746, new_n2806);
xor_4  g00458(new_n2633, new_n2632, new_n2807);
and_5  g00459(new_n2807, new_n2806, new_n2808);
xor_4  g00460(new_n2807, new_n2806, new_n2809_1);
xor_4  g00461(new_n2755, new_n2753, new_n2810);
xor_4  g00462(new_n2630, new_n2629, new_n2811);
nand_5 g00463(new_n2811, new_n2810, new_n2812);
xnor_4 g00464(new_n2628, n23541, new_n2813);
xor_4  g00465(new_n2752, new_n2751, new_n2814);
nor_5  g00466(new_n2814, new_n2813, new_n2815);
xor_4  g00467(new_n2811, new_n2810, new_n2816_1);
not_10 g00468(new_n2816_1, new_n2817);
or_5   g00469(new_n2817, new_n2815, new_n2818);
and_5  g00470(new_n2818, new_n2812, new_n2819);
and_5  g00471(new_n2819, new_n2809_1, new_n2820);
nor_5  g00472(new_n2820, new_n2808, new_n2821);
nand_5 g00473(new_n2821, new_n2805, new_n2822);
and_5  g00474(new_n2822, new_n2804, new_n2823);
or_5   g00475(new_n2823, new_n2800, new_n2824);
and_5  g00476(new_n2824, new_n2797, new_n2825);
and_5  g00477(new_n2825, new_n2794, new_n2826_1);
nor_5  g00478(new_n2826_1, new_n2793, new_n2827);
nand_5 g00479(new_n2827, new_n2790, new_n2828);
and_5  g00480(new_n2828, new_n2789, new_n2829);
or_5   g00481(new_n2829, new_n2785, new_n2830);
and_5  g00482(new_n2830, new_n2783_1, new_n2831);
and_5  g00483(new_n2831, new_n2779_1, new_n2832);
nor_5  g00484(new_n2832, new_n2778, new_n2833);
xnor_4 g00485(new_n2833, new_n2775, n108);
xnor_4 g00486(n22379, n767, new_n2835);
not_10 g00487(new_n2835, new_n2836);
not_10 g00488(n1662, new_n2837);
or_5   g00489(n7330, new_n2837, new_n2838);
xnor_4 g00490(n7330, n1662, new_n2839);
not_10 g00491(new_n2839, new_n2840);
not_10 g00492(n12875, new_n2841);
or_5   g00493(n22492, new_n2841, new_n2842);
xnor_4 g00494(n22492, n12875, new_n2843);
not_10 g00495(new_n2843, new_n2844);
not_10 g00496(n2035, new_n2845);
or_5   g00497(n12821, new_n2845, new_n2846);
xnor_4 g00498(n12821, n2035, new_n2847);
not_10 g00499(new_n2847, new_n2848);
not_10 g00500(n5213, new_n2849);
or_5   g00501(new_n2849, n3468, new_n2850);
xnor_4 g00502(n5213, n3468, new_n2851);
not_10 g00503(new_n2851, new_n2852);
not_10 g00504(n4665, new_n2853_1);
or_5   g00505(n18558, new_n2853_1, new_n2854);
xnor_4 g00506(n18558, n4665, new_n2855);
not_10 g00507(n7149, new_n2856);
or_5   g00508(n19005, new_n2856, new_n2857);
not_10 g00509(n19005, new_n2858_1);
or_5   g00510(new_n2858_1, n7149, new_n2859);
not_10 g00511(n4326, new_n2860_1);
and_5  g00512(n14148, new_n2860_1, new_n2861);
not_10 g00513(n14148, new_n2862);
and_5  g00514(new_n2862, n4326, new_n2863);
not_10 g00515(new_n2863, new_n2864);
not_10 g00516(n5438, new_n2865);
and_5  g00517(new_n2865, n1152, new_n2866);
and_5  g00518(new_n2866, new_n2864, new_n2867);
nor_5  g00519(new_n2867, new_n2861, new_n2868);
not_10 g00520(new_n2868, new_n2869);
nand_5 g00521(new_n2869, new_n2859, new_n2870);
and_5  g00522(new_n2870, new_n2857, new_n2871);
nand_5 g00523(new_n2871, new_n2855, new_n2872);
and_5  g00524(new_n2872, new_n2854, new_n2873);
or_5   g00525(new_n2873, new_n2852, new_n2874);
and_5  g00526(new_n2874, new_n2850, new_n2875);
or_5   g00527(new_n2875, new_n2848, new_n2876);
and_5  g00528(new_n2876, new_n2846, new_n2877);
or_5   g00529(new_n2877, new_n2844, new_n2878);
and_5  g00530(new_n2878, new_n2842, new_n2879);
or_5   g00531(new_n2879, new_n2840, new_n2880);
and_5  g00532(new_n2880, new_n2838, new_n2881);
xor_4  g00533(new_n2881, new_n2836, new_n2882);
xnor_4 g00534(n10763, n6814, new_n2883);
or_5   g00535(n19701, n7437, new_n2884);
xnor_4 g00536(n19701, n7437, new_n2885);
or_5   g00537(n23529, n20700, new_n2886_1);
xnor_4 g00538(n23529, n20700, new_n2887_1);
or_5   g00539(n24620, n7099, new_n2888);
xnor_4 g00540(n24620, n7099, new_n2889);
or_5   g00541(n12811, n5211, new_n2890);
xnor_4 g00542(n12811, n5211, new_n2891);
or_5   g00543(n12956, n1118, new_n2892);
xnor_4 g00544(n12956, n1118, new_n2893);
or_5   g00545(n25974, n18295, new_n2894);
xnor_4 g00546(n25974, n18295, new_n2895);
or_5   g00547(n6502, n1630, new_n2896);
and_5  g00548(n15780, n1451, new_n2897);
xnor_4 g00549(n6502, n1630, new_n2898);
or_5   g00550(new_n2898, new_n2897, new_n2899);
and_5  g00551(new_n2899, new_n2896, new_n2900);
or_5   g00552(new_n2900, new_n2895, new_n2901);
and_5  g00553(new_n2901, new_n2894, new_n2902);
or_5   g00554(new_n2902, new_n2893, new_n2903);
and_5  g00555(new_n2903, new_n2892, new_n2904);
or_5   g00556(new_n2904, new_n2891, new_n2905);
and_5  g00557(new_n2905, new_n2890, new_n2906);
or_5   g00558(new_n2906, new_n2889, new_n2907);
and_5  g00559(new_n2907, new_n2888, new_n2908);
or_5   g00560(new_n2908, new_n2887_1, new_n2909);
and_5  g00561(new_n2909, new_n2886_1, new_n2910);
or_5   g00562(new_n2910, new_n2885, new_n2911);
and_5  g00563(new_n2911, new_n2884, new_n2912);
xor_4  g00564(new_n2912, new_n2883, new_n2913);
xor_4  g00565(n27089, n12657, new_n2914);
not_10 g00566(new_n2914, new_n2915);
or_5   g00567(n17077, n11841, new_n2916);
xor_4  g00568(n17077, n11841, new_n2917);
not_10 g00569(new_n2917, new_n2918);
or_5   g00570(n26510, n10710, new_n2919);
xor_4  g00571(n26510, n10710, new_n2920);
not_10 g00572(new_n2920, new_n2921);
or_5   g00573(n23068, n20929, new_n2922);
xor_4  g00574(n23068, n20929, new_n2923);
not_10 g00575(new_n2923, new_n2924);
or_5   g00576(n19514, n8006, new_n2925);
xor_4  g00577(n19514, n8006, new_n2926);
not_10 g00578(new_n2926, new_n2927);
or_5   g00579(n25074, n10053, new_n2928);
xor_4  g00580(n25074, n10053, new_n2929_1);
not_10 g00581(new_n2929_1, new_n2930);
or_5   g00582(n16396, n8399, new_n2931);
xor_4  g00583(n16396, n8399, new_n2932);
not_10 g00584(new_n2932, new_n2933);
or_5   g00585(n9507, n9399, new_n2934);
nand_5 g00586(n26979, n2088, new_n2935);
xor_4  g00587(n9507, n9399, new_n2936);
nand_5 g00588(new_n2936, new_n2935, new_n2937);
and_5  g00589(new_n2937, new_n2934, new_n2938);
or_5   g00590(new_n2938, new_n2933, new_n2939);
and_5  g00591(new_n2939, new_n2931, new_n2940);
or_5   g00592(new_n2940, new_n2930, new_n2941);
and_5  g00593(new_n2941, new_n2928, new_n2942);
or_5   g00594(new_n2942, new_n2927, new_n2943);
and_5  g00595(new_n2943, new_n2925, new_n2944_1);
or_5   g00596(new_n2944_1, new_n2924, new_n2945);
and_5  g00597(new_n2945, new_n2922, new_n2946);
or_5   g00598(new_n2946, new_n2921, new_n2947);
and_5  g00599(new_n2947, new_n2919, new_n2948_1);
or_5   g00600(new_n2948_1, new_n2918, new_n2949);
and_5  g00601(new_n2949, new_n2916, new_n2950);
xor_4  g00602(new_n2950, new_n2915, new_n2951);
xor_4  g00603(new_n2951, new_n2913, new_n2952);
xor_4  g00604(new_n2910, new_n2885, new_n2953);
xor_4  g00605(new_n2948_1, new_n2918, new_n2954);
not_10 g00606(new_n2954, new_n2955);
or_5   g00607(new_n2955, new_n2953, new_n2956);
xnor_4 g00608(new_n2954, new_n2953, new_n2957);
xor_4  g00609(new_n2908, new_n2887_1, new_n2958);
xor_4  g00610(new_n2946, new_n2921, new_n2959);
not_10 g00611(new_n2959, new_n2960);
nand_5 g00612(new_n2960, new_n2958, new_n2961_1);
xnor_4 g00613(new_n2959, new_n2958, new_n2962);
not_10 g00614(new_n2962, new_n2963);
xor_4  g00615(new_n2906, new_n2889, new_n2964);
xor_4  g00616(new_n2944_1, new_n2924, new_n2965);
not_10 g00617(new_n2965, new_n2966);
nand_5 g00618(new_n2966, new_n2964, new_n2967);
xnor_4 g00619(new_n2965, new_n2964, new_n2968);
not_10 g00620(new_n2968, new_n2969);
xor_4  g00621(new_n2904, new_n2891, new_n2970);
xor_4  g00622(new_n2942, new_n2927, new_n2971_1);
not_10 g00623(new_n2971_1, new_n2972);
nand_5 g00624(new_n2972, new_n2970, new_n2973);
xnor_4 g00625(new_n2971_1, new_n2970, new_n2974);
not_10 g00626(new_n2974, new_n2975);
xor_4  g00627(new_n2902, new_n2893, new_n2976);
xor_4  g00628(new_n2940, new_n2930, new_n2977);
not_10 g00629(new_n2977, new_n2978_1);
nand_5 g00630(new_n2978_1, new_n2976, new_n2979_1);
xnor_4 g00631(new_n2977, new_n2976, new_n2980);
xor_4  g00632(new_n2900, new_n2895, new_n2981);
xor_4  g00633(new_n2938, new_n2933, new_n2982);
not_10 g00634(new_n2982, new_n2983);
or_5   g00635(new_n2983, new_n2981, new_n2984);
xnor_4 g00636(new_n2982, new_n2981, new_n2985_1);
xor_4  g00637(n6502, n1630, new_n2986);
xnor_4 g00638(new_n2986, new_n2897, new_n2987);
not_10 g00639(new_n2987, new_n2988);
xor_4  g00640(new_n2936, new_n2935, new_n2989);
or_5   g00641(new_n2989, new_n2988, new_n2990);
xor_4  g00642(n15780, n1451, new_n2991);
xnor_4 g00643(n26979, n2088, new_n2992);
nor_5  g00644(new_n2992, new_n2991, new_n2993);
xor_4  g00645(new_n2989, new_n2988, new_n2994);
nand_5 g00646(new_n2994, new_n2993, new_n2995);
and_5  g00647(new_n2995, new_n2990, new_n2996);
nand_5 g00648(new_n2996, new_n2985_1, new_n2997);
and_5  g00649(new_n2997, new_n2984, new_n2998);
nand_5 g00650(new_n2998, new_n2980, new_n2999_1);
and_5  g00651(new_n2999_1, new_n2979_1, new_n3000);
or_5   g00652(new_n3000, new_n2975, new_n3001);
and_5  g00653(new_n3001, new_n2973, new_n3002);
or_5   g00654(new_n3002, new_n2969, new_n3003);
and_5  g00655(new_n3003, new_n2967, new_n3004);
or_5   g00656(new_n3004, new_n2963, new_n3005);
and_5  g00657(new_n3005, new_n2961_1, new_n3006);
nand_5 g00658(new_n3006, new_n2957, new_n3007);
and_5  g00659(new_n3007, new_n2956, new_n3008);
xor_4  g00660(new_n3008, new_n2952, new_n3009);
xor_4  g00661(new_n3009, new_n2882, new_n3010_1);
not_10 g00662(new_n3010_1, new_n3011);
xor_4  g00663(new_n2879, new_n2840, new_n3012);
xor_4  g00664(new_n3006, new_n2957, new_n3013);
nor_5  g00665(new_n3013, new_n3012, new_n3014);
xor_4  g00666(new_n3013, new_n3012, new_n3015);
not_10 g00667(new_n3015, new_n3016);
xor_4  g00668(new_n2877, new_n2844, new_n3017_1);
not_10 g00669(new_n3017_1, new_n3018_1);
xor_4  g00670(new_n3004, new_n2963, new_n3019);
and_5  g00671(new_n3019, new_n3018_1, new_n3020_1);
xor_4  g00672(new_n3019, new_n3018_1, new_n3021);
not_10 g00673(new_n3021, new_n3022);
xor_4  g00674(new_n2875, new_n2848, new_n3023);
not_10 g00675(new_n3023, new_n3024);
xor_4  g00676(new_n3002, new_n2969, new_n3025);
and_5  g00677(new_n3025, new_n3024, new_n3026);
xor_4  g00678(new_n3025, new_n3024, new_n3027);
not_10 g00679(new_n3027, new_n3028);
xor_4  g00680(new_n2873, new_n2852, new_n3029);
not_10 g00681(new_n3029, new_n3030_1);
xor_4  g00682(new_n3000, new_n2975, new_n3031);
and_5  g00683(new_n3031, new_n3030_1, new_n3032);
xor_4  g00684(new_n3031, new_n3030_1, new_n3033);
not_10 g00685(new_n3033, new_n3034);
xor_4  g00686(new_n2998, new_n2980, new_n3035);
not_10 g00687(new_n3035, new_n3036);
xor_4  g00688(new_n2871, new_n2855, new_n3037);
nor_5  g00689(new_n3037, new_n3036, new_n3038);
xor_4  g00690(new_n3037, new_n3036, new_n3039);
xor_4  g00691(new_n2996, new_n2985_1, new_n3040);
not_10 g00692(new_n3040, new_n3041);
xnor_4 g00693(n19005, n7149, new_n3042);
xor_4  g00694(new_n3042, new_n2869, new_n3043);
and_5  g00695(new_n3043, new_n3041, new_n3044);
xor_4  g00696(new_n3043, new_n3041, new_n3045);
xnor_4 g00697(n5438, n1152, new_n3046);
xor_4  g00698(n26979, n2088, new_n3047);
xnor_4 g00699(new_n3047, new_n2991, new_n3048);
nor_5  g00700(new_n3048, new_n3046, new_n3049);
not_10 g00701(new_n3049, new_n3050);
xnor_4 g00702(n14148, n4326, new_n3051);
xor_4  g00703(new_n3051, new_n2866, new_n3052);
and_5  g00704(new_n3052, new_n3050, new_n3053);
not_10 g00705(new_n3053, new_n3054);
xor_4  g00706(new_n2994, new_n2993, new_n3055);
xor_4  g00707(new_n3052, new_n3050, new_n3056);
and_5  g00708(new_n3056, new_n3055, new_n3057);
not_10 g00709(new_n3057, new_n3058);
and_5  g00710(new_n3058, new_n3054, new_n3059);
not_10 g00711(new_n3059, new_n3060);
and_5  g00712(new_n3060, new_n3045, new_n3061);
nor_5  g00713(new_n3061, new_n3044, new_n3062);
not_10 g00714(new_n3062, new_n3063);
and_5  g00715(new_n3063, new_n3039, new_n3064);
nor_5  g00716(new_n3064, new_n3038, new_n3065);
nor_5  g00717(new_n3065, new_n3034, new_n3066);
nor_5  g00718(new_n3066, new_n3032, new_n3067_1);
nor_5  g00719(new_n3067_1, new_n3028, new_n3068);
nor_5  g00720(new_n3068, new_n3026, new_n3069);
nor_5  g00721(new_n3069, new_n3022, new_n3070);
nor_5  g00722(new_n3070, new_n3020_1, new_n3071);
nor_5  g00723(new_n3071, new_n3016, new_n3072);
nor_5  g00724(new_n3072, new_n3014, new_n3073);
xnor_4 g00725(new_n3073, new_n3011, n142);
not_10 g00726(n5025, new_n3075);
xor_4  g00727(n7335, n4319, new_n3076_1);
not_10 g00728(new_n3076_1, new_n3077);
or_5   g00729(n23463, n5696, new_n3078);
xor_4  g00730(n23463, n5696, new_n3079);
not_10 g00731(new_n3079, new_n3080);
or_5   g00732(n13367, n13074, new_n3081);
xor_4  g00733(n13367, n13074, new_n3082);
not_10 g00734(new_n3082, new_n3083);
or_5   g00735(n10739, n932, new_n3084);
xor_4  g00736(n10739, n932, new_n3085);
not_10 g00737(new_n3085, new_n3086);
or_5   g00738(n21753, n6691, new_n3087);
xor_4  g00739(n21753, n6691, new_n3088);
not_10 g00740(new_n3088, new_n3089_1);
or_5   g00741(n21832, n3260, new_n3090);
xor_4  g00742(n21832, n3260, new_n3091);
not_10 g00743(new_n3091, new_n3092);
or_5   g00744(n26913, n20489, new_n3093);
xor_4  g00745(n26913, n20489, new_n3094);
not_10 g00746(new_n3094, new_n3095);
or_5   g00747(n16223, n2355, new_n3096);
xor_4  g00748(n16223, n2355, new_n3097);
not_10 g00749(new_n3097, new_n3098);
or_5   g00750(n19494, n11121, new_n3099);
nand_5 g00751(n16217, n2387, new_n3100);
xor_4  g00752(n19494, n11121, new_n3101);
nand_5 g00753(new_n3101, new_n3100, new_n3102);
and_5  g00754(new_n3102, new_n3099, new_n3103);
or_5   g00755(new_n3103, new_n3098, new_n3104);
and_5  g00756(new_n3104, new_n3096, new_n3105);
or_5   g00757(new_n3105, new_n3095, new_n3106);
and_5  g00758(new_n3106, new_n3093, new_n3107);
or_5   g00759(new_n3107, new_n3092, new_n3108);
and_5  g00760(new_n3108, new_n3090, new_n3109);
or_5   g00761(new_n3109, new_n3089_1, new_n3110);
and_5  g00762(new_n3110, new_n3087, new_n3111);
or_5   g00763(new_n3111, new_n3086, new_n3112);
and_5  g00764(new_n3112, new_n3084, new_n3113);
or_5   g00765(new_n3113, new_n3083, new_n3114);
and_5  g00766(new_n3114, new_n3081, new_n3115);
or_5   g00767(new_n3115, new_n3080, new_n3116);
and_5  g00768(new_n3116, new_n3078, new_n3117);
xor_4  g00769(new_n3117, new_n3077, new_n3118);
not_10 g00770(new_n3118, new_n3119);
nand_5 g00771(new_n3119, new_n3075, new_n3120);
xor_4  g00772(new_n3119, n5025, new_n3121);
xor_4  g00773(new_n3115, new_n3080, new_n3122);
or_5   g00774(new_n3122, n6485, new_n3123);
not_10 g00775(new_n3122, new_n3124);
xor_4  g00776(new_n3124, n6485, new_n3125_1);
xor_4  g00777(new_n3113, new_n3083, new_n3126_1);
or_5   g00778(new_n3126_1, n26036, new_n3127);
not_10 g00779(new_n3126_1, new_n3128);
xor_4  g00780(new_n3128, n26036, new_n3129);
xor_4  g00781(new_n3111, new_n3086, new_n3130);
or_5   g00782(new_n3130, n19770, new_n3131);
not_10 g00783(new_n3130, new_n3132);
xor_4  g00784(new_n3132, n19770, new_n3133);
xor_4  g00785(new_n3109, new_n3089_1, new_n3134);
or_5   g00786(new_n3134, n8782, new_n3135);
not_10 g00787(new_n3134, new_n3136_1);
xor_4  g00788(new_n3136_1, n8782, new_n3137);
xor_4  g00789(new_n3107, new_n3092, new_n3138);
or_5   g00790(new_n3138, n8678, new_n3139);
not_10 g00791(new_n3138, new_n3140);
xor_4  g00792(new_n3140, n8678, new_n3141);
xor_4  g00793(new_n3105, new_n3095, new_n3142);
or_5   g00794(new_n3142, n1432, new_n3143);
not_10 g00795(new_n3142, new_n3144);
xor_4  g00796(new_n3144, n1432, new_n3145);
not_10 g00797(n21599, new_n3146);
xor_4  g00798(new_n3103, new_n3098, new_n3147);
not_10 g00799(new_n3147, new_n3148);
nand_5 g00800(new_n3148, new_n3146, new_n3149);
xor_4  g00801(new_n3148, n21599, new_n3150);
not_10 g00802(n25336, new_n3151);
not_10 g00803(n11424, new_n3152);
xor_4  g00804(n16217, n2387, new_n3153);
and_5  g00805(new_n3153, new_n3152, new_n3154);
nand_5 g00806(new_n3154, new_n3151, new_n3155);
xor_4  g00807(new_n3154, n25336, new_n3156);
xor_4  g00808(new_n3101, new_n3100, new_n3157);
or_5   g00809(new_n3157, new_n3156, new_n3158);
and_5  g00810(new_n3158, new_n3155, new_n3159);
or_5   g00811(new_n3159, new_n3150, new_n3160);
and_5  g00812(new_n3160, new_n3149, new_n3161_1);
or_5   g00813(new_n3161_1, new_n3145, new_n3162);
and_5  g00814(new_n3162, new_n3143, new_n3163);
or_5   g00815(new_n3163, new_n3141, new_n3164_1);
and_5  g00816(new_n3164_1, new_n3139, new_n3165);
or_5   g00817(new_n3165, new_n3137, new_n3166);
and_5  g00818(new_n3166, new_n3135, new_n3167);
or_5   g00819(new_n3167, new_n3133, new_n3168);
and_5  g00820(new_n3168, new_n3131, new_n3169);
or_5   g00821(new_n3169, new_n3129, new_n3170);
and_5  g00822(new_n3170, new_n3127, new_n3171);
or_5   g00823(new_n3171, new_n3125_1, new_n3172);
and_5  g00824(new_n3172, new_n3123, new_n3173);
or_5   g00825(new_n3173, new_n3121, new_n3174);
and_5  g00826(new_n3174, new_n3120, new_n3175);
nor_5  g00827(n7335, n4319, new_n3176);
not_10 g00828(new_n3176, new_n3177);
nor_5  g00829(new_n3117, new_n3077, new_n3178);
not_10 g00830(new_n3178, new_n3179);
and_5  g00831(new_n3179, new_n3177, new_n3180);
not_10 g00832(new_n3180, new_n3181);
and_5  g00833(new_n3181, new_n3175, new_n3182);
not_10 g00834(n3425, new_n3183);
not_10 g00835(n9967, new_n3184);
not_10 g00836(n20946, new_n3185);
not_10 g00837(n7751, new_n3186);
not_10 g00838(n26823, new_n3187);
not_10 g00839(n4812, new_n3188);
not_10 g00840(n24278, new_n3189);
not_10 g00841(n24618, new_n3190);
nor_5  g00842(n12315, n3952, new_n3191);
and_5  g00843(new_n3191, new_n3190, new_n3192);
and_5  g00844(new_n3192, new_n3189, new_n3193);
and_5  g00845(new_n3193, new_n3188, new_n3194);
and_5  g00846(new_n3194, new_n3187, new_n3195);
and_5  g00847(new_n3195, new_n3186, new_n3196);
and_5  g00848(new_n3196, new_n3185, new_n3197);
and_5  g00849(new_n3197, new_n3184, new_n3198);
xor_4  g00850(new_n3198, new_n3183, new_n3199);
not_10 g00851(new_n3199, new_n3200);
xor_4  g00852(new_n3173, new_n3121, new_n3201);
nor_5  g00853(new_n3201, new_n3200, new_n3202);
and_5  g00854(new_n3198, new_n3183, new_n3203);
not_10 g00855(new_n3203, new_n3204);
xor_4  g00856(new_n3201, new_n3199, new_n3205);
xor_4  g00857(new_n3197, new_n3184, new_n3206);
xor_4  g00858(new_n3171, new_n3125_1, new_n3207);
not_10 g00859(new_n3207, new_n3208_1);
nand_5 g00860(new_n3208_1, new_n3206, new_n3209);
xnor_4 g00861(new_n3208_1, new_n3206, new_n3210);
xor_4  g00862(new_n3196, new_n3185, new_n3211);
not_10 g00863(new_n3211, new_n3212);
xor_4  g00864(new_n3169, new_n3129, new_n3213);
or_5   g00865(new_n3213, new_n3212, new_n3214);
xor_4  g00866(new_n3213, new_n3211, new_n3215);
xor_4  g00867(new_n3195, new_n3186, new_n3216);
not_10 g00868(new_n3216, new_n3217);
xor_4  g00869(new_n3167, new_n3133, new_n3218);
or_5   g00870(new_n3218, new_n3217, new_n3219_1);
xor_4  g00871(new_n3218, new_n3216, new_n3220);
xor_4  g00872(new_n3194, new_n3187, new_n3221);
not_10 g00873(new_n3221, new_n3222);
xor_4  g00874(new_n3165, new_n3137, new_n3223);
or_5   g00875(new_n3223, new_n3222, new_n3224);
xor_4  g00876(new_n3223, new_n3221, new_n3225);
xor_4  g00877(new_n3193, new_n3188, new_n3226);
not_10 g00878(new_n3226, new_n3227);
xor_4  g00879(new_n3163, new_n3141, new_n3228_1);
or_5   g00880(new_n3228_1, new_n3227, new_n3229);
xor_4  g00881(new_n3228_1, new_n3226, new_n3230);
xor_4  g00882(new_n3192, new_n3189, new_n3231);
not_10 g00883(new_n3231, new_n3232);
xor_4  g00884(new_n3161_1, new_n3145, new_n3233);
or_5   g00885(new_n3233, new_n3232, new_n3234);
xor_4  g00886(new_n3233, new_n3231, new_n3235_1);
xor_4  g00887(new_n3191, new_n3190, new_n3236);
not_10 g00888(new_n3236, new_n3237);
xor_4  g00889(new_n3159, new_n3150, new_n3238);
or_5   g00890(new_n3238, new_n3237, new_n3239);
xor_4  g00891(new_n3238, new_n3236, new_n3240);
not_10 g00892(n3952, new_n3241);
xor_4  g00893(new_n3153, new_n3152, new_n3242);
not_10 g00894(new_n3242, new_n3243);
and_5  g00895(new_n3243, n12315, new_n3244_1);
nand_5 g00896(new_n3244_1, new_n3241, new_n3245);
xnor_4 g00897(new_n3157, new_n3156, new_n3246);
xor_4  g00898(n12315, n3952, new_n3247);
or_5   g00899(new_n3247, new_n3244_1, new_n3248);
and_5  g00900(new_n3248, new_n3245, new_n3249);
nand_5 g00901(new_n3249, new_n3246, new_n3250);
and_5  g00902(new_n3250, new_n3245, new_n3251);
or_5   g00903(new_n3251, new_n3240, new_n3252);
and_5  g00904(new_n3252, new_n3239, new_n3253_1);
or_5   g00905(new_n3253_1, new_n3235_1, new_n3254);
and_5  g00906(new_n3254, new_n3234, new_n3255);
or_5   g00907(new_n3255, new_n3230, new_n3256);
and_5  g00908(new_n3256, new_n3229, new_n3257);
or_5   g00909(new_n3257, new_n3225, new_n3258);
and_5  g00910(new_n3258, new_n3224, new_n3259);
or_5   g00911(new_n3259, new_n3220, new_n3260_1);
and_5  g00912(new_n3260_1, new_n3219_1, new_n3261);
or_5   g00913(new_n3261, new_n3215, new_n3262);
and_5  g00914(new_n3262, new_n3214, new_n3263_1);
or_5   g00915(new_n3263_1, new_n3210, new_n3264);
and_5  g00916(new_n3264, new_n3209, new_n3265);
or_5   g00917(new_n3265, new_n3205, new_n3266);
and_5  g00918(new_n3266, new_n3204, new_n3267);
not_10 g00919(new_n3267, new_n3268);
nor_5  g00920(new_n3268, new_n3202, new_n3269);
and_5  g00921(new_n3269, new_n3182, new_n3270);
or_5   g00922(n7593, n5101, new_n3271);
xor_4  g00923(n7593, n5101, new_n3272);
not_10 g00924(new_n3272, new_n3273);
or_5   g00925(n16507, n337, new_n3274);
xor_4  g00926(n16507, n337, new_n3275);
not_10 g00927(new_n3275, new_n3276);
or_5   g00928(n22470, n3228, new_n3277);
xor_4  g00929(n22470, n3228, new_n3278);
not_10 g00930(new_n3278, new_n3279_1);
or_5   g00931(n19116, n5302, new_n3280);
xnor_4 g00932(n19116, n5302, new_n3281);
or_5   g00933(n25738, n6861, new_n3282);
xor_4  g00934(n25738, n6861, new_n3283);
not_10 g00935(new_n3283, new_n3284);
or_5   g00936(n21471, n19357, new_n3285);
xor_4  g00937(n21471, n19357, new_n3286);
not_10 g00938(new_n3286, new_n3287);
or_5   g00939(n18737, n2328, new_n3288);
xor_4  g00940(n18737, n2328, new_n3289_1);
not_10 g00941(new_n3289_1, new_n3290);
or_5   g00942(n15053, n14603, new_n3291);
xor_4  g00943(n15053, n14603, new_n3292);
not_10 g00944(new_n3292, new_n3293);
or_5   g00945(n25471, n20794, new_n3294);
and_5  g00946(n23333, n16502, new_n3295);
not_10 g00947(new_n3295, new_n3296);
xor_4  g00948(n25471, n20794, new_n3297);
nand_5 g00949(new_n3297, new_n3296, new_n3298);
and_5  g00950(new_n3298, new_n3294, new_n3299);
or_5   g00951(new_n3299, new_n3293, new_n3300);
and_5  g00952(new_n3300, new_n3291, new_n3301_1);
or_5   g00953(new_n3301_1, new_n3290, new_n3302);
and_5  g00954(new_n3302, new_n3288, new_n3303);
or_5   g00955(new_n3303, new_n3287, new_n3304);
and_5  g00956(new_n3304, new_n3285, new_n3305);
or_5   g00957(new_n3305, new_n3284, new_n3306_1);
and_5  g00958(new_n3306_1, new_n3282, new_n3307);
or_5   g00959(new_n3307, new_n3281, new_n3308);
and_5  g00960(new_n3308, new_n3280, new_n3309);
or_5   g00961(new_n3309, new_n3279_1, new_n3310);
and_5  g00962(new_n3310, new_n3277, new_n3311);
or_5   g00963(new_n3311, new_n3276, new_n3312);
and_5  g00964(new_n3312, new_n3274, new_n3313);
or_5   g00965(new_n3313, new_n3273, new_n3314);
and_5  g00966(new_n3314, new_n3271, new_n3315);
xnor_4 g00967(new_n3180, new_n3175, new_n3316_1);
xor_4  g00968(new_n3316_1, new_n3269, new_n3317);
and_5  g00969(new_n3317, new_n3315, new_n3318);
or_5   g00970(new_n3317, new_n3315, new_n3319);
xor_4  g00971(new_n3265, new_n3205, new_n3320_1);
not_10 g00972(new_n3320_1, new_n3321);
xor_4  g00973(new_n3313, new_n3273, new_n3322);
and_5  g00974(new_n3322, new_n3321, new_n3323);
not_10 g00975(new_n3322, new_n3324_1);
xor_4  g00976(new_n3324_1, new_n3321, new_n3325);
xor_4  g00977(new_n3263_1, new_n3210, new_n3326);
not_10 g00978(new_n3326, new_n3327);
xor_4  g00979(new_n3311, new_n3276, new_n3328);
and_5  g00980(new_n3328, new_n3327, new_n3329);
not_10 g00981(new_n3328, new_n3330);
xor_4  g00982(new_n3330, new_n3327, new_n3331);
xor_4  g00983(new_n3261, new_n3215, new_n3332_1);
not_10 g00984(new_n3332_1, new_n3333);
xor_4  g00985(new_n3309, new_n3279_1, new_n3334);
and_5  g00986(new_n3334, new_n3333, new_n3335);
not_10 g00987(new_n3334, new_n3336);
xor_4  g00988(new_n3336, new_n3333, new_n3337);
xor_4  g00989(new_n3259, new_n3220, new_n3338);
not_10 g00990(new_n3338, new_n3339);
xor_4  g00991(new_n3307, new_n3281, new_n3340_1);
and_5  g00992(new_n3340_1, new_n3339, new_n3341);
xnor_4 g00993(new_n3340_1, new_n3339, new_n3342);
xor_4  g00994(new_n3257, new_n3225, new_n3343_1);
not_10 g00995(new_n3343_1, new_n3344);
xor_4  g00996(new_n3305, new_n3284, new_n3345);
and_5  g00997(new_n3345, new_n3344, new_n3346);
not_10 g00998(new_n3345, new_n3347);
xor_4  g00999(new_n3347, new_n3344, new_n3348);
xor_4  g01000(new_n3255, new_n3230, new_n3349_1);
not_10 g01001(new_n3349_1, new_n3350);
xor_4  g01002(new_n3303, new_n3287, new_n3351);
and_5  g01003(new_n3351, new_n3350, new_n3352);
not_10 g01004(new_n3351, new_n3353);
xor_4  g01005(new_n3353, new_n3350, new_n3354);
xor_4  g01006(new_n3253_1, new_n3235_1, new_n3355);
not_10 g01007(new_n3355, new_n3356);
xor_4  g01008(new_n3301_1, new_n3290, new_n3357);
and_5  g01009(new_n3357, new_n3356, new_n3358);
not_10 g01010(new_n3357, new_n3359);
xor_4  g01011(new_n3359, new_n3356, new_n3360);
xor_4  g01012(new_n3251, new_n3240, new_n3361);
not_10 g01013(new_n3361, new_n3362);
xor_4  g01014(new_n3299, new_n3293, new_n3363);
and_5  g01015(new_n3363, new_n3362, new_n3364);
not_10 g01016(new_n3363, new_n3365);
xor_4  g01017(new_n3365, new_n3362, new_n3366_1);
xor_4  g01018(n23333, n16502, new_n3367);
xor_4  g01019(new_n3243, n12315, new_n3368);
and_5  g01020(new_n3368, new_n3367, new_n3369);
xnor_4 g01021(new_n3297, new_n3295, new_n3370);
not_10 g01022(new_n3370, new_n3371);
nor_5  g01023(new_n3371, new_n3369, new_n3372);
xor_4  g01024(new_n3249, new_n3246, new_n3373);
not_10 g01025(new_n3373, new_n3374);
and_5  g01026(new_n3369, new_n3297, new_n3375);
nor_5  g01027(new_n3375, new_n3372, new_n3376);
and_5  g01028(new_n3376, new_n3374, new_n3377);
nor_5  g01029(new_n3377, new_n3372, new_n3378);
nor_5  g01030(new_n3378, new_n3366_1, new_n3379);
nor_5  g01031(new_n3379, new_n3364, new_n3380);
nor_5  g01032(new_n3380, new_n3360, new_n3381);
nor_5  g01033(new_n3381, new_n3358, new_n3382);
nor_5  g01034(new_n3382, new_n3354, new_n3383);
nor_5  g01035(new_n3383, new_n3352, new_n3384);
nor_5  g01036(new_n3384, new_n3348, new_n3385);
nor_5  g01037(new_n3385, new_n3346, new_n3386);
nor_5  g01038(new_n3386, new_n3342, new_n3387);
nor_5  g01039(new_n3387, new_n3341, new_n3388);
nor_5  g01040(new_n3388, new_n3337, new_n3389);
nor_5  g01041(new_n3389, new_n3335, new_n3390_1);
nor_5  g01042(new_n3390_1, new_n3331, new_n3391);
nor_5  g01043(new_n3391, new_n3329, new_n3392);
nor_5  g01044(new_n3392, new_n3325, new_n3393);
nor_5  g01045(new_n3393, new_n3323, new_n3394);
and_5  g01046(new_n3394, new_n3319, new_n3395);
nor_5  g01047(new_n3395, new_n3318, new_n3396);
not_10 g01048(new_n3396, new_n3397);
nand_5 g01049(new_n3397, new_n3270, new_n3398);
not_10 g01050(new_n3182, new_n3399);
or_5   g01051(new_n3269, new_n3399, new_n3400);
nor_5  g01052(new_n3181, new_n3175, new_n3401);
nand_5 g01053(new_n3401, new_n3269, new_n3402);
and_5  g01054(new_n3402, new_n3400, new_n3403);
and_5  g01055(new_n3403, new_n3397, new_n3404);
or_5   g01056(new_n3404, new_n3270, new_n3405);
and_5  g01057(new_n3405, new_n3398, n175);
not_10 g01058(n26180, new_n3407);
not_10 g01059(n25494, new_n3408);
not_10 g01060(n8856, new_n3409);
not_10 g01061(n14130, new_n3410);
not_10 g01062(n16482, new_n3411);
not_10 g01063(n9942, new_n3412);
not_10 g01064(n25643, new_n3413);
not_10 g01065(n9557, new_n3414);
not_10 g01066(n3136, new_n3415);
nor_5  g01067(n20138, n9251, new_n3416);
and_5  g01068(new_n3416, new_n2361_1, new_n3417);
and_5  g01069(new_n3417, new_n3415, new_n3418);
and_5  g01070(new_n3418, new_n3414, new_n3419);
and_5  g01071(new_n3419, new_n3413, new_n3420);
and_5  g01072(new_n3420, new_n3412, new_n3421);
and_5  g01073(new_n3421, new_n3411, new_n3422);
and_5  g01074(new_n3422, new_n3410, new_n3423);
xor_4  g01075(new_n3423, new_n3409, new_n3424);
xor_4  g01076(new_n3424, new_n3408, new_n3425_1);
xor_4  g01077(new_n3422, new_n3410, new_n3426_1);
nor_5  g01078(new_n3426_1, n10117, new_n3427);
xnor_4 g01079(new_n3426_1, n10117, new_n3428);
xor_4  g01080(new_n3421, new_n3411, new_n3429);
or_5   g01081(new_n3429, n13460, new_n3430);
xnor_4 g01082(new_n3429, n13460, new_n3431);
xor_4  g01083(new_n3420, new_n3412, new_n3432);
or_5   g01084(new_n3432, n6104, new_n3433);
xnor_4 g01085(new_n3432, n6104, new_n3434);
xor_4  g01086(new_n3419, new_n3413, new_n3435);
or_5   g01087(new_n3435, n4119, new_n3436);
not_10 g01088(n4119, new_n3437);
xor_4  g01089(new_n3435, new_n3437, new_n3438);
xor_4  g01090(new_n3418, new_n3414, new_n3439);
or_5   g01091(new_n3439, n14510, new_n3440);
xor_4  g01092(new_n3439, n14510, new_n3441);
not_10 g01093(new_n3441, new_n3442);
xor_4  g01094(new_n3417, new_n3415, new_n3443);
or_5   g01095(new_n3443, n13263, new_n3444);
xor_4  g01096(new_n3416, new_n2361_1, new_n3445);
nor_5  g01097(new_n3445, n20455, new_n3446);
xor_4  g01098(new_n3445, n20455, new_n3447);
not_10 g01099(new_n3447, new_n3448);
xor_4  g01100(n20138, n9251, new_n3449);
or_5   g01101(new_n3449, n1639, new_n3450);
and_5  g01102(n16968, n9251, new_n3451_1);
not_10 g01103(new_n3451_1, new_n3452);
xor_4  g01104(new_n3449, n1639, new_n3453);
nand_5 g01105(new_n3453, new_n3452, new_n3454);
and_5  g01106(new_n3454, new_n3450, new_n3455);
nor_5  g01107(new_n3455, new_n3448, new_n3456);
or_5   g01108(new_n3456, new_n3446, new_n3457);
xor_4  g01109(new_n3443, n13263, new_n3458);
nand_5 g01110(new_n3458, new_n3457, new_n3459_1);
and_5  g01111(new_n3459_1, new_n3444, new_n3460_1);
or_5   g01112(new_n3460_1, new_n3442, new_n3461);
and_5  g01113(new_n3461, new_n3440, new_n3462);
or_5   g01114(new_n3462, new_n3438, new_n3463);
and_5  g01115(new_n3463, new_n3436, new_n3464);
or_5   g01116(new_n3464, new_n3434, new_n3465);
and_5  g01117(new_n3465, new_n3433, new_n3466);
or_5   g01118(new_n3466, new_n3431, new_n3467);
and_5  g01119(new_n3467, new_n3430, new_n3468_1);
nor_5  g01120(new_n3468_1, new_n3428, new_n3469);
nor_5  g01121(new_n3469, new_n3427, new_n3470);
xor_4  g01122(new_n3470, new_n3425_1, new_n3471);
xor_4  g01123(new_n3471, new_n3407, new_n3472);
not_10 g01124(new_n3472, new_n3473);
not_10 g01125(n24004, new_n3474);
xor_4  g01126(new_n3468_1, new_n3428, new_n3475);
nand_5 g01127(new_n3475, new_n3474, new_n3476);
xor_4  g01128(new_n3475, new_n3474, new_n3477);
not_10 g01129(new_n3477, new_n3478);
not_10 g01130(n12871, new_n3479);
xor_4  g01131(new_n3466, new_n3431, new_n3480_1);
nand_5 g01132(new_n3480_1, new_n3479, new_n3481);
xor_4  g01133(new_n3480_1, new_n3479, new_n3482);
not_10 g01134(new_n3482, new_n3483);
not_10 g01135(n23304, new_n3484);
xor_4  g01136(new_n3464, new_n3434, new_n3485);
nand_5 g01137(new_n3485, new_n3484, new_n3486);
xor_4  g01138(new_n3485, new_n3484, new_n3487);
not_10 g01139(new_n3487, new_n3488);
not_10 g01140(n19361, new_n3489);
xor_4  g01141(new_n3462, new_n3438, new_n3490);
nand_5 g01142(new_n3490, new_n3489, new_n3491);
xor_4  g01143(new_n3490, new_n3489, new_n3492);
not_10 g01144(new_n3492, new_n3493);
xor_4  g01145(new_n3460_1, new_n3442, new_n3494);
not_10 g01146(new_n3494, new_n3495);
or_5   g01147(new_n3495, n1437, new_n3496);
xor_4  g01148(new_n3495, n1437, new_n3497);
not_10 g01149(new_n3497, new_n3498);
not_10 g01150(n4722, new_n3499);
xor_4  g01151(new_n3458, new_n3457, new_n3500);
nand_5 g01152(new_n3500, new_n3499, new_n3501);
xor_4  g01153(new_n3500, new_n3499, new_n3502_1);
xor_4  g01154(new_n3455, new_n3448, new_n3503);
not_10 g01155(new_n3503, new_n3504);
nand_5 g01156(new_n3504, n14633, new_n3505);
xor_4  g01157(new_n3504, n14633, new_n3506_1);
xor_4  g01158(new_n3453, new_n3452, new_n3507);
not_10 g01159(new_n3507, new_n3508);
nand_5 g01160(new_n3508, n8721, new_n3509);
xor_4  g01161(n16968, n9251, new_n3510);
and_5  g01162(new_n3510, n18578, new_n3511);
xor_4  g01163(new_n3508, n8721, new_n3512);
nand_5 g01164(new_n3512, new_n3511, new_n3513);
nand_5 g01165(new_n3513, new_n3509, new_n3514);
nand_5 g01166(new_n3514, new_n3506_1, new_n3515);
and_5  g01167(new_n3515, new_n3505, new_n3516_1);
nand_5 g01168(new_n3516_1, new_n3502_1, new_n3517);
and_5  g01169(new_n3517, new_n3501, new_n3518);
or_5   g01170(new_n3518, new_n3498, new_n3519);
and_5  g01171(new_n3519, new_n3496, new_n3520);
or_5   g01172(new_n3520, new_n3493, new_n3521);
and_5  g01173(new_n3521, new_n3491, new_n3522);
or_5   g01174(new_n3522, new_n3488, new_n3523);
and_5  g01175(new_n3523, new_n3486, new_n3524);
or_5   g01176(new_n3524, new_n3483, new_n3525);
and_5  g01177(new_n3525, new_n3481, new_n3526);
or_5   g01178(new_n3526, new_n3478, new_n3527);
and_5  g01179(new_n3527, new_n3476, new_n3528_1);
xor_4  g01180(new_n3528_1, new_n3473, new_n3529);
not_10 g01181(new_n3529, new_n3530);
xnor_4 g01182(n3506, n2743, new_n3531);
not_10 g01183(new_n3531, new_n3532);
not_10 g01184(n7026, new_n3533);
or_5   g01185(n14899, new_n3533, new_n3534);
xnor_4 g01186(n14899, n7026, new_n3535);
not_10 g01187(new_n3535, new_n3536);
not_10 g01188(n13719, new_n3537);
or_5   g01189(n18444, new_n3537, new_n3538);
xnor_4 g01190(n18444, n13719, new_n3539);
not_10 g01191(new_n3539, new_n3540);
not_10 g01192(n442, new_n3541_1);
or_5   g01193(n24638, new_n3541_1, new_n3542);
xnor_4 g01194(n24638, n442, new_n3543);
not_10 g01195(new_n3543, new_n3544);
not_10 g01196(n9172, new_n3545);
or_5   g01197(n21674, new_n3545, new_n3546);
xnor_4 g01198(n21674, n9172, new_n3547);
not_10 g01199(new_n3547, new_n3548);
not_10 g01200(n4913, new_n3549);
or_5   g01201(n17251, new_n3549, new_n3550);
xnor_4 g01202(n17251, n4913, new_n3551);
not_10 g01203(new_n3551, new_n3552);
not_10 g01204(n604, new_n3553);
or_5   g01205(n14790, new_n3553, new_n3554);
xnor_4 g01206(n14790, n604, new_n3555_1);
not_10 g01207(n10096, new_n3556);
or_5   g01208(n16824, new_n3556, new_n3557);
not_10 g01209(n16824, new_n3558);
or_5   g01210(new_n3558, n10096, new_n3559);
not_10 g01211(n16521, new_n3560);
and_5  g01212(n16994, new_n3560, new_n3561_1);
nor_5  g01213(n16994, new_n3560, new_n3562);
not_10 g01214(new_n3562, new_n3563_1);
not_10 g01215(n7139, new_n3564);
and_5  g01216(n9246, new_n3564, new_n3565);
and_5  g01217(new_n3565, new_n3563_1, new_n3566);
nor_5  g01218(new_n3566, new_n3561_1, new_n3567);
not_10 g01219(new_n3567, new_n3568);
nand_5 g01220(new_n3568, new_n3559, new_n3569);
and_5  g01221(new_n3569, new_n3557, new_n3570_1);
nand_5 g01222(new_n3570_1, new_n3555_1, new_n3571);
and_5  g01223(new_n3571, new_n3554, new_n3572);
or_5   g01224(new_n3572, new_n3552, new_n3573);
and_5  g01225(new_n3573, new_n3550, new_n3574);
or_5   g01226(new_n3574, new_n3548, new_n3575);
and_5  g01227(new_n3575, new_n3546, new_n3576);
or_5   g01228(new_n3576, new_n3544, new_n3577);
and_5  g01229(new_n3577, new_n3542, new_n3578);
or_5   g01230(new_n3578, new_n3540, new_n3579);
and_5  g01231(new_n3579, new_n3538, new_n3580);
or_5   g01232(new_n3580, new_n3536, new_n3581);
and_5  g01233(new_n3581, new_n3534, new_n3582_1);
xor_4  g01234(new_n3582_1, new_n3532, new_n3583);
not_10 g01235(n9259, new_n3584);
not_10 g01236(n21489, new_n3585);
not_10 g01237(n20213, new_n3586);
not_10 g01238(n13912, new_n3587);
not_10 g01239(n7670, new_n3588);
not_10 g01240(n9598, new_n3589);
not_10 g01241(n22290, new_n3590);
not_10 g01242(n11273, new_n3591);
nor_5  g01243(n25565, n21993, new_n3592);
and_5  g01244(new_n3592, new_n3591, new_n3593);
and_5  g01245(new_n3593, new_n3590, new_n3594);
and_5  g01246(new_n3594, new_n3589, new_n3595);
and_5  g01247(new_n3595, new_n3588, new_n3596);
and_5  g01248(new_n3596, new_n3587, new_n3597);
and_5  g01249(new_n3597, new_n3586, new_n3598);
and_5  g01250(new_n3598, new_n3585, new_n3599);
xor_4  g01251(new_n3599, new_n3584, new_n3600);
xnor_4 g01252(new_n3600, new_n3583, new_n3601);
xor_4  g01253(new_n3580, new_n3536, new_n3602);
xor_4  g01254(new_n3598, new_n3585, new_n3603);
nand_5 g01255(new_n3603, new_n3602, new_n3604);
xor_4  g01256(new_n3603, new_n3602, new_n3605);
xor_4  g01257(new_n3578, new_n3540, new_n3606);
xor_4  g01258(new_n3597, new_n3586, new_n3607);
or_5   g01259(new_n3607, new_n3606, new_n3608);
xnor_4 g01260(new_n3607, new_n3606, new_n3609);
xor_4  g01261(new_n3576, new_n3544, new_n3610);
xor_4  g01262(new_n3596, new_n3587, new_n3611);
or_5   g01263(new_n3611, new_n3610, new_n3612);
xnor_4 g01264(new_n3611, new_n3610, new_n3613);
xor_4  g01265(new_n3574, new_n3548, new_n3614);
xor_4  g01266(new_n3595, new_n3588, new_n3615);
or_5   g01267(new_n3615, new_n3614, new_n3616);
xnor_4 g01268(new_n3615, new_n3614, new_n3617_1);
xor_4  g01269(new_n3594, new_n3589, new_n3618_1);
xor_4  g01270(new_n3572, new_n3552, new_n3619);
or_5   g01271(new_n3619, new_n3618_1, new_n3620);
not_10 g01272(new_n3619, new_n3621);
xor_4  g01273(new_n3621, new_n3618_1, new_n3622);
xor_4  g01274(new_n3593, new_n3590, new_n3623);
xor_4  g01275(new_n3570_1, new_n3555_1, new_n3624);
or_5   g01276(new_n3624, new_n3623, new_n3625);
xor_4  g01277(new_n3592, new_n3591, new_n3626);
not_10 g01278(new_n3626, new_n3627);
xnor_4 g01279(n16824, n10096, new_n3628);
xor_4  g01280(new_n3628, new_n3568, new_n3629);
and_5  g01281(new_n3629, new_n3627, new_n3630);
xor_4  g01282(new_n3629, new_n3626, new_n3631);
xor_4  g01283(n25565, n21993, new_n3632);
not_10 g01284(new_n3632, new_n3633);
xnor_4 g01285(n16994, n16521, new_n3634);
xor_4  g01286(new_n3634, new_n3565, new_n3635);
nand_5 g01287(new_n3635, new_n3633, new_n3636);
not_10 g01288(n21993, new_n3637);
xnor_4 g01289(n9246, n7139, new_n3638);
nor_5  g01290(new_n3638, new_n3637, new_n3639);
not_10 g01291(new_n3639, new_n3640);
xnor_4 g01292(new_n3635, new_n3632, new_n3641);
nand_5 g01293(new_n3641, new_n3640, new_n3642_1);
and_5  g01294(new_n3642_1, new_n3636, new_n3643);
nor_5  g01295(new_n3643, new_n3631, new_n3644);
or_5   g01296(new_n3644, new_n3630, new_n3645);
not_10 g01297(new_n3624, new_n3646);
xnor_4 g01298(new_n3646, new_n3623, new_n3647);
nand_5 g01299(new_n3647, new_n3645, new_n3648);
and_5  g01300(new_n3648, new_n3625, new_n3649_1);
or_5   g01301(new_n3649_1, new_n3622, new_n3650);
and_5  g01302(new_n3650, new_n3620, new_n3651);
or_5   g01303(new_n3651, new_n3617_1, new_n3652);
and_5  g01304(new_n3652, new_n3616, new_n3653);
or_5   g01305(new_n3653, new_n3613, new_n3654);
and_5  g01306(new_n3654, new_n3612, new_n3655);
or_5   g01307(new_n3655, new_n3609, new_n3656);
and_5  g01308(new_n3656, new_n3608, new_n3657);
nand_5 g01309(new_n3657, new_n3605, new_n3658);
and_5  g01310(new_n3658, new_n3604, new_n3659);
xor_4  g01311(new_n3659, new_n3601, new_n3660);
xor_4  g01312(new_n3660, new_n3530, new_n3661);
xor_4  g01313(new_n3526, new_n3478, new_n3662);
not_10 g01314(new_n3662, new_n3663);
xor_4  g01315(new_n3657, new_n3605, new_n3664);
or_5   g01316(new_n3664, new_n3663, new_n3665_1);
xor_4  g01317(new_n3664, new_n3663, new_n3666);
xor_4  g01318(new_n3524, new_n3483, new_n3667);
xor_4  g01319(new_n3655, new_n3609, new_n3668);
nand_5 g01320(new_n3668, new_n3667, new_n3669);
xor_4  g01321(new_n3668, new_n3667, new_n3670);
not_10 g01322(new_n3670, new_n3671);
xor_4  g01323(new_n3522, new_n3488, new_n3672);
xor_4  g01324(new_n3653, new_n3613, new_n3673);
nand_5 g01325(new_n3673, new_n3672, new_n3674);
xor_4  g01326(new_n3673, new_n3672, new_n3675);
not_10 g01327(new_n3675, new_n3676);
xor_4  g01328(new_n3520, new_n3493, new_n3677);
xor_4  g01329(new_n3651, new_n3617_1, new_n3678);
nand_5 g01330(new_n3678, new_n3677, new_n3679_1);
xor_4  g01331(new_n3678, new_n3677, new_n3680);
not_10 g01332(new_n3680, new_n3681);
xnor_4 g01333(new_n3518, new_n3497, new_n3682);
xor_4  g01334(new_n3649_1, new_n3622, new_n3683);
nand_5 g01335(new_n3683, new_n3682, new_n3684);
not_10 g01336(new_n3682, new_n3685);
xnor_4 g01337(new_n3683, new_n3685, new_n3686);
xor_4  g01338(new_n3516_1, new_n3502_1, new_n3687);
xor_4  g01339(new_n3647, new_n3645, new_n3688);
nand_5 g01340(new_n3688, new_n3687, new_n3689);
not_10 g01341(new_n3687, new_n3690);
xnor_4 g01342(new_n3688, new_n3690, new_n3691);
and_5  g01343(new_n3513, new_n3509, new_n3692);
xnor_4 g01344(new_n3692, new_n3506_1, new_n3693);
not_10 g01345(new_n3693, new_n3694);
xor_4  g01346(new_n3643, new_n3631, new_n3695);
nand_5 g01347(new_n3695, new_n3694, new_n3696);
xor_4  g01348(new_n3695, new_n3694, new_n3697);
not_10 g01349(new_n3697, new_n3698);
xor_4  g01350(new_n3641, new_n3640, new_n3699);
not_10 g01351(new_n3699, new_n3700);
xor_4  g01352(new_n3512, new_n3511, new_n3701);
or_5   g01353(new_n3701, new_n3700, new_n3702);
xor_4  g01354(new_n3510, n18578, new_n3703);
xor_4  g01355(new_n3638, new_n3637, new_n3704);
nand_5 g01356(new_n3704, new_n3703, new_n3705);
xor_4  g01357(new_n3701, new_n3700, new_n3706);
nand_5 g01358(new_n3706, new_n3705, new_n3707);
and_5  g01359(new_n3707, new_n3702, new_n3708);
or_5   g01360(new_n3708, new_n3698, new_n3709);
nand_5 g01361(new_n3709, new_n3696, new_n3710_1);
nand_5 g01362(new_n3710_1, new_n3691, new_n3711);
nand_5 g01363(new_n3711, new_n3689, new_n3712);
nand_5 g01364(new_n3712, new_n3686, new_n3713);
and_5  g01365(new_n3713, new_n3684, new_n3714);
or_5   g01366(new_n3714, new_n3681, new_n3715);
and_5  g01367(new_n3715, new_n3679_1, new_n3716);
or_5   g01368(new_n3716, new_n3676, new_n3717);
and_5  g01369(new_n3717, new_n3674, new_n3718);
or_5   g01370(new_n3718, new_n3671, new_n3719);
nand_5 g01371(new_n3719, new_n3669, new_n3720);
nand_5 g01372(new_n3720, new_n3666, new_n3721);
nand_5 g01373(new_n3721, new_n3665_1, new_n3722);
xnor_4 g01374(new_n3722, new_n3661, n235);
not_10 g01375(n19327, new_n3724);
not_10 g01376(n2113, new_n3725_1);
not_10 g01377(n21134, new_n3726);
not_10 g01378(n6369, new_n3727);
not_10 g01379(n25797, new_n3728);
not_10 g01380(n15967, new_n3729);
nor_5  g01381(n25435, n13319, new_n3730);
and_5  g01382(new_n3730, new_n3729, new_n3731);
and_5  g01383(new_n3731, new_n3728, new_n3732);
and_5  g01384(new_n3732, new_n3727, new_n3733_1);
and_5  g01385(new_n3733_1, new_n3726, new_n3734);
xor_4  g01386(new_n3734, new_n3725_1, new_n3735);
xor_4  g01387(new_n3735, new_n3724, new_n3736);
xor_4  g01388(new_n3733_1, new_n3726, new_n3737);
or_5   g01389(new_n3737, n22597, new_n3738);
not_10 g01390(n22597, new_n3739);
xor_4  g01391(new_n3737, new_n3739, new_n3740_1);
xor_4  g01392(new_n3732, new_n3727, new_n3741);
or_5   g01393(new_n3741, n26107, new_n3742);
xor_4  g01394(new_n3741, n26107, new_n3743);
not_10 g01395(new_n3743, new_n3744);
xor_4  g01396(new_n3731, new_n3728, new_n3745);
or_5   g01397(new_n3745, n342, new_n3746);
xor_4  g01398(new_n3730, new_n3729, new_n3747);
nor_5  g01399(new_n3747, n26553, new_n3748);
xor_4  g01400(new_n3747, n26553, new_n3749);
not_10 g01401(new_n3749, new_n3750);
xor_4  g01402(n25435, n13319, new_n3751);
or_5   g01403(new_n3751, n4964, new_n3752);
and_5  g01404(n25435, n7876, new_n3753);
not_10 g01405(new_n3753, new_n3754);
xor_4  g01406(new_n3751, n4964, new_n3755_1);
nand_5 g01407(new_n3755_1, new_n3754, new_n3756);
and_5  g01408(new_n3756, new_n3752, new_n3757);
nor_5  g01409(new_n3757, new_n3750, new_n3758_1);
or_5   g01410(new_n3758_1, new_n3748, new_n3759);
xor_4  g01411(new_n3745, n342, new_n3760_1);
nand_5 g01412(new_n3760_1, new_n3759, new_n3761);
and_5  g01413(new_n3761, new_n3746, new_n3762);
or_5   g01414(new_n3762, new_n3744, new_n3763);
and_5  g01415(new_n3763, new_n3742, new_n3764);
or_5   g01416(new_n3764, new_n3740_1, new_n3765);
and_5  g01417(new_n3765, new_n3738, new_n3766);
xor_4  g01418(new_n3766, new_n3736, new_n3767);
xor_4  g01419(new_n3767, n25749, new_n3768);
not_10 g01420(n3161, new_n3769);
xor_4  g01421(new_n3764, new_n3740_1, new_n3770);
or_5   g01422(new_n3770, new_n3769, new_n3771);
xor_4  g01423(new_n3770, n3161, new_n3772);
xor_4  g01424(new_n3762, new_n3744, new_n3773);
not_10 g01425(new_n3773, new_n3774);
nand_5 g01426(new_n3774, n9003, new_n3775);
not_10 g01427(n9003, new_n3776);
xor_4  g01428(new_n3774, new_n3776, new_n3777);
not_10 g01429(n4957, new_n3778);
xor_4  g01430(new_n3760_1, new_n3759, new_n3779);
or_5   g01431(new_n3779, new_n3778, new_n3780);
xor_4  g01432(new_n3779, n4957, new_n3781_1);
xor_4  g01433(new_n3757, new_n3750, new_n3782);
not_10 g01434(new_n3782, new_n3783);
nand_5 g01435(new_n3783, n7524, new_n3784);
not_10 g01436(n7524, new_n3785_1);
xor_4  g01437(new_n3783, new_n3785_1, new_n3786);
xor_4  g01438(new_n3755_1, new_n3754, new_n3787);
not_10 g01439(new_n3787, new_n3788);
nand_5 g01440(new_n3788, n15743, new_n3789);
xor_4  g01441(n25435, n7876, new_n3790);
and_5  g01442(new_n3790, n20658, new_n3791);
xor_4  g01443(new_n3788, n15743, new_n3792);
nand_5 g01444(new_n3792, new_n3791, new_n3793);
and_5  g01445(new_n3793, new_n3789, new_n3794_1);
or_5   g01446(new_n3794_1, new_n3786, new_n3795_1);
and_5  g01447(new_n3795_1, new_n3784, new_n3796);
or_5   g01448(new_n3796, new_n3781_1, new_n3797);
and_5  g01449(new_n3797, new_n3780, new_n3798);
or_5   g01450(new_n3798, new_n3777, new_n3799);
and_5  g01451(new_n3799, new_n3775, new_n3800);
or_5   g01452(new_n3800, new_n3772, new_n3801);
and_5  g01453(new_n3801, new_n3771, new_n3802);
xor_4  g01454(new_n3802, new_n3768, new_n3803);
xnor_4 g01455(n26510, n22332, new_n3804);
not_10 g01456(new_n3804, new_n3805);
not_10 g01457(n18907, new_n3806);
or_5   g01458(n23068, new_n3806, new_n3807);
xnor_4 g01459(n23068, n18907, new_n3808);
not_10 g01460(new_n3808, new_n3809);
not_10 g01461(n2731, new_n3810);
or_5   g01462(n19514, new_n3810, new_n3811);
xnor_4 g01463(n19514, n2731, new_n3812);
not_10 g01464(new_n3812, new_n3813);
not_10 g01465(n19911, new_n3814);
or_5   g01466(new_n3814, n10053, new_n3815);
xnor_4 g01467(n19911, n10053, new_n3816);
not_10 g01468(n8399, new_n3817);
or_5   g01469(n13708, new_n3817, new_n3818);
not_10 g01470(n13708, new_n3819);
or_5   g01471(new_n3819, n8399, new_n3820);
not_10 g01472(n18409, new_n3821);
and_5  g01473(new_n3821, n9507, new_n3822);
not_10 g01474(n9507, new_n3823);
and_5  g01475(n18409, new_n3823, new_n3824);
not_10 g01476(new_n3824, new_n3825);
not_10 g01477(n5704, new_n3826);
and_5  g01478(n26979, new_n3826, new_n3827);
and_5  g01479(new_n3827, new_n3825, new_n3828_1);
nor_5  g01480(new_n3828_1, new_n3822, new_n3829);
not_10 g01481(new_n3829, new_n3830);
nand_5 g01482(new_n3830, new_n3820, new_n3831);
and_5  g01483(new_n3831, new_n3818, new_n3832);
nand_5 g01484(new_n3832, new_n3816, new_n3833);
and_5  g01485(new_n3833, new_n3815, new_n3834);
or_5   g01486(new_n3834, new_n3813, new_n3835);
and_5  g01487(new_n3835, new_n3811, new_n3836);
or_5   g01488(new_n3836, new_n3809, new_n3837);
and_5  g01489(new_n3837, new_n3807, new_n3838);
xor_4  g01490(new_n3838, new_n3805, new_n3839);
not_10 g01491(new_n3839, new_n3840);
not_10 g01492(n4325, new_n3841);
not_10 g01493(n5337, new_n3842_1);
not_10 g01494(n626, new_n3843);
not_10 g01495(n1204, new_n3844);
not_10 g01496(n19618, new_n3845);
nor_5  g01497(n22043, n12121, new_n3846);
and_5  g01498(new_n3846, new_n3845, new_n3847);
and_5  g01499(new_n3847, new_n3844, new_n3848);
and_5  g01500(new_n3848, new_n3843, new_n3849);
and_5  g01501(new_n3849, new_n3842_1, new_n3850_1);
xor_4  g01502(new_n3850_1, new_n3841, new_n3851);
xnor_4 g01503(new_n3851, new_n3840, new_n3852);
not_10 g01504(new_n3852, new_n3853);
xor_4  g01505(new_n3836, new_n3809, new_n3854);
xor_4  g01506(new_n3849, new_n3842_1, new_n3855);
or_5   g01507(new_n3855, new_n3854, new_n3856);
not_10 g01508(new_n3854, new_n3857);
xnor_4 g01509(new_n3855, new_n3857, new_n3858);
not_10 g01510(new_n3858, new_n3859);
xor_4  g01511(new_n3834, new_n3813, new_n3860);
xor_4  g01512(new_n3848, new_n3843, new_n3861);
or_5   g01513(new_n3861, new_n3860, new_n3862);
not_10 g01514(new_n3860, new_n3863);
xnor_4 g01515(new_n3861, new_n3863, new_n3864);
not_10 g01516(new_n3864, new_n3865);
xor_4  g01517(new_n3847, new_n3844, new_n3866);
xor_4  g01518(new_n3832, new_n3816, new_n3867);
or_5   g01519(new_n3867, new_n3866, new_n3868);
xor_4  g01520(new_n3867, new_n3866, new_n3869_1);
not_10 g01521(new_n3869_1, new_n3870);
xor_4  g01522(new_n3846, new_n3845, new_n3871_1);
not_10 g01523(new_n3871_1, new_n3872);
xnor_4 g01524(n13708, n8399, new_n3873);
xor_4  g01525(new_n3873, new_n3830, new_n3874);
nand_5 g01526(new_n3874, new_n3872, new_n3875);
xor_4  g01527(new_n3874, new_n3872, new_n3876);
xnor_4 g01528(n22043, n12121, new_n3877);
xnor_4 g01529(n18409, n9507, new_n3878);
xor_4  g01530(new_n3878, new_n3827, new_n3879);
or_5   g01531(new_n3879, new_n3877, new_n3880);
not_10 g01532(n12121, new_n3881);
xnor_4 g01533(n26979, n5704, new_n3882);
nor_5  g01534(new_n3882, new_n3881, new_n3883);
xor_4  g01535(new_n3879, new_n3877, new_n3884);
nand_5 g01536(new_n3884, new_n3883, new_n3885);
and_5  g01537(new_n3885, new_n3880, new_n3886);
nand_5 g01538(new_n3886, new_n3876, new_n3887);
and_5  g01539(new_n3887, new_n3875, new_n3888);
or_5   g01540(new_n3888, new_n3870, new_n3889);
and_5  g01541(new_n3889, new_n3868, new_n3890);
or_5   g01542(new_n3890, new_n3865, new_n3891_1);
and_5  g01543(new_n3891_1, new_n3862, new_n3892);
or_5   g01544(new_n3892, new_n3859, new_n3893);
and_5  g01545(new_n3893, new_n3856, new_n3894);
xor_4  g01546(new_n3894, new_n3853, new_n3895);
xnor_4 g01547(new_n3895, new_n3803, new_n3896);
xor_4  g01548(new_n3892, new_n3859, new_n3897);
not_10 g01549(new_n3897, new_n3898);
xor_4  g01550(new_n3800, new_n3772, new_n3899);
or_5   g01551(new_n3899, new_n3898, new_n3900);
xor_4  g01552(new_n3899, new_n3898, new_n3901);
xor_4  g01553(new_n3890, new_n3865, new_n3902);
not_10 g01554(new_n3902, new_n3903);
xor_4  g01555(new_n3798, new_n3777, new_n3904);
or_5   g01556(new_n3904, new_n3903, new_n3905);
xor_4  g01557(new_n3904, new_n3903, new_n3906);
xor_4  g01558(new_n3888, new_n3870, new_n3907);
not_10 g01559(new_n3907, new_n3908);
xor_4  g01560(new_n3796, new_n3781_1, new_n3909_1);
or_5   g01561(new_n3909_1, new_n3908, new_n3910);
xor_4  g01562(new_n3909_1, new_n3908, new_n3911);
xor_4  g01563(new_n3886, new_n3876, new_n3912);
not_10 g01564(new_n3912, new_n3913);
xor_4  g01565(new_n3794_1, new_n3786, new_n3914);
or_5   g01566(new_n3914, new_n3913, new_n3915);
xor_4  g01567(new_n3914, new_n3913, new_n3916);
xor_4  g01568(new_n3884, new_n3883, new_n3917);
xor_4  g01569(new_n3792, new_n3791, new_n3918_1);
or_5   g01570(new_n3918_1, new_n3917, new_n3919);
xor_4  g01571(new_n3790, n20658, new_n3920);
xor_4  g01572(new_n3882, new_n3881, new_n3921);
and_5  g01573(new_n3921, new_n3920, new_n3922);
xor_4  g01574(new_n3918_1, new_n3917, new_n3923);
not_10 g01575(new_n3923, new_n3924);
or_5   g01576(new_n3924, new_n3922, new_n3925_1);
nand_5 g01577(new_n3925_1, new_n3919, new_n3926);
nand_5 g01578(new_n3926, new_n3916, new_n3927);
nand_5 g01579(new_n3927, new_n3915, new_n3928);
nand_5 g01580(new_n3928, new_n3911, new_n3929);
nand_5 g01581(new_n3929, new_n3910, new_n3930);
nand_5 g01582(new_n3930, new_n3906, new_n3931);
nand_5 g01583(new_n3931, new_n3905, new_n3932_1);
nand_5 g01584(new_n3932_1, new_n3901, new_n3933);
and_5  g01585(new_n3933, new_n3900, new_n3934_1);
xor_4  g01586(new_n3934_1, new_n3896, n242);
not_10 g01587(n19477, new_n3936);
not_10 g01588(n11223, new_n3937);
not_10 g01589(n5115, new_n3938);
not_10 g01590(n26572, new_n3939);
nor_5  g01591(n21398, n11667, new_n3940);
and_5  g01592(new_n3940, new_n3939, new_n3941);
and_5  g01593(new_n3941, new_n3938, new_n3942);
and_5  g01594(new_n3942, new_n3937, new_n3943);
xor_4  g01595(new_n3943, new_n3936, new_n3944);
xor_4  g01596(new_n3944, n11011, new_n3945_1);
not_10 g01597(new_n3945_1, new_n3946);
xor_4  g01598(new_n3942, new_n3937, new_n3947);
or_5   g01599(new_n3947, n16029, new_n3948);
xor_4  g01600(new_n3947, n16029, new_n3949);
xor_4  g01601(new_n3941, new_n3938, new_n3950);
nand_5 g01602(new_n3950, n16476, new_n3951);
xor_4  g01603(new_n3950, n16476, new_n3952_1);
xor_4  g01604(new_n3940, new_n3939, new_n3953);
or_5   g01605(new_n3953, n11615, new_n3954);
xor_4  g01606(new_n3953, n11615, new_n3955);
not_10 g01607(new_n3955, new_n3956);
xor_4  g01608(n21398, n11667, new_n3957);
or_5   g01609(new_n3957, n22433, new_n3958);
and_5  g01610(n21398, n14090, new_n3959_1);
not_10 g01611(new_n3959_1, new_n3960);
xor_4  g01612(new_n3957, n22433, new_n3961);
nand_5 g01613(new_n3961, new_n3960, new_n3962_1);
and_5  g01614(new_n3962_1, new_n3958, new_n3963);
or_5   g01615(new_n3963, new_n3956, new_n3964);
and_5  g01616(new_n3964, new_n3954, new_n3965);
nand_5 g01617(new_n3965, new_n3952_1, new_n3966);
and_5  g01618(new_n3966, new_n3951, new_n3967);
nand_5 g01619(new_n3967, new_n3949, new_n3968);
and_5  g01620(new_n3968, new_n3948, new_n3969);
xor_4  g01621(new_n3969, new_n3946, new_n3970);
not_10 g01622(new_n3970, new_n3971_1);
xor_4  g01623(new_n3971_1, n13677, new_n3972);
xor_4  g01624(new_n3967, new_n3949, new_n3973);
not_10 g01625(new_n3973, new_n3974);
or_5   g01626(new_n3974, n18926, new_n3975);
xor_4  g01627(new_n3965, new_n3952_1, new_n3976);
and_5  g01628(new_n3976, n5451, new_n3977);
not_10 g01629(n5451, new_n3978);
xor_4  g01630(new_n3976, new_n3978, new_n3979);
xor_4  g01631(new_n3963, new_n3956, new_n3980);
not_10 g01632(new_n3980, new_n3981);
nand_5 g01633(new_n3981, n5330, new_n3982);
xor_4  g01634(new_n3981, n5330, new_n3983_1);
xor_4  g01635(new_n3961, new_n3960, new_n3984_1);
not_10 g01636(new_n3984_1, new_n3985);
nand_5 g01637(new_n3985, n7657, new_n3986);
and_5  g01638(new_n2554, n25926, new_n3987);
xor_4  g01639(new_n3985, n7657, new_n3988);
nand_5 g01640(new_n3988, new_n3987, new_n3989);
nand_5 g01641(new_n3989, new_n3986, new_n3990);
nand_5 g01642(new_n3990, new_n3983_1, new_n3991);
and_5  g01643(new_n3991, new_n3982, new_n3992);
nor_5  g01644(new_n3992, new_n3979, new_n3993);
nor_5  g01645(new_n3993, new_n3977, new_n3994);
xor_4  g01646(new_n3974, n18926, new_n3995);
nand_5 g01647(new_n3995, new_n3994, new_n3996);
nand_5 g01648(new_n3996, new_n3975, new_n3997);
xor_4  g01649(new_n3997, new_n3972, new_n3998);
not_10 g01650(new_n3998, new_n3999);
not_10 g01651(n12398, new_n4000_1);
not_10 g01652(n19789, new_n4001);
not_10 g01653(n20169, new_n4002);
not_10 g01654(n8285, new_n4003);
nor_5  g01655(n21687, n6729, new_n4004);
and_5  g01656(new_n4004, new_n4003, new_n4005);
and_5  g01657(new_n4005, new_n4002, new_n4006);
and_5  g01658(new_n4006, new_n4001, new_n4007);
xor_4  g01659(new_n4007, new_n4000_1, new_n4008);
not_10 g01660(n20151, new_n4009);
not_10 g01661(n25694, new_n4010_1);
not_10 g01662(n15424, new_n4011);
not_10 g01663(n1949, new_n4012);
not_10 g01664(n9323, new_n4013);
nor_5  g01665(n19922, n10792, new_n4014_1);
and_5  g01666(new_n4014_1, new_n4013, new_n4015);
and_5  g01667(new_n4015, new_n4012, new_n4016);
and_5  g01668(new_n4016, new_n4011, new_n4017);
xor_4  g01669(new_n4017, new_n4010_1, new_n4018);
xor_4  g01670(new_n4018, new_n4009, new_n4019);
xor_4  g01671(new_n4016, new_n4011, new_n4020);
nand_5 g01672(new_n4020, n7693, new_n4021);
xor_4  g01673(new_n4015, new_n4012, new_n4022);
and_5  g01674(new_n4022, n10405, new_n4023);
not_10 g01675(new_n4023, new_n4024);
xor_4  g01676(new_n4022, n10405, new_n4025);
xor_4  g01677(new_n4014_1, new_n4013, new_n4026);
or_5   g01678(new_n4026, n11302, new_n4027);
xor_4  g01679(new_n4026, n11302, new_n4028);
not_10 g01680(new_n4028, new_n4029);
xor_4  g01681(n19922, n10792, new_n4030);
or_5   g01682(new_n4030, n17090, new_n4031);
nand_5 g01683(n19922, n6773, new_n4032);
xor_4  g01684(new_n4030, n17090, new_n4033);
nand_5 g01685(new_n4033, new_n4032, new_n4034);
and_5  g01686(new_n4034, new_n4031, new_n4035);
or_5   g01687(new_n4035, new_n4029, new_n4036);
and_5  g01688(new_n4036, new_n4027, new_n4037);
and_5  g01689(new_n4037, new_n4025, new_n4038);
not_10 g01690(new_n4038, new_n4039);
and_5  g01691(new_n4039, new_n4024, new_n4040);
not_10 g01692(n7693, new_n4041);
xor_4  g01693(new_n4020, new_n4041, new_n4042);
or_5   g01694(new_n4042, new_n4040, new_n4043);
and_5  g01695(new_n4043, new_n4021, new_n4044);
xor_4  g01696(new_n4044, new_n4019, new_n4045);
xnor_4 g01697(new_n4045, new_n4008, new_n4046);
xor_4  g01698(new_n4006, new_n4001, new_n4047);
xor_4  g01699(new_n4020, n7693, new_n4048);
xnor_4 g01700(new_n4048, new_n4040, new_n4049);
nand_5 g01701(new_n4049, new_n4047, new_n4050);
xor_4  g01702(new_n4049, new_n4047, new_n4051);
xor_4  g01703(new_n4037, new_n4025, new_n4052);
xor_4  g01704(new_n4005, new_n4002, new_n4053);
or_5   g01705(new_n4053, new_n4052, new_n4054);
not_10 g01706(new_n4052, new_n4055);
xnor_4 g01707(new_n4053, new_n4055, new_n4056);
xor_4  g01708(new_n4035, new_n4029, new_n4057);
not_10 g01709(new_n4057, new_n4058);
xor_4  g01710(new_n4004, new_n4003, new_n4059);
nand_5 g01711(new_n4059, new_n4058, new_n4060);
xnor_4 g01712(new_n4059, new_n4058, new_n4061);
xnor_4 g01713(n21687, n6729, new_n4062);
xor_4  g01714(new_n4033, new_n4032, new_n4063);
or_5   g01715(new_n4063, new_n4062, new_n4064);
and_5  g01716(new_n2552, n21687, new_n4065);
xor_4  g01717(new_n4063, new_n4062, new_n4066);
nand_5 g01718(new_n4066, new_n4065, new_n4067);
and_5  g01719(new_n4067, new_n4064, new_n4068);
or_5   g01720(new_n4068, new_n4061, new_n4069);
and_5  g01721(new_n4069, new_n4060, new_n4070);
nand_5 g01722(new_n4070, new_n4056, new_n4071_1);
and_5  g01723(new_n4071_1, new_n4054, new_n4072);
nand_5 g01724(new_n4072, new_n4051, new_n4073);
and_5  g01725(new_n4073, new_n4050, new_n4074);
xor_4  g01726(new_n4074, new_n4046, new_n4075);
xor_4  g01727(new_n4075, new_n3999, new_n4076);
xor_4  g01728(new_n4072, new_n4051, new_n4077);
not_10 g01729(new_n4077, new_n4078);
xor_4  g01730(new_n3995, new_n3994, new_n4079);
and_5  g01731(new_n4079, new_n4078, new_n4080);
not_10 g01732(new_n4080, new_n4081);
not_10 g01733(new_n4079, new_n4082);
xnor_4 g01734(new_n4082, new_n4078, new_n4083);
xor_4  g01735(new_n4070, new_n4056, new_n4084);
not_10 g01736(new_n4084, new_n4085_1);
xor_4  g01737(new_n3992, new_n3979, new_n4086);
nor_5  g01738(new_n4086, new_n4085_1, new_n4087);
not_10 g01739(new_n4087, new_n4088_1);
xor_4  g01740(new_n4086, new_n4085_1, new_n4089_1);
xor_4  g01741(new_n3990, new_n3983_1, new_n4090);
xor_4  g01742(new_n4068, new_n4061, new_n4091);
nor_5  g01743(new_n4091, new_n4090, new_n4092);
xor_4  g01744(new_n4091, new_n4090, new_n4093);
not_10 g01745(new_n4093, new_n4094);
xor_4  g01746(new_n4066, new_n4065, new_n4095);
xor_4  g01747(new_n3988, new_n3987, new_n4096);
nor_5  g01748(new_n4096, new_n4095, new_n4097);
and_5  g01749(new_n2555_1, new_n2553_1, new_n4098);
xor_4  g01750(new_n4096, new_n4095, new_n4099);
not_10 g01751(new_n4099, new_n4100_1);
nor_5  g01752(new_n4100_1, new_n4098, new_n4101);
nor_5  g01753(new_n4101, new_n4097, new_n4102);
nor_5  g01754(new_n4102, new_n4094, new_n4103_1);
nor_5  g01755(new_n4103_1, new_n4092, new_n4104);
not_10 g01756(new_n4104, new_n4105);
and_5  g01757(new_n4105, new_n4089_1, new_n4106);
not_10 g01758(new_n4106, new_n4107);
and_5  g01759(new_n4107, new_n4088_1, new_n4108);
not_10 g01760(new_n4108, new_n4109);
and_5  g01761(new_n4109, new_n4083, new_n4110);
not_10 g01762(new_n4110, new_n4111);
and_5  g01763(new_n4111, new_n4081, new_n4112);
xor_4  g01764(new_n4112, new_n4076, n243);
xnor_4 g01765(n24786, n11302, new_n4114);
or_5   g01766(n27120, n17090, new_n4115);
nand_5 g01767(n23065, n6773, new_n4116);
xor_4  g01768(n27120, n17090, new_n4117);
nand_5 g01769(new_n4117, new_n4116, new_n4118);
and_5  g01770(new_n4118, new_n4115, new_n4119_1);
xor_4  g01771(new_n4119_1, new_n4114, new_n4120);
xor_4  g01772(n20036, n1689, new_n4121);
not_10 g01773(n11192, new_n4122);
and_5  g01774(n22274, new_n4122, new_n4123_1);
or_5   g01775(n22274, new_n4122, new_n4124);
not_10 g01776(n9380, new_n4125);
and_5  g01777(n24129, new_n4125, new_n4126);
and_5  g01778(new_n4126, new_n4124, new_n4127);
nor_5  g01779(new_n4127, new_n4123_1, new_n4128);
xor_4  g01780(new_n4128, new_n4121, new_n4129);
xor_4  g01781(new_n4129, new_n4120, new_n4130);
xor_4  g01782(new_n4117, new_n4116, new_n4131);
xnor_4 g01783(n22274, n11192, new_n4132);
xor_4  g01784(new_n4132, new_n4126, new_n4133);
or_5   g01785(new_n4133, new_n4131, new_n4134_1);
xor_4  g01786(n23065, n6773, new_n4135);
not_10 g01787(new_n4135, new_n4136);
xnor_4 g01788(n24129, n9380, new_n4137);
nor_5  g01789(new_n4137, new_n4136, new_n4138);
xor_4  g01790(new_n4133, new_n4131, new_n4139);
nand_5 g01791(new_n4139, new_n4138, new_n4140);
and_5  g01792(new_n4140, new_n4134_1, new_n4141);
xor_4  g01793(new_n4141, new_n4130, new_n4142);
not_10 g01794(new_n4142, new_n4143);
xnor_4 g01795(n5330, n919, new_n4144);
or_5   g01796(n25316, n7657, new_n4145);
nand_5 g01797(n25926, n20385, new_n4146_1);
xor_4  g01798(n25316, n7657, new_n4147);
nand_5 g01799(new_n4147, new_n4146_1, new_n4148);
and_5  g01800(new_n4148, new_n4145, new_n4149);
xor_4  g01801(new_n4149, new_n4144, new_n4150_1);
xor_4  g01802(new_n4150_1, new_n4143, new_n4151_1);
xor_4  g01803(new_n4139, new_n4138, new_n4152_1);
xor_4  g01804(new_n4147, new_n4146_1, new_n4153_1);
nor_5  g01805(new_n4153_1, new_n4152_1, new_n4154);
not_10 g01806(new_n4154, new_n4155);
xor_4  g01807(n25926, n20385, new_n4156);
xnor_4 g01808(new_n4137, new_n4135, new_n4157);
not_10 g01809(new_n4157, new_n4158);
and_5  g01810(new_n4158, new_n4156, new_n4159);
xor_4  g01811(new_n4153_1, new_n4152_1, new_n4160);
and_5  g01812(new_n4160, new_n4159, new_n4161);
not_10 g01813(new_n4161, new_n4162);
and_5  g01814(new_n4162, new_n4155, new_n4163);
xor_4  g01815(new_n4163, new_n4151_1, n248);
not_10 g01816(n19905, new_n4165_1);
not_10 g01817(n17035, new_n4166);
not_10 g01818(n14684, new_n4167);
nor_5  g01819(n24732, n6631, new_n4168);
and_5  g01820(new_n4168, new_n4167, new_n4169);
and_5  g01821(new_n4169, new_n4166, new_n4170);
xor_4  g01822(new_n4170, new_n4165_1, new_n4171);
xor_4  g01823(new_n4171, n6369, new_n4172_1);
xor_4  g01824(new_n4169, new_n4166, new_n4173_1);
nand_5 g01825(new_n4173_1, n25797, new_n4174);
xor_4  g01826(new_n4173_1, n25797, new_n4175);
xor_4  g01827(new_n4168, new_n4167, new_n4176_1);
or_5   g01828(new_n4176_1, n15967, new_n4177);
xor_4  g01829(new_n4176_1, new_n3729, new_n4178);
xor_4  g01830(n24732, n6631, new_n4179);
or_5   g01831(new_n4179, n13319, new_n4180);
and_5  g01832(n25435, n24732, new_n4181);
not_10 g01833(new_n4181, new_n4182);
xor_4  g01834(new_n4179, n13319, new_n4183);
nand_5 g01835(new_n4183, new_n4182, new_n4184);
and_5  g01836(new_n4184, new_n4180, new_n4185);
or_5   g01837(new_n4185, new_n4178, new_n4186_1);
and_5  g01838(new_n4186_1, new_n4177, new_n4187);
nand_5 g01839(new_n4187, new_n4175, new_n4188);
and_5  g01840(new_n4188, new_n4174, new_n4189);
xor_4  g01841(new_n4189, new_n4172_1, new_n4190);
not_10 g01842(new_n4190, new_n4191);
not_10 g01843(n3468, new_n4192);
not_10 g01844(n18558, new_n4193);
nor_5  g01845(n14148, n1152, new_n4194);
and_5  g01846(new_n4194, new_n2856, new_n4195);
and_5  g01847(new_n4195, new_n4193, new_n4196);
xor_4  g01848(new_n4196, new_n4192, new_n4197);
xor_4  g01849(new_n4197, n19514, new_n4198);
not_10 g01850(new_n4198, new_n4199);
xor_4  g01851(new_n4195, new_n4193, new_n4200);
nand_5 g01852(new_n4200, n10053, new_n4201);
xor_4  g01853(new_n4200, n10053, new_n4202);
not_10 g01854(new_n4202, new_n4203);
xor_4  g01855(new_n4194, new_n2856, new_n4204_1);
nand_5 g01856(new_n4204_1, n8399, new_n4205_1);
xor_4  g01857(new_n4204_1, n8399, new_n4206);
not_10 g01858(new_n4206, new_n4207);
xor_4  g01859(n14148, n1152, new_n4208);
nand_5 g01860(new_n4208, n9507, new_n4209);
and_5  g01861(n26979, n1152, new_n4210);
xor_4  g01862(new_n4208, n9507, new_n4211);
nand_5 g01863(new_n4211, new_n4210, new_n4212);
and_5  g01864(new_n4212, new_n4209, new_n4213);
or_5   g01865(new_n4213, new_n4207, new_n4214);
and_5  g01866(new_n4214, new_n4205_1, new_n4215_1);
or_5   g01867(new_n4215_1, new_n4203, new_n4216);
and_5  g01868(new_n4216, new_n4201, new_n4217);
xor_4  g01869(new_n4217, new_n4199, new_n4218);
not_10 g01870(new_n4218, new_n4219);
not_10 g01871(n13668, new_n4220);
not_10 g01872(n21276, new_n4221_1);
not_10 g01873(n26748, new_n4222);
nor_5  g01874(n10057, n8920, new_n4223);
and_5  g01875(new_n4223, new_n4222, new_n4224_1);
and_5  g01876(new_n4224_1, new_n4221_1, new_n4225);
xor_4  g01877(new_n4225, new_n4220, new_n4226);
xor_4  g01878(new_n4226, n626, new_n4227);
not_10 g01879(new_n4227, new_n4228);
xor_4  g01880(new_n4224_1, new_n4221_1, new_n4229);
nand_5 g01881(new_n4229, n1204, new_n4230);
xor_4  g01882(new_n4229, n1204, new_n4231_1);
not_10 g01883(new_n4231_1, new_n4232);
xor_4  g01884(new_n4223, new_n4222, new_n4233);
nand_5 g01885(new_n4233, n19618, new_n4234);
xor_4  g01886(new_n4233, n19618, new_n4235);
xor_4  g01887(n10057, n8920, new_n4236);
or_5   g01888(new_n4236, n22043, new_n4237);
nand_5 g01889(n12121, n8920, new_n4238);
xor_4  g01890(new_n4236, n22043, new_n4239);
nand_5 g01891(new_n4239, new_n4238, new_n4240);
and_5  g01892(new_n4240, new_n4237, new_n4241);
nand_5 g01893(new_n4241, new_n4235, new_n4242);
and_5  g01894(new_n4242, new_n4234, new_n4243);
or_5   g01895(new_n4243, new_n4232, new_n4244);
and_5  g01896(new_n4244, new_n4230, new_n4245);
xor_4  g01897(new_n4245, new_n4228, new_n4246);
not_10 g01898(new_n4246, new_n4247);
xnor_4 g01899(new_n4247, new_n4219, new_n4248);
xor_4  g01900(new_n4215_1, new_n4203, new_n4249);
not_10 g01901(new_n4249, new_n4250);
xor_4  g01902(new_n4243, new_n4232, new_n4251);
not_10 g01903(new_n4251, new_n4252);
or_5   g01904(new_n4252, new_n4250, new_n4253);
xnor_4 g01905(new_n4252, new_n4250, new_n4254);
xor_4  g01906(new_n4241, new_n4235, new_n4255);
not_10 g01907(new_n4255, new_n4256_1);
xor_4  g01908(new_n4211, new_n4210, new_n4257);
not_10 g01909(new_n4257, new_n4258);
xor_4  g01910(new_n4239, new_n4238, new_n4259);
or_5   g01911(new_n4259, new_n4258, new_n4260);
xor_4  g01912(n12121, n8920, new_n4261);
xor_4  g01913(n26979, n1152, new_n4262);
and_5  g01914(new_n4262, new_n4261, new_n4263);
xor_4  g01915(new_n4259, new_n4258, new_n4264);
nand_5 g01916(new_n4264, new_n4263, new_n4265);
and_5  g01917(new_n4265, new_n4260, new_n4266_1);
or_5   g01918(new_n4266_1, new_n4256_1, new_n4267);
xor_4  g01919(new_n4213, new_n4207, new_n4268);
xor_4  g01920(new_n4266_1, new_n4256_1, new_n4269);
nand_5 g01921(new_n4269, new_n4268, new_n4270);
and_5  g01922(new_n4270, new_n4267, new_n4271);
or_5   g01923(new_n4271, new_n4254, new_n4272_1);
and_5  g01924(new_n4272_1, new_n4253, new_n4273);
xor_4  g01925(new_n4273, new_n4248, new_n4274);
xor_4  g01926(new_n4274, new_n4191, new_n4275);
xor_4  g01927(new_n4187, new_n4175, new_n4276);
xor_4  g01928(new_n4271, new_n4254, new_n4277);
and_5  g01929(new_n4277, new_n4276, new_n4278);
not_10 g01930(new_n4276, new_n4279);
xor_4  g01931(new_n4277, new_n4279, new_n4280);
xor_4  g01932(new_n4269, new_n4268, new_n4281);
not_10 g01933(new_n4281, new_n4282);
xor_4  g01934(new_n4185, new_n4178, new_n4283);
or_5   g01935(new_n4283, new_n4282, new_n4284);
xor_4  g01936(new_n4283, new_n4282, new_n4285);
xor_4  g01937(new_n4264, new_n4263, new_n4286);
or_5   g01938(new_n4286, new_n4183, new_n4287);
not_10 g01939(new_n4286, new_n4288);
xor_4  g01940(new_n4183, new_n4182, new_n4289);
nor_5  g01941(new_n4289, new_n4288, new_n4290);
xor_4  g01942(n25435, n24732, new_n4291);
xor_4  g01943(new_n4262, new_n4261, new_n4292);
and_5  g01944(new_n4292, new_n4291, new_n4293);
or_5   g01945(new_n4293, new_n4290, new_n4294);
and_5  g01946(new_n4294, new_n4287, new_n4295);
nand_5 g01947(new_n4295, new_n4285, new_n4296);
and_5  g01948(new_n4296, new_n4284, new_n4297);
nor_5  g01949(new_n4297, new_n4280, new_n4298);
nor_5  g01950(new_n4298, new_n4278, new_n4299);
xnor_4 g01951(new_n4299, new_n4275, n266);
not_10 g01952(n21839, new_n4301);
nor_5  g01953(n22270, new_n4301, new_n4302);
xor_4  g01954(n22270, n21839, new_n4303);
not_10 g01955(n27089, new_n4304);
or_5   g01956(new_n4304, n8806, new_n4305);
xor_4  g01957(n27089, n8806, new_n4306_1);
not_10 g01958(n11841, new_n4307);
or_5   g01959(new_n4307, n2479, new_n4308);
xor_4  g01960(n11841, n2479, new_n4309);
not_10 g01961(n10710, new_n4310);
or_5   g01962(new_n4310, n9372, new_n4311);
xor_4  g01963(n10710, n9372, new_n4312);
not_10 g01964(n20929, new_n4313);
or_5   g01965(new_n4313, n6596, new_n4314);
xor_4  g01966(n20929, n6596, new_n4315);
not_10 g01967(n8006, new_n4316);
or_5   g01968(n15289, new_n4316, new_n4317);
xor_4  g01969(n15289, n8006, new_n4318);
not_10 g01970(n25074, new_n4319_1);
or_5   g01971(new_n4319_1, n6556, new_n4320);
xnor_4 g01972(n25074, n6556, new_n4321);
not_10 g01973(n16396, new_n4322);
and_5  g01974(n22871, new_n4322, new_n4323);
or_5   g01975(n22871, new_n4322, new_n4324);
not_10 g01976(n9399, new_n4325_1);
and_5  g01977(n14275, new_n4325_1, new_n4326_1);
nor_5  g01978(n14275, new_n4325_1, new_n4327);
not_10 g01979(new_n4327, new_n4328);
not_10 g01980(n2088, new_n4329);
and_5  g01981(n25023, new_n4329, new_n4330);
and_5  g01982(new_n4330, new_n4328, new_n4331);
nor_5  g01983(new_n4331, new_n4326_1, new_n4332);
not_10 g01984(new_n4332, new_n4333);
and_5  g01985(new_n4333, new_n4324, new_n4334);
nor_5  g01986(new_n4334, new_n4323, new_n4335);
nand_5 g01987(new_n4335, new_n4321, new_n4336);
and_5  g01988(new_n4336, new_n4320, new_n4337);
or_5   g01989(new_n4337, new_n4318, new_n4338);
and_5  g01990(new_n4338, new_n4317, new_n4339);
or_5   g01991(new_n4339, new_n4315, new_n4340_1);
and_5  g01992(new_n4340_1, new_n4314, new_n4341);
or_5   g01993(new_n4341, new_n4312, new_n4342);
and_5  g01994(new_n4342, new_n4311, new_n4343);
or_5   g01995(new_n4343, new_n4309, new_n4344);
and_5  g01996(new_n4344, new_n4308, new_n4345);
or_5   g01997(new_n4345, new_n4306_1, new_n4346);
and_5  g01998(new_n4346, new_n4305, new_n4347);
nor_5  g01999(new_n4347, new_n4303, new_n4348);
nor_5  g02000(new_n4348, new_n4302, new_n4349);
xor_4  g02001(new_n4347, new_n4303, new_n4350);
or_5   g02002(new_n4350, n23272, new_n4351);
xor_4  g02003(new_n4350, n23272, new_n4352);
not_10 g02004(new_n4352, new_n4353);
xor_4  g02005(new_n4345, new_n4306_1, new_n4354);
or_5   g02006(new_n4354, n11481, new_n4355);
xor_4  g02007(new_n4354, n11481, new_n4356);
not_10 g02008(new_n4356, new_n4357);
xor_4  g02009(new_n4343, new_n4309, new_n4358);
or_5   g02010(new_n4358, n16439, new_n4359);
not_10 g02011(n16439, new_n4360);
xor_4  g02012(new_n4358, new_n4360, new_n4361);
xor_4  g02013(new_n4341, new_n4312, new_n4362);
or_5   g02014(new_n4362, n15241, new_n4363);
not_10 g02015(n15241, new_n4364);
xor_4  g02016(new_n4362, new_n4364, new_n4365);
xor_4  g02017(new_n4339, new_n4315, new_n4366);
or_5   g02018(new_n4366, n7678, new_n4367);
not_10 g02019(n7678, new_n4368);
xor_4  g02020(new_n4366, new_n4368, new_n4369);
xor_4  g02021(new_n4337, new_n4318, new_n4370);
or_5   g02022(new_n4370, n3785, new_n4371);
xor_4  g02023(new_n4370, n3785, new_n4372);
not_10 g02024(new_n4372, new_n4373);
xor_4  g02025(new_n4335, new_n4321, new_n4374_1);
or_5   g02026(new_n4374_1, n20250, new_n4375);
xor_4  g02027(new_n4374_1, n20250, new_n4376_1);
not_10 g02028(n5822, new_n4377);
xnor_4 g02029(n22871, n16396, new_n4378);
xor_4  g02030(new_n4378, new_n4333, new_n4379);
or_5   g02031(new_n4379, new_n4377, new_n4380);
nand_5 g02032(new_n4379, new_n4377, new_n4381);
not_10 g02033(n26443, new_n4382);
xnor_4 g02034(n14275, n9399, new_n4383);
xor_4  g02035(new_n4383, new_n4330, new_n4384);
and_5  g02036(new_n4384, new_n4382, new_n4385);
not_10 g02037(n1681, new_n4386);
xnor_4 g02038(n25023, n2088, new_n4387);
nor_5  g02039(new_n4387, new_n4386, new_n4388);
not_10 g02040(new_n4388, new_n4389);
xor_4  g02041(new_n4384, new_n4382, new_n4390);
and_5  g02042(new_n4390, new_n4389, new_n4391);
nor_5  g02043(new_n4391, new_n4385, new_n4392);
nand_5 g02044(new_n4392, new_n4381, new_n4393);
and_5  g02045(new_n4393, new_n4380, new_n4394);
nand_5 g02046(new_n4394, new_n4376_1, new_n4395);
and_5  g02047(new_n4395, new_n4375, new_n4396);
or_5   g02048(new_n4396, new_n4373, new_n4397);
and_5  g02049(new_n4397, new_n4371, new_n4398);
or_5   g02050(new_n4398, new_n4369, new_n4399);
and_5  g02051(new_n4399, new_n4367, new_n4400);
or_5   g02052(new_n4400, new_n4365, new_n4401_1);
and_5  g02053(new_n4401_1, new_n4363, new_n4402);
or_5   g02054(new_n4402, new_n4361, new_n4403);
and_5  g02055(new_n4403, new_n4359, new_n4404);
or_5   g02056(new_n4404, new_n4357, new_n4405);
and_5  g02057(new_n4405, new_n4355, new_n4406);
or_5   g02058(new_n4406, new_n4353, new_n4407);
and_5  g02059(new_n4407, new_n4351, new_n4408);
and_5  g02060(new_n4408, new_n4349, new_n4409_1);
not_10 g02061(n9396, new_n4410);
not_10 g02062(n1999, new_n4411);
not_10 g02063(n25168, new_n4412);
not_10 g02064(n9318, new_n4413);
and_5  g02065(new_n3943, new_n3936, new_n4414);
and_5  g02066(new_n4414, new_n4413, new_n4415);
and_5  g02067(new_n4415, new_n4412, new_n4416);
and_5  g02068(new_n4416, new_n4411, new_n4417);
and_5  g02069(new_n4417, new_n4410, new_n4418);
xor_4  g02070(new_n4417, new_n4410, new_n4419);
nor_5  g02071(new_n4419, n18880, new_n4420);
xor_4  g02072(new_n4416, new_n4411, new_n4421);
nor_5  g02073(new_n4421, n25475, new_n4422);
xor_4  g02074(new_n4421, n25475, new_n4423);
not_10 g02075(new_n4423, new_n4424_1);
xor_4  g02076(new_n4415, new_n4412, new_n4425);
or_5   g02077(new_n4425, n23849, new_n4426_1);
xor_4  g02078(new_n4425, n23849, new_n4427);
not_10 g02079(new_n4427, new_n4428);
xor_4  g02080(new_n4414, new_n4413, new_n4429);
or_5   g02081(new_n4429, n12446, new_n4430);
nor_5  g02082(new_n3944, n11011, new_n4431);
not_10 g02083(new_n4431, new_n4432_1);
nor_5  g02084(new_n3969, new_n3946, new_n4433);
not_10 g02085(new_n4433, new_n4434);
and_5  g02086(new_n4434, new_n4432_1, new_n4435);
not_10 g02087(n12446, new_n4436);
xor_4  g02088(new_n4429, new_n4436, new_n4437);
or_5   g02089(new_n4437, new_n4435, new_n4438);
and_5  g02090(new_n4438, new_n4430, new_n4439);
or_5   g02091(new_n4439, new_n4428, new_n4440);
and_5  g02092(new_n4440, new_n4426_1, new_n4441_1);
nor_5  g02093(new_n4441_1, new_n4424_1, new_n4442);
nor_5  g02094(new_n4442, new_n4422, new_n4443);
and_5  g02095(new_n4419, n18880, new_n4444);
nor_5  g02096(new_n4444, new_n4443, new_n4445);
nor_5  g02097(new_n4445, new_n4420, new_n4446);
nor_5  g02098(new_n4446, new_n4418, new_n4447);
not_10 g02099(new_n4447, new_n4448);
not_10 g02100(n18105, new_n4449);
not_10 g02101(n24196, new_n4450);
not_10 g02102(n16376, new_n4451_1);
not_10 g02103(n25381, new_n4452);
not_10 g02104(n12587, new_n4453);
not_10 g02105(n268, new_n4454);
not_10 g02106(n24879, new_n4455);
not_10 g02107(n6785, new_n4456);
nor_5  g02108(n24032, n22843, new_n4457);
and_5  g02109(new_n4457, new_n4456, new_n4458);
and_5  g02110(new_n4458, new_n4455, new_n4459);
and_5  g02111(new_n4459, new_n4454, new_n4460);
and_5  g02112(new_n4460, new_n4453, new_n4461);
and_5  g02113(new_n4461, new_n4452, new_n4462);
and_5  g02114(new_n4462, new_n4451_1, new_n4463);
and_5  g02115(new_n4463, new_n4450, new_n4464);
xor_4  g02116(new_n4464, new_n4449, new_n4465);
xor_4  g02117(new_n4419, n18880, new_n4466);
xnor_4 g02118(new_n4466, new_n4443, new_n4467);
not_10 g02119(new_n4467, new_n4468);
nand_5 g02120(new_n4468, new_n4465, new_n4469);
nand_5 g02121(new_n4464, new_n4449, new_n4470);
xor_4  g02122(new_n4468, new_n4465, new_n4471);
xor_4  g02123(new_n4463, new_n4450, new_n4472);
xor_4  g02124(new_n4441_1, new_n4424_1, new_n4473);
not_10 g02125(new_n4473, new_n4474);
or_5   g02126(new_n4474, new_n4472, new_n4475);
xor_4  g02127(new_n4474, new_n4472, new_n4476_1);
not_10 g02128(new_n4476_1, new_n4477);
xor_4  g02129(new_n4462, new_n4451_1, new_n4478_1);
xor_4  g02130(new_n4439, new_n4428, new_n4479);
not_10 g02131(new_n4479, new_n4480);
or_5   g02132(new_n4480, new_n4478_1, new_n4481);
xnor_4 g02133(new_n4479, new_n4478_1, new_n4482);
not_10 g02134(new_n4482, new_n4483);
xor_4  g02135(new_n4461, new_n4452, new_n4484);
not_10 g02136(new_n4484, new_n4485);
xor_4  g02137(new_n4437, new_n4435, new_n4486);
nand_5 g02138(new_n4486, new_n4485, new_n4487);
xor_4  g02139(new_n4486, new_n4485, new_n4488);
not_10 g02140(new_n4488, new_n4489);
xor_4  g02141(new_n4460, new_n4453, new_n4490);
or_5   g02142(new_n4490, new_n3971_1, new_n4491);
xor_4  g02143(new_n4490, new_n3971_1, new_n4492);
xor_4  g02144(new_n4459, new_n4454, new_n4493);
or_5   g02145(new_n4493, new_n3974, new_n4494);
xor_4  g02146(new_n4458, new_n4455, new_n4495);
nor_5  g02147(new_n4495, new_n3976, new_n4496);
xor_4  g02148(new_n4495, new_n3976, new_n4497);
xor_4  g02149(new_n4457, new_n4456, new_n4498);
nand_5 g02150(new_n4498, new_n3981, new_n4499);
xor_4  g02151(new_n4498, new_n3981, new_n4500);
xor_4  g02152(n24032, n22843, new_n4501);
or_5   g02153(new_n4501, new_n3985, new_n4502);
nand_5 g02154(new_n2554, n22843, new_n4503);
xor_4  g02155(new_n4501, new_n3985, new_n4504);
nand_5 g02156(new_n4504, new_n4503, new_n4505);
and_5  g02157(new_n4505, new_n4502, new_n4506);
nand_5 g02158(new_n4506, new_n4500, new_n4507);
and_5  g02159(new_n4507, new_n4499, new_n4508);
and_5  g02160(new_n4508, new_n4497, new_n4509);
or_5   g02161(new_n4509, new_n4496, new_n4510);
xor_4  g02162(new_n4493, new_n3974, new_n4511);
nand_5 g02163(new_n4511, new_n4510, new_n4512);
nand_5 g02164(new_n4512, new_n4494, new_n4513);
nand_5 g02165(new_n4513, new_n4492, new_n4514_1);
and_5  g02166(new_n4514_1, new_n4491, new_n4515);
or_5   g02167(new_n4515, new_n4489, new_n4516);
and_5  g02168(new_n4516, new_n4487, new_n4517);
or_5   g02169(new_n4517, new_n4483, new_n4518);
and_5  g02170(new_n4518, new_n4481, new_n4519);
or_5   g02171(new_n4519, new_n4477, new_n4520);
and_5  g02172(new_n4520, new_n4475, new_n4521);
nand_5 g02173(new_n4521, new_n4471, new_n4522);
and_5  g02174(new_n4522, new_n4470, new_n4523);
and_5  g02175(new_n4523, new_n4469, new_n4524);
and_5  g02176(new_n4524, new_n4448, new_n4525);
xor_4  g02177(new_n4525, new_n4409_1, new_n4526);
xor_4  g02178(new_n4408, new_n4349, new_n4527);
not_10 g02179(new_n4527, new_n4528);
xnor_4 g02180(new_n4524, new_n4447, new_n4529_1);
and_5  g02181(new_n4529_1, new_n4528, new_n4530);
xor_4  g02182(new_n4529_1, new_n4528, new_n4531);
not_10 g02183(new_n4531, new_n4532);
xor_4  g02184(new_n4521, new_n4471, new_n4533);
not_10 g02185(new_n4533, new_n4534);
xor_4  g02186(new_n4406, new_n4353, new_n4535);
and_5  g02187(new_n4535, new_n4534, new_n4536);
not_10 g02188(new_n4536, new_n4537);
not_10 g02189(new_n4535, new_n4538);
xnor_4 g02190(new_n4538, new_n4534, new_n4539);
xor_4  g02191(new_n4519, new_n4477, new_n4540);
not_10 g02192(new_n4540, new_n4541);
xor_4  g02193(new_n4404, new_n4357, new_n4542);
not_10 g02194(new_n4542, new_n4543);
nor_5  g02195(new_n4543, new_n4541, new_n4544);
not_10 g02196(new_n4544, new_n4545);
xor_4  g02197(new_n4543, new_n4541, new_n4546);
xnor_4 g02198(new_n4517, new_n4482, new_n4547);
xor_4  g02199(new_n4402, new_n4361, new_n4548);
and_5  g02200(new_n4548, new_n4547, new_n4549);
xor_4  g02201(new_n4548, new_n4547, new_n4550);
not_10 g02202(new_n4550, new_n4551);
xor_4  g02203(new_n4515, new_n4489, new_n4552_1);
xor_4  g02204(new_n4400, new_n4365, new_n4553);
and_5  g02205(new_n4553, new_n4552_1, new_n4554);
xor_4  g02206(new_n4553, new_n4552_1, new_n4555);
not_10 g02207(new_n4555, new_n4556);
xor_4  g02208(new_n4513, new_n4492, new_n4557);
xor_4  g02209(new_n4398, new_n4369, new_n4558);
and_5  g02210(new_n4558, new_n4557, new_n4559);
xor_4  g02211(new_n4558, new_n4557, new_n4560);
not_10 g02212(new_n4560, new_n4561);
xor_4  g02213(new_n4396, new_n4373, new_n4562);
xor_4  g02214(new_n4511, new_n4510, new_n4563);
and_5  g02215(new_n4563, new_n4562, new_n4564);
xor_4  g02216(new_n4563, new_n4562, new_n4565);
not_10 g02217(new_n4565, new_n4566);
xor_4  g02218(new_n4508, new_n4497, new_n4567);
xor_4  g02219(new_n4394, new_n4376_1, new_n4568);
and_5  g02220(new_n4568, new_n4567, new_n4569);
not_10 g02221(new_n4569, new_n4570);
xor_4  g02222(new_n4568, new_n4567, new_n4571);
xor_4  g02223(new_n4506, new_n4500, new_n4572);
xor_4  g02224(new_n4379, new_n4377, new_n4573);
xor_4  g02225(new_n4573, new_n4392, new_n4574);
and_5  g02226(new_n4574, new_n4572, new_n4575);
xor_4  g02227(new_n4390, new_n4389, new_n4576);
xor_4  g02228(new_n4504, new_n4503, new_n4577);
nand_5 g02229(new_n4577, new_n4576, new_n4578);
xor_4  g02230(new_n2554, n22843, new_n4579);
xor_4  g02231(new_n4387, new_n4386, new_n4580);
nand_5 g02232(new_n4580, new_n4579, new_n4581);
not_10 g02233(new_n4576, new_n4582);
xnor_4 g02234(new_n4577, new_n4582, new_n4583);
nand_5 g02235(new_n4583, new_n4581, new_n4584);
and_5  g02236(new_n4584, new_n4578, new_n4585);
not_10 g02237(new_n4574, new_n4586);
xnor_4 g02238(new_n4586, new_n4572, new_n4587);
and_5  g02239(new_n4587, new_n4585, new_n4588_1);
nor_5  g02240(new_n4588_1, new_n4575, new_n4589);
and_5  g02241(new_n4589, new_n4571, new_n4590_1);
not_10 g02242(new_n4590_1, new_n4591);
and_5  g02243(new_n4591, new_n4570, new_n4592);
nor_5  g02244(new_n4592, new_n4566, new_n4593);
nor_5  g02245(new_n4593, new_n4564, new_n4594);
nor_5  g02246(new_n4594, new_n4561, new_n4595_1);
nor_5  g02247(new_n4595_1, new_n4559, new_n4596);
nor_5  g02248(new_n4596, new_n4556, new_n4597);
nor_5  g02249(new_n4597, new_n4554, new_n4598);
nor_5  g02250(new_n4598, new_n4551, new_n4599);
nor_5  g02251(new_n4599, new_n4549, new_n4600);
not_10 g02252(new_n4600, new_n4601);
and_5  g02253(new_n4601, new_n4546, new_n4602);
not_10 g02254(new_n4602, new_n4603);
and_5  g02255(new_n4603, new_n4545, new_n4604);
not_10 g02256(new_n4604, new_n4605);
and_5  g02257(new_n4605, new_n4539, new_n4606);
not_10 g02258(new_n4606, new_n4607);
and_5  g02259(new_n4607, new_n4537, new_n4608);
nor_5  g02260(new_n4608, new_n4532, new_n4609);
nor_5  g02261(new_n4609, new_n4530, new_n4610);
xor_4  g02262(new_n4610, new_n4526, n298);
xor_4  g02263(n21735, n20604, new_n4612);
not_10 g02264(n16158, new_n4613);
nand_5 g02265(n24085, new_n4613, new_n4614);
xnor_4 g02266(n24085, n16158, new_n4615);
not_10 g02267(new_n4615, new_n4616);
not_10 g02268(n14071, new_n4617);
or_5   g02269(new_n4617, n5752, new_n4618);
xnor_4 g02270(n14071, n5752, new_n4619);
not_10 g02271(n18171, new_n4620);
or_5   g02272(new_n4620, n1738, new_n4621);
nand_5 g02273(new_n4620, n1738, new_n4622);
not_10 g02274(n12152, new_n4623);
and_5  g02275(n25073, new_n4623, new_n4624_1);
nor_5  g02276(n25073, new_n4623, new_n4625);
not_10 g02277(new_n4625, new_n4626);
not_10 g02278(n19107, new_n4627);
and_5  g02279(n22309, new_n4627, new_n4628);
and_5  g02280(new_n4628, new_n4626, new_n4629);
nor_5  g02281(new_n4629, new_n4624_1, new_n4630);
not_10 g02282(new_n4630, new_n4631);
nand_5 g02283(new_n4631, new_n4622, new_n4632);
and_5  g02284(new_n4632, new_n4621, new_n4633);
nand_5 g02285(new_n4633, new_n4619, new_n4634);
and_5  g02286(new_n4634, new_n4618, new_n4635);
or_5   g02287(new_n4635, new_n4616, new_n4636);
and_5  g02288(new_n4636, new_n4614, new_n4637);
xor_4  g02289(new_n4637, new_n4612, new_n4638);
xnor_4 g02290(n4119, n1525, new_n4639);
not_10 g02291(new_n4639, new_n4640);
not_10 g02292(n16988, new_n4641);
or_5   g02293(new_n4641, n14510, new_n4642);
xnor_4 g02294(n16988, n14510, new_n4643);
not_10 g02295(new_n4643, new_n4644);
not_10 g02296(n21779, new_n4645);
or_5   g02297(new_n4645, n13263, new_n4646_1);
xnor_4 g02298(n21779, n13263, new_n4647);
not_10 g02299(n20455, new_n4648);
or_5   g02300(new_n4648, n5376, new_n4649);
not_10 g02301(n5376, new_n4650);
or_5   g02302(n20455, new_n4650, new_n4651);
not_10 g02303(n1639, new_n4652);
nor_5  g02304(n5128, new_n4652, new_n4653);
and_5  g02305(n5128, new_n4652, new_n4654);
not_10 g02306(n16968, new_n4655);
nor_5  g02307(n23120, new_n4655, new_n4656);
not_10 g02308(new_n4656, new_n4657);
nor_5  g02309(new_n4657, new_n4654, new_n4658);
nor_5  g02310(new_n4658, new_n4653, new_n4659);
not_10 g02311(new_n4659, new_n4660);
nand_5 g02312(new_n4660, new_n4651, new_n4661);
and_5  g02313(new_n4661, new_n4649, new_n4662);
nand_5 g02314(new_n4662, new_n4647, new_n4663);
and_5  g02315(new_n4663, new_n4646_1, new_n4664);
or_5   g02316(new_n4664, new_n4644, new_n4665_1);
and_5  g02317(new_n4665_1, new_n4642, new_n4666);
xor_4  g02318(new_n4666, new_n4640, new_n4667);
not_10 g02319(new_n4667, new_n4668);
xor_4  g02320(n12626, n4272, new_n4669);
not_10 g02321(n24319, new_n4670);
or_5   g02322(new_n4670, n6971, new_n4671);
xnor_4 g02323(n24319, n6971, new_n4672);
not_10 g02324(new_n4672, new_n4673);
not_10 g02325(n7460, new_n4674_1);
or_5   g02326(n22068, new_n4674_1, new_n4675);
xnor_4 g02327(n22068, n7460, new_n4676);
not_10 g02328(n9460, new_n4677);
or_5   g02329(new_n4677, n196, new_n4678);
nand_5 g02330(new_n4677, n196, new_n4679);
not_10 g02331(n11749, new_n4680);
and_5  g02332(n14954, new_n4680, new_n4681);
nor_5  g02333(n14954, new_n4680, new_n4682);
not_10 g02334(n13424, new_n4683);
and_5  g02335(n23831, new_n4683, new_n4684);
not_10 g02336(new_n4684, new_n4685);
nor_5  g02337(new_n4685, new_n4682, new_n4686);
nor_5  g02338(new_n4686, new_n4681, new_n4687);
not_10 g02339(new_n4687, new_n4688);
nand_5 g02340(new_n4688, new_n4679, new_n4689);
and_5  g02341(new_n4689, new_n4678, new_n4690);
nand_5 g02342(new_n4690, new_n4676, new_n4691);
and_5  g02343(new_n4691, new_n4675, new_n4692);
or_5   g02344(new_n4692, new_n4673, new_n4693_1);
and_5  g02345(new_n4693_1, new_n4671, new_n4694);
xor_4  g02346(new_n4694, new_n4669, new_n4695);
xor_4  g02347(new_n4695, new_n4668, new_n4696);
xor_4  g02348(new_n4664, new_n4644, new_n4697);
not_10 g02349(new_n4697, new_n4698);
xor_4  g02350(new_n4692, new_n4673, new_n4699);
not_10 g02351(new_n4699, new_n4700);
or_5   g02352(new_n4700, new_n4698, new_n4701);
xor_4  g02353(new_n4700, new_n4698, new_n4702);
xor_4  g02354(new_n4662, new_n4647, new_n4703);
xor_4  g02355(new_n4690, new_n4676, new_n4704);
or_5   g02356(new_n4704, new_n4703, new_n4705);
xor_4  g02357(new_n4704, new_n4703, new_n4706);
not_10 g02358(new_n4706, new_n4707);
xnor_4 g02359(n20455, n5376, new_n4708);
xor_4  g02360(new_n4708, new_n4660, new_n4709);
xnor_4 g02361(n9460, n196, new_n4710);
xor_4  g02362(new_n4710, new_n4688, new_n4711);
nand_5 g02363(new_n4711, new_n4709, new_n4712);
xor_4  g02364(new_n4711, new_n4709, new_n4713);
xnor_4 g02365(n5128, n1639, new_n4714);
xnor_4 g02366(new_n4714, new_n4657, new_n4715);
xnor_4 g02367(n14954, n11749, new_n4716);
xnor_4 g02368(new_n4716, new_n4685, new_n4717);
or_5   g02369(new_n4717, new_n4715, new_n4718);
xnor_4 g02370(n23120, n16968, new_n4719);
xnor_4 g02371(n23831, n13424, new_n4720);
nor_5  g02372(new_n4720, new_n4719, new_n4721);
xor_4  g02373(new_n4717, new_n4715, new_n4722_1);
nand_5 g02374(new_n4722_1, new_n4721, new_n4723);
and_5  g02375(new_n4723, new_n4718, new_n4724);
nand_5 g02376(new_n4724, new_n4713, new_n4725);
and_5  g02377(new_n4725, new_n4712, new_n4726);
or_5   g02378(new_n4726, new_n4707, new_n4727);
and_5  g02379(new_n4727, new_n4705, new_n4728);
nand_5 g02380(new_n4728, new_n4702, new_n4729);
and_5  g02381(new_n4729, new_n4701, new_n4730);
xor_4  g02382(new_n4730, new_n4696, new_n4731_1);
xor_4  g02383(new_n4731_1, new_n4638, new_n4732);
xor_4  g02384(new_n4635, new_n4616, new_n4733);
xor_4  g02385(new_n4728, new_n4702, new_n4734);
or_5   g02386(new_n4734, new_n4733, new_n4735);
xor_4  g02387(new_n4734, new_n4733, new_n4736);
not_10 g02388(new_n4736, new_n4737);
xor_4  g02389(new_n4726, new_n4707, new_n4738);
xnor_4 g02390(new_n4633, new_n4619, new_n4739);
nand_5 g02391(new_n4739, new_n4738, new_n4740);
xor_4  g02392(new_n4724, new_n4713, new_n4741);
xnor_4 g02393(n18171, n1738, new_n4742);
xor_4  g02394(new_n4742, new_n4631, new_n4743);
nand_5 g02395(new_n4743, new_n4741, new_n4744);
not_10 g02396(new_n4741, new_n4745_1);
xnor_4 g02397(new_n4743, new_n4745_1, new_n4746);
xnor_4 g02398(n22309, n19107, new_n4747_1);
xor_4  g02399(new_n4720, new_n4719, new_n4748);
not_10 g02400(new_n4748, new_n4749);
nor_5  g02401(new_n4749, new_n4747_1, new_n4750);
xnor_4 g02402(n25073, n12152, new_n4751);
xnor_4 g02403(new_n4751, new_n4628, new_n4752);
or_5   g02404(new_n4752, new_n4750, new_n4753);
xor_4  g02405(new_n4722_1, new_n4721, new_n4754);
xor_4  g02406(new_n4751, new_n4628, new_n4755);
xnor_4 g02407(new_n4755, new_n4750, new_n4756);
not_10 g02408(new_n4756, new_n4757);
or_5   g02409(new_n4757, new_n4754, new_n4758);
nand_5 g02410(new_n4758, new_n4753, new_n4759);
nand_5 g02411(new_n4759, new_n4746, new_n4760);
and_5  g02412(new_n4760, new_n4744, new_n4761);
xor_4  g02413(new_n4739, new_n4738, new_n4762);
not_10 g02414(new_n4762, new_n4763);
or_5   g02415(new_n4763, new_n4761, new_n4764);
and_5  g02416(new_n4764, new_n4740, new_n4765);
or_5   g02417(new_n4765, new_n4737, new_n4766_1);
and_5  g02418(new_n4766_1, new_n4735, new_n4767);
xor_4  g02419(new_n4767, new_n4732, n317);
nor_5  g02420(n9934, n3506, new_n4769);
not_10 g02421(new_n4769, new_n4770_1);
xor_4  g02422(n9934, n3506, new_n4771);
not_10 g02423(new_n4771, new_n4772);
or_5   g02424(n18496, n14899, new_n4773);
xor_4  g02425(n18496, n14899, new_n4774);
not_10 g02426(new_n4774, new_n4775);
or_5   g02427(n26224, n18444, new_n4776);
xor_4  g02428(n26224, n18444, new_n4777_1);
not_10 g02429(new_n4777_1, new_n4778);
or_5   g02430(n24638, n19327, new_n4779);
xor_4  g02431(n24638, n19327, new_n4780);
not_10 g02432(new_n4780, new_n4781);
or_5   g02433(n22597, n21674, new_n4782);
xor_4  g02434(n22597, n21674, new_n4783);
not_10 g02435(new_n4783, new_n4784);
or_5   g02436(n26107, n17251, new_n4785_1);
xor_4  g02437(n26107, n17251, new_n4786);
not_10 g02438(new_n4786, new_n4787);
or_5   g02439(n14790, n342, new_n4788);
xor_4  g02440(n14790, n342, new_n4789);
not_10 g02441(new_n4789, new_n4790);
or_5   g02442(n26553, n10096, new_n4791);
xnor_4 g02443(n26553, n10096, new_n4792);
or_5   g02444(n16994, n4964, new_n4793);
and_5  g02445(n9246, n7876, new_n4794);
not_10 g02446(new_n4794, new_n4795);
xor_4  g02447(n16994, n4964, new_n4796);
nand_5 g02448(new_n4796, new_n4795, new_n4797);
and_5  g02449(new_n4797, new_n4793, new_n4798);
or_5   g02450(new_n4798, new_n4792, new_n4799);
and_5  g02451(new_n4799, new_n4791, new_n4800);
or_5   g02452(new_n4800, new_n4790, new_n4801);
and_5  g02453(new_n4801, new_n4788, new_n4802);
or_5   g02454(new_n4802, new_n4787, new_n4803);
and_5  g02455(new_n4803, new_n4785_1, new_n4804_1);
or_5   g02456(new_n4804_1, new_n4784, new_n4805);
and_5  g02457(new_n4805, new_n4782, new_n4806);
or_5   g02458(new_n4806, new_n4781, new_n4807);
and_5  g02459(new_n4807, new_n4779, new_n4808);
or_5   g02460(new_n4808, new_n4778, new_n4809);
and_5  g02461(new_n4809, new_n4776, new_n4810_1);
or_5   g02462(new_n4810_1, new_n4775, new_n4811);
and_5  g02463(new_n4811, new_n4773, new_n4812_1);
nor_5  g02464(new_n4812_1, new_n4772, new_n4813);
not_10 g02465(new_n4813, new_n4814_1);
and_5  g02466(new_n4814_1, new_n4770_1, new_n4815);
xor_4  g02467(n9554, n2979, new_n4816);
not_10 g02468(new_n4816, new_n4817);
or_5   g02469(n26408, n647, new_n4818);
xor_4  g02470(n26408, n647, new_n4819);
not_10 g02471(new_n4819, new_n4820);
or_5   g02472(n20409, n18227, new_n4821);
xor_4  g02473(n20409, n18227, new_n4822);
not_10 g02474(new_n4822, new_n4823);
or_5   g02475(n25749, n7377, new_n4824);
xor_4  g02476(n25749, n7377, new_n4825);
not_10 g02477(new_n4825, new_n4826);
or_5   g02478(n11630, n3161, new_n4827);
xnor_4 g02479(n11630, n3161, new_n4828);
or_5   g02480(n13453, n9003, new_n4829);
xnor_4 g02481(n13453, n9003, new_n4830);
or_5   g02482(n7421, n4957, new_n4831);
xor_4  g02483(n7421, n4957, new_n4832);
not_10 g02484(new_n4832, new_n4833);
or_5   g02485(n19680, n7524, new_n4834);
xor_4  g02486(n19680, n7524, new_n4835);
not_10 g02487(new_n4835, new_n4836);
or_5   g02488(n15743, n2809, new_n4837);
and_5  g02489(n20658, n15508, new_n4838);
xnor_4 g02490(n15743, n2809, new_n4839);
or_5   g02491(new_n4839, new_n4838, new_n4840);
and_5  g02492(new_n4840, new_n4837, new_n4841);
or_5   g02493(new_n4841, new_n4836, new_n4842);
and_5  g02494(new_n4842, new_n4834, new_n4843);
or_5   g02495(new_n4843, new_n4833, new_n4844);
and_5  g02496(new_n4844, new_n4831, new_n4845);
or_5   g02497(new_n4845, new_n4830, new_n4846);
and_5  g02498(new_n4846, new_n4829, new_n4847);
or_5   g02499(new_n4847, new_n4828, new_n4848);
and_5  g02500(new_n4848, new_n4827, new_n4849);
or_5   g02501(new_n4849, new_n4826, new_n4850_1);
and_5  g02502(new_n4850_1, new_n4824, new_n4851);
or_5   g02503(new_n4851, new_n4823, new_n4852);
and_5  g02504(new_n4852, new_n4821, new_n4853);
or_5   g02505(new_n4853, new_n4820, new_n4854);
and_5  g02506(new_n4854, new_n4818, new_n4855);
xor_4  g02507(new_n4855, new_n4817, new_n4856);
not_10 g02508(new_n4856, new_n4857);
and_5  g02509(new_n4857, n9259, new_n4858_1);
not_10 g02510(new_n4858_1, new_n4859);
xor_4  g02511(new_n4857, new_n3584, new_n4860);
xor_4  g02512(new_n4853, new_n4820, new_n4861);
not_10 g02513(new_n4861, new_n4862);
nand_5 g02514(new_n4862, n21489, new_n4863);
xor_4  g02515(new_n4862, new_n3585, new_n4864);
xor_4  g02516(new_n4851, new_n4823, new_n4865);
not_10 g02517(new_n4865, new_n4866);
nand_5 g02518(new_n4866, n20213, new_n4867);
xor_4  g02519(new_n4866, new_n3586, new_n4868);
xor_4  g02520(new_n4849, new_n4826, new_n4869);
not_10 g02521(new_n4869, new_n4870);
nand_5 g02522(new_n4870, n13912, new_n4871);
xor_4  g02523(new_n4870, new_n3587, new_n4872);
xor_4  g02524(new_n4847, new_n4828, new_n4873);
or_5   g02525(new_n4873, new_n3588, new_n4874);
xor_4  g02526(new_n4873, n7670, new_n4875);
xor_4  g02527(new_n4845, new_n4830, new_n4876);
or_5   g02528(new_n4876, new_n3589, new_n4877);
xor_4  g02529(new_n4876, n9598, new_n4878);
xor_4  g02530(new_n4843, new_n4833, new_n4879);
not_10 g02531(new_n4879, new_n4880);
nand_5 g02532(new_n4880, n22290, new_n4881);
xor_4  g02533(new_n4880, new_n3590, new_n4882);
xor_4  g02534(new_n4841, new_n4836, new_n4883);
not_10 g02535(new_n4883, new_n4884);
nand_5 g02536(new_n4884, n11273, new_n4885);
xor_4  g02537(n15743, n2809, new_n4886);
xnor_4 g02538(new_n4886, new_n4838, new_n4887);
not_10 g02539(new_n4887, new_n4888);
or_5   g02540(new_n4888, n25565, new_n4889);
xor_4  g02541(n20658, n15508, new_n4890);
and_5  g02542(new_n4890, n21993, new_n4891_1);
not_10 g02543(new_n4891_1, new_n4892);
xor_4  g02544(new_n4888, n25565, new_n4893);
nand_5 g02545(new_n4893, new_n4892, new_n4894);
and_5  g02546(new_n4894, new_n4889, new_n4895);
xor_4  g02547(new_n4884, n11273, new_n4896);
nand_5 g02548(new_n4896, new_n4895, new_n4897);
and_5  g02549(new_n4897, new_n4885, new_n4898);
or_5   g02550(new_n4898, new_n4882, new_n4899);
and_5  g02551(new_n4899, new_n4881, new_n4900);
or_5   g02552(new_n4900, new_n4878, new_n4901);
and_5  g02553(new_n4901, new_n4877, new_n4902);
or_5   g02554(new_n4902, new_n4875, new_n4903);
and_5  g02555(new_n4903, new_n4874, new_n4904);
or_5   g02556(new_n4904, new_n4872, new_n4905);
and_5  g02557(new_n4905, new_n4871, new_n4906);
or_5   g02558(new_n4906, new_n4868, new_n4907);
and_5  g02559(new_n4907, new_n4867, new_n4908);
or_5   g02560(new_n4908, new_n4864, new_n4909);
and_5  g02561(new_n4909, new_n4863, new_n4910);
nor_5  g02562(new_n4910, new_n4860, new_n4911);
not_10 g02563(new_n4911, new_n4912);
and_5  g02564(new_n4912, new_n4859, new_n4913_1);
or_5   g02565(n9554, n2979, new_n4914);
or_5   g02566(new_n4855, new_n4817, new_n4915);
and_5  g02567(new_n4915, new_n4914, new_n4916);
xnor_4 g02568(new_n4916, new_n4913_1, new_n4917);
not_10 g02569(new_n4917, new_n4918);
not_10 g02570(n3740, new_n4919);
xor_4  g02571(new_n4910, new_n4860, new_n4920);
and_5  g02572(new_n4920, new_n4919, new_n4921);
xor_4  g02573(new_n4920, new_n4919, new_n4922);
not_10 g02574(n2858, new_n4923);
xor_4  g02575(new_n4908, new_n4864, new_n4924);
or_5   g02576(new_n4924, new_n4923, new_n4925_1);
xor_4  g02577(new_n4924, n2858, new_n4926);
not_10 g02578(n2659, new_n4927);
xor_4  g02579(new_n4906, new_n4868, new_n4928);
or_5   g02580(new_n4928, new_n4927, new_n4929);
xor_4  g02581(new_n4928, n2659, new_n4930);
not_10 g02582(n24327, new_n4931);
xor_4  g02583(new_n4904, new_n4872, new_n4932);
or_5   g02584(new_n4932, new_n4931, new_n4933);
xor_4  g02585(new_n4932, n24327, new_n4934);
not_10 g02586(n22198, new_n4935);
xor_4  g02587(new_n4902, new_n4875, new_n4936);
or_5   g02588(new_n4936, new_n4935, new_n4937);
xor_4  g02589(new_n4936, n22198, new_n4938);
not_10 g02590(n20826, new_n4939_1);
xor_4  g02591(new_n4900, new_n4878, new_n4940);
or_5   g02592(new_n4940, new_n4939_1, new_n4941);
xor_4  g02593(new_n4940, n20826, new_n4942);
not_10 g02594(n7305, new_n4943);
xor_4  g02595(new_n4898, new_n4882, new_n4944);
or_5   g02596(new_n4944, new_n4943, new_n4945);
not_10 g02597(n25872, new_n4946);
xor_4  g02598(new_n4896, new_n4895, new_n4947_1);
nand_5 g02599(new_n4947_1, new_n4946, new_n4948);
xor_4  g02600(new_n4947_1, new_n4946, new_n4949);
xor_4  g02601(new_n4893, new_n4892, new_n4950);
nand_5 g02602(new_n4950, n20259, new_n4951);
not_10 g02603(n3925, new_n4952_1);
xor_4  g02604(new_n4890, n21993, new_n4953);
nand_5 g02605(new_n4953, new_n4952_1, new_n4954);
xor_4  g02606(new_n4950, n20259, new_n4955);
nand_5 g02607(new_n4955, new_n4954, new_n4956);
and_5  g02608(new_n4956, new_n4951, new_n4957_1);
nand_5 g02609(new_n4957_1, new_n4949, new_n4958);
and_5  g02610(new_n4958, new_n4948, new_n4959);
xor_4  g02611(new_n4944, new_n4943, new_n4960);
nand_5 g02612(new_n4960, new_n4959, new_n4961);
and_5  g02613(new_n4961, new_n4945, new_n4962);
or_5   g02614(new_n4962, new_n4942, new_n4963);
and_5  g02615(new_n4963, new_n4941, new_n4964_1);
or_5   g02616(new_n4964_1, new_n4938, new_n4965);
and_5  g02617(new_n4965, new_n4937, new_n4966_1);
or_5   g02618(new_n4966_1, new_n4934, new_n4967_1);
and_5  g02619(new_n4967_1, new_n4933, new_n4968);
or_5   g02620(new_n4968, new_n4930, new_n4969);
and_5  g02621(new_n4969, new_n4929, new_n4970);
or_5   g02622(new_n4970, new_n4926, new_n4971);
and_5  g02623(new_n4971, new_n4925_1, new_n4972_1);
and_5  g02624(new_n4972_1, new_n4922, new_n4973);
nor_5  g02625(new_n4973, new_n4921, new_n4974);
xor_4  g02626(new_n4974, new_n4918, new_n4975);
xor_4  g02627(new_n4975, new_n4815, new_n4976);
xor_4  g02628(new_n4812_1, new_n4772, new_n4977);
xor_4  g02629(new_n4972_1, new_n4922, new_n4978);
and_5  g02630(new_n4978, new_n4977, new_n4979);
xor_4  g02631(new_n4978, new_n4977, new_n4980);
not_10 g02632(new_n4980, new_n4981);
xor_4  g02633(new_n4810_1, new_n4775, new_n4982);
not_10 g02634(new_n4982, new_n4983);
xor_4  g02635(new_n4970, new_n4926, new_n4984);
nor_5  g02636(new_n4984, new_n4983, new_n4985);
xor_4  g02637(new_n4984, new_n4983, new_n4986);
not_10 g02638(new_n4986, new_n4987);
xor_4  g02639(new_n4808, new_n4778, new_n4988);
not_10 g02640(new_n4988, new_n4989);
xor_4  g02641(new_n4968, new_n4930, new_n4990);
nor_5  g02642(new_n4990, new_n4989, new_n4991);
xor_4  g02643(new_n4990, new_n4989, new_n4992);
not_10 g02644(new_n4992, new_n4993);
xor_4  g02645(new_n4806, new_n4781, new_n4994);
not_10 g02646(new_n4994, new_n4995);
xor_4  g02647(new_n4966_1, new_n4934, new_n4996);
nor_5  g02648(new_n4996, new_n4995, new_n4997);
xor_4  g02649(new_n4996, new_n4995, new_n4998);
not_10 g02650(new_n4998, new_n4999);
xor_4  g02651(new_n4804_1, new_n4784, new_n5000);
not_10 g02652(new_n5000, new_n5001);
xor_4  g02653(new_n4964_1, new_n4938, new_n5002);
nor_5  g02654(new_n5002, new_n5001, new_n5003);
xor_4  g02655(new_n5002, new_n5001, new_n5004);
not_10 g02656(new_n5004, new_n5005);
xor_4  g02657(new_n4802, new_n4787, new_n5006);
not_10 g02658(new_n5006, new_n5007);
xor_4  g02659(new_n4962, new_n4942, new_n5008);
nor_5  g02660(new_n5008, new_n5007, new_n5009);
xor_4  g02661(new_n5008, new_n5007, new_n5010);
not_10 g02662(new_n5010, new_n5011_1);
xor_4  g02663(new_n4800, new_n4790, new_n5012);
not_10 g02664(new_n5012, new_n5013);
xor_4  g02665(new_n4960, new_n4959, new_n5014);
nor_5  g02666(new_n5014, new_n5013, new_n5015);
xor_4  g02667(new_n5014, new_n5013, new_n5016);
not_10 g02668(new_n5016, new_n5017);
xor_4  g02669(new_n4957_1, new_n4949, new_n5018);
xor_4  g02670(new_n4798, new_n4792, new_n5019);
and_5  g02671(new_n5019, new_n5018, new_n5020_1);
not_10 g02672(new_n5020_1, new_n5021);
xor_4  g02673(new_n5019, new_n5018, new_n5022);
xor_4  g02674(new_n4953, n3925, new_n5023);
xor_4  g02675(n9246, n7876, new_n5024_1);
and_5  g02676(new_n5024_1, new_n5023, new_n5025_1);
and_5  g02677(new_n5025_1, new_n4796, new_n5026_1);
xor_4  g02678(new_n4955, new_n4954, new_n5027);
not_10 g02679(new_n5025_1, new_n5028);
xnor_4 g02680(new_n4796, new_n4794, new_n5029);
and_5  g02681(new_n5029, new_n5028, new_n5030);
nor_5  g02682(new_n5030, new_n5026_1, new_n5031_1);
and_5  g02683(new_n5031_1, new_n5027, new_n5032);
nor_5  g02684(new_n5032, new_n5026_1, new_n5033);
and_5  g02685(new_n5033, new_n5022, new_n5034);
not_10 g02686(new_n5034, new_n5035);
and_5  g02687(new_n5035, new_n5021, new_n5036);
nor_5  g02688(new_n5036, new_n5017, new_n5037);
nor_5  g02689(new_n5037, new_n5015, new_n5038);
nor_5  g02690(new_n5038, new_n5011_1, new_n5039);
nor_5  g02691(new_n5039, new_n5009, new_n5040);
nor_5  g02692(new_n5040, new_n5005, new_n5041);
nor_5  g02693(new_n5041, new_n5003, new_n5042);
nor_5  g02694(new_n5042, new_n4999, new_n5043);
nor_5  g02695(new_n5043, new_n4997, new_n5044);
nor_5  g02696(new_n5044, new_n4993, new_n5045);
nor_5  g02697(new_n5045, new_n4991, new_n5046_1);
nor_5  g02698(new_n5046_1, new_n4987, new_n5047);
nor_5  g02699(new_n5047, new_n4985, new_n5048);
nor_5  g02700(new_n5048, new_n4981, new_n5049);
nor_5  g02701(new_n5049, new_n4979, new_n5050);
xor_4  g02702(new_n5050, new_n4976, n332);
xnor_4 g02703(n18295, n16223, new_n5052);
or_5   g02704(n19494, n6502, new_n5053);
nand_5 g02705(n15780, n2387, new_n5054);
xor_4  g02706(n19494, n6502, new_n5055);
nand_5 g02707(new_n5055, new_n5054, new_n5056);
and_5  g02708(new_n5056, new_n5053, new_n5057);
xor_4  g02709(new_n5057, new_n5052, new_n5058);
xor_4  g02710(new_n5058, n8381, new_n5059);
not_10 g02711(new_n5059, new_n5060_1);
not_10 g02712(n20235, new_n5061);
not_10 g02713(n12495, new_n5062_1);
xor_4  g02714(n15780, n2387, new_n5063);
and_5  g02715(new_n5063, new_n5062_1, new_n5064_1);
nand_5 g02716(new_n5064_1, new_n5061, new_n5065);
xor_4  g02717(new_n5064_1, n20235, new_n5066);
xor_4  g02718(new_n5055, new_n5054, new_n5067);
or_5   g02719(new_n5067, new_n5066, new_n5068);
and_5  g02720(new_n5068, new_n5065, new_n5069);
xor_4  g02721(new_n5069, new_n5060_1, new_n5070);
not_10 g02722(new_n5070, new_n5071);
not_10 g02723(n23146, new_n5072);
not_10 g02724(n21654, new_n5073);
and_5  g02725(new_n5073, n16502, new_n5074);
xnor_4 g02726(n25471, n23842, new_n5075);
xor_4  g02727(new_n5075, new_n5074, new_n5076);
nor_5  g02728(new_n5076, new_n5072, new_n5077_1);
not_10 g02729(n17968, new_n5078);
xnor_4 g02730(n21654, n16502, new_n5079);
nor_5  g02731(new_n5079, new_n5078, new_n5080);
not_10 g02732(new_n5080, new_n5081);
xor_4  g02733(new_n5076, n23146, new_n5082_1);
nor_5  g02734(new_n5082_1, new_n5081, new_n5083);
or_5   g02735(new_n5083, new_n5077_1, new_n5084);
not_10 g02736(n11184, new_n5085);
xor_4  g02737(n15053, n3828, new_n5086);
not_10 g02738(n25471, new_n5087);
or_5   g02739(new_n5087, n23842, new_n5088);
nand_5 g02740(new_n5075, new_n5074, new_n5089);
and_5  g02741(new_n5089, new_n5088, new_n5090);
xor_4  g02742(new_n5090, new_n5086, new_n5091);
xor_4  g02743(new_n5091, new_n5085, new_n5092);
xor_4  g02744(new_n5092, new_n5084, new_n5093);
xor_4  g02745(new_n5093, new_n5071, new_n5094);
not_10 g02746(new_n5094, new_n5095);
xor_4  g02747(new_n5082_1, new_n5081, new_n5096);
not_10 g02748(new_n5096, new_n5097);
xor_4  g02749(new_n5067, new_n5066, new_n5098_1);
nand_5 g02750(new_n5098_1, new_n5097, new_n5099);
xor_4  g02751(new_n5063, n12495, new_n5100);
xor_4  g02752(new_n5079, new_n5078, new_n5101_1);
nand_5 g02753(new_n5101_1, new_n5100, new_n5102);
xor_4  g02754(new_n5098_1, new_n5097, new_n5103);
nand_5 g02755(new_n5103, new_n5102, new_n5104);
and_5  g02756(new_n5104, new_n5099, new_n5105);
xnor_4 g02757(new_n5105, new_n5095, n357);
xor_4  g02758(n22309, n9251, new_n5107);
and_5  g02759(n22309, n9251, new_n5108);
xnor_4 g02760(n25073, n20138, new_n5109);
xnor_4 g02761(new_n5109, new_n5108, new_n5110);
nor_5  g02762(new_n5110, new_n5107, new_n5111);
not_10 g02763(new_n5111, new_n5112);
xor_4  g02764(n18171, n6385, new_n5113);
not_10 g02765(new_n5113, new_n5114);
nor_5  g02766(n25073, n20138, new_n5115_1);
nor_5  g02767(new_n5109, new_n5108, new_n5116);
nor_5  g02768(new_n5116, new_n5115_1, new_n5117);
xor_4  g02769(new_n5117, new_n5114, new_n5118);
not_10 g02770(new_n5118, new_n5119);
nor_5  g02771(new_n5119, new_n5112, new_n5120_1);
xor_4  g02772(n5752, n3136, new_n5121);
not_10 g02773(new_n5121, new_n5122);
or_5   g02774(n18171, n6385, new_n5123);
or_5   g02775(new_n5117, new_n5114, new_n5124);
and_5  g02776(new_n5124, new_n5123, new_n5125);
xor_4  g02777(new_n5125, new_n5122, new_n5126);
and_5  g02778(new_n5126, new_n5120_1, new_n5127);
xor_4  g02779(n16158, n9557, new_n5128_1);
not_10 g02780(new_n5128_1, new_n5129);
or_5   g02781(n5752, n3136, new_n5130);
or_5   g02782(new_n5125, new_n5122, new_n5131_1);
and_5  g02783(new_n5131_1, new_n5130, new_n5132);
xor_4  g02784(new_n5132, new_n5129, new_n5133);
and_5  g02785(new_n5133, new_n5127, new_n5134);
xor_4  g02786(n25643, n20604, new_n5135);
not_10 g02787(new_n5135, new_n5136);
or_5   g02788(n16158, n9557, new_n5137);
or_5   g02789(new_n5132, new_n5129, new_n5138);
and_5  g02790(new_n5138, new_n5137, new_n5139);
xor_4  g02791(new_n5139, new_n5136, new_n5140_1);
not_10 g02792(new_n5140_1, new_n5141);
xnor_4 g02793(new_n5141, new_n5134, new_n5142);
xnor_4 g02794(new_n5142, new_n3134, new_n5143);
not_10 g02795(new_n5143, new_n5144);
not_10 g02796(new_n5133, new_n5145);
xnor_4 g02797(new_n5145, new_n5127, new_n5146);
or_5   g02798(new_n5146, new_n3140, new_n5147);
xnor_4 g02799(new_n5146, new_n3138, new_n5148);
not_10 g02800(new_n5148, new_n5149);
not_10 g02801(new_n5126, new_n5150);
xnor_4 g02802(new_n5150, new_n5120_1, new_n5151);
or_5   g02803(new_n5151, new_n3144, new_n5152);
xor_4  g02804(new_n5151, new_n3144, new_n5153);
xor_4  g02805(new_n5119, new_n5112, new_n5154);
nand_5 g02806(new_n5154, new_n3148, new_n5155);
nand_5 g02807(new_n5107, new_n3153, new_n5156);
and_5  g02808(new_n5156, new_n3157, new_n5157);
nor_5  g02809(n22309, n9251, new_n5158_1);
not_10 g02810(new_n5116, new_n5159);
nor_5  g02811(new_n5159, new_n5158_1, new_n5160);
nor_5  g02812(new_n5160, new_n5111, new_n5161);
not_10 g02813(new_n5161, new_n5162);
not_10 g02814(new_n5157, new_n5163);
not_10 g02815(new_n3101, new_n5164);
or_5   g02816(new_n5156, new_n5164, new_n5165);
and_5  g02817(new_n5165, new_n5163, new_n5166);
and_5  g02818(new_n5166, new_n5162, new_n5167);
nor_5  g02819(new_n5167, new_n5157, new_n5168_1);
xor_4  g02820(new_n5154, new_n3148, new_n5169);
nand_5 g02821(new_n5169, new_n5168_1, new_n5170);
and_5  g02822(new_n5170, new_n5155, new_n5171);
nand_5 g02823(new_n5171, new_n5153, new_n5172);
and_5  g02824(new_n5172, new_n5152, new_n5173);
or_5   g02825(new_n5173, new_n5149, new_n5174);
and_5  g02826(new_n5174, new_n5147, new_n5175);
xor_4  g02827(new_n5175, new_n5144, new_n5176);
not_10 g02828(new_n5176, new_n5177);
xor_4  g02829(n5255, n4119, new_n5178);
not_10 g02830(n21649, new_n5179);
or_5   g02831(new_n5179, n14510, new_n5180);
xnor_4 g02832(n21649, n14510, new_n5181);
not_10 g02833(new_n5181, new_n5182);
not_10 g02834(n18274, new_n5183);
or_5   g02835(new_n5183, n13263, new_n5184_1);
xnor_4 g02836(n18274, n13263, new_n5185);
or_5   g02837(new_n4648, n3828, new_n5186);
not_10 g02838(n3828, new_n5187);
or_5   g02839(n20455, new_n5187, new_n5188);
not_10 g02840(n23842, new_n5189);
and_5  g02841(new_n5189, n1639, new_n5190);
and_5  g02842(n23842, new_n4652, new_n5191);
not_10 g02843(new_n5191, new_n5192);
and_5  g02844(new_n5073, n16968, new_n5193);
and_5  g02845(new_n5193, new_n5192, new_n5194);
nor_5  g02846(new_n5194, new_n5190, new_n5195);
not_10 g02847(new_n5195, new_n5196);
nand_5 g02848(new_n5196, new_n5188, new_n5197);
and_5  g02849(new_n5197, new_n5186, new_n5198);
nand_5 g02850(new_n5198, new_n5185, new_n5199);
and_5  g02851(new_n5199, new_n5184_1, new_n5200);
or_5   g02852(new_n5200, new_n5182, new_n5201);
and_5  g02853(new_n5201, new_n5180, new_n5202);
xor_4  g02854(new_n5202, new_n5178, new_n5203);
xor_4  g02855(new_n5203, new_n5177, new_n5204);
xor_4  g02856(new_n5200, new_n5182, new_n5205);
xor_4  g02857(new_n5173, new_n5149, new_n5206);
not_10 g02858(new_n5206, new_n5207);
or_5   g02859(new_n5207, new_n5205, new_n5208);
xor_4  g02860(new_n5207, new_n5205, new_n5209);
xor_4  g02861(new_n5171, new_n5153, new_n5210);
not_10 g02862(new_n5210, new_n5211_1);
xor_4  g02863(new_n5198, new_n5185, new_n5212);
or_5   g02864(new_n5212, new_n5211_1, new_n5213_1);
xor_4  g02865(new_n5212, new_n5211_1, new_n5214);
xor_4  g02866(new_n5169, new_n5168_1, new_n5215);
not_10 g02867(new_n5215, new_n5216);
xnor_4 g02868(n20455, n3828, new_n5217);
xor_4  g02869(new_n5217, new_n5196, new_n5218);
nand_5 g02870(new_n5218, new_n5216, new_n5219);
xor_4  g02871(new_n5218, new_n5216, new_n5220);
not_10 g02872(new_n5220, new_n5221);
xnor_4 g02873(n21654, n16968, new_n5222);
xor_4  g02874(new_n5107, new_n3153, new_n5223);
not_10 g02875(new_n5223, new_n5224);
nor_5  g02876(new_n5224, new_n5222, new_n5225);
xnor_4 g02877(n23842, n1639, new_n5226_1);
xnor_4 g02878(new_n5226_1, new_n5193, new_n5227);
or_5   g02879(new_n5227, new_n5225, new_n5228_1);
xor_4  g02880(new_n5166, new_n5161, new_n5229);
xor_4  g02881(new_n5226_1, new_n5193, new_n5230);
xnor_4 g02882(new_n5230, new_n5225, new_n5231);
not_10 g02883(new_n5231, new_n5232);
or_5   g02884(new_n5232, new_n5229, new_n5233);
and_5  g02885(new_n5233, new_n5228_1, new_n5234);
or_5   g02886(new_n5234, new_n5221, new_n5235);
nand_5 g02887(new_n5235, new_n5219, new_n5236);
nand_5 g02888(new_n5236, new_n5214, new_n5237);
nand_5 g02889(new_n5237, new_n5213_1, new_n5238);
nand_5 g02890(new_n5238, new_n5209, new_n5239);
and_5  g02891(new_n5239, new_n5208, new_n5240);
xor_4  g02892(new_n5240, new_n5204, n422);
not_10 g02893(n337, new_n5242);
not_10 g02894(n3228, new_n5243);
not_10 g02895(n5302, new_n5244);
not_10 g02896(n25738, new_n5245);
not_10 g02897(n21471, new_n5246);
not_10 g02898(n18737, new_n5247);
not_10 g02899(n14603, new_n5248);
nor_5  g02900(n23333, n20794, new_n5249);
and_5  g02901(new_n5249, new_n5248, new_n5250);
and_5  g02902(new_n5250, new_n5247, new_n5251);
and_5  g02903(new_n5251, new_n5246, new_n5252);
and_5  g02904(new_n5252, new_n5245, new_n5253);
and_5  g02905(new_n5253, new_n5244, new_n5254);
and_5  g02906(new_n5254, new_n5243, new_n5255_1);
xor_4  g02907(new_n5255_1, new_n5242, new_n5256_1);
xor_4  g02908(new_n5256_1, n6485, new_n5257);
xor_4  g02909(new_n5254, new_n5243, new_n5258);
or_5   g02910(new_n5258, n26036, new_n5259);
xor_4  g02911(new_n5258, n26036, new_n5260);
not_10 g02912(new_n5260, new_n5261);
xor_4  g02913(new_n5253, new_n5244, new_n5262);
or_5   g02914(new_n5262, n19770, new_n5263);
xor_4  g02915(new_n5262, n19770, new_n5264);
not_10 g02916(new_n5264, new_n5265_1);
xor_4  g02917(new_n5252, new_n5245, new_n5266);
or_5   g02918(new_n5266, n8782, new_n5267);
xor_4  g02919(new_n5266, n8782, new_n5268);
not_10 g02920(new_n5268, new_n5269);
xor_4  g02921(new_n5251, new_n5246, new_n5270);
or_5   g02922(new_n5270, n8678, new_n5271);
xor_4  g02923(new_n5270, n8678, new_n5272);
not_10 g02924(new_n5272, new_n5273_1);
xor_4  g02925(new_n5250, new_n5247, new_n5274_1);
or_5   g02926(new_n5274_1, n1432, new_n5275);
xor_4  g02927(new_n5249, new_n5248, new_n5276);
nor_5  g02928(new_n5276, n21599, new_n5277);
xor_4  g02929(new_n5276, new_n3146, new_n5278);
xor_4  g02930(n23333, n20794, new_n5279);
or_5   g02931(new_n5279, n25336, new_n5280);
nand_5 g02932(n23333, n11424, new_n5281);
xor_4  g02933(new_n5279, n25336, new_n5282);
nand_5 g02934(new_n5282, new_n5281, new_n5283);
and_5  g02935(new_n5283, new_n5280, new_n5284);
nor_5  g02936(new_n5284, new_n5278, new_n5285);
or_5   g02937(new_n5285, new_n5277, new_n5286);
xor_4  g02938(new_n5274_1, n1432, new_n5287);
nand_5 g02939(new_n5287, new_n5286, new_n5288);
and_5  g02940(new_n5288, new_n5275, new_n5289);
or_5   g02941(new_n5289, new_n5273_1, new_n5290);
and_5  g02942(new_n5290, new_n5271, new_n5291);
or_5   g02943(new_n5291, new_n5269, new_n5292);
and_5  g02944(new_n5292, new_n5267, new_n5293);
or_5   g02945(new_n5293, new_n5265_1, new_n5294);
and_5  g02946(new_n5294, new_n5263, new_n5295);
or_5   g02947(new_n5295, new_n5261, new_n5296);
and_5  g02948(new_n5296, new_n5259, new_n5297);
xor_4  g02949(new_n5297, new_n5257, new_n5298);
xor_4  g02950(n22379, n9967, new_n5299);
not_10 g02951(new_n5299, new_n5300_1);
or_5   g02952(n20946, n1662, new_n5301);
xor_4  g02953(n20946, n1662, new_n5302_1);
not_10 g02954(new_n5302_1, new_n5303);
or_5   g02955(n12875, n7751, new_n5304);
xor_4  g02956(n12875, n7751, new_n5305);
not_10 g02957(new_n5305, new_n5306);
or_5   g02958(n26823, n2035, new_n5307);
xor_4  g02959(n26823, n2035, new_n5308);
not_10 g02960(new_n5308, new_n5309);
or_5   g02961(n5213, n4812, new_n5310);
xor_4  g02962(n5213, n4812, new_n5311);
not_10 g02963(new_n5311, new_n5312);
or_5   g02964(n24278, n4665, new_n5313);
xor_4  g02965(n24278, n4665, new_n5314);
not_10 g02966(new_n5314, new_n5315);
or_5   g02967(n24618, n19005, new_n5316);
xor_4  g02968(n24618, n19005, new_n5317);
not_10 g02969(new_n5317, new_n5318);
or_5   g02970(n4326, n3952, new_n5319);
and_5  g02971(n12315, n5438, new_n5320);
xnor_4 g02972(n4326, n3952, new_n5321);
or_5   g02973(new_n5321, new_n5320, new_n5322);
and_5  g02974(new_n5322, new_n5319, new_n5323);
or_5   g02975(new_n5323, new_n5318, new_n5324);
and_5  g02976(new_n5324, new_n5316, new_n5325_1);
or_5   g02977(new_n5325_1, new_n5315, new_n5326);
and_5  g02978(new_n5326, new_n5313, new_n5327);
or_5   g02979(new_n5327, new_n5312, new_n5328);
and_5  g02980(new_n5328, new_n5310, new_n5329);
or_5   g02981(new_n5329, new_n5309, new_n5330_1);
and_5  g02982(new_n5330_1, new_n5307, new_n5331);
or_5   g02983(new_n5331, new_n5306, new_n5332);
and_5  g02984(new_n5332, new_n5304, new_n5333);
or_5   g02985(new_n5333, new_n5303, new_n5334);
and_5  g02986(new_n5334, new_n5301, new_n5335);
xor_4  g02987(new_n5335, new_n5300_1, new_n5336);
not_10 g02988(new_n5336, new_n5337_1);
xnor_4 g02989(n10763, n5696, new_n5338);
or_5   g02990(n13367, n7437, new_n5339);
xor_4  g02991(n13367, n7437, new_n5340);
not_10 g02992(new_n5340, new_n5341);
or_5   g02993(n20700, n932, new_n5342);
xor_4  g02994(n20700, n932, new_n5343);
not_10 g02995(new_n5343, new_n5344);
or_5   g02996(n7099, n6691, new_n5345);
xor_4  g02997(n7099, n6691, new_n5346);
not_10 g02998(new_n5346, new_n5347);
or_5   g02999(n12811, n3260, new_n5348);
xnor_4 g03000(n12811, n3260, new_n5349);
or_5   g03001(n20489, n1118, new_n5350);
xor_4  g03002(n20489, n1118, new_n5351_1);
not_10 g03003(new_n5351_1, new_n5352);
or_5   g03004(n25974, n2355, new_n5353_1);
xor_4  g03005(n25974, n2355, new_n5354);
not_10 g03006(new_n5354, new_n5355);
or_5   g03007(n11121, n1630, new_n5356);
nand_5 g03008(n16217, n1451, new_n5357);
xor_4  g03009(n11121, n1630, new_n5358);
nand_5 g03010(new_n5358, new_n5357, new_n5359);
and_5  g03011(new_n5359, new_n5356, new_n5360);
or_5   g03012(new_n5360, new_n5355, new_n5361);
and_5  g03013(new_n5361, new_n5353_1, new_n5362);
or_5   g03014(new_n5362, new_n5352, new_n5363);
and_5  g03015(new_n5363, new_n5350, new_n5364);
or_5   g03016(new_n5364, new_n5349, new_n5365);
and_5  g03017(new_n5365, new_n5348, new_n5366);
or_5   g03018(new_n5366, new_n5347, new_n5367);
and_5  g03019(new_n5367, new_n5345, new_n5368);
or_5   g03020(new_n5368, new_n5344, new_n5369);
and_5  g03021(new_n5369, new_n5342, new_n5370);
or_5   g03022(new_n5370, new_n5341, new_n5371);
and_5  g03023(new_n5371, new_n5339, new_n5372);
xor_4  g03024(new_n5372, new_n5338, new_n5373);
xnor_4 g03025(new_n5373, new_n5337_1, new_n5374);
xor_4  g03026(new_n5370, new_n5341, new_n5375);
xor_4  g03027(new_n5333, new_n5303, new_n5376_1);
not_10 g03028(new_n5376_1, new_n5377);
or_5   g03029(new_n5377, new_n5375, new_n5378);
xor_4  g03030(new_n5377, new_n5375, new_n5379);
xor_4  g03031(new_n5368, new_n5344, new_n5380);
xor_4  g03032(new_n5331, new_n5306, new_n5381);
not_10 g03033(new_n5381, new_n5382);
nand_5 g03034(new_n5382, new_n5380, new_n5383);
xnor_4 g03035(new_n5382, new_n5380, new_n5384);
xor_4  g03036(new_n5366, new_n5346, new_n5385);
xor_4  g03037(new_n5329, new_n5309, new_n5386_1);
or_5   g03038(new_n5386_1, new_n5385, new_n5387);
xor_4  g03039(new_n5362, new_n5352, new_n5388);
xor_4  g03040(new_n5325_1, new_n5315, new_n5389);
not_10 g03041(new_n5389, new_n5390);
and_5  g03042(new_n5390, new_n5388, new_n5391);
xnor_4 g03043(new_n5390, new_n5388, new_n5392);
xor_4  g03044(new_n5360, new_n5354, new_n5393);
xor_4  g03045(new_n5323, new_n5318, new_n5394);
or_5   g03046(new_n5394, new_n5393, new_n5395);
xor_4  g03047(new_n5321, new_n5320, new_n5396);
not_10 g03048(new_n5396, new_n5397);
xor_4  g03049(new_n5358, new_n5357, new_n5398);
and_5  g03050(new_n5398, new_n5397, new_n5399_1);
xor_4  g03051(n12315, n5438, new_n5400_1);
xnor_4 g03052(n16217, n1451, new_n5401);
and_5  g03053(new_n5401, new_n5400_1, new_n5402);
xor_4  g03054(new_n5398, new_n5397, new_n5403_1);
and_5  g03055(new_n5403_1, new_n5402, new_n5404);
or_5   g03056(new_n5404, new_n5399_1, new_n5405);
not_10 g03057(new_n5394, new_n5406);
xnor_4 g03058(new_n5406, new_n5393, new_n5407);
nand_5 g03059(new_n5407, new_n5405, new_n5408);
and_5  g03060(new_n5408, new_n5395, new_n5409);
nor_5  g03061(new_n5409, new_n5392, new_n5410);
or_5   g03062(new_n5410, new_n5391, new_n5411);
xor_4  g03063(new_n5364, new_n5349, new_n5412);
or_5   g03064(new_n5412, new_n5411, new_n5413);
xor_4  g03065(new_n5412, new_n5411, new_n5414);
xor_4  g03066(new_n5327, new_n5312, new_n5415);
nand_5 g03067(new_n5415, new_n5414, new_n5416);
and_5  g03068(new_n5416, new_n5413, new_n5417);
not_10 g03069(new_n5386_1, new_n5418);
xnor_4 g03070(new_n5418, new_n5385, new_n5419);
nand_5 g03071(new_n5419, new_n5417, new_n5420);
and_5  g03072(new_n5420, new_n5387, new_n5421);
or_5   g03073(new_n5421, new_n5384, new_n5422);
and_5  g03074(new_n5422, new_n5383, new_n5423);
nand_5 g03075(new_n5423, new_n5379, new_n5424);
and_5  g03076(new_n5424, new_n5378, new_n5425);
xor_4  g03077(new_n5425, new_n5374, new_n5426);
xor_4  g03078(new_n5426, new_n5298, new_n5427);
xor_4  g03079(new_n5295, new_n5261, new_n5428);
xor_4  g03080(new_n5423, new_n5379, new_n5429);
not_10 g03081(new_n5429, new_n5430_1);
nand_5 g03082(new_n5430_1, new_n5428, new_n5431);
xor_4  g03083(new_n5430_1, new_n5428, new_n5432);
xor_4  g03084(new_n5293, new_n5265_1, new_n5433);
xor_4  g03085(new_n5421, new_n5384, new_n5434);
nand_5 g03086(new_n5434, new_n5433, new_n5435);
xor_4  g03087(new_n5434, new_n5433, new_n5436);
not_10 g03088(new_n5436, new_n5437);
xor_4  g03089(new_n5291, new_n5269, new_n5438_1);
xor_4  g03090(new_n5419, new_n5417, new_n5439_1);
nand_5 g03091(new_n5439_1, new_n5438_1, new_n5440);
xor_4  g03092(new_n5439_1, new_n5438_1, new_n5441);
not_10 g03093(new_n5441, new_n5442);
xor_4  g03094(new_n5289, new_n5273_1, new_n5443_1);
not_10 g03095(new_n5443_1, new_n5444);
xor_4  g03096(new_n5415, new_n5414, new_n5445);
or_5   g03097(new_n5445, new_n5444, new_n5446);
xor_4  g03098(new_n5445, new_n5444, new_n5447);
not_10 g03099(new_n5447, new_n5448);
xor_4  g03100(new_n5409, new_n5392, new_n5449);
xor_4  g03101(new_n5287, new_n5286, new_n5450);
nand_5 g03102(new_n5450, new_n5449, new_n5451_1);
xor_4  g03103(new_n5450, new_n5449, new_n5452);
xor_4  g03104(new_n5284, new_n5278, new_n5453);
xor_4  g03105(new_n5407, new_n5405, new_n5454);
nor_5  g03106(new_n5454, new_n5453, new_n5455);
xor_4  g03107(new_n5454, new_n5453, new_n5456);
xor_4  g03108(new_n5403_1, new_n5402, new_n5457);
not_10 g03109(new_n5457, new_n5458);
or_5   g03110(new_n5458, new_n5282, new_n5459);
xor_4  g03111(new_n5282, new_n5281, new_n5460);
nor_5  g03112(new_n5460, new_n5457, new_n5461);
xnor_4 g03113(n23333, n11424, new_n5462);
xor_4  g03114(new_n5401, new_n5400_1, new_n5463);
nor_5  g03115(new_n5463, new_n5462, new_n5464);
or_5   g03116(new_n5464, new_n5461, new_n5465);
and_5  g03117(new_n5465, new_n5459, new_n5466);
and_5  g03118(new_n5466, new_n5456, new_n5467);
nor_5  g03119(new_n5467, new_n5455, new_n5468);
nand_5 g03120(new_n5468, new_n5452, new_n5469);
and_5  g03121(new_n5469, new_n5451_1, new_n5470);
or_5   g03122(new_n5470, new_n5448, new_n5471);
and_5  g03123(new_n5471, new_n5446, new_n5472_1);
or_5   g03124(new_n5472_1, new_n5442, new_n5473);
and_5  g03125(new_n5473, new_n5440, new_n5474);
or_5   g03126(new_n5474, new_n5437, new_n5475);
nand_5 g03127(new_n5475, new_n5435, new_n5476);
nand_5 g03128(new_n5476, new_n5432, new_n5477);
and_5  g03129(new_n5477, new_n5431, new_n5478);
xor_4  g03130(new_n5478, new_n5427, n431);
not_10 g03131(n8614, new_n5480);
and_5  g03132(n23895, new_n5480, new_n5481);
xnor_4 g03133(n23895, n8614, new_n5482);
not_10 g03134(new_n5482, new_n5483);
not_10 g03135(n17351, new_n5484);
or_5   g03136(new_n5484, n15182, new_n5485_1);
xnor_4 g03137(n17351, n15182, new_n5486);
not_10 g03138(new_n5486, new_n5487);
not_10 g03139(n11736, new_n5488);
or_5   g03140(n27037, new_n5488, new_n5489);
xnor_4 g03141(n27037, n11736, new_n5490);
not_10 g03142(new_n5490, new_n5491);
not_10 g03143(n23200, new_n5492);
or_5   g03144(new_n5492, n8964, new_n5493);
xnor_4 g03145(n23200, n8964, new_n5494);
not_10 g03146(new_n5494, new_n5495);
not_10 g03147(n17959, new_n5496);
or_5   g03148(n20151, new_n5496, new_n5497);
xnor_4 g03149(n20151, n17959, new_n5498);
not_10 g03150(new_n5498, new_n5499);
not_10 g03151(n7566, new_n5500);
or_5   g03152(n7693, new_n5500, new_n5501);
xnor_4 g03153(n7693, n7566, new_n5502);
not_10 g03154(new_n5502, new_n5503);
not_10 g03155(n7731, new_n5504);
or_5   g03156(n10405, new_n5504, new_n5505);
xnor_4 g03157(n10405, n7731, new_n5506);
not_10 g03158(n11302, new_n5507);
or_5   g03159(n12341, new_n5507, new_n5508);
not_10 g03160(n12341, new_n5509);
or_5   g03161(new_n5509, n11302, new_n5510);
not_10 g03162(n20986, new_n5511);
and_5  g03163(new_n5511, n17090, new_n5512);
not_10 g03164(n17090, new_n5513);
and_5  g03165(n20986, new_n5513, new_n5514);
not_10 g03166(new_n5514, new_n5515);
not_10 g03167(n12384, new_n5516);
and_5  g03168(new_n5516, n6773, new_n5517_1);
and_5  g03169(new_n5517_1, new_n5515, new_n5518);
nor_5  g03170(new_n5518, new_n5512, new_n5519);
not_10 g03171(new_n5519, new_n5520);
nand_5 g03172(new_n5520, new_n5510, new_n5521_1);
and_5  g03173(new_n5521_1, new_n5508, new_n5522);
nand_5 g03174(new_n5522, new_n5506, new_n5523);
and_5  g03175(new_n5523, new_n5505, new_n5524_1);
or_5   g03176(new_n5524_1, new_n5503, new_n5525);
and_5  g03177(new_n5525, new_n5501, new_n5526);
or_5   g03178(new_n5526, new_n5499, new_n5527);
and_5  g03179(new_n5527, new_n5497, new_n5528);
or_5   g03180(new_n5528, new_n5495, new_n5529);
and_5  g03181(new_n5529, new_n5493, new_n5530);
or_5   g03182(new_n5530, new_n5491, new_n5531);
and_5  g03183(new_n5531, new_n5489, new_n5532_1);
or_5   g03184(new_n5532_1, new_n5487, new_n5533);
and_5  g03185(new_n5533, new_n5485_1, new_n5534);
nor_5  g03186(new_n5534, new_n5483, new_n5535);
nor_5  g03187(new_n5535, new_n5481, new_n5536);
not_10 g03188(n18880, new_n5537);
and_5  g03189(new_n5537, n13494, new_n5538);
not_10 g03190(new_n5538, new_n5539);
xor_4  g03191(n18880, n13494, new_n5540);
not_10 g03192(n25345, new_n5541);
or_5   g03193(n25475, new_n5541, new_n5542);
xnor_4 g03194(n25475, n25345, new_n5543);
not_10 g03195(new_n5543, new_n5544);
not_10 g03196(n9655, new_n5545);
or_5   g03197(n23849, new_n5545, new_n5546);
xnor_4 g03198(n23849, n9655, new_n5547);
not_10 g03199(new_n5547, new_n5548);
not_10 g03200(n13490, new_n5549);
or_5   g03201(new_n5549, n12446, new_n5550);
xnor_4 g03202(n13490, n12446, new_n5551);
not_10 g03203(new_n5551, new_n5552);
not_10 g03204(n22660, new_n5553);
or_5   g03205(new_n5553, n11011, new_n5554);
xnor_4 g03206(n22660, n11011, new_n5555);
not_10 g03207(new_n5555, new_n5556);
not_10 g03208(n1777, new_n5557);
or_5   g03209(n16029, new_n5557, new_n5558);
xnor_4 g03210(n16029, n1777, new_n5559);
not_10 g03211(new_n5559, new_n5560);
not_10 g03212(n8745, new_n5561);
or_5   g03213(n16476, new_n5561, new_n5562);
xnor_4 g03214(n16476, n8745, new_n5563);
not_10 g03215(n11615, new_n5564_1);
or_5   g03216(n15636, new_n5564_1, new_n5565);
and_5  g03217(n15636, new_n5564_1, new_n5566);
not_10 g03218(n20077, new_n5567);
and_5  g03219(n22433, new_n5567, new_n5568);
or_5   g03220(n22433, new_n5567, new_n5569);
not_10 g03221(n6794, new_n5570);
and_5  g03222(n14090, new_n5570, new_n5571);
and_5  g03223(new_n5571, new_n5569, new_n5572);
nor_5  g03224(new_n5572, new_n5568, new_n5573);
or_5   g03225(new_n5573, new_n5566, new_n5574);
and_5  g03226(new_n5574, new_n5565, new_n5575);
nand_5 g03227(new_n5575, new_n5563, new_n5576);
and_5  g03228(new_n5576, new_n5562, new_n5577);
or_5   g03229(new_n5577, new_n5560, new_n5578);
and_5  g03230(new_n5578, new_n5558, new_n5579_1);
or_5   g03231(new_n5579_1, new_n5556, new_n5580);
and_5  g03232(new_n5580, new_n5554, new_n5581);
or_5   g03233(new_n5581, new_n5552, new_n5582);
and_5  g03234(new_n5582, new_n5550, new_n5583);
or_5   g03235(new_n5583, new_n5548, new_n5584);
and_5  g03236(new_n5584, new_n5546, new_n5585);
or_5   g03237(new_n5585, new_n5544, new_n5586);
and_5  g03238(new_n5586, new_n5542, new_n5587);
nor_5  g03239(new_n5587, new_n5540, new_n5588);
not_10 g03240(new_n5588, new_n5589);
and_5  g03241(new_n5589, new_n5539, new_n5590);
xor_4  g03242(new_n5587, new_n5540, new_n5591);
not_10 g03243(n26797, new_n5592);
not_10 g03244(n23913, new_n5593_1);
not_10 g03245(n22554, new_n5594);
not_10 g03246(n20429, new_n5595);
not_10 g03247(n3909, new_n5596);
not_10 g03248(n23974, new_n5597);
not_10 g03249(n2146, new_n5598);
nor_5  g03250(n22173, n583, new_n5599);
and_5  g03251(new_n5599, new_n5598, new_n5600);
and_5  g03252(new_n5600, new_n5597, new_n5601);
and_5  g03253(new_n5601, new_n5596, new_n5602);
and_5  g03254(new_n5602, new_n5595, new_n5603_1);
and_5  g03255(new_n5603_1, new_n5594, new_n5604);
and_5  g03256(new_n5604, new_n5593_1, new_n5605_1);
xor_4  g03257(new_n5605_1, new_n5592, new_n5606);
nor_5  g03258(new_n5606, n10201, new_n5607);
not_10 g03259(n10201, new_n5608);
xor_4  g03260(new_n5606, new_n5608, new_n5609_1);
xor_4  g03261(new_n5604, new_n5593_1, new_n5610);
or_5   g03262(new_n5610, n10593, new_n5611);
not_10 g03263(n10593, new_n5612);
xor_4  g03264(new_n5610, new_n5612, new_n5613);
xor_4  g03265(new_n5603_1, new_n5594, new_n5614);
or_5   g03266(new_n5614, n18290, new_n5615);
not_10 g03267(n18290, new_n5616);
xor_4  g03268(new_n5614, new_n5616, new_n5617);
xor_4  g03269(new_n5602, new_n5595, new_n5618);
or_5   g03270(new_n5618, n11580, new_n5619);
not_10 g03271(n11580, new_n5620);
xor_4  g03272(new_n5618, new_n5620, new_n5621);
xor_4  g03273(new_n5601, new_n5596, new_n5622);
or_5   g03274(new_n5622, n15884, new_n5623);
not_10 g03275(n15884, new_n5624);
xor_4  g03276(new_n5622, new_n5624, new_n5625);
xor_4  g03277(new_n5600, new_n5597, new_n5626);
or_5   g03278(new_n5626, n6356, new_n5627);
xor_4  g03279(new_n5599, new_n5598, new_n5628);
nor_5  g03280(new_n5628, n27104, new_n5629);
xor_4  g03281(new_n5628, n27104, new_n5630);
not_10 g03282(new_n5630, new_n5631);
xor_4  g03283(n22173, n583, new_n5632);
or_5   g03284(new_n5632, n27188, new_n5633);
nand_5 g03285(n6611, n583, new_n5634_1);
xor_4  g03286(new_n5632, n27188, new_n5635);
nand_5 g03287(new_n5635, new_n5634_1, new_n5636);
and_5  g03288(new_n5636, new_n5633, new_n5637);
nor_5  g03289(new_n5637, new_n5631, new_n5638);
or_5   g03290(new_n5638, new_n5629, new_n5639);
xor_4  g03291(new_n5626, n6356, new_n5640);
nand_5 g03292(new_n5640, new_n5639, new_n5641);
and_5  g03293(new_n5641, new_n5627, new_n5642);
or_5   g03294(new_n5642, new_n5625, new_n5643_1);
and_5  g03295(new_n5643_1, new_n5623, new_n5644);
or_5   g03296(new_n5644, new_n5621, new_n5645);
and_5  g03297(new_n5645, new_n5619, new_n5646);
or_5   g03298(new_n5646, new_n5617, new_n5647);
and_5  g03299(new_n5647, new_n5615, new_n5648);
or_5   g03300(new_n5648, new_n5613, new_n5649);
and_5  g03301(new_n5649, new_n5611, new_n5650);
nor_5  g03302(new_n5650, new_n5609_1, new_n5651);
nor_5  g03303(new_n5651, new_n5607, new_n5652);
not_10 g03304(n12702, new_n5653);
and_5  g03305(new_n5605_1, new_n5592, new_n5654);
xor_4  g03306(new_n5654, new_n5653, new_n5655);
xor_4  g03307(new_n5655, n12650, new_n5656);
xor_4  g03308(new_n5656, new_n5652, new_n5657);
nor_5  g03309(new_n5657, new_n5591, new_n5658);
xor_4  g03310(new_n5657, new_n5591, new_n5659);
not_10 g03311(new_n5659, new_n5660);
xor_4  g03312(new_n5585, new_n5544, new_n5661);
not_10 g03313(new_n5661, new_n5662);
xor_4  g03314(new_n5650, new_n5609_1, new_n5663);
nand_5 g03315(new_n5663, new_n5662, new_n5664);
xnor_4 g03316(new_n5663, new_n5661, new_n5665);
not_10 g03317(new_n5665, new_n5666);
xor_4  g03318(new_n5583, new_n5548, new_n5667);
not_10 g03319(new_n5667, new_n5668);
xor_4  g03320(new_n5648, new_n5613, new_n5669);
nand_5 g03321(new_n5669, new_n5668, new_n5670);
xor_4  g03322(new_n5669, new_n5667, new_n5671);
xor_4  g03323(new_n5581, new_n5552, new_n5672);
not_10 g03324(new_n5672, new_n5673);
xor_4  g03325(new_n5646, new_n5617, new_n5674);
nand_5 g03326(new_n5674, new_n5673, new_n5675);
xor_4  g03327(new_n5674, new_n5672, new_n5676);
xor_4  g03328(new_n5579_1, new_n5556, new_n5677);
not_10 g03329(new_n5677, new_n5678);
xor_4  g03330(new_n5644, new_n5621, new_n5679);
nand_5 g03331(new_n5679, new_n5678, new_n5680_1);
xnor_4 g03332(new_n5679, new_n5677, new_n5681);
not_10 g03333(new_n5681, new_n5682);
xor_4  g03334(new_n5577, new_n5560, new_n5683);
not_10 g03335(new_n5683, new_n5684);
xor_4  g03336(new_n5642, new_n5625, new_n5685);
nand_5 g03337(new_n5685, new_n5684, new_n5686);
xor_4  g03338(new_n5685, new_n5683, new_n5687_1);
xor_4  g03339(new_n5575, new_n5563, new_n5688);
not_10 g03340(new_n5688, new_n5689);
xor_4  g03341(new_n5640, new_n5639, new_n5690);
nand_5 g03342(new_n5690, new_n5689, new_n5691);
xnor_4 g03343(new_n5690, new_n5688, new_n5692);
xor_4  g03344(new_n5637, new_n5631, new_n5693);
not_10 g03345(new_n5693, new_n5694);
xnor_4 g03346(n15636, n11615, new_n5695);
xnor_4 g03347(new_n5695, new_n5573, new_n5696_1);
not_10 g03348(new_n5696_1, new_n5697);
nand_5 g03349(new_n5697, new_n5694, new_n5698);
xor_4  g03350(new_n5697, new_n5694, new_n5699);
xor_4  g03351(new_n5635, new_n5634_1, new_n5700_1);
xnor_4 g03352(n22433, n20077, new_n5701);
xor_4  g03353(new_n5701, new_n5571, new_n5702);
or_5   g03354(new_n5702, new_n5700_1, new_n5703);
xnor_4 g03355(n14090, n6794, new_n5704_1);
not_10 g03356(new_n5704_1, new_n5705);
xor_4  g03357(n6611, n583, new_n5706);
and_5  g03358(new_n5706, new_n5705, new_n5707);
xor_4  g03359(new_n5702, new_n5700_1, new_n5708);
nand_5 g03360(new_n5708, new_n5707, new_n5709);
nand_5 g03361(new_n5709, new_n5703, new_n5710);
nand_5 g03362(new_n5710, new_n5699, new_n5711);
and_5  g03363(new_n5711, new_n5698, new_n5712);
nand_5 g03364(new_n5712, new_n5692, new_n5713);
and_5  g03365(new_n5713, new_n5691, new_n5714);
or_5   g03366(new_n5714, new_n5687_1, new_n5715);
and_5  g03367(new_n5715, new_n5686, new_n5716);
or_5   g03368(new_n5716, new_n5682, new_n5717);
and_5  g03369(new_n5717, new_n5680_1, new_n5718);
or_5   g03370(new_n5718, new_n5676, new_n5719);
and_5  g03371(new_n5719, new_n5675, new_n5720);
or_5   g03372(new_n5720, new_n5671, new_n5721);
and_5  g03373(new_n5721, new_n5670, new_n5722);
or_5   g03374(new_n5722, new_n5666, new_n5723);
and_5  g03375(new_n5723, new_n5664, new_n5724);
nor_5  g03376(new_n5724, new_n5660, new_n5725);
or_5   g03377(new_n5725, new_n5658, new_n5726);
nand_5 g03378(new_n5654, new_n5653, new_n5727);
nand_5 g03379(new_n5655, n12650, new_n5728);
or_5   g03380(new_n5655, n12650, new_n5729);
nand_5 g03381(new_n5729, new_n5652, new_n5730);
and_5  g03382(new_n5730, new_n5728, new_n5731);
and_5  g03383(new_n5731, new_n5727, new_n5732_1);
nor_5  g03384(new_n5732_1, new_n5726, new_n5733);
and_5  g03385(new_n5733, new_n5590, new_n5734);
not_10 g03386(new_n5734, new_n5735);
not_10 g03387(new_n5590, new_n5736);
and_5  g03388(new_n5732_1, new_n5726, new_n5737);
and_5  g03389(new_n5737, new_n5736, new_n5738);
not_10 g03390(new_n5738, new_n5739);
and_5  g03391(new_n5739, new_n5735, new_n5740);
xor_4  g03392(new_n5740, new_n5536, new_n5741);
xor_4  g03393(new_n5732_1, new_n5726, new_n5742_1);
xnor_4 g03394(new_n5742_1, new_n5590, new_n5743);
and_5  g03395(new_n5743, new_n5536, new_n5744);
nor_5  g03396(new_n5743, new_n5536, new_n5745);
not_10 g03397(new_n5745, new_n5746);
xor_4  g03398(new_n5534, new_n5483, new_n5747);
not_10 g03399(new_n5747, new_n5748);
xor_4  g03400(new_n5724, new_n5660, new_n5749);
and_5  g03401(new_n5749, new_n5748, new_n5750);
xor_4  g03402(new_n5749, new_n5748, new_n5751);
not_10 g03403(new_n5751, new_n5752_1);
xor_4  g03404(new_n5532_1, new_n5487, new_n5753);
not_10 g03405(new_n5753, new_n5754);
xor_4  g03406(new_n5722, new_n5666, new_n5755);
and_5  g03407(new_n5755, new_n5754, new_n5756);
xor_4  g03408(new_n5755, new_n5754, new_n5757);
not_10 g03409(new_n5757, new_n5758);
xor_4  g03410(new_n5530, new_n5491, new_n5759);
not_10 g03411(new_n5759, new_n5760);
xor_4  g03412(new_n5720, new_n5671, new_n5761);
and_5  g03413(new_n5761, new_n5760, new_n5762);
xor_4  g03414(new_n5761, new_n5760, new_n5763);
not_10 g03415(new_n5763, new_n5764);
xor_4  g03416(new_n5528, new_n5495, new_n5765_1);
not_10 g03417(new_n5765_1, new_n5766);
xor_4  g03418(new_n5718, new_n5676, new_n5767);
and_5  g03419(new_n5767, new_n5766, new_n5768);
xor_4  g03420(new_n5767, new_n5766, new_n5769);
not_10 g03421(new_n5769, new_n5770);
xor_4  g03422(new_n5526, new_n5499, new_n5771);
not_10 g03423(new_n5771, new_n5772);
xor_4  g03424(new_n5716, new_n5682, new_n5773);
and_5  g03425(new_n5773, new_n5772, new_n5774);
xor_4  g03426(new_n5773, new_n5772, new_n5775);
not_10 g03427(new_n5775, new_n5776_1);
xor_4  g03428(new_n5524_1, new_n5503, new_n5777);
not_10 g03429(new_n5777, new_n5778);
xor_4  g03430(new_n5714, new_n5687_1, new_n5779);
and_5  g03431(new_n5779, new_n5778, new_n5780);
xor_4  g03432(new_n5779, new_n5778, new_n5781);
not_10 g03433(new_n5781, new_n5782_1);
xor_4  g03434(new_n5712, new_n5692, new_n5783);
not_10 g03435(new_n5783, new_n5784);
xor_4  g03436(new_n5522, new_n5506, new_n5785);
nor_5  g03437(new_n5785, new_n5784, new_n5786);
xor_4  g03438(new_n5785, new_n5784, new_n5787);
xor_4  g03439(new_n5710, new_n5699, new_n5788);
not_10 g03440(new_n5788, new_n5789);
xnor_4 g03441(n12341, n11302, new_n5790);
xor_4  g03442(new_n5790, new_n5520, new_n5791);
and_5  g03443(new_n5791, new_n5789, new_n5792);
not_10 g03444(new_n5792, new_n5793);
xor_4  g03445(new_n5791, new_n5789, new_n5794);
xor_4  g03446(new_n5706, new_n5704_1, new_n5795);
xnor_4 g03447(n12384, n6773, new_n5796);
nor_5  g03448(new_n5796, new_n5795, new_n5797);
not_10 g03449(new_n5797, new_n5798);
xnor_4 g03450(n20986, n17090, new_n5799);
xor_4  g03451(new_n5799, new_n5517_1, new_n5800);
and_5  g03452(new_n5800, new_n5798, new_n5801);
xor_4  g03453(new_n5708, new_n5707, new_n5802);
not_10 g03454(new_n5802, new_n5803);
xor_4  g03455(new_n5800, new_n5798, new_n5804);
and_5  g03456(new_n5804, new_n5803, new_n5805);
nor_5  g03457(new_n5805, new_n5801, new_n5806);
not_10 g03458(new_n5806, new_n5807);
and_5  g03459(new_n5807, new_n5794, new_n5808);
not_10 g03460(new_n5808, new_n5809);
and_5  g03461(new_n5809, new_n5793, new_n5810);
not_10 g03462(new_n5810, new_n5811);
and_5  g03463(new_n5811, new_n5787, new_n5812);
nor_5  g03464(new_n5812, new_n5786, new_n5813);
nor_5  g03465(new_n5813, new_n5782_1, new_n5814);
nor_5  g03466(new_n5814, new_n5780, new_n5815);
nor_5  g03467(new_n5815, new_n5776_1, new_n5816);
nor_5  g03468(new_n5816, new_n5774, new_n5817);
nor_5  g03469(new_n5817, new_n5770, new_n5818);
nor_5  g03470(new_n5818, new_n5768, new_n5819);
nor_5  g03471(new_n5819, new_n5764, new_n5820);
nor_5  g03472(new_n5820, new_n5762, new_n5821);
nor_5  g03473(new_n5821, new_n5758, new_n5822_1);
nor_5  g03474(new_n5822_1, new_n5756, new_n5823);
nor_5  g03475(new_n5823, new_n5752_1, new_n5824);
nor_5  g03476(new_n5824, new_n5750, new_n5825);
and_5  g03477(new_n5825, new_n5746, new_n5826);
nor_5  g03478(new_n5826, new_n5744, new_n5827);
xor_4  g03479(new_n5827, new_n5741, n457);
xnor_4 g03480(n24323, n1681, new_n5829);
xor_4  g03481(n13781, n2088, new_n5830);
xnor_4 g03482(new_n5830, new_n5829, new_n5831);
and_5  g03483(new_n5831, new_n5705, new_n5832);
xnor_4 g03484(new_n5832, new_n5702, new_n5833_1);
not_10 g03485(new_n5829, new_n5834_1);
and_5  g03486(new_n5830, new_n5834_1, new_n5835);
nor_5  g03487(n24323, new_n4386, new_n5836);
xnor_4 g03488(n26443, n25877, new_n5837);
xor_4  g03489(new_n5837, new_n5836, new_n5838);
not_10 g03490(new_n5838, new_n5839);
xor_4  g03491(new_n5839, new_n5835, new_n5840_1);
xor_4  g03492(n9399, n2088, new_n5841_1);
and_5  g03493(n13781, n2088, new_n5842_1);
or_5   g03494(new_n5842_1, n11486, new_n5843);
nand_5 g03495(n13781, n11486, new_n5844);
or_5   g03496(new_n5844, new_n4329, new_n5845);
and_5  g03497(new_n5845, new_n5843, new_n5846);
xnor_4 g03498(new_n5846, new_n5841_1, new_n5847);
xnor_4 g03499(new_n5847, new_n5840_1, new_n5848);
not_10 g03500(new_n5848, new_n5849);
xnor_4 g03501(new_n5849, new_n5833_1, n463);
xor_4  g03502(n12121, n6775, new_n5851);
xor_4  g03503(new_n5851, n8920, new_n5852);
xor_4  g03504(new_n2991, n5438, new_n5853);
xor_4  g03505(new_n5853, new_n5852, n491);
xor_4  g03506(new_n5810, new_n5787, n496);
xor_4  g03507(n25926, n12384, new_n5856);
xor_4  g03508(new_n5856, n6773, new_n5857);
not_10 g03509(n16167, new_n5858);
xor_4  g03510(new_n5704_1, new_n5858, new_n5859);
and_5  g03511(new_n5859, new_n5857, new_n5860);
nor_5  g03512(new_n5704_1, new_n5858, new_n5861);
not_10 g03513(new_n5861, new_n5862);
not_10 g03514(new_n5702, new_n5863);
xor_4  g03515(new_n5863, n18745, new_n5864);
xor_4  g03516(new_n5864, new_n5862, new_n5865);
not_10 g03517(new_n5865, new_n5866);
and_5  g03518(n25926, n12384, new_n5867);
xor_4  g03519(n25926, n7657, new_n5868);
xor_4  g03520(new_n5868, n20986, new_n5869);
xor_4  g03521(new_n5869, new_n5867, new_n5870);
not_10 g03522(new_n5870, new_n5871);
nand_5 g03523(new_n5856, n6773, new_n5872);
or_5   g03524(new_n5872, n17090, new_n5873);
nor_5  g03525(n17090, n6773, new_n5874);
nand_5 g03526(n17090, n6773, new_n5875);
nor_5  g03527(new_n5875, new_n5856, new_n5876);
nor_5  g03528(new_n5876, new_n5874, new_n5877);
and_5  g03529(new_n5877, new_n5873, new_n5878);
xor_4  g03530(new_n5878, new_n5871, new_n5879);
xnor_4 g03531(new_n5879, new_n5866, new_n5880);
xor_4  g03532(new_n5880, new_n5860, n498);
xnor_4 g03533(n25872, n19618, new_n5882_1);
or_5   g03534(n22043, n20259, new_n5883);
nand_5 g03535(n12121, n3925, new_n5884);
xor_4  g03536(n22043, n20259, new_n5885);
nand_5 g03537(new_n5885, new_n5884, new_n5886);
and_5  g03538(new_n5886, new_n5883, new_n5887);
xor_4  g03539(new_n5887, new_n5882_1, new_n5888);
xnor_4 g03540(new_n5888, new_n4884, new_n5889);
xor_4  g03541(new_n5885, new_n5884, new_n5890);
or_5   g03542(new_n5890, new_n4888, new_n5891);
xnor_4 g03543(n12121, n3925, new_n5892);
nand_5 g03544(new_n5892, new_n4890, new_n5893);
xnor_4 g03545(new_n5890, new_n4887, new_n5894);
nand_5 g03546(new_n5894, new_n5893, new_n5895);
and_5  g03547(new_n5895, new_n5891, new_n5896);
xor_4  g03548(new_n5896, new_n5889, new_n5897);
xnor_4 g03549(new_n5897, new_n3782, new_n5898);
xor_4  g03550(new_n5894, new_n5893, new_n5899);
or_5   g03551(new_n5899, new_n3755_1, new_n5900);
and_5  g03552(new_n5899, new_n3788, new_n5901);
not_10 g03553(new_n3790, new_n5902);
xor_4  g03554(new_n5892, new_n4890, new_n5903_1);
nor_5  g03555(new_n5903_1, new_n5902, new_n5904_1);
or_5   g03556(new_n5904_1, new_n5901, new_n5905);
and_5  g03557(new_n5905, new_n5900, new_n5906);
xor_4  g03558(new_n5906, new_n5898, n521);
xor_4  g03559(new_n5796, new_n5795, n548);
xor_4  g03560(new_n4297, new_n4280, n554);
not_10 g03561(n2979, new_n5910);
not_10 g03562(n647, new_n5911_1);
not_10 g03563(n20409, new_n5912);
not_10 g03564(n25749, new_n5913);
nor_5  g03565(n20658, n15743, new_n5914);
and_5  g03566(new_n5914, new_n3785_1, new_n5915);
and_5  g03567(new_n5915, new_n3778, new_n5916);
and_5  g03568(new_n5916, new_n3776, new_n5917);
and_5  g03569(new_n5917, new_n3769, new_n5918);
and_5  g03570(new_n5918, new_n5913, new_n5919);
and_5  g03571(new_n5919, new_n5912, new_n5920);
and_5  g03572(new_n5920, new_n5911_1, new_n5921);
xor_4  g03573(new_n5921, new_n5910, new_n5922);
xor_4  g03574(n9259, n6456, new_n5923);
not_10 g03575(new_n5923, new_n5924);
or_5   g03576(n21489, n4085, new_n5925);
xor_4  g03577(n21489, n4085, new_n5926);
not_10 g03578(new_n5926, new_n5927);
or_5   g03579(n26725, n20213, new_n5928);
xor_4  g03580(n26725, n20213, new_n5929);
not_10 g03581(new_n5929, new_n5930);
or_5   g03582(n13912, n11980, new_n5931);
xor_4  g03583(n13912, n11980, new_n5932);
not_10 g03584(new_n5932, new_n5933);
or_5   g03585(n7670, n3253, new_n5934);
xor_4  g03586(n7670, n3253, new_n5935);
not_10 g03587(new_n5935, new_n5936_1);
or_5   g03588(n9598, n7759, new_n5937);
xor_4  g03589(n9598, n7759, new_n5938);
not_10 g03590(new_n5938, new_n5939);
or_5   g03591(n22290, n12562, new_n5940);
xor_4  g03592(n22290, n12562, new_n5941);
not_10 g03593(new_n5941, new_n5942);
or_5   g03594(n11273, n7949, new_n5943_1);
xor_4  g03595(n11273, n7949, new_n5944);
not_10 g03596(new_n5944, new_n5945);
or_5   g03597(n25565, n24374, new_n5946);
nand_5 g03598(n21993, n14575, new_n5947);
xor_4  g03599(n25565, n24374, new_n5948);
nand_5 g03600(new_n5948, new_n5947, new_n5949);
and_5  g03601(new_n5949, new_n5946, new_n5950);
or_5   g03602(new_n5950, new_n5945, new_n5951);
and_5  g03603(new_n5951, new_n5943_1, new_n5952);
or_5   g03604(new_n5952, new_n5942, new_n5953);
and_5  g03605(new_n5953, new_n5940, new_n5954);
or_5   g03606(new_n5954, new_n5939, new_n5955);
and_5  g03607(new_n5955, new_n5937, new_n5956);
or_5   g03608(new_n5956, new_n5936_1, new_n5957);
and_5  g03609(new_n5957, new_n5934, new_n5958);
or_5   g03610(new_n5958, new_n5933, new_n5959);
and_5  g03611(new_n5959, new_n5931, new_n5960);
or_5   g03612(new_n5960, new_n5930, new_n5961);
and_5  g03613(new_n5961, new_n5928, new_n5962);
or_5   g03614(new_n5962, new_n5927, new_n5963);
and_5  g03615(new_n5963, new_n5925, new_n5964_1);
xor_4  g03616(new_n5964_1, new_n5924, new_n5965);
not_10 g03617(new_n5965, new_n5966);
xnor_4 g03618(new_n5966, new_n5922, new_n5967);
not_10 g03619(new_n5967, new_n5968);
xor_4  g03620(new_n5920, new_n5911_1, new_n5969);
xor_4  g03621(new_n5962, new_n5927, new_n5970);
nand_5 g03622(new_n5970, new_n5969, new_n5971);
not_10 g03623(new_n5970, new_n5972);
xnor_4 g03624(new_n5972, new_n5969, new_n5973);
xor_4  g03625(new_n5919, new_n5912, new_n5974);
xor_4  g03626(new_n5960, new_n5930, new_n5975);
or_5   g03627(new_n5975, new_n5974, new_n5976);
not_10 g03628(new_n5975, new_n5977);
xnor_4 g03629(new_n5977, new_n5974, new_n5978);
not_10 g03630(new_n5978, new_n5979);
xor_4  g03631(new_n5918, new_n5913, new_n5980_1);
xor_4  g03632(new_n5958, new_n5933, new_n5981);
or_5   g03633(new_n5981, new_n5980_1, new_n5982);
not_10 g03634(new_n5981, new_n5983);
xnor_4 g03635(new_n5983, new_n5980_1, new_n5984);
not_10 g03636(new_n5984, new_n5985);
xor_4  g03637(new_n5917, new_n3769, new_n5986);
xor_4  g03638(new_n5956, new_n5936_1, new_n5987);
or_5   g03639(new_n5987, new_n5986, new_n5988);
not_10 g03640(new_n5987, new_n5989);
xnor_4 g03641(new_n5989, new_n5986, new_n5990);
not_10 g03642(new_n5990, new_n5991);
xor_4  g03643(new_n5916, new_n3776, new_n5992);
xor_4  g03644(new_n5954, new_n5939, new_n5993);
or_5   g03645(new_n5993, new_n5992, new_n5994);
not_10 g03646(new_n5993, new_n5995);
xnor_4 g03647(new_n5995, new_n5992, new_n5996);
not_10 g03648(new_n5996, new_n5997);
xor_4  g03649(new_n5915, new_n3778, new_n5998);
xor_4  g03650(new_n5952, new_n5942, new_n5999);
or_5   g03651(new_n5999, new_n5998, new_n6000);
not_10 g03652(new_n5999, new_n6001);
xnor_4 g03653(new_n6001, new_n5998, new_n6002);
xor_4  g03654(new_n5914, new_n3785_1, new_n6003);
xor_4  g03655(new_n5950, new_n5945, new_n6004);
nand_5 g03656(new_n6004, new_n6003, new_n6005);
not_10 g03657(new_n6004, new_n6006);
xnor_4 g03658(new_n6006, new_n6003, new_n6007);
not_10 g03659(n20658, new_n6008);
xor_4  g03660(n21993, n14575, new_n6009);
and_5  g03661(new_n6009, new_n6008, new_n6010);
not_10 g03662(new_n6010, new_n6011);
or_5   g03663(new_n6011, n15743, new_n6012_1);
xnor_4 g03664(new_n5948, new_n5947, new_n6013);
xor_4  g03665(n20658, n15743, new_n6014);
nand_5 g03666(new_n6014, new_n6011, new_n6015);
and_5  g03667(new_n6015, new_n6012_1, new_n6016);
nand_5 g03668(new_n6016, new_n6013, new_n6017);
and_5  g03669(new_n6017, new_n6012_1, new_n6018);
nand_5 g03670(new_n6018, new_n6007, new_n6019);
and_5  g03671(new_n6019, new_n6005, new_n6020);
nand_5 g03672(new_n6020, new_n6002, new_n6021);
and_5  g03673(new_n6021, new_n6000, new_n6022_1);
or_5   g03674(new_n6022_1, new_n5997, new_n6023);
and_5  g03675(new_n6023, new_n5994, new_n6024);
or_5   g03676(new_n6024, new_n5991, new_n6025);
and_5  g03677(new_n6025, new_n5988, new_n6026);
or_5   g03678(new_n6026, new_n5985, new_n6027);
and_5  g03679(new_n6027, new_n5982, new_n6028);
or_5   g03680(new_n6028, new_n5979, new_n6029);
and_5  g03681(new_n6029, new_n5976, new_n6030);
nand_5 g03682(new_n6030, new_n5973, new_n6031_1);
and_5  g03683(new_n6031_1, new_n5971, new_n6032);
xor_4  g03684(new_n6032, new_n5968, new_n6033);
not_10 g03685(new_n6033, new_n6034);
not_10 g03686(n8526, new_n6035);
xnor_4 g03687(n21784, n3582, new_n6036);
or_5   g03688(n5521, n2145, new_n6037);
xnor_4 g03689(n5521, n2145, new_n6038);
or_5   g03690(n11926, n5031, new_n6039);
xnor_4 g03691(n11926, n5031, new_n6040);
or_5   g03692(n11044, n4325, new_n6041);
xnor_4 g03693(n11044, n4325, new_n6042);
or_5   g03694(n5337, n2421, new_n6043);
xnor_4 g03695(n5337, n2421, new_n6044_1);
or_5   g03696(n987, n626, new_n6045);
xnor_4 g03697(n987, n626, new_n6046_1);
or_5   g03698(n20478, n1204, new_n6047);
xnor_4 g03699(n20478, n1204, new_n6048);
or_5   g03700(n26882, n19618, new_n6049);
xnor_4 g03701(n26882, n19618, new_n6050);
or_5   g03702(n22619, n22043, new_n6051);
nand_5 g03703(n12121, n6775, new_n6052);
xor_4  g03704(n22619, n22043, new_n6053);
nand_5 g03705(new_n6053, new_n6052, new_n6054);
and_5  g03706(new_n6054, new_n6051, new_n6055);
or_5   g03707(new_n6055, new_n6050, new_n6056);
and_5  g03708(new_n6056, new_n6049, new_n6057);
or_5   g03709(new_n6057, new_n6048, new_n6058);
and_5  g03710(new_n6058, new_n6047, new_n6059);
or_5   g03711(new_n6059, new_n6046_1, new_n6060);
and_5  g03712(new_n6060, new_n6045, new_n6061);
or_5   g03713(new_n6061, new_n6044_1, new_n6062);
and_5  g03714(new_n6062, new_n6043, new_n6063);
or_5   g03715(new_n6063, new_n6042, new_n6064);
and_5  g03716(new_n6064, new_n6041, new_n6065);
or_5   g03717(new_n6065, new_n6040, new_n6066);
and_5  g03718(new_n6066, new_n6039, new_n6067);
or_5   g03719(new_n6067, new_n6038, new_n6068);
and_5  g03720(new_n6068, new_n6037, new_n6069);
xor_4  g03721(new_n6069, new_n6036, new_n6070);
xor_4  g03722(new_n6070, new_n6035, new_n6071);
not_10 g03723(new_n6071, new_n6072);
not_10 g03724(n2816, new_n6073);
xor_4  g03725(new_n6067, new_n6038, new_n6074);
or_5   g03726(new_n6074, new_n6073, new_n6075);
xor_4  g03727(new_n6074, new_n6073, new_n6076);
not_10 g03728(new_n6076, new_n6077);
not_10 g03729(n20359, new_n6078);
xor_4  g03730(new_n6065, new_n6040, new_n6079);
or_5   g03731(new_n6079, new_n6078, new_n6080);
xor_4  g03732(new_n6079, new_n6078, new_n6081);
not_10 g03733(new_n6081, new_n6082);
not_10 g03734(n4409, new_n6083);
xor_4  g03735(new_n6063, new_n6042, new_n6084_1);
or_5   g03736(new_n6084_1, new_n6083, new_n6085);
xor_4  g03737(new_n6084_1, new_n6083, new_n6086);
not_10 g03738(new_n6086, new_n6087);
not_10 g03739(n3570, new_n6088);
xor_4  g03740(new_n6061, new_n6044_1, new_n6089);
or_5   g03741(new_n6089, new_n6088, new_n6090);
xor_4  g03742(new_n6089, new_n6088, new_n6091);
not_10 g03743(new_n6091, new_n6092);
xor_4  g03744(new_n6059, new_n6046_1, new_n6093);
or_5   g03745(new_n6093, new_n4220, new_n6094);
xor_4  g03746(new_n6093, new_n4220, new_n6095);
not_10 g03747(new_n6095, new_n6096);
xor_4  g03748(new_n6057, new_n6048, new_n6097);
or_5   g03749(new_n6097, new_n4221_1, new_n6098);
xor_4  g03750(new_n6097, new_n4221_1, new_n6099);
not_10 g03751(new_n6099, new_n6100);
xor_4  g03752(new_n6055, new_n6050, new_n6101);
or_5   g03753(new_n6101, new_n4222, new_n6102);
not_10 g03754(n10057, new_n6103);
xor_4  g03755(new_n6053, new_n6052, new_n6104_1);
and_5  g03756(new_n6104_1, new_n6103, new_n6105_1);
and_5  g03757(new_n5851, n8920, new_n6106);
not_10 g03758(new_n6106, new_n6107);
xor_4  g03759(new_n6104_1, new_n6103, new_n6108);
and_5  g03760(new_n6108, new_n6107, new_n6109);
nor_5  g03761(new_n6109, new_n6105_1, new_n6110);
xor_4  g03762(new_n6101, new_n4222, new_n6111);
nand_5 g03763(new_n6111, new_n6110, new_n6112);
and_5  g03764(new_n6112, new_n6102, new_n6113);
or_5   g03765(new_n6113, new_n6100, new_n6114);
and_5  g03766(new_n6114, new_n6098, new_n6115);
or_5   g03767(new_n6115, new_n6096, new_n6116);
and_5  g03768(new_n6116, new_n6094, new_n6117);
or_5   g03769(new_n6117, new_n6092, new_n6118);
and_5  g03770(new_n6118, new_n6090, new_n6119);
or_5   g03771(new_n6119, new_n6087, new_n6120);
and_5  g03772(new_n6120, new_n6085, new_n6121);
or_5   g03773(new_n6121, new_n6082, new_n6122);
and_5  g03774(new_n6122, new_n6080, new_n6123);
or_5   g03775(new_n6123, new_n6077, new_n6124);
and_5  g03776(new_n6124, new_n6075, new_n6125);
xor_4  g03777(new_n6125, new_n6072, new_n6126);
xnor_4 g03778(new_n6126, new_n6034, new_n6127);
xor_4  g03779(new_n6123, new_n6077, new_n6128);
xor_4  g03780(new_n6030, new_n5973, new_n6129);
nor_5  g03781(new_n6129, new_n6128, new_n6130);
xor_4  g03782(new_n6129, new_n6128, new_n6131);
not_10 g03783(new_n6131, new_n6132);
xor_4  g03784(new_n6028, new_n5979, new_n6133);
not_10 g03785(new_n6133, new_n6134);
xor_4  g03786(new_n6121, new_n6082, new_n6135);
nor_5  g03787(new_n6135, new_n6134, new_n6136);
xor_4  g03788(new_n6135, new_n6134, new_n6137);
xor_4  g03789(new_n6026, new_n5985, new_n6138);
not_10 g03790(new_n6138, new_n6139);
xor_4  g03791(new_n6119, new_n6087, new_n6140);
nor_5  g03792(new_n6140, new_n6139, new_n6141);
xor_4  g03793(new_n6140, new_n6139, new_n6142);
xor_4  g03794(new_n6024, new_n5991, new_n6143);
not_10 g03795(new_n6143, new_n6144);
xor_4  g03796(new_n6117, new_n6092, new_n6145);
nor_5  g03797(new_n6145, new_n6144, new_n6146);
xor_4  g03798(new_n6145, new_n6144, new_n6147);
xnor_4 g03799(new_n6022_1, new_n5996, new_n6148);
not_10 g03800(new_n6148, new_n6149);
xor_4  g03801(new_n6115, new_n6096, new_n6150);
nor_5  g03802(new_n6150, new_n6149, new_n6151);
xor_4  g03803(new_n6150, new_n6149, new_n6152);
xor_4  g03804(new_n6020, new_n6002, new_n6153);
not_10 g03805(new_n6153, new_n6154);
xor_4  g03806(new_n6113, new_n6100, new_n6155);
nor_5  g03807(new_n6155, new_n6154, new_n6156);
xor_4  g03808(new_n6155, new_n6154, new_n6157);
xor_4  g03809(new_n6018, new_n6007, new_n6158);
not_10 g03810(new_n6158, new_n6159);
xor_4  g03811(new_n6111, new_n6110, new_n6160_1);
not_10 g03812(new_n6160_1, new_n6161);
and_5  g03813(new_n6161, new_n6159, new_n6162);
xor_4  g03814(new_n6161, new_n6159, new_n6163);
xor_4  g03815(new_n6108, new_n6107, new_n6164);
xor_4  g03816(new_n6016, new_n6013, new_n6165);
nor_5  g03817(new_n6165, new_n6164, new_n6166);
not_10 g03818(new_n5852, new_n6167);
xor_4  g03819(new_n6009, new_n6008, new_n6168);
nor_5  g03820(new_n6168, new_n6167, new_n6169);
xor_4  g03821(new_n6165, new_n6164, new_n6170);
and_5  g03822(new_n6170, new_n6169, new_n6171_1);
nor_5  g03823(new_n6171_1, new_n6166, new_n6172);
and_5  g03824(new_n6172, new_n6163, new_n6173);
nor_5  g03825(new_n6173, new_n6162, new_n6174);
not_10 g03826(new_n6174, new_n6175);
and_5  g03827(new_n6175, new_n6157, new_n6176);
nor_5  g03828(new_n6176, new_n6156, new_n6177);
not_10 g03829(new_n6177, new_n6178);
and_5  g03830(new_n6178, new_n6152, new_n6179);
nor_5  g03831(new_n6179, new_n6151, new_n6180);
not_10 g03832(new_n6180, new_n6181);
and_5  g03833(new_n6181, new_n6147, new_n6182);
nor_5  g03834(new_n6182, new_n6146, new_n6183_1);
not_10 g03835(new_n6183_1, new_n6184);
and_5  g03836(new_n6184, new_n6142, new_n6185);
nor_5  g03837(new_n6185, new_n6141, new_n6186);
not_10 g03838(new_n6186, new_n6187);
and_5  g03839(new_n6187, new_n6137, new_n6188);
nor_5  g03840(new_n6188, new_n6136, new_n6189_1);
nor_5  g03841(new_n6189_1, new_n6132, new_n6190);
nor_5  g03842(new_n6190, new_n6130, new_n6191);
xor_4  g03843(new_n6191, new_n6127, n567);
nor_5  g03844(n10250, n1831, new_n6193);
xnor_4 g03845(n10250, n1831, new_n6194);
or_5   g03846(n13137, n7674, new_n6195);
xor_4  g03847(n13137, n7674, new_n6196);
not_10 g03848(new_n6196, new_n6197);
or_5   g03849(n18452, n6397, new_n6198);
xor_4  g03850(n18452, n6397, new_n6199);
not_10 g03851(new_n6199, new_n6200);
or_5   g03852(n21317, n19196, new_n6201);
xor_4  g03853(n21317, n19196, new_n6202);
not_10 g03854(new_n6202, new_n6203);
or_5   g03855(n23586, n12398, new_n6204_1);
xor_4  g03856(n23586, n12398, new_n6205);
not_10 g03857(new_n6205, new_n6206);
or_5   g03858(n21226, n19789, new_n6207);
xor_4  g03859(n21226, n19789, new_n6208);
not_10 g03860(new_n6208, new_n6209);
or_5   g03861(n20169, n4426, new_n6210);
xnor_4 g03862(n20169, n4426, new_n6211);
or_5   g03863(n20036, n8285, new_n6212);
xor_4  g03864(n20036, n8285, new_n6213);
not_10 g03865(new_n6213, new_n6214);
or_5   g03866(n11192, n6729, new_n6215);
nand_5 g03867(n21687, n9380, new_n6216);
xor_4  g03868(n11192, n6729, new_n6217);
nand_5 g03869(new_n6217, new_n6216, new_n6218_1);
and_5  g03870(new_n6218_1, new_n6215, new_n6219);
or_5   g03871(new_n6219, new_n6214, new_n6220);
and_5  g03872(new_n6220, new_n6212, new_n6221);
or_5   g03873(new_n6221, new_n6211, new_n6222);
and_5  g03874(new_n6222, new_n6210, new_n6223_1);
or_5   g03875(new_n6223_1, new_n6209, new_n6224);
and_5  g03876(new_n6224, new_n6207, new_n6225);
or_5   g03877(new_n6225, new_n6206, new_n6226);
and_5  g03878(new_n6226, new_n6204_1, new_n6227);
or_5   g03879(new_n6227, new_n6203, new_n6228);
and_5  g03880(new_n6228, new_n6201, new_n6229);
or_5   g03881(new_n6229, new_n6200, new_n6230);
and_5  g03882(new_n6230, new_n6198, new_n6231);
or_5   g03883(new_n6231, new_n6197, new_n6232);
and_5  g03884(new_n6232, new_n6195, new_n6233_1);
nor_5  g03885(new_n6233_1, new_n6194, new_n6234);
or_5   g03886(new_n6234, new_n6193, new_n6235);
not_10 g03887(n3320, new_n6236);
not_10 g03888(n1288, new_n6237);
not_10 g03889(n1752, new_n6238);
not_10 g03890(n13110, new_n6239);
and_5  g03891(new_n4017, new_n4010_1, new_n6240);
and_5  g03892(new_n6240, new_n6239, new_n6241);
and_5  g03893(new_n6241, new_n6238, new_n6242);
and_5  g03894(new_n6242, new_n6237, new_n6243);
xor_4  g03895(new_n6243, new_n6236, new_n6244);
not_10 g03896(new_n6244, new_n6245_1);
nor_5  g03897(new_n6245_1, new_n5480, new_n6246);
not_10 g03898(new_n6246, new_n6247);
and_5  g03899(new_n6243, new_n6236, new_n6248_1);
and_5  g03900(new_n6245_1, new_n5480, new_n6249);
xor_4  g03901(new_n6242, new_n6237, new_n6250);
nor_5  g03902(new_n6250, n15182, new_n6251);
xor_4  g03903(new_n6250, n15182, new_n6252);
not_10 g03904(new_n6252, new_n6253);
xor_4  g03905(new_n6241, new_n6238, new_n6254);
or_5   g03906(new_n6254, n27037, new_n6255);
xor_4  g03907(new_n6254, n27037, new_n6256_1);
xor_4  g03908(new_n6240, new_n6239, new_n6257);
nand_5 g03909(new_n6257, n8964, new_n6258);
not_10 g03910(n8964, new_n6259);
xor_4  g03911(new_n6257, new_n6259, new_n6260);
nand_5 g03912(new_n4018, n20151, new_n6261);
or_5   g03913(new_n4044, new_n4019, new_n6262);
and_5  g03914(new_n6262, new_n6261, new_n6263);
or_5   g03915(new_n6263, new_n6260, new_n6264);
and_5  g03916(new_n6264, new_n6258, new_n6265);
nand_5 g03917(new_n6265, new_n6256_1, new_n6266);
and_5  g03918(new_n6266, new_n6255, new_n6267);
nor_5  g03919(new_n6267, new_n6253, new_n6268);
nor_5  g03920(new_n6268, new_n6251, new_n6269);
not_10 g03921(new_n6269, new_n6270);
nor_5  g03922(new_n6270, new_n6249, new_n6271_1);
nor_5  g03923(new_n6271_1, new_n6248_1, new_n6272);
and_5  g03924(new_n6272, new_n6247, new_n6273);
not_10 g03925(new_n6273, new_n6274);
and_5  g03926(new_n6274, new_n6235, new_n6275);
xnor_4 g03927(new_n6273, new_n6235, new_n6276_1);
xor_4  g03928(new_n6233_1, new_n6194, new_n6277);
not_10 g03929(new_n6277, new_n6278);
or_5   g03930(new_n6249, new_n6246, new_n6279);
xor_4  g03931(new_n6279, new_n6270, new_n6280);
nand_5 g03932(new_n6280, new_n6278, new_n6281);
xor_4  g03933(new_n6267, new_n6253, new_n6282);
not_10 g03934(new_n6282, new_n6283);
xor_4  g03935(new_n6231, new_n6197, new_n6284);
not_10 g03936(new_n6284, new_n6285);
nor_5  g03937(new_n6285, new_n6283, new_n6286);
xor_4  g03938(new_n6285, new_n6283, new_n6287);
not_10 g03939(new_n6287, new_n6288);
xor_4  g03940(new_n6265, new_n6256_1, new_n6289);
not_10 g03941(new_n6289, new_n6290);
xor_4  g03942(new_n6229, new_n6200, new_n6291);
not_10 g03943(new_n6291, new_n6292);
or_5   g03944(new_n6292, new_n6290, new_n6293);
xor_4  g03945(new_n6292, new_n6290, new_n6294);
xor_4  g03946(new_n6227, new_n6203, new_n6295);
not_10 g03947(new_n6295, new_n6296);
xor_4  g03948(new_n6263, new_n6260, new_n6297);
nand_5 g03949(new_n6297, new_n6296, new_n6298);
xor_4  g03950(new_n6225, new_n6206, new_n6299);
not_10 g03951(new_n6299, new_n6300);
or_5   g03952(new_n6300, new_n4045, new_n6301);
xor_4  g03953(new_n6300, new_n4045, new_n6302);
not_10 g03954(new_n6302, new_n6303);
xor_4  g03955(new_n6223_1, new_n6209, new_n6304);
not_10 g03956(new_n6304, new_n6305);
xor_4  g03957(new_n6221, new_n6211, new_n6306);
nand_5 g03958(new_n6306, new_n4055, new_n6307);
xor_4  g03959(new_n6219, new_n6214, new_n6308_1);
not_10 g03960(new_n6308_1, new_n6309);
and_5  g03961(new_n6309, new_n4058, new_n6310);
xor_4  g03962(new_n6308_1, new_n4058, new_n6311_1);
xor_4  g03963(new_n6217, new_n6216, new_n6312);
or_5   g03964(new_n6312, new_n4063, new_n6313);
xor_4  g03965(n21687, n9380, new_n6314);
and_5  g03966(new_n6314, new_n2552, new_n6315);
xor_4  g03967(new_n6312, new_n4063, new_n6316);
nand_5 g03968(new_n6316, new_n6315, new_n6317);
and_5  g03969(new_n6317, new_n6313, new_n6318);
nor_5  g03970(new_n6318, new_n6311_1, new_n6319);
nor_5  g03971(new_n6319, new_n6310, new_n6320);
xor_4  g03972(new_n6306, new_n4055, new_n6321);
nand_5 g03973(new_n6321, new_n6320, new_n6322);
and_5  g03974(new_n6322, new_n6307, new_n6323_1);
or_5   g03975(new_n6323_1, new_n6305, new_n6324);
not_10 g03976(new_n4049, new_n6325);
xnor_4 g03977(new_n6323_1, new_n6304, new_n6326);
nand_5 g03978(new_n6326, new_n6325, new_n6327);
and_5  g03979(new_n6327, new_n6324, new_n6328);
or_5   g03980(new_n6328, new_n6303, new_n6329);
and_5  g03981(new_n6329, new_n6301, new_n6330_1);
xor_4  g03982(new_n6297, new_n6296, new_n6331);
nand_5 g03983(new_n6331, new_n6330_1, new_n6332);
and_5  g03984(new_n6332, new_n6298, new_n6333);
nand_5 g03985(new_n6333, new_n6294, new_n6334);
and_5  g03986(new_n6334, new_n6293, new_n6335);
nor_5  g03987(new_n6335, new_n6288, new_n6336);
or_5   g03988(new_n6336, new_n6286, new_n6337);
xor_4  g03989(new_n6280, new_n6278, new_n6338);
not_10 g03990(new_n6338, new_n6339_1);
or_5   g03991(new_n6339_1, new_n6337, new_n6340);
and_5  g03992(new_n6340, new_n6281, new_n6341);
and_5  g03993(new_n6341, new_n6276_1, new_n6342);
nor_5  g03994(new_n6342, new_n6275, new_n6343);
xor_4  g03995(new_n6341, new_n6276_1, new_n6344);
or_5   g03996(n15766, n6105, new_n6345);
xor_4  g03997(n15766, n6105, new_n6346);
not_10 g03998(new_n6346, new_n6347);
or_5   g03999(n25629, n3795, new_n6348);
xor_4  g04000(n25629, n3795, new_n6349);
not_10 g04001(new_n6349, new_n6350);
or_5   g04002(n25464, n7692, new_n6351);
xor_4  g04003(n25464, n7692, new_n6352);
not_10 g04004(new_n6352, new_n6353);
or_5   g04005(n23039, n4590, new_n6354_1);
xor_4  g04006(n23039, n4590, new_n6355);
not_10 g04007(new_n6355, new_n6356_1);
or_5   g04008(n26752, n13677, new_n6357);
xor_4  g04009(n26752, n13677, new_n6358);
not_10 g04010(new_n6358, new_n6359);
or_5   g04011(n18926, n6513, new_n6360);
xor_4  g04012(n18926, n6513, new_n6361);
nand_5 g04013(n5451, n3918, new_n6362);
or_5   g04014(n5451, n3918, new_n6363);
nor_5  g04015(n5330, n919, new_n6364);
nor_5  g04016(new_n4149, new_n4144, new_n6365);
nor_5  g04017(new_n6365, new_n6364, new_n6366);
nand_5 g04018(new_n6366, new_n6363, new_n6367);
and_5  g04019(new_n6367, new_n6362, new_n6368);
nand_5 g04020(new_n6368, new_n6361, new_n6369_1);
and_5  g04021(new_n6369_1, new_n6360, new_n6370);
or_5   g04022(new_n6370, new_n6359, new_n6371);
and_5  g04023(new_n6371, new_n6357, new_n6372);
or_5   g04024(new_n6372, new_n6356_1, new_n6373);
and_5  g04025(new_n6373, new_n6354_1, new_n6374);
or_5   g04026(new_n6374, new_n6353, new_n6375_1);
and_5  g04027(new_n6375_1, new_n6351, new_n6376);
or_5   g04028(new_n6376, new_n6350, new_n6377);
and_5  g04029(new_n6377, new_n6348, new_n6378);
or_5   g04030(new_n6378, new_n6347, new_n6379_1);
and_5  g04031(new_n6379_1, new_n6345, new_n6380);
and_5  g04032(new_n6380, new_n6344, new_n6381_1);
xor_4  g04033(new_n6380, new_n6344, new_n6382);
not_10 g04034(new_n6382, new_n6383_1);
xor_4  g04035(new_n6378, new_n6347, new_n6384);
xnor_4 g04036(new_n6338, new_n6337, new_n6385_1);
nor_5  g04037(new_n6385_1, new_n6384, new_n6386);
xor_4  g04038(new_n6385_1, new_n6384, new_n6387);
not_10 g04039(new_n6387, new_n6388);
xnor_4 g04040(new_n6335, new_n6287, new_n6389);
not_10 g04041(new_n6389, new_n6390);
xor_4  g04042(new_n6376, new_n6350, new_n6391);
nor_5  g04043(new_n6391, new_n6390, new_n6392);
xor_4  g04044(new_n6391, new_n6390, new_n6393);
xor_4  g04045(new_n6333, new_n6294, new_n6394);
not_10 g04046(new_n6394, new_n6395);
xor_4  g04047(new_n6374, new_n6353, new_n6396);
nor_5  g04048(new_n6396, new_n6395, new_n6397_1);
xor_4  g04049(new_n6396, new_n6395, new_n6398);
xor_4  g04050(new_n6372, new_n6356_1, new_n6399);
xor_4  g04051(new_n6331, new_n6330_1, new_n6400);
nor_5  g04052(new_n6400, new_n6399, new_n6401);
xor_4  g04053(new_n6400, new_n6399, new_n6402);
not_10 g04054(new_n6402, new_n6403);
xor_4  g04055(new_n6328, new_n6303, new_n6404);
xor_4  g04056(new_n6370, new_n6359, new_n6405);
not_10 g04057(new_n6405, new_n6406);
and_5  g04058(new_n6406, new_n6404, new_n6407_1);
xor_4  g04059(new_n6406, new_n6404, new_n6408);
not_10 g04060(new_n6408, new_n6409);
xnor_4 g04061(new_n6326, new_n4049, new_n6410);
not_10 g04062(new_n6410, new_n6411);
xor_4  g04063(new_n6368, new_n6361, new_n6412);
nor_5  g04064(new_n6412, new_n6411, new_n6413);
xor_4  g04065(new_n6412, new_n6411, new_n6414);
xor_4  g04066(new_n6321, new_n6320, new_n6415);
xor_4  g04067(n5451, n3918, new_n6416);
xor_4  g04068(new_n6416, new_n6366, new_n6417);
and_5  g04069(new_n6417, new_n6415, new_n6418);
xor_4  g04070(new_n6417, new_n6415, new_n6419);
not_10 g04071(new_n6419, new_n6420);
xor_4  g04072(new_n6318, new_n6311_1, new_n6421);
nor_5  g04073(new_n6421, new_n4150_1, new_n6422);
xor_4  g04074(new_n6421, new_n4150_1, new_n6423);
not_10 g04075(new_n6423, new_n6424);
xor_4  g04076(new_n6316, new_n6315, new_n6425);
nor_5  g04077(new_n6425, new_n4153_1, new_n6426);
not_10 g04078(new_n6426, new_n6427_1);
xor_4  g04079(new_n6314, new_n2552, new_n6428);
not_10 g04080(new_n6428, new_n6429);
and_5  g04081(new_n6429, new_n4156, new_n6430);
xor_4  g04082(new_n6425, new_n4153_1, new_n6431_1);
and_5  g04083(new_n6431_1, new_n6430, new_n6432);
not_10 g04084(new_n6432, new_n6433);
and_5  g04085(new_n6433, new_n6427_1, new_n6434);
nor_5  g04086(new_n6434, new_n6424, new_n6435);
nor_5  g04087(new_n6435, new_n6422, new_n6436);
nor_5  g04088(new_n6436, new_n6420, new_n6437_1);
nor_5  g04089(new_n6437_1, new_n6418, new_n6438);
not_10 g04090(new_n6438, new_n6439);
and_5  g04091(new_n6439, new_n6414, new_n6440);
nor_5  g04092(new_n6440, new_n6413, new_n6441);
nor_5  g04093(new_n6441, new_n6409, new_n6442);
nor_5  g04094(new_n6442, new_n6407_1, new_n6443);
nor_5  g04095(new_n6443, new_n6403, new_n6444);
nor_5  g04096(new_n6444, new_n6401, new_n6445);
not_10 g04097(new_n6445, new_n6446);
and_5  g04098(new_n6446, new_n6398, new_n6447);
nor_5  g04099(new_n6447, new_n6397_1, new_n6448);
not_10 g04100(new_n6448, new_n6449);
and_5  g04101(new_n6449, new_n6393, new_n6450);
nor_5  g04102(new_n6450, new_n6392, new_n6451);
nor_5  g04103(new_n6451, new_n6388, new_n6452);
nor_5  g04104(new_n6452, new_n6386, new_n6453);
nor_5  g04105(new_n6453, new_n6383_1, new_n6454);
nor_5  g04106(new_n6454, new_n6381_1, new_n6455);
nor_5  g04107(new_n6455, new_n6343, n588);
xnor_4 g04108(n19803, n18584, new_n6457_1);
not_10 g04109(new_n6457_1, new_n6458);
not_10 g04110(n12626, new_n6459);
or_5   g04111(new_n6459, n4272, new_n6460);
or_5   g04112(new_n4694, new_n4669, new_n6461);
and_5  g04113(new_n6461, new_n6460, new_n6462);
xor_4  g04114(new_n6462, new_n6458, new_n6463);
xnor_4 g04115(n16911, n7773, new_n6464);
not_10 g04116(new_n6464, new_n6465_1);
not_10 g04117(n376, new_n6466);
or_5   g04118(n7721, new_n6466, new_n6467);
xnor_4 g04119(n7721, n376, new_n6468);
not_10 g04120(new_n6468, new_n6469);
not_10 g04121(n5517, new_n6470_1);
or_5   g04122(n21981, new_n6470_1, new_n6471);
xnor_4 g04123(n21981, n5517, new_n6472);
not_10 g04124(new_n6472, new_n6473);
not_10 g04125(n12113, new_n6474);
or_5   g04126(n12917, new_n6474, new_n6475);
xnor_4 g04127(n12917, n12113, new_n6476_1);
not_10 g04128(n21898, new_n6477);
or_5   g04129(new_n6477, n10614, new_n6478);
nand_5 g04130(new_n6477, n10614, new_n6479);
not_10 g04131(n11266, new_n6480);
and_5  g04132(new_n6480, n9926, new_n6481);
nor_5  g04133(new_n6480, n9926, new_n6482);
not_10 g04134(n2646, new_n6483);
and_5  g04135(n22072, new_n6483, new_n6484);
not_10 g04136(new_n6484, new_n6485_1);
nor_5  g04137(new_n6485_1, new_n6482, new_n6486);
nor_5  g04138(new_n6486, new_n6481, new_n6487);
not_10 g04139(new_n6487, new_n6488);
nand_5 g04140(new_n6488, new_n6479, new_n6489);
and_5  g04141(new_n6489, new_n6478, new_n6490);
nand_5 g04142(new_n6490, new_n6476_1, new_n6491);
and_5  g04143(new_n6491, new_n6475, new_n6492);
or_5   g04144(new_n6492, new_n6473, new_n6493);
and_5  g04145(new_n6493, new_n6471, new_n6494);
or_5   g04146(new_n6494, new_n6469, new_n6495);
and_5  g04147(new_n6495, new_n6467, new_n6496);
xor_4  g04148(new_n6496, new_n6465_1, new_n6497);
not_10 g04149(new_n6497, new_n6498);
not_10 g04150(n1742, new_n6499);
not_10 g04151(n16818, new_n6500);
not_10 g04152(n1269, new_n6501);
not_10 g04153(n14576, new_n6502_1);
not_10 g04154(n2985, new_n6503);
not_10 g04155(n5605, new_n6504);
nor_5  g04156(n15652, n4939, new_n6505);
and_5  g04157(new_n6505, new_n6504, new_n6506_1);
and_5  g04158(new_n6506_1, new_n6503, new_n6507);
and_5  g04159(new_n6507, new_n6502_1, new_n6508);
and_5  g04160(new_n6508, new_n6501, new_n6509);
xor_4  g04161(new_n6509, new_n6500, new_n6510);
not_10 g04162(new_n6510, new_n6511);
nor_5  g04163(new_n6511, new_n6499, new_n6512);
and_5  g04164(new_n6511, new_n6499, new_n6513_1);
or_5   g04165(new_n6513_1, new_n6512, new_n6514_1);
not_10 g04166(n4858, new_n6515);
xor_4  g04167(new_n6508, new_n6501, new_n6516);
not_10 g04168(new_n6516, new_n6517);
and_5  g04169(new_n6517, new_n6515, new_n6518);
xor_4  g04170(new_n6517, n4858, new_n6519);
not_10 g04171(n8244, new_n6520);
xor_4  g04172(new_n6507, new_n6502_1, new_n6521);
not_10 g04173(new_n6521, new_n6522);
nand_5 g04174(new_n6522, new_n6520, new_n6523);
xor_4  g04175(new_n6522, n8244, new_n6524);
not_10 g04176(n9493, new_n6525);
xor_4  g04177(new_n6506_1, new_n6503, new_n6526);
not_10 g04178(new_n6526, new_n6527);
nand_5 g04179(new_n6527, new_n6525, new_n6528);
not_10 g04180(n15167, new_n6529);
xor_4  g04181(new_n6505, new_n6504, new_n6530);
not_10 g04182(new_n6530, new_n6531);
and_5  g04183(new_n6531, new_n6529, new_n6532);
xor_4  g04184(new_n6531, new_n6529, new_n6533);
not_10 g04185(new_n6533, new_n6534);
xor_4  g04186(n15652, n4939, new_n6535);
or_5   g04187(new_n6535, n21095, new_n6536);
and_5  g04188(n8656, n4939, new_n6537);
not_10 g04189(new_n6537, new_n6538);
xor_4  g04190(new_n6535, n21095, new_n6539);
nand_5 g04191(new_n6539, new_n6538, new_n6540);
and_5  g04192(new_n6540, new_n6536, new_n6541);
nor_5  g04193(new_n6541, new_n6534, new_n6542_1);
or_5   g04194(new_n6542_1, new_n6532, new_n6543);
xor_4  g04195(new_n6527, new_n6525, new_n6544);
nand_5 g04196(new_n6544, new_n6543, new_n6545);
and_5  g04197(new_n6545, new_n6528, new_n6546);
or_5   g04198(new_n6546, new_n6524, new_n6547);
and_5  g04199(new_n6547, new_n6523, new_n6548);
nor_5  g04200(new_n6548, new_n6519, new_n6549);
nor_5  g04201(new_n6549, new_n6518, new_n6550);
xor_4  g04202(new_n6550, new_n6514_1, new_n6551);
xnor_4 g04203(new_n6551, new_n6498, new_n6552);
xor_4  g04204(new_n6494, new_n6469, new_n6553);
not_10 g04205(new_n6553, new_n6554);
xor_4  g04206(new_n6548, new_n6519, new_n6555);
or_5   g04207(new_n6555, new_n6554, new_n6556_1);
xnor_4 g04208(new_n6555, new_n6553, new_n6557);
xor_4  g04209(new_n6492, new_n6473, new_n6558_1);
not_10 g04210(new_n6558_1, new_n6559);
xor_4  g04211(new_n6546, new_n6524, new_n6560_1);
nand_5 g04212(new_n6560_1, new_n6559, new_n6561);
xnor_4 g04213(new_n6560_1, new_n6558_1, new_n6562);
xor_4  g04214(new_n6490, new_n6476_1, new_n6563);
not_10 g04215(new_n6563, new_n6564);
xor_4  g04216(new_n6544, new_n6543, new_n6565);
or_5   g04217(new_n6565, new_n6564, new_n6566);
xor_4  g04218(new_n6541, new_n6534, new_n6567_1);
xnor_4 g04219(n21898, n10614, new_n6568);
xor_4  g04220(new_n6568, new_n6488, new_n6569);
and_5  g04221(new_n6569, new_n6567_1, new_n6570);
xnor_4 g04222(new_n6569, new_n6567_1, new_n6571);
xor_4  g04223(n8656, n4939, new_n6572);
not_10 g04224(new_n6572, new_n6573);
xnor_4 g04225(n22072, n2646, new_n6574);
nor_5  g04226(new_n6574, new_n6573, new_n6575);
not_10 g04227(new_n6575, new_n6576_1);
xnor_4 g04228(n11266, n9926, new_n6577);
xnor_4 g04229(new_n6577, new_n6485_1, new_n6578);
nand_5 g04230(new_n6578, new_n6576_1, new_n6579);
xor_4  g04231(new_n6539, new_n6538, new_n6580);
xnor_4 g04232(new_n6578, new_n6575, new_n6581);
nand_5 g04233(new_n6581, new_n6580, new_n6582);
and_5  g04234(new_n6582, new_n6579, new_n6583);
nor_5  g04235(new_n6583, new_n6571, new_n6584);
nor_5  g04236(new_n6584, new_n6570, new_n6585);
xnor_4 g04237(new_n6565, new_n6563, new_n6586);
nand_5 g04238(new_n6586, new_n6585, new_n6587_1);
and_5  g04239(new_n6587_1, new_n6566, new_n6588);
nand_5 g04240(new_n6588, new_n6562, new_n6589);
and_5  g04241(new_n6589, new_n6561, new_n6590_1);
nand_5 g04242(new_n6590_1, new_n6557, new_n6591);
and_5  g04243(new_n6591, new_n6556_1, new_n6592);
xor_4  g04244(new_n6592, new_n6552, new_n6593);
xor_4  g04245(new_n6593, new_n6463, new_n6594);
xor_4  g04246(new_n6590_1, new_n6557, new_n6595);
or_5   g04247(new_n6595, new_n4695, new_n6596_1);
xor_4  g04248(new_n6595, new_n4695, new_n6597);
not_10 g04249(new_n6597, new_n6598);
xor_4  g04250(new_n6588, new_n6562, new_n6599);
not_10 g04251(new_n6599, new_n6600);
or_5   g04252(new_n6600, new_n4699, new_n6601);
xor_4  g04253(new_n6600, new_n4699, new_n6602);
xor_4  g04254(new_n6586, new_n6585, new_n6603);
or_5   g04255(new_n6603, new_n4704, new_n6604);
not_10 g04256(new_n6603, new_n6605);
xnor_4 g04257(new_n6605, new_n4704, new_n6606);
xor_4  g04258(new_n6583, new_n6571, new_n6607);
nand_5 g04259(new_n6607, new_n4711, new_n6608);
xor_4  g04260(new_n6607, new_n4711, new_n6609);
not_10 g04261(new_n6609, new_n6610);
xnor_4 g04262(new_n6574, new_n6572, new_n6611_1);
not_10 g04263(new_n6611_1, new_n6612_1);
nor_5  g04264(new_n6612_1, new_n4720, new_n6613);
not_10 g04265(new_n6613, new_n6614);
nand_5 g04266(new_n6614, new_n4717, new_n6615);
xor_4  g04267(new_n6581, new_n6580, new_n6616);
xnor_4 g04268(new_n6613, new_n4717, new_n6617);
nand_5 g04269(new_n6617, new_n6616, new_n6618);
and_5  g04270(new_n6618, new_n6615, new_n6619);
or_5   g04271(new_n6619, new_n6610, new_n6620);
nand_5 g04272(new_n6620, new_n6608, new_n6621);
nand_5 g04273(new_n6621, new_n6606, new_n6622);
nand_5 g04274(new_n6622, new_n6604, new_n6623);
nand_5 g04275(new_n6623, new_n6602, new_n6624);
and_5  g04276(new_n6624, new_n6601, new_n6625);
or_5   g04277(new_n6625, new_n6598, new_n6626);
and_5  g04278(new_n6626, new_n6596_1, new_n6627);
xor_4  g04279(new_n6627, new_n6594, n597);
not_10 g04280(new_n5859, new_n6629);
not_10 g04281(n14230, new_n6630_1);
xor_4  g04282(n25926, n9646, new_n6631_1);
xor_4  g04283(new_n6631_1, new_n6630_1, new_n6632);
xor_4  g04284(new_n6632, new_n6629, n637);
not_10 g04285(n7421, new_n6634_1);
xnor_4 g04286(n25797, n10611, new_n6635);
or_5   g04287(n15967, n2783, new_n6636);
xnor_4 g04288(n15967, n2783, new_n6637);
or_5   g04289(n15490, n13319, new_n6638);
nand_5 g04290(n25435, n18, new_n6639);
xor_4  g04291(n15490, n13319, new_n6640);
nand_5 g04292(new_n6640, new_n6639, new_n6641);
and_5  g04293(new_n6641, new_n6638, new_n6642);
or_5   g04294(new_n6642, new_n6637, new_n6643);
and_5  g04295(new_n6643, new_n6636, new_n6644);
xor_4  g04296(new_n6644, new_n6635, new_n6645);
xor_4  g04297(new_n6645, new_n6634_1, new_n6646);
not_10 g04298(new_n6646, new_n6647);
not_10 g04299(n19680, new_n6648);
xor_4  g04300(new_n6642, new_n6637, new_n6649);
or_5   g04301(new_n6649, new_n6648, new_n6650);
xor_4  g04302(new_n6649, new_n6648, new_n6651);
not_10 g04303(n2809, new_n6652_1);
xor_4  g04304(new_n6640, new_n6639, new_n6653);
nand_5 g04305(new_n6653, new_n6652_1, new_n6654);
xor_4  g04306(n25435, n18, new_n6655_1);
and_5  g04307(new_n6655_1, n15508, new_n6656);
not_10 g04308(new_n6656, new_n6657);
xor_4  g04309(new_n6653, new_n6652_1, new_n6658);
nand_5 g04310(new_n6658, new_n6657, new_n6659_1);
and_5  g04311(new_n6659_1, new_n6654, new_n6660);
nand_5 g04312(new_n6660, new_n6651, new_n6661);
and_5  g04313(new_n6661, new_n6650, new_n6662);
xor_4  g04314(new_n6662, new_n6647, new_n6663);
not_10 g04315(n20250, new_n6664);
xnor_4 g04316(n18157, n11056, new_n6665);
or_5   g04317(n15271, n12161, new_n6666);
xnor_4 g04318(n15271, n12161, new_n6667);
or_5   g04319(n25877, n5026, new_n6668);
nand_5 g04320(n24323, n8581, new_n6669_1);
xor_4  g04321(n25877, n5026, new_n6670);
nand_5 g04322(new_n6670, new_n6669_1, new_n6671_1);
and_5  g04323(new_n6671_1, new_n6668, new_n6672);
or_5   g04324(new_n6672, new_n6667, new_n6673_1);
and_5  g04325(new_n6673_1, new_n6666, new_n6674_1);
xor_4  g04326(new_n6674_1, new_n6665, new_n6675);
xor_4  g04327(new_n6675, new_n6664, new_n6676);
not_10 g04328(new_n6676, new_n6677);
xor_4  g04329(new_n6672, new_n6667, new_n6678);
nand_5 g04330(new_n6678, new_n4377, new_n6679);
xor_4  g04331(new_n6670, new_n6669_1, new_n6680);
and_5  g04332(new_n6680, new_n4382, new_n6681);
xor_4  g04333(n24323, n8581, new_n6682);
nand_5 g04334(new_n6682, n1681, new_n6683);
xor_4  g04335(new_n6680, new_n4382, new_n6684_1);
and_5  g04336(new_n6684_1, new_n6683, new_n6685);
or_5   g04337(new_n6685, new_n6681, new_n6686);
xor_4  g04338(new_n6678, new_n4377, new_n6687);
nand_5 g04339(new_n6687, new_n6686, new_n6688);
and_5  g04340(new_n6688, new_n6679, new_n6689);
xor_4  g04341(new_n6689, new_n6677, new_n6690);
xor_4  g04342(new_n6690, new_n6663, new_n6691_1);
xor_4  g04343(new_n6660, new_n6651, new_n6692);
xor_4  g04344(new_n6687, new_n6686, new_n6693);
nor_5  g04345(new_n6693, new_n6692, new_n6694);
xor_4  g04346(new_n6693, new_n6692, new_n6695);
xor_4  g04347(new_n6658, new_n6657, new_n6696);
not_10 g04348(new_n6696, new_n6697);
xor_4  g04349(new_n6684_1, new_n6683, new_n6698);
nand_5 g04350(new_n6698, new_n6697, new_n6699);
xor_4  g04351(new_n6655_1, n15508, new_n6700);
not_10 g04352(new_n6700, new_n6701);
xor_4  g04353(new_n6682, n1681, new_n6702);
nor_5  g04354(new_n6702, new_n6701, new_n6703);
xor_4  g04355(new_n6698, new_n6697, new_n6704);
nand_5 g04356(new_n6704, new_n6703, new_n6705);
and_5  g04357(new_n6705, new_n6699, new_n6706_1);
and_5  g04358(new_n6706_1, new_n6695, new_n6707_1);
nor_5  g04359(new_n6707_1, new_n6694, new_n6708);
xnor_4 g04360(new_n6708, new_n6691_1, n646);
nor_5  g04361(n19494, n2387, new_n6710);
and_5  g04362(new_n6710, new_n2363_1, new_n6711);
and_5  g04363(new_n6711, new_n2358, new_n6712);
xor_4  g04364(new_n6712, new_n2354, new_n6713);
xor_4  g04365(new_n2461, new_n5500, new_n6714);
nand_5 g04366(new_n2466, n7731, new_n6715);
xor_4  g04367(new_n2466, new_n5504, new_n6716);
nand_5 g04368(new_n2472, n12341, new_n6717);
xor_4  g04369(new_n2472, n12341, new_n6718);
and_5  g04370(new_n2475, new_n5516, new_n6719);
nand_5 g04371(new_n6719, new_n5511, new_n6720);
xor_4  g04372(new_n6719, new_n5511, new_n6721);
nand_5 g04373(new_n6721, new_n2478, new_n6722);
and_5  g04374(new_n6722, new_n6720, new_n6723);
nand_5 g04375(new_n6723, new_n6718, new_n6724);
and_5  g04376(new_n6724, new_n6717, new_n6725);
or_5   g04377(new_n6725, new_n6716, new_n6726);
and_5  g04378(new_n6726, new_n6715, new_n6727);
xor_4  g04379(new_n6727, new_n6714, new_n6728);
xnor_4 g04380(new_n6728, new_n6713, new_n6729_1);
xor_4  g04381(new_n6711, new_n2358, new_n6730);
xor_4  g04382(new_n6725, new_n6716, new_n6731);
nand_5 g04383(new_n6731, new_n6730, new_n6732);
not_10 g04384(new_n6731, new_n6733);
xor_4  g04385(new_n6733, new_n6730, new_n6734);
xor_4  g04386(new_n2475, new_n5516, new_n6735);
not_10 g04387(new_n6735, new_n6736_1);
and_5  g04388(new_n6736_1, n2387, new_n6737);
nand_5 g04389(new_n6737, new_n2365, new_n6738);
xnor_4 g04390(new_n6721, new_n2478, new_n6739);
xor_4  g04391(n19494, n2387, new_n6740);
or_5   g04392(new_n6740, new_n6737, new_n6741);
and_5  g04393(new_n6741, new_n6738, new_n6742);
nand_5 g04394(new_n6742, new_n6739, new_n6743);
nand_5 g04395(new_n6743, new_n6738, new_n6744);
xor_4  g04396(new_n6710, new_n2363_1, new_n6745);
nand_5 g04397(new_n6745, new_n6744, new_n6746);
xor_4  g04398(new_n6723, new_n6718, new_n6747);
xor_4  g04399(new_n6745, new_n6744, new_n6748);
nand_5 g04400(new_n6748, new_n6747, new_n6749);
and_5  g04401(new_n6749, new_n6746, new_n6750);
or_5   g04402(new_n6750, new_n6734, new_n6751);
and_5  g04403(new_n6751, new_n6732, new_n6752);
xor_4  g04404(new_n6752, new_n6729_1, new_n6753);
xnor_4 g04405(new_n6753, new_n3351, new_n6754);
xor_4  g04406(new_n6750, new_n6734, new_n6755);
or_5   g04407(new_n6755, new_n3359, new_n6756);
xor_4  g04408(new_n6748, new_n6747, new_n6757);
and_5  g04409(new_n6757, new_n3365, new_n6758);
xor_4  g04410(new_n6757, new_n3365, new_n6759);
xor_4  g04411(new_n6736_1, n2387, new_n6760);
and_5  g04412(new_n6760, new_n3367, new_n6761);
nor_5  g04413(new_n6761, new_n3371, new_n6762);
xnor_4 g04414(new_n6742, new_n6739, new_n6763);
and_5  g04415(new_n6761, new_n3297, new_n6764);
nor_5  g04416(new_n6764, new_n6762, new_n6765);
and_5  g04417(new_n6765, new_n6763, new_n6766);
nor_5  g04418(new_n6766, new_n6762, new_n6767);
and_5  g04419(new_n6767, new_n6759, new_n6768);
or_5   g04420(new_n6768, new_n6758, new_n6769);
xnor_4 g04421(new_n6755, new_n3357, new_n6770);
not_10 g04422(new_n6770, new_n6771);
or_5   g04423(new_n6771, new_n6769, new_n6772);
and_5  g04424(new_n6772, new_n6756, new_n6773_1);
xor_4  g04425(new_n6773_1, new_n6754, n696);
xnor_4 g04426(n25475, n23697, new_n6775_1);
or_5   g04427(n23849, n2289, new_n6776);
xnor_4 g04428(n23849, n2289, new_n6777);
or_5   g04429(n12446, n1112, new_n6778);
xnor_4 g04430(n12446, n1112, new_n6779);
or_5   g04431(n20179, n11011, new_n6780);
xnor_4 g04432(n20179, n11011, new_n6781);
or_5   g04433(n19228, n16029, new_n6782);
xnor_4 g04434(n19228, n16029, new_n6783);
or_5   g04435(n16476, n15539, new_n6784);
xnor_4 g04436(n16476, n15539, new_n6785_1);
or_5   g04437(n11615, n8052, new_n6786);
xnor_4 g04438(n11615, n8052, new_n6787);
or_5   g04439(n22433, n10158, new_n6788);
nand_5 g04440(n18962, n14090, new_n6789);
xor_4  g04441(n22433, n10158, new_n6790_1);
nand_5 g04442(new_n6790_1, new_n6789, new_n6791_1);
and_5  g04443(new_n6791_1, new_n6788, new_n6792);
or_5   g04444(new_n6792, new_n6787, new_n6793);
and_5  g04445(new_n6793, new_n6786, new_n6794_1);
or_5   g04446(new_n6794_1, new_n6785_1, new_n6795);
and_5  g04447(new_n6795, new_n6784, new_n6796);
or_5   g04448(new_n6796, new_n6783, new_n6797);
and_5  g04449(new_n6797, new_n6782, new_n6798);
or_5   g04450(new_n6798, new_n6781, new_n6799);
and_5  g04451(new_n6799, new_n6780, new_n6800);
or_5   g04452(new_n6800, new_n6779, new_n6801);
and_5  g04453(new_n6801, new_n6778, new_n6802_1);
or_5   g04454(new_n6802_1, new_n6777, new_n6803);
and_5  g04455(new_n6803, new_n6776, new_n6804);
xor_4  g04456(new_n6804, new_n6775_1, new_n6805);
xor_4  g04457(new_n6805, new_n5541, new_n6806);
not_10 g04458(new_n6806, new_n6807);
xor_4  g04459(new_n6802_1, new_n6777, new_n6808);
or_5   g04460(new_n6808, new_n5545, new_n6809);
xor_4  g04461(new_n6808, n9655, new_n6810);
xor_4  g04462(new_n6800, new_n6779, new_n6811);
or_5   g04463(new_n6811, new_n5549, new_n6812);
xor_4  g04464(new_n6811, n13490, new_n6813);
xor_4  g04465(new_n6798, new_n6781, new_n6814_1);
or_5   g04466(new_n6814_1, new_n5553, new_n6815);
xor_4  g04467(new_n6796, new_n6783, new_n6816);
nand_5 g04468(new_n6816, new_n5557, new_n6817);
xor_4  g04469(new_n6816, new_n5557, new_n6818);
not_10 g04470(new_n6818, new_n6819);
xor_4  g04471(new_n6794_1, new_n6785_1, new_n6820);
nand_5 g04472(new_n6820, new_n5561, new_n6821);
xor_4  g04473(new_n6820, new_n5561, new_n6822);
not_10 g04474(n15636, new_n6823);
xor_4  g04475(new_n6792, new_n6787, new_n6824);
or_5   g04476(new_n6824, new_n6823, new_n6825);
xor_4  g04477(new_n6824, new_n6823, new_n6826_1);
xor_4  g04478(n18962, n14090, new_n6827);
and_5  g04479(new_n6827, n6794, new_n6828);
or_5   g04480(new_n6828, n20077, new_n6829);
xor_4  g04481(new_n6790_1, new_n6789, new_n6830);
xor_4  g04482(new_n6828, n20077, new_n6831);
nand_5 g04483(new_n6831, new_n6830, new_n6832);
and_5  g04484(new_n6832, new_n6829, new_n6833);
nand_5 g04485(new_n6833, new_n6826_1, new_n6834);
and_5  g04486(new_n6834, new_n6825, new_n6835_1);
nand_5 g04487(new_n6835_1, new_n6822, new_n6836);
and_5  g04488(new_n6836, new_n6821, new_n6837);
or_5   g04489(new_n6837, new_n6819, new_n6838);
and_5  g04490(new_n6838, new_n6817, new_n6839);
xor_4  g04491(new_n6814_1, new_n5553, new_n6840);
nand_5 g04492(new_n6840, new_n6839, new_n6841);
and_5  g04493(new_n6841, new_n6815, new_n6842);
or_5   g04494(new_n6842, new_n6813, new_n6843);
and_5  g04495(new_n6843, new_n6812, new_n6844);
or_5   g04496(new_n6844, new_n6810, new_n6845);
and_5  g04497(new_n6845, new_n6809, new_n6846);
xor_4  g04498(new_n6846, new_n6807, new_n6847);
xor_4  g04499(n21915, n15182, new_n6848);
not_10 g04500(new_n6848, new_n6849);
or_5   g04501(n27037, n13775, new_n6850);
xor_4  g04502(n27037, n13775, new_n6851);
not_10 g04503(new_n6851, new_n6852);
or_5   g04504(n8964, n1293, new_n6853_1);
xor_4  g04505(n8964, n1293, new_n6854);
not_10 g04506(new_n6854, new_n6855);
or_5   g04507(n20151, n19042, new_n6856);
xor_4  g04508(n20151, n19042, new_n6857);
not_10 g04509(new_n6857, new_n6858);
or_5   g04510(n19472, n7693, new_n6859);
xor_4  g04511(n19472, n7693, new_n6860);
nand_5 g04512(n25370, n10405, new_n6861_1);
or_5   g04513(n25370, n10405, new_n6862_1);
nor_5  g04514(n24786, n11302, new_n6863_1);
nor_5  g04515(new_n4119_1, new_n4114, new_n6864);
nor_5  g04516(new_n6864, new_n6863_1, new_n6865);
nand_5 g04517(new_n6865, new_n6862_1, new_n6866);
and_5  g04518(new_n6866, new_n6861_1, new_n6867_1);
nand_5 g04519(new_n6867_1, new_n6860, new_n6868);
and_5  g04520(new_n6868, new_n6859, new_n6869);
or_5   g04521(new_n6869, new_n6858, new_n6870);
and_5  g04522(new_n6870, new_n6856, new_n6871);
or_5   g04523(new_n6871, new_n6855, new_n6872);
and_5  g04524(new_n6872, new_n6853_1, new_n6873);
or_5   g04525(new_n6873, new_n6852, new_n6874);
and_5  g04526(new_n6874, new_n6850, new_n6875);
xor_4  g04527(new_n6875, new_n6849, new_n6876);
not_10 g04528(new_n6876, new_n6877);
xor_4  g04529(new_n6877, new_n5484, new_n6878);
xor_4  g04530(new_n6873, new_n6852, new_n6879);
not_10 g04531(new_n6879, new_n6880);
nand_5 g04532(new_n6880, n11736, new_n6881);
xor_4  g04533(new_n6880, n11736, new_n6882);
not_10 g04534(new_n6882, new_n6883);
xor_4  g04535(new_n6871, new_n6855, new_n6884);
not_10 g04536(new_n6884, new_n6885);
nand_5 g04537(new_n6885, n23200, new_n6886);
xor_4  g04538(new_n6885, n23200, new_n6887);
not_10 g04539(new_n6887, new_n6888);
xor_4  g04540(new_n6869, new_n6858, new_n6889);
not_10 g04541(new_n6889, new_n6890);
nand_5 g04542(new_n6890, n17959, new_n6891);
xor_4  g04543(new_n6890, n17959, new_n6892);
not_10 g04544(new_n6892, new_n6893);
xor_4  g04545(new_n6867_1, new_n6860, new_n6894);
not_10 g04546(new_n6894, new_n6895);
nand_5 g04547(new_n6895, n7566, new_n6896);
xor_4  g04548(new_n6895, new_n5500, new_n6897);
xor_4  g04549(n25370, n10405, new_n6898);
xor_4  g04550(new_n6898, new_n6865, new_n6899);
not_10 g04551(new_n6899, new_n6900);
or_5   g04552(new_n6900, new_n5504, new_n6901);
xor_4  g04553(new_n6900, n7731, new_n6902);
or_5   g04554(new_n4120, new_n5509, new_n6903);
and_5  g04555(new_n4131, new_n5511, new_n6904);
and_5  g04556(new_n4135, n12384, new_n6905);
not_10 g04557(new_n6905, new_n6906);
xor_4  g04558(new_n4131, new_n5511, new_n6907);
and_5  g04559(new_n6907, new_n6906, new_n6908);
nor_5  g04560(new_n6908, new_n6904, new_n6909);
xor_4  g04561(new_n4120, new_n5509, new_n6910);
nand_5 g04562(new_n6910, new_n6909, new_n6911);
and_5  g04563(new_n6911, new_n6903, new_n6912);
or_5   g04564(new_n6912, new_n6902, new_n6913);
and_5  g04565(new_n6913, new_n6901, new_n6914);
or_5   g04566(new_n6914, new_n6897, new_n6915);
and_5  g04567(new_n6915, new_n6896, new_n6916);
or_5   g04568(new_n6916, new_n6893, new_n6917);
and_5  g04569(new_n6917, new_n6891, new_n6918);
or_5   g04570(new_n6918, new_n6888, new_n6919);
and_5  g04571(new_n6919, new_n6886, new_n6920);
or_5   g04572(new_n6920, new_n6883, new_n6921);
and_5  g04573(new_n6921, new_n6881, new_n6922);
xor_4  g04574(new_n6922, new_n6878, new_n6923);
xnor_4 g04575(new_n6923, new_n6847, new_n6924);
not_10 g04576(new_n6924, new_n6925);
xor_4  g04577(new_n6920, new_n6883, new_n6926);
not_10 g04578(new_n6926, new_n6927);
xor_4  g04579(new_n6844, new_n6810, new_n6928);
and_5  g04580(new_n6928, new_n6927, new_n6929);
not_10 g04581(new_n6929, new_n6930);
xor_4  g04582(new_n6928, new_n6927, new_n6931);
xor_4  g04583(new_n6918, new_n6888, new_n6932);
not_10 g04584(new_n6932, new_n6933);
xor_4  g04585(new_n6842, new_n6813, new_n6934);
and_5  g04586(new_n6934, new_n6933, new_n6935);
not_10 g04587(new_n6935, new_n6936);
xor_4  g04588(new_n6934, new_n6933, new_n6937);
xnor_4 g04589(new_n6916, new_n6892, new_n6938);
not_10 g04590(new_n6938, new_n6939);
xor_4  g04591(new_n6840, new_n6839, new_n6940);
and_5  g04592(new_n6940, new_n6939, new_n6941);
not_10 g04593(new_n6941, new_n6942);
xor_4  g04594(new_n6940, new_n6939, new_n6943);
xor_4  g04595(new_n6837, new_n6819, new_n6944);
xor_4  g04596(new_n6914, new_n6897, new_n6945);
nor_5  g04597(new_n6945, new_n6944, new_n6946);
xor_4  g04598(new_n6945, new_n6944, new_n6947);
not_10 g04599(new_n6947, new_n6948);
xor_4  g04600(new_n6835_1, new_n6822, new_n6949);
xor_4  g04601(new_n6912, new_n6902, new_n6950);
nor_5  g04602(new_n6950, new_n6949, new_n6951);
xor_4  g04603(new_n6950, new_n6949, new_n6952);
not_10 g04604(new_n6952, new_n6953);
xor_4  g04605(new_n6910, new_n6909, new_n6954);
not_10 g04606(new_n6954, new_n6955);
xor_4  g04607(new_n6833, new_n6826_1, new_n6956);
and_5  g04608(new_n6956, new_n6955, new_n6957);
not_10 g04609(new_n6957, new_n6958);
not_10 g04610(new_n6956, new_n6959);
xnor_4 g04611(new_n6959, new_n6955, new_n6960);
xor_4  g04612(new_n6907, new_n6906, new_n6961);
not_10 g04613(new_n6961, new_n6962);
xor_4  g04614(new_n6831, new_n6830, new_n6963);
nor_5  g04615(new_n6963, new_n6962, new_n6964);
not_10 g04616(new_n6964, new_n6965_1);
xor_4  g04617(new_n6827, n6794, new_n6966);
not_10 g04618(new_n6966, new_n6967_1);
xor_4  g04619(new_n4135, n12384, new_n6968);
nor_5  g04620(new_n6968, new_n6967_1, new_n6969);
xor_4  g04621(new_n6963, new_n6962, new_n6970);
and_5  g04622(new_n6970, new_n6969, new_n6971_1);
not_10 g04623(new_n6971_1, new_n6972);
and_5  g04624(new_n6972, new_n6965_1, new_n6973);
not_10 g04625(new_n6973, new_n6974);
and_5  g04626(new_n6974, new_n6960, new_n6975_1);
not_10 g04627(new_n6975_1, new_n6976);
and_5  g04628(new_n6976, new_n6958, new_n6977);
nor_5  g04629(new_n6977, new_n6953, new_n6978);
nor_5  g04630(new_n6978, new_n6951, new_n6979);
nor_5  g04631(new_n6979, new_n6948, new_n6980);
nor_5  g04632(new_n6980, new_n6946, new_n6981);
not_10 g04633(new_n6981, new_n6982);
and_5  g04634(new_n6982, new_n6943, new_n6983_1);
not_10 g04635(new_n6983_1, new_n6984);
and_5  g04636(new_n6984, new_n6942, new_n6985_1);
not_10 g04637(new_n6985_1, new_n6986);
and_5  g04638(new_n6986, new_n6937, new_n6987);
not_10 g04639(new_n6987, new_n6988);
and_5  g04640(new_n6988, new_n6936, new_n6989);
not_10 g04641(new_n6989, new_n6990);
and_5  g04642(new_n6990, new_n6931, new_n6991);
not_10 g04643(new_n6991, new_n6992);
and_5  g04644(new_n6992, new_n6930, new_n6993);
xnor_4 g04645(new_n6993, new_n6925, n723);
xnor_4 g04646(n26986, n2272, new_n6995);
not_10 g04647(new_n6995, new_n6996);
not_10 g04648(n21287, new_n6997);
nand_5 g04649(n25331, new_n6997, new_n6998_1);
xnor_4 g04650(n25331, n21287, new_n6999);
not_10 g04651(new_n6999, new_n7000);
not_10 g04652(n4256, new_n7001);
nand_5 g04653(n18483, new_n7001, new_n7002);
xnor_4 g04654(n18483, n4256, new_n7003);
not_10 g04655(new_n7003, new_n7004);
not_10 g04656(n22332, new_n7005);
nand_5 g04657(new_n7005, n21934, new_n7006);
xnor_4 g04658(n22332, n21934, new_n7007);
not_10 g04659(new_n7007, new_n7008);
nand_5 g04660(new_n3806, n18901, new_n7009);
xnor_4 g04661(n18907, n18901, new_n7010);
not_10 g04662(new_n7010, new_n7011);
nand_5 g04663(n4376, new_n3810, new_n7012);
xnor_4 g04664(n4376, n2731, new_n7013);
not_10 g04665(new_n7013, new_n7014);
nand_5 g04666(new_n3814, n14570, new_n7015);
xnor_4 g04667(n19911, n14570, new_n7016);
or_5   g04668(n23775, new_n3819, new_n7017);
nand_5 g04669(n23775, new_n3819, new_n7018);
nor_5  g04670(new_n3821, n8259, new_n7019);
and_5  g04671(new_n3821, n8259, new_n7020);
not_10 g04672(new_n7020, new_n7021);
not_10 g04673(n11479, new_n7022);
and_5  g04674(new_n7022, n5704, new_n7023);
and_5  g04675(new_n7023, new_n7021, new_n7024);
nor_5  g04676(new_n7024, new_n7019, new_n7025);
not_10 g04677(new_n7025, new_n7026_1);
nand_5 g04678(new_n7026_1, new_n7018, new_n7027);
and_5  g04679(new_n7027, new_n7017, new_n7028);
nand_5 g04680(new_n7028, new_n7016, new_n7029);
and_5  g04681(new_n7029, new_n7015, new_n7030);
or_5   g04682(new_n7030, new_n7014, new_n7031);
and_5  g04683(new_n7031, new_n7012, new_n7032_1);
or_5   g04684(new_n7032_1, new_n7011, new_n7033);
and_5  g04685(new_n7033, new_n7009, new_n7034);
or_5   g04686(new_n7034, new_n7008, new_n7035);
and_5  g04687(new_n7035, new_n7006, new_n7036);
or_5   g04688(new_n7036, new_n7004, new_n7037);
and_5  g04689(new_n7037, new_n7002, new_n7038_1);
or_5   g04690(new_n7038_1, new_n7000, new_n7039);
and_5  g04691(new_n7039, new_n6998_1, new_n7040);
xor_4  g04692(new_n7040, new_n6996, new_n7041);
not_10 g04693(new_n7041, new_n7042);
xor_4  g04694(n1255, n468, new_n7043);
not_10 g04695(new_n7043, new_n7044);
or_5   g04696(n9512, n5400, new_n7045);
xor_4  g04697(n9512, n5400, new_n7046);
not_10 g04698(new_n7046, new_n7047);
or_5   g04699(n23923, n16608, new_n7048);
xnor_4 g04700(n23923, n16608, new_n7049);
or_5   g04701(n21735, n329, new_n7050);
xnor_4 g04702(n21735, n329, new_n7051);
or_5   g04703(n24170, n24085, new_n7052);
xnor_4 g04704(n24170, n24085, new_n7053);
or_5   g04705(n14071, n2409, new_n7054);
xnor_4 g04706(n14071, n2409, new_n7055);
or_5   g04707(n8869, n1738, new_n7056);
xnor_4 g04708(n8869, n1738, new_n7057_1);
or_5   g04709(n12152, n10372, new_n7058);
nand_5 g04710(n19107, n7428, new_n7059);
xor_4  g04711(n12152, n10372, new_n7060);
nand_5 g04712(new_n7060, new_n7059, new_n7061);
and_5  g04713(new_n7061, new_n7058, new_n7062);
or_5   g04714(new_n7062, new_n7057_1, new_n7063);
and_5  g04715(new_n7063, new_n7056, new_n7064);
or_5   g04716(new_n7064, new_n7055, new_n7065);
and_5  g04717(new_n7065, new_n7054, new_n7066);
or_5   g04718(new_n7066, new_n7053, new_n7067);
and_5  g04719(new_n7067, new_n7052, new_n7068);
or_5   g04720(new_n7068, new_n7051, new_n7069);
and_5  g04721(new_n7069, new_n7050, new_n7070);
or_5   g04722(new_n7070, new_n7049, new_n7071);
and_5  g04723(new_n7071, new_n7048, new_n7072);
or_5   g04724(new_n7072, new_n7047, new_n7073);
and_5  g04725(new_n7073, new_n7045, new_n7074);
xor_4  g04726(new_n7074, new_n7044, new_n7075);
not_10 g04727(new_n7075, new_n7076);
xnor_4 g04728(n14130, n12861, new_n7077);
or_5   g04729(n16482, n13333, new_n7078);
xnor_4 g04730(n16482, n13333, new_n7079_1);
or_5   g04731(n9942, n2210, new_n7080);
xor_4  g04732(n9942, n2210, new_n7081);
not_10 g04733(new_n7081, new_n7082);
or_5   g04734(n25643, n20604, new_n7083);
or_5   g04735(new_n5139, new_n5136, new_n7084);
and_5  g04736(new_n7084, new_n7083, new_n7085);
or_5   g04737(new_n7085, new_n7082, new_n7086);
and_5  g04738(new_n7086, new_n7080, new_n7087);
or_5   g04739(new_n7087, new_n7079_1, new_n7088);
and_5  g04740(new_n7088, new_n7078, new_n7089);
xor_4  g04741(new_n7089, new_n7077, new_n7090);
nor_5  g04742(new_n7090, new_n7076, new_n7091);
xor_4  g04743(new_n7090, new_n7075, new_n7092);
xor_4  g04744(new_n7072, new_n7047, new_n7093);
not_10 g04745(new_n7093, new_n7094);
xor_4  g04746(new_n7087, new_n7079_1, new_n7095);
or_5   g04747(new_n7095, new_n7094, new_n7096);
xor_4  g04748(new_n7095, new_n7093, new_n7097);
xor_4  g04749(new_n7085, new_n7082, new_n7098);
not_10 g04750(new_n7098, new_n7099_1);
xor_4  g04751(new_n7070, new_n7049, new_n7100);
nand_5 g04752(new_n7100, new_n7099_1, new_n7101);
xor_4  g04753(new_n7100, new_n7099_1, new_n7102);
not_10 g04754(new_n7102, new_n7103);
xor_4  g04755(new_n7068, new_n7051, new_n7104);
nand_5 g04756(new_n7104, new_n5141, new_n7105);
xnor_4 g04757(new_n7104, new_n5141, new_n7106);
xor_4  g04758(new_n7066, new_n7053, new_n7107);
nand_5 g04759(new_n7107, new_n5145, new_n7108);
xnor_4 g04760(new_n7107, new_n5145, new_n7109);
xor_4  g04761(new_n7064, new_n7055, new_n7110);
nand_5 g04762(new_n7110, new_n5150, new_n7111);
xor_4  g04763(new_n7110, new_n5150, new_n7112);
xor_4  g04764(new_n7062, new_n7057_1, new_n7113);
nand_5 g04765(new_n7113, new_n5119, new_n7114);
xnor_4 g04766(new_n7113, new_n5119, new_n7115);
xor_4  g04767(new_n7060, new_n7059, new_n7116);
nand_5 g04768(new_n7116, new_n5110, new_n7117);
xnor_4 g04769(n19107, n7428, new_n7118);
and_5  g04770(new_n7118, new_n5107, new_n7119);
xor_4  g04771(new_n7116, new_n5110, new_n7120);
nand_5 g04772(new_n7120, new_n7119, new_n7121);
and_5  g04773(new_n7121, new_n7117, new_n7122);
or_5   g04774(new_n7122, new_n7115, new_n7123);
nand_5 g04775(new_n7123, new_n7114, new_n7124);
nand_5 g04776(new_n7124, new_n7112, new_n7125);
and_5  g04777(new_n7125, new_n7111, new_n7126);
or_5   g04778(new_n7126, new_n7109, new_n7127);
and_5  g04779(new_n7127, new_n7108, new_n7128);
or_5   g04780(new_n7128, new_n7106, new_n7129);
and_5  g04781(new_n7129, new_n7105, new_n7130);
or_5   g04782(new_n7130, new_n7103, new_n7131);
and_5  g04783(new_n7131, new_n7101, new_n7132);
or_5   g04784(new_n7132, new_n7097, new_n7133);
and_5  g04785(new_n7133, new_n7096, new_n7134);
nor_5  g04786(new_n7134, new_n7092, new_n7135);
or_5   g04787(new_n7135, new_n7091, new_n7136);
xor_4  g04788(n22442, n22253, new_n7137);
or_5   g04789(n1255, n468, new_n7138);
or_5   g04790(new_n7074, new_n7044, new_n7139_1);
and_5  g04791(new_n7139_1, new_n7138, new_n7140);
xor_4  g04792(new_n7140, new_n7137, new_n7141);
xnor_4 g04793(n8856, n8305, new_n7142);
or_5   g04794(n14130, n12861, new_n7143);
or_5   g04795(new_n7089, new_n7077, new_n7144);
and_5  g04796(new_n7144, new_n7143, new_n7145);
xor_4  g04797(new_n7145, new_n7142, new_n7146);
xor_4  g04798(new_n7146, new_n7141, new_n7147);
xor_4  g04799(new_n7147, new_n7136, new_n7148);
and_5  g04800(new_n7148, new_n7042, new_n7149_1);
xor_4  g04801(new_n7148, new_n7042, new_n7150);
not_10 g04802(new_n7150, new_n7151);
xor_4  g04803(new_n7038_1, new_n7000, new_n7152);
not_10 g04804(new_n7152, new_n7153);
xor_4  g04805(new_n7134, new_n7092, new_n7154);
and_5  g04806(new_n7154, new_n7153, new_n7155);
xor_4  g04807(new_n7154, new_n7153, new_n7156);
not_10 g04808(new_n7156, new_n7157);
xor_4  g04809(new_n7036, new_n7004, new_n7158);
not_10 g04810(new_n7158, new_n7159);
xor_4  g04811(new_n7132, new_n7097, new_n7160);
and_5  g04812(new_n7160, new_n7159, new_n7161);
xor_4  g04813(new_n7160, new_n7159, new_n7162);
not_10 g04814(new_n7162, new_n7163);
xor_4  g04815(new_n7034, new_n7008, new_n7164);
xnor_4 g04816(new_n7130, new_n7102, new_n7165);
not_10 g04817(new_n7165, new_n7166);
nor_5  g04818(new_n7166, new_n7164, new_n7167);
xor_4  g04819(new_n7166, new_n7164, new_n7168);
xor_4  g04820(new_n7032_1, new_n7011, new_n7169);
not_10 g04821(new_n7169, new_n7170);
xor_4  g04822(new_n7128, new_n7106, new_n7171);
and_5  g04823(new_n7171, new_n7170, new_n7172);
xor_4  g04824(new_n7171, new_n7170, new_n7173);
not_10 g04825(new_n7173, new_n7174);
xor_4  g04826(new_n7030, new_n7014, new_n7175);
not_10 g04827(new_n7175, new_n7176);
xor_4  g04828(new_n7126, new_n7109, new_n7177);
and_5  g04829(new_n7177, new_n7176, new_n7178);
xor_4  g04830(new_n7177, new_n7176, new_n7179);
not_10 g04831(new_n7179, new_n7180);
xor_4  g04832(new_n7124, new_n7112, new_n7181);
not_10 g04833(new_n7181, new_n7182);
xor_4  g04834(new_n7028, new_n7016, new_n7183);
nor_5  g04835(new_n7183, new_n7182, new_n7184);
not_10 g04836(new_n7184, new_n7185);
xor_4  g04837(new_n7122, new_n7115, new_n7186);
xnor_4 g04838(n23775, n13708, new_n7187);
xor_4  g04839(new_n7187, new_n7026_1, new_n7188);
and_5  g04840(new_n7188, new_n7186, new_n7189);
not_10 g04841(new_n7189, new_n7190_1);
xor_4  g04842(new_n7188, new_n7186, new_n7191);
xor_4  g04843(new_n7118, new_n5107, new_n7192);
xnor_4 g04844(n11479, n5704, new_n7193);
or_5   g04845(new_n7193, new_n7192, new_n7194);
xnor_4 g04846(n18409, n8259, new_n7195);
xor_4  g04847(new_n7195, new_n7023, new_n7196);
nor_5  g04848(new_n7196, new_n7194, new_n7197);
xnor_4 g04849(new_n7120, new_n7119, new_n7198);
xor_4  g04850(new_n7196, new_n7194, new_n7199);
and_5  g04851(new_n7199, new_n7198, new_n7200);
nor_5  g04852(new_n7200, new_n7197, new_n7201);
and_5  g04853(new_n7201, new_n7191, new_n7202);
not_10 g04854(new_n7202, new_n7203);
and_5  g04855(new_n7203, new_n7190_1, new_n7204);
not_10 g04856(new_n7204, new_n7205);
xor_4  g04857(new_n7183, new_n7182, new_n7206);
and_5  g04858(new_n7206, new_n7205, new_n7207);
not_10 g04859(new_n7207, new_n7208);
and_5  g04860(new_n7208, new_n7185, new_n7209);
nor_5  g04861(new_n7209, new_n7180, new_n7210);
nor_5  g04862(new_n7210, new_n7178, new_n7211);
nor_5  g04863(new_n7211, new_n7174, new_n7212);
nor_5  g04864(new_n7212, new_n7172, new_n7213);
not_10 g04865(new_n7213, new_n7214);
and_5  g04866(new_n7214, new_n7168, new_n7215);
nor_5  g04867(new_n7215, new_n7167, new_n7216);
nor_5  g04868(new_n7216, new_n7163, new_n7217);
nor_5  g04869(new_n7217, new_n7161, new_n7218);
nor_5  g04870(new_n7218, new_n7157, new_n7219);
nor_5  g04871(new_n7219, new_n7155, new_n7220);
nor_5  g04872(new_n7220, new_n7151, new_n7221);
nor_5  g04873(new_n7221, new_n7149_1, new_n7222);
not_10 g04874(n26986, new_n7223);
and_5  g04875(new_n7223, n2272, new_n7224);
not_10 g04876(new_n7224, new_n7225);
nor_5  g04877(new_n7040, new_n6996, new_n7226);
not_10 g04878(new_n7226, new_n7227);
and_5  g04879(new_n7227, new_n7225, new_n7228);
nor_5  g04880(n22442, n22253, new_n7229_1);
not_10 g04881(new_n7137, new_n7230_1);
nor_5  g04882(new_n7140, new_n7230_1, new_n7231);
or_5   g04883(new_n7231, new_n7229_1, new_n7232);
nor_5  g04884(n8856, n8305, new_n7233_1);
not_10 g04885(new_n7233_1, new_n7234);
or_5   g04886(new_n7145, new_n7142, new_n7235);
and_5  g04887(new_n7235, new_n7234, new_n7236_1);
xor_4  g04888(new_n7236_1, new_n7232, new_n7237);
or_5   g04889(new_n7146, new_n7141, new_n7238);
nand_5 g04890(new_n7147, new_n7136, new_n7239);
and_5  g04891(new_n7239, new_n7238, new_n7240);
xor_4  g04892(new_n7240, new_n7237, new_n7241);
xor_4  g04893(new_n7241, new_n7228, new_n7242);
xor_4  g04894(new_n7242, new_n7222, n735);
xor_4  g04895(n21138, n14230, new_n7244);
not_10 g04896(new_n7244, new_n7245);
xor_4  g04897(new_n6827, n19234, new_n7246);
not_10 g04898(new_n7246, new_n7247);
xor_4  g04899(new_n7247, n26167, new_n7248);
xor_4  g04900(new_n7248, new_n7245, n779);
not_10 g04901(n17458, new_n7250);
and_5  g04902(new_n7250, n8526, new_n7251);
xnor_4 g04903(n17458, n8526, new_n7252);
not_10 g04904(new_n7252, new_n7253_1);
or_5   g04905(new_n6073, n1222, new_n7254);
xnor_4 g04906(n2816, n1222, new_n7255);
not_10 g04907(new_n7255, new_n7256_1);
or_5   g04908(n25240, new_n6078, new_n7257);
xnor_4 g04909(n25240, n20359, new_n7258);
not_10 g04910(new_n7258, new_n7259);
or_5   g04911(n10125, new_n6083, new_n7260);
xor_4  g04912(n10125, n4409, new_n7261);
or_5   g04913(n8067, new_n6088, new_n7262);
xor_4  g04914(n8067, n3570, new_n7263);
or_5   g04915(n20923, new_n4220, new_n7264);
xor_4  g04916(n20923, n13668, new_n7265);
or_5   g04917(new_n4221_1, n18157, new_n7266);
xnor_4 g04918(n21276, n18157, new_n7267);
not_10 g04919(n12161, new_n7268_1);
or_5   g04920(n26748, new_n7268_1, new_n7269);
and_5  g04921(n26748, new_n7268_1, new_n7270);
and_5  g04922(new_n6103, n5026, new_n7271);
not_10 g04923(n5026, new_n7272);
and_5  g04924(n10057, new_n7272, new_n7273);
not_10 g04925(n8581, new_n7274);
or_5   g04926(n8920, new_n7274, new_n7275);
or_5   g04927(new_n7275, new_n7273, new_n7276);
not_10 g04928(new_n7276, new_n7277_1);
nor_5  g04929(new_n7277_1, new_n7271, new_n7278);
or_5   g04930(new_n7278, new_n7270, new_n7279);
and_5  g04931(new_n7279, new_n7269, new_n7280_1);
nand_5 g04932(new_n7280_1, new_n7267, new_n7281);
and_5  g04933(new_n7281, new_n7266, new_n7282);
or_5   g04934(new_n7282, new_n7265, new_n7283);
and_5  g04935(new_n7283, new_n7264, new_n7284);
or_5   g04936(new_n7284, new_n7263, new_n7285);
and_5  g04937(new_n7285, new_n7262, new_n7286);
or_5   g04938(new_n7286, new_n7261, new_n7287);
and_5  g04939(new_n7287, new_n7260, new_n7288);
or_5   g04940(new_n7288, new_n7259, new_n7289);
and_5  g04941(new_n7289, new_n7257, new_n7290);
or_5   g04942(new_n7290, new_n7256_1, new_n7291);
and_5  g04943(new_n7291, new_n7254, new_n7292);
nor_5  g04944(new_n7292, new_n7253_1, new_n7293);
nor_5  g04945(new_n7293, new_n7251, new_n7294);
not_10 g04946(n19282, new_n7295);
and_5  g04947(n26986, new_n7295, new_n7296);
xor_4  g04948(n26986, n19282, new_n7297);
or_5   g04949(new_n6997, n12657, new_n7298_1);
xor_4  g04950(n21287, n12657, new_n7299);
or_5   g04951(n17077, new_n7001, new_n7300);
xor_4  g04952(n17077, n4256, new_n7301);
or_5   g04953(n26510, new_n7005, new_n7302);
or_5   g04954(new_n3838, new_n3805, new_n7303);
and_5  g04955(new_n7303, new_n7302, new_n7304);
or_5   g04956(new_n7304, new_n7301, new_n7305_1);
and_5  g04957(new_n7305_1, new_n7300, new_n7306);
or_5   g04958(new_n7306, new_n7299, new_n7307);
and_5  g04959(new_n7307, new_n7298_1, new_n7308_1);
nor_5  g04960(new_n7308_1, new_n7297, new_n7309);
nor_5  g04961(new_n7309, new_n7296, new_n7310);
xor_4  g04962(new_n7310, new_n7294, new_n7311);
xor_4  g04963(new_n7292, new_n7253_1, new_n7312);
xor_4  g04964(new_n7308_1, new_n7297, new_n7313_1);
nand_5 g04965(new_n7313_1, new_n7312, new_n7314);
xor_4  g04966(new_n7313_1, new_n7312, new_n7315);
xor_4  g04967(new_n7290, new_n7256_1, new_n7316);
xor_4  g04968(new_n7306, new_n7299, new_n7317);
or_5   g04969(new_n7317, new_n7316, new_n7318);
xor_4  g04970(new_n7317, new_n7316, new_n7319);
not_10 g04971(new_n7319, new_n7320);
xor_4  g04972(new_n7288, new_n7259, new_n7321);
xor_4  g04973(new_n7304, new_n7301, new_n7322);
or_5   g04974(new_n7322, new_n7321, new_n7323);
xor_4  g04975(new_n7322, new_n7321, new_n7324);
not_10 g04976(new_n7324, new_n7325);
xor_4  g04977(new_n7286, new_n7261, new_n7326);
or_5   g04978(new_n7326, new_n3839, new_n7327);
xnor_4 g04979(new_n7326, new_n3840, new_n7328);
not_10 g04980(new_n7328, new_n7329);
xor_4  g04981(new_n7284, new_n7263, new_n7330_1);
or_5   g04982(new_n7330_1, new_n3854, new_n7331);
xnor_4 g04983(new_n7330_1, new_n3857, new_n7332);
not_10 g04984(new_n7332, new_n7333);
xor_4  g04985(new_n7282, new_n7265, new_n7334);
or_5   g04986(new_n7334, new_n3860, new_n7335_1);
xnor_4 g04987(new_n7334, new_n3863, new_n7336);
not_10 g04988(new_n7336, new_n7337);
xor_4  g04989(new_n7280_1, new_n7267, new_n7338);
or_5   g04990(new_n7338, new_n3867, new_n7339_1);
xor_4  g04991(new_n7338, new_n3867, new_n7340);
not_10 g04992(new_n7340, new_n7341);
xnor_4 g04993(n26748, n12161, new_n7342);
xor_4  g04994(new_n7342, new_n7278, new_n7343);
not_10 g04995(new_n7343, new_n7344);
nand_5 g04996(new_n7344, new_n3874, new_n7345);
xnor_4 g04997(new_n7343, new_n3874, new_n7346_1);
xnor_4 g04998(n10057, n5026, new_n7347);
xnor_4 g04999(new_n7347, new_n7275, new_n7348);
or_5   g05000(new_n7348, new_n3879, new_n7349_1);
xnor_4 g05001(n8920, n8581, new_n7350);
nor_5  g05002(new_n7350, new_n3882, new_n7351);
xor_4  g05003(new_n7348, new_n3879, new_n7352);
nand_5 g05004(new_n7352, new_n7351, new_n7353);
and_5  g05005(new_n7353, new_n7349_1, new_n7354);
nand_5 g05006(new_n7354, new_n7346_1, new_n7355);
and_5  g05007(new_n7355, new_n7345, new_n7356);
or_5   g05008(new_n7356, new_n7341, new_n7357);
and_5  g05009(new_n7357, new_n7339_1, new_n7358);
or_5   g05010(new_n7358, new_n7337, new_n7359);
and_5  g05011(new_n7359, new_n7335_1, new_n7360);
or_5   g05012(new_n7360, new_n7333, new_n7361);
and_5  g05013(new_n7361, new_n7331, new_n7362);
or_5   g05014(new_n7362, new_n7329, new_n7363_1);
and_5  g05015(new_n7363_1, new_n7327, new_n7364);
or_5   g05016(new_n7364, new_n7325, new_n7365);
and_5  g05017(new_n7365, new_n7323, new_n7366);
or_5   g05018(new_n7366, new_n7320, new_n7367);
and_5  g05019(new_n7367, new_n7318, new_n7368);
nand_5 g05020(new_n7368, new_n7315, new_n7369);
and_5  g05021(new_n7369, new_n7314, new_n7370);
xnor_4 g05022(new_n7370, new_n7311, new_n7371);
or_5   g05023(n11898, new_n5910, new_n7372);
xnor_4 g05024(n11898, n2979, new_n7373);
not_10 g05025(new_n7373, new_n7374);
or_5   g05026(n19941, new_n5911_1, new_n7375);
xnor_4 g05027(n19941, n647, new_n7376);
not_10 g05028(new_n7376, new_n7377_1);
or_5   g05029(new_n5912, n1099, new_n7378);
xnor_4 g05030(n20409, n1099, new_n7379);
not_10 g05031(new_n7379, new_n7380);
or_5   g05032(new_n5913, n2113, new_n7381);
xnor_4 g05033(n25749, n2113, new_n7382);
not_10 g05034(new_n7382, new_n7383);
or_5   g05035(n21134, new_n3769, new_n7384);
xnor_4 g05036(n21134, n3161, new_n7385);
not_10 g05037(new_n7385, new_n7386);
or_5   g05038(new_n3776, n6369, new_n7387);
xnor_4 g05039(n9003, n6369, new_n7388);
not_10 g05040(new_n7388, new_n7389);
or_5   g05041(n25797, new_n3778, new_n7390_1);
xnor_4 g05042(n25797, n4957, new_n7391);
or_5   g05043(new_n3729, n7524, new_n7392);
or_5   g05044(n15967, new_n3785_1, new_n7393);
not_10 g05045(n15743, new_n7394);
and_5  g05046(new_n7394, n13319, new_n7395);
nor_5  g05047(new_n7394, n13319, new_n7396);
not_10 g05048(new_n7396, new_n7397);
and_5  g05049(n25435, new_n6008, new_n7398);
and_5  g05050(new_n7398, new_n7397, new_n7399);
nor_5  g05051(new_n7399, new_n7395, new_n7400);
not_10 g05052(new_n7400, new_n7401);
nand_5 g05053(new_n7401, new_n7393, new_n7402);
and_5  g05054(new_n7402, new_n7392, new_n7403_1);
nand_5 g05055(new_n7403_1, new_n7391, new_n7404);
and_5  g05056(new_n7404, new_n7390_1, new_n7405);
or_5   g05057(new_n7405, new_n7389, new_n7406);
and_5  g05058(new_n7406, new_n7387, new_n7407);
or_5   g05059(new_n7407, new_n7386, new_n7408_1);
and_5  g05060(new_n7408_1, new_n7384, new_n7409);
or_5   g05061(new_n7409, new_n7383, new_n7410);
and_5  g05062(new_n7410, new_n7381, new_n7411);
or_5   g05063(new_n7411, new_n7380, new_n7412);
and_5  g05064(new_n7412, new_n7378, new_n7413);
or_5   g05065(new_n7413, new_n7377_1, new_n7414);
and_5  g05066(new_n7414, new_n7375, new_n7415);
or_5   g05067(new_n7415, new_n7374, new_n7416);
and_5  g05068(new_n7416, new_n7372, new_n7417);
xor_4  g05069(new_n7417, new_n7371, new_n7418);
xor_4  g05070(new_n7415, new_n7374, new_n7419);
xor_4  g05071(new_n7368, new_n7315, new_n7420);
nor_5  g05072(new_n7420, new_n7419, new_n7421_1);
xor_4  g05073(new_n7420, new_n7419, new_n7422);
not_10 g05074(new_n7422, new_n7423);
xor_4  g05075(new_n7413, new_n7377_1, new_n7424);
xor_4  g05076(new_n7366, new_n7320, new_n7425);
not_10 g05077(new_n7425, new_n7426);
nor_5  g05078(new_n7426, new_n7424, new_n7427);
not_10 g05079(new_n7427, new_n7428_1);
xor_4  g05080(new_n7426, new_n7424, new_n7429);
xor_4  g05081(new_n7411, new_n7380, new_n7430);
xor_4  g05082(new_n7364, new_n7325, new_n7431);
not_10 g05083(new_n7431, new_n7432_1);
nor_5  g05084(new_n7432_1, new_n7430, new_n7433);
not_10 g05085(new_n7433, new_n7434);
xor_4  g05086(new_n7432_1, new_n7430, new_n7435);
xor_4  g05087(new_n7409, new_n7383, new_n7436);
xor_4  g05088(new_n7362, new_n7329, new_n7437_1);
not_10 g05089(new_n7437_1, new_n7438);
nor_5  g05090(new_n7438, new_n7436, new_n7439);
not_10 g05091(new_n7439, new_n7440);
xor_4  g05092(new_n7438, new_n7436, new_n7441);
xor_4  g05093(new_n7407, new_n7386, new_n7442);
xor_4  g05094(new_n7360, new_n7333, new_n7443);
not_10 g05095(new_n7443, new_n7444);
nor_5  g05096(new_n7444, new_n7442, new_n7445);
not_10 g05097(new_n7445, new_n7446);
xor_4  g05098(new_n7444, new_n7442, new_n7447);
xor_4  g05099(new_n7405, new_n7389, new_n7448);
xor_4  g05100(new_n7358, new_n7337, new_n7449);
not_10 g05101(new_n7449, new_n7450);
nor_5  g05102(new_n7450, new_n7448, new_n7451);
not_10 g05103(new_n7451, new_n7452);
xor_4  g05104(new_n7450, new_n7448, new_n7453);
xor_4  g05105(new_n7356, new_n7341, new_n7454);
not_10 g05106(new_n7454, new_n7455);
xor_4  g05107(new_n7403_1, new_n7391, new_n7456);
nor_5  g05108(new_n7456, new_n7455, new_n7457);
not_10 g05109(new_n7457, new_n7458);
xor_4  g05110(new_n7354, new_n7346_1, new_n7459);
xnor_4 g05111(n15967, n7524, new_n7460_1);
xor_4  g05112(new_n7460_1, new_n7401, new_n7461);
and_5  g05113(new_n7461, new_n7459, new_n7462);
not_10 g05114(new_n7459, new_n7463);
xnor_4 g05115(new_n7461, new_n7463, new_n7464);
xnor_4 g05116(n25435, n20658, new_n7465);
xor_4  g05117(new_n7350, new_n3882, new_n7466);
not_10 g05118(new_n7466, new_n7467);
nor_5  g05119(new_n7467, new_n7465, new_n7468);
xnor_4 g05120(n15743, n13319, new_n7469);
xnor_4 g05121(new_n7469, new_n7398, new_n7470);
nor_5  g05122(new_n7470, new_n7468, new_n7471);
xor_4  g05123(new_n7352, new_n7351, new_n7472);
not_10 g05124(new_n7472, new_n7473);
xor_4  g05125(new_n7470, new_n7468, new_n7474);
and_5  g05126(new_n7474, new_n7473, new_n7475_1);
nor_5  g05127(new_n7475_1, new_n7471, new_n7476);
not_10 g05128(new_n7476, new_n7477_1);
and_5  g05129(new_n7477_1, new_n7464, new_n7478);
nor_5  g05130(new_n7478, new_n7462, new_n7479);
not_10 g05131(new_n7479, new_n7480);
xor_4  g05132(new_n7456, new_n7455, new_n7481);
and_5  g05133(new_n7481, new_n7480, new_n7482);
not_10 g05134(new_n7482, new_n7483);
and_5  g05135(new_n7483, new_n7458, new_n7484);
not_10 g05136(new_n7484, new_n7485);
and_5  g05137(new_n7485, new_n7453, new_n7486);
not_10 g05138(new_n7486, new_n7487);
and_5  g05139(new_n7487, new_n7452, new_n7488);
not_10 g05140(new_n7488, new_n7489);
and_5  g05141(new_n7489, new_n7447, new_n7490);
not_10 g05142(new_n7490, new_n7491);
and_5  g05143(new_n7491, new_n7446, new_n7492);
not_10 g05144(new_n7492, new_n7493);
and_5  g05145(new_n7493, new_n7441, new_n7494);
not_10 g05146(new_n7494, new_n7495);
and_5  g05147(new_n7495, new_n7440, new_n7496);
not_10 g05148(new_n7496, new_n7497);
and_5  g05149(new_n7497, new_n7435, new_n7498);
not_10 g05150(new_n7498, new_n7499);
and_5  g05151(new_n7499, new_n7434, new_n7500);
not_10 g05152(new_n7500, new_n7501);
and_5  g05153(new_n7501, new_n7429, new_n7502);
not_10 g05154(new_n7502, new_n7503);
and_5  g05155(new_n7503, new_n7428_1, new_n7504);
nor_5  g05156(new_n7504, new_n7423, new_n7505);
nor_5  g05157(new_n7505, new_n7421_1, new_n7506);
xor_4  g05158(new_n7506, new_n7418, n809);
and_5  g05159(new_n7295, n2978, new_n7508);
xnor_4 g05160(n19282, n2978, new_n7509);
not_10 g05161(new_n7509, new_n7510);
not_10 g05162(n23697, new_n7511);
or_5   g05163(new_n7511, n12657, new_n7512);
xnor_4 g05164(n23697, n12657, new_n7513);
not_10 g05165(new_n7513, new_n7514_1);
not_10 g05166(n2289, new_n7515);
or_5   g05167(n17077, new_n7515, new_n7516);
xnor_4 g05168(n17077, n2289, new_n7517);
not_10 g05169(new_n7517, new_n7518);
not_10 g05170(n1112, new_n7519);
or_5   g05171(n26510, new_n7519, new_n7520);
xor_4  g05172(n26510, n1112, new_n7521);
not_10 g05173(n20179, new_n7522);
or_5   g05174(n23068, new_n7522, new_n7523);
xor_4  g05175(n23068, n20179, new_n7524_1);
not_10 g05176(n19228, new_n7525);
or_5   g05177(n19514, new_n7525, new_n7526);
xor_4  g05178(n19514, n19228, new_n7527);
not_10 g05179(n15539, new_n7528);
or_5   g05180(new_n7528, n10053, new_n7529);
xnor_4 g05181(n15539, n10053, new_n7530);
or_5   g05182(new_n3817, n8052, new_n7531);
not_10 g05183(n8052, new_n7532);
or_5   g05184(n8399, new_n7532, new_n7533);
not_10 g05185(n10158, new_n7534);
and_5  g05186(new_n7534, n9507, new_n7535);
and_5  g05187(n10158, new_n3823, new_n7536);
not_10 g05188(new_n7536, new_n7537);
not_10 g05189(n18962, new_n7538);
and_5  g05190(n26979, new_n7538, new_n7539);
and_5  g05191(new_n7539, new_n7537, new_n7540);
nor_5  g05192(new_n7540, new_n7535, new_n7541);
not_10 g05193(new_n7541, new_n7542);
nand_5 g05194(new_n7542, new_n7533, new_n7543);
and_5  g05195(new_n7543, new_n7531, new_n7544);
nand_5 g05196(new_n7544, new_n7530, new_n7545);
and_5  g05197(new_n7545, new_n7529, new_n7546);
or_5   g05198(new_n7546, new_n7527, new_n7547);
and_5  g05199(new_n7547, new_n7526, new_n7548);
or_5   g05200(new_n7548, new_n7524_1, new_n7549);
and_5  g05201(new_n7549, new_n7523, new_n7550);
or_5   g05202(new_n7550, new_n7521, new_n7551);
and_5  g05203(new_n7551, new_n7520, new_n7552);
or_5   g05204(new_n7552, new_n7518, new_n7553);
and_5  g05205(new_n7553, new_n7516, new_n7554);
or_5   g05206(new_n7554, new_n7514_1, new_n7555);
and_5  g05207(new_n7555, new_n7512, new_n7556);
nor_5  g05208(new_n7556, new_n7510, new_n7557);
nor_5  g05209(new_n7557, new_n7508, new_n7558_1);
nor_5  g05210(n26986, n22626, new_n7559);
and_5  g05211(new_n2426, new_n2421_1, new_n7560);
not_10 g05212(new_n7560, new_n7561);
xor_4  g05213(n4256, n1654, new_n7562);
not_10 g05214(new_n7562, new_n7563);
or_5   g05215(n22332, n13783, new_n7564);
or_5   g05216(new_n2425, new_n2422, new_n7565);
and_5  g05217(new_n7565, new_n7564, new_n7566_1);
xor_4  g05218(new_n7566_1, new_n7563, new_n7567);
not_10 g05219(new_n7567, new_n7568);
nor_5  g05220(new_n7568, new_n7561, new_n7569_1);
not_10 g05221(new_n7569_1, new_n7570);
xor_4  g05222(n21287, n14440, new_n7571);
not_10 g05223(new_n7571, new_n7572_1);
or_5   g05224(n4256, n1654, new_n7573);
or_5   g05225(new_n7566_1, new_n7563, new_n7574);
and_5  g05226(new_n7574, new_n7573, new_n7575_1);
xor_4  g05227(new_n7575_1, new_n7572_1, new_n7576);
not_10 g05228(new_n7576, new_n7577);
nor_5  g05229(new_n7577, new_n7570, new_n7578);
not_10 g05230(new_n7578, new_n7579);
xor_4  g05231(n26986, n22626, new_n7580);
not_10 g05232(new_n7580, new_n7581);
or_5   g05233(n21287, n14440, new_n7582);
or_5   g05234(new_n7575_1, new_n7572_1, new_n7583);
and_5  g05235(new_n7583, new_n7582, new_n7584);
xor_4  g05236(new_n7584, new_n7581, new_n7585_1);
not_10 g05237(new_n7585_1, new_n7586);
nor_5  g05238(new_n7586, new_n7579, new_n7587);
and_5  g05239(new_n7587, new_n7559, new_n7588_1);
nor_5  g05240(new_n7584, new_n7581, new_n7589);
or_5   g05241(new_n7589, new_n7559, new_n7590);
nor_5  g05242(new_n7590, new_n7587, new_n7591);
nor_5  g05243(new_n7591, new_n7588_1, new_n7592);
nor_5  g05244(n13494, n3425, new_n7593_1);
not_10 g05245(new_n7593_1, new_n7594);
xnor_4 g05246(n13494, n3425, new_n7595);
or_5   g05247(n25345, n9967, new_n7596);
xor_4  g05248(n25345, n9967, new_n7597);
nand_5 g05249(n20946, n9655, new_n7598_1);
or_5   g05250(n20946, n9655, new_n7599);
nor_5  g05251(n13490, n7751, new_n7600);
nor_5  g05252(new_n2450, new_n2429, new_n7601);
nor_5  g05253(new_n7601, new_n7600, new_n7602);
nand_5 g05254(new_n7602, new_n7599, new_n7603);
and_5  g05255(new_n7603, new_n7598_1, new_n7604);
nand_5 g05256(new_n7604, new_n7597, new_n7605);
and_5  g05257(new_n7605, new_n7596, new_n7606);
nor_5  g05258(new_n7606, new_n7595, new_n7607_1);
not_10 g05259(new_n7607_1, new_n7608);
and_5  g05260(new_n7608, new_n7594, new_n7609);
and_5  g05261(new_n7609, new_n7592, new_n7610_1);
nor_5  g05262(new_n7609, new_n7592, new_n7611);
xor_4  g05263(new_n7586, new_n7579, new_n7612);
xnor_4 g05264(new_n7606, new_n7595, new_n7613);
nor_5  g05265(new_n7613, new_n7612, new_n7614);
xor_4  g05266(new_n7606, new_n7595, new_n7615);
xnor_4 g05267(new_n7615, new_n7612, new_n7616_1);
not_10 g05268(new_n7616_1, new_n7617);
xor_4  g05269(new_n7577, new_n7570, new_n7618);
xnor_4 g05270(new_n7604, new_n7597, new_n7619);
or_5   g05271(new_n7619, new_n7618, new_n7620);
xor_4  g05272(new_n7604, new_n7597, new_n7621);
xnor_4 g05273(new_n7621, new_n7618, new_n7622);
not_10 g05274(new_n7622, new_n7623);
xor_4  g05275(new_n7568, new_n7561, new_n7624);
xor_4  g05276(n20946, n9655, new_n7625);
xor_4  g05277(new_n7625, new_n7602, new_n7626);
or_5   g05278(new_n7626, new_n7624, new_n7627);
xor_4  g05279(new_n7626, new_n7624, new_n7628);
not_10 g05280(new_n7628, new_n7629);
nand_5 g05281(new_n2451, new_n2428, new_n7630_1);
not_10 g05282(new_n2452, new_n7631);
or_5   g05283(new_n2500, new_n7631, new_n7632);
and_5  g05284(new_n7632, new_n7630_1, new_n7633);
or_5   g05285(new_n7633, new_n7629, new_n7634);
and_5  g05286(new_n7634, new_n7627, new_n7635);
or_5   g05287(new_n7635, new_n7623, new_n7636);
and_5  g05288(new_n7636, new_n7620, new_n7637);
nor_5  g05289(new_n7637, new_n7617, new_n7638);
nor_5  g05290(new_n7638, new_n7614, new_n7639);
not_10 g05291(new_n7639, new_n7640);
nor_5  g05292(new_n7640, new_n7611, new_n7641);
nor_5  g05293(new_n7641, new_n7588_1, new_n7642);
not_10 g05294(new_n7642, new_n7643_1);
nor_5  g05295(new_n7643_1, new_n7610_1, new_n7644);
xor_4  g05296(new_n7644, new_n7558_1, new_n7645);
xnor_4 g05297(new_n7609, new_n7592, new_n7646);
xor_4  g05298(new_n7646, new_n7640, new_n7647_1);
nor_5  g05299(new_n7647_1, new_n7558_1, new_n7648);
xor_4  g05300(new_n7647_1, new_n7558_1, new_n7649);
not_10 g05301(new_n7649, new_n7650);
xor_4  g05302(new_n7556, new_n7510, new_n7651);
xor_4  g05303(new_n7637, new_n7617, new_n7652);
not_10 g05304(new_n7652, new_n7653);
nor_5  g05305(new_n7653, new_n7651, new_n7654);
xor_4  g05306(new_n7653, new_n7651, new_n7655);
xor_4  g05307(new_n7554, new_n7514_1, new_n7656);
xor_4  g05308(new_n7635, new_n7623, new_n7657_1);
not_10 g05309(new_n7657_1, new_n7658);
nor_5  g05310(new_n7658, new_n7656, new_n7659);
xor_4  g05311(new_n7658, new_n7656, new_n7660);
xor_4  g05312(new_n7552, new_n7518, new_n7661);
xor_4  g05313(new_n7633, new_n7629, new_n7662);
not_10 g05314(new_n7662, new_n7663);
nor_5  g05315(new_n7663, new_n7661, new_n7664);
xor_4  g05316(new_n7663, new_n7661, new_n7665);
not_10 g05317(new_n2501, new_n7666);
xor_4  g05318(new_n7550, new_n7521, new_n7667);
nor_5  g05319(new_n7667, new_n7666, new_n7668);
xnor_4 g05320(new_n7667, new_n2501, new_n7669);
not_10 g05321(new_n7669, new_n7670_1);
xor_4  g05322(new_n7548, new_n7524_1, new_n7671);
nor_5  g05323(new_n7671, new_n2506, new_n7672);
not_10 g05324(new_n7672, new_n7673);
xor_4  g05325(new_n7671, new_n2506, new_n7674_1);
not_10 g05326(new_n7674_1, new_n7675);
xor_4  g05327(new_n7546, new_n7527, new_n7676);
nor_5  g05328(new_n7676, new_n2512, new_n7677);
not_10 g05329(new_n7677, new_n7678_1);
xor_4  g05330(new_n7676, new_n2512, new_n7679_1);
not_10 g05331(new_n7679_1, new_n7680);
xor_4  g05332(new_n7544, new_n7530, new_n7681);
nor_5  g05333(new_n7681, new_n2517, new_n7682);
not_10 g05334(new_n7682, new_n7683);
xor_4  g05335(new_n7681, new_n2517, new_n7684);
xnor_4 g05336(n8399, n8052, new_n7685);
xor_4  g05337(new_n7685, new_n7542, new_n7686_1);
and_5  g05338(new_n7686_1, new_n2520, new_n7687);
not_10 g05339(new_n7687, new_n7688);
xnor_4 g05340(new_n7686_1, new_n2524, new_n7689);
xnor_4 g05341(n26979, n18962, new_n7690);
nor_5  g05342(new_n7690, new_n2528, new_n7691);
xnor_4 g05343(n10158, n9507, new_n7692_1);
xnor_4 g05344(new_n7692_1, new_n7539, new_n7693_1);
nor_5  g05345(new_n7693_1, new_n7691, new_n7694);
not_10 g05346(new_n7694, new_n7695);
xor_4  g05347(new_n7693_1, new_n7691, new_n7696);
and_5  g05348(new_n7696, new_n2533_1, new_n7697);
not_10 g05349(new_n7697, new_n7698_1);
and_5  g05350(new_n7698_1, new_n7695, new_n7699);
not_10 g05351(new_n7699, new_n7700);
and_5  g05352(new_n7700, new_n7689, new_n7701);
not_10 g05353(new_n7701, new_n7702);
and_5  g05354(new_n7702, new_n7688, new_n7703);
not_10 g05355(new_n7703, new_n7704);
and_5  g05356(new_n7704, new_n7684, new_n7705);
not_10 g05357(new_n7705, new_n7706);
and_5  g05358(new_n7706, new_n7683, new_n7707);
nor_5  g05359(new_n7707, new_n7680, new_n7708_1);
not_10 g05360(new_n7708_1, new_n7709);
and_5  g05361(new_n7709, new_n7678_1, new_n7710);
nor_5  g05362(new_n7710, new_n7675, new_n7711);
not_10 g05363(new_n7711, new_n7712);
and_5  g05364(new_n7712, new_n7673, new_n7713);
nor_5  g05365(new_n7713, new_n7670_1, new_n7714);
nor_5  g05366(new_n7714, new_n7668, new_n7715);
not_10 g05367(new_n7715, new_n7716);
and_5  g05368(new_n7716, new_n7665, new_n7717);
nor_5  g05369(new_n7717, new_n7664, new_n7718);
not_10 g05370(new_n7718, new_n7719);
and_5  g05371(new_n7719, new_n7660, new_n7720);
nor_5  g05372(new_n7720, new_n7659, new_n7721_1);
not_10 g05373(new_n7721_1, new_n7722);
and_5  g05374(new_n7722, new_n7655, new_n7723);
nor_5  g05375(new_n7723, new_n7654, new_n7724);
nor_5  g05376(new_n7724, new_n7650, new_n7725);
nor_5  g05377(new_n7725, new_n7648, new_n7726);
xor_4  g05378(new_n7726, new_n7645, n819);
not_10 g05379(n22626, new_n7728);
and_5  g05380(new_n7728, n8856, new_n7729);
not_10 g05381(new_n7729, new_n7730);
xnor_4 g05382(n22626, n8856, new_n7731_1);
not_10 g05383(new_n7731_1, new_n7732);
or_5   g05384(n14440, new_n3410, new_n7733);
xnor_4 g05385(n14440, n14130, new_n7734);
not_10 g05386(new_n7734, new_n7735);
or_5   g05387(new_n3411, n1654, new_n7736);
xnor_4 g05388(n16482, n1654, new_n7737);
not_10 g05389(new_n7737, new_n7738);
or_5   g05390(n13783, new_n3412, new_n7739);
xnor_4 g05391(n13783, n9942, new_n7740);
not_10 g05392(new_n7740, new_n7741);
or_5   g05393(n26660, new_n3413, new_n7742);
xnor_4 g05394(n26660, n25643, new_n7743);
not_10 g05395(new_n7743, new_n7744);
or_5   g05396(new_n3414, n3018, new_n7745);
xnor_4 g05397(n9557, n3018, new_n7746);
not_10 g05398(new_n7746, new_n7747);
or_5   g05399(n3480, new_n3415, new_n7748);
xnor_4 g05400(n3480, n3136, new_n7749);
not_10 g05401(n16722, new_n7750);
or_5   g05402(new_n7750, n6385, new_n7751_1);
or_5   g05403(n16722, new_n2361_1, new_n7752);
and_5  g05404(new_n2367, n11486, new_n7753);
not_10 g05405(n11486, new_n7754);
and_5  g05406(n20138, new_n7754, new_n7755);
not_10 g05407(new_n7755, new_n7756);
not_10 g05408(n13781, new_n7757);
nor_5  g05409(new_n7757, n9251, new_n7758);
and_5  g05410(new_n7758, new_n7756, new_n7759_1);
nor_5  g05411(new_n7759_1, new_n7753, new_n7760);
not_10 g05412(new_n7760, new_n7761);
nand_5 g05413(new_n7761, new_n7752, new_n7762);
and_5  g05414(new_n7762, new_n7751_1, new_n7763);
nand_5 g05415(new_n7763, new_n7749, new_n7764);
and_5  g05416(new_n7764, new_n7748, new_n7765);
or_5   g05417(new_n7765, new_n7747, new_n7766);
and_5  g05418(new_n7766, new_n7745, new_n7767);
or_5   g05419(new_n7767, new_n7744, new_n7768);
and_5  g05420(new_n7768, new_n7742, new_n7769_1);
or_5   g05421(new_n7769_1, new_n7741, new_n7770);
and_5  g05422(new_n7770, new_n7739, new_n7771);
or_5   g05423(new_n7771, new_n7738, new_n7772);
and_5  g05424(new_n7772, new_n7736, new_n7773_1);
or_5   g05425(new_n7773_1, new_n7735, new_n7774);
and_5  g05426(new_n7774, new_n7733, new_n7775);
nor_5  g05427(new_n7775, new_n7732, new_n7776);
not_10 g05428(new_n7776, new_n7777);
and_5  g05429(new_n7777, new_n7730, new_n7778);
not_10 g05430(n25120, new_n7779);
and_5  g05431(new_n7779, n3582, new_n7780_1);
xor_4  g05432(n25120, n3582, new_n7781);
not_10 g05433(n2145, new_n7782);
or_5   g05434(n8363, new_n7782, new_n7783);
xor_4  g05435(n8363, n2145, new_n7784);
not_10 g05436(n5031, new_n7785);
or_5   g05437(n14680, new_n7785, new_n7786);
xnor_4 g05438(n14680, n5031, new_n7787);
not_10 g05439(new_n7787, new_n7788_1);
not_10 g05440(n11044, new_n7789);
or_5   g05441(n17250, new_n7789, new_n7790);
xor_4  g05442(n17250, n11044, new_n7791);
not_10 g05443(n2421, new_n7792);
or_5   g05444(n23160, new_n7792, new_n7793);
xor_4  g05445(n23160, n2421, new_n7794_1);
not_10 g05446(n987, new_n7795);
or_5   g05447(n16524, new_n7795, new_n7796);
xor_4  g05448(n16524, n987, new_n7797);
not_10 g05449(n20478, new_n7798);
or_5   g05450(new_n7798, n11056, new_n7799);
xnor_4 g05451(n20478, n11056, new_n7800);
not_10 g05452(n15271, new_n7801);
or_5   g05453(n26882, new_n7801, new_n7802);
not_10 g05454(n26882, new_n7803);
or_5   g05455(new_n7803, n15271, new_n7804);
not_10 g05456(n22619, new_n7805);
and_5  g05457(n25877, new_n7805, new_n7806);
nor_5  g05458(n25877, new_n7805, new_n7807);
not_10 g05459(n6775, new_n7808);
and_5  g05460(n24323, new_n7808, new_n7809);
not_10 g05461(new_n7809, new_n7810);
nor_5  g05462(new_n7810, new_n7807, new_n7811_1);
nor_5  g05463(new_n7811_1, new_n7806, new_n7812);
not_10 g05464(new_n7812, new_n7813);
nand_5 g05465(new_n7813, new_n7804, new_n7814);
and_5  g05466(new_n7814, new_n7802, new_n7815);
nand_5 g05467(new_n7815, new_n7800, new_n7816);
and_5  g05468(new_n7816, new_n7799, new_n7817);
or_5   g05469(new_n7817, new_n7797, new_n7818);
and_5  g05470(new_n7818, new_n7796, new_n7819);
or_5   g05471(new_n7819, new_n7794_1, new_n7820);
and_5  g05472(new_n7820, new_n7793, new_n7821);
or_5   g05473(new_n7821, new_n7791, new_n7822);
and_5  g05474(new_n7822, new_n7790, new_n7823);
or_5   g05475(new_n7823, new_n7788_1, new_n7824);
and_5  g05476(new_n7824, new_n7786, new_n7825);
or_5   g05477(new_n7825, new_n7784, new_n7826);
and_5  g05478(new_n7826, new_n7783, new_n7827);
nor_5  g05479(new_n7827, new_n7781, new_n7828);
nor_5  g05480(new_n7828, new_n7780_1, new_n7829);
xor_4  g05481(new_n7829, new_n7778, new_n7830_1);
not_10 g05482(new_n7830_1, new_n7831);
xor_4  g05483(new_n7827, new_n7781, new_n7832);
xor_4  g05484(new_n7775, new_n7732, new_n7833);
or_5   g05485(new_n7833, new_n7832, new_n7834_1);
xor_4  g05486(new_n7833, new_n7832, new_n7835);
not_10 g05487(new_n7835, new_n7836);
xor_4  g05488(new_n7825, new_n7784, new_n7837);
xor_4  g05489(new_n7773_1, new_n7735, new_n7838);
or_5   g05490(new_n7838, new_n7837, new_n7839);
xor_4  g05491(new_n7838, new_n7837, new_n7840);
not_10 g05492(new_n7840, new_n7841_1);
xor_4  g05493(new_n7823, new_n7788_1, new_n7842);
not_10 g05494(new_n7842, new_n7843);
xor_4  g05495(new_n7771, new_n7738, new_n7844);
not_10 g05496(new_n7844, new_n7845);
nand_5 g05497(new_n7845, new_n7843, new_n7846);
xor_4  g05498(new_n7845, new_n7843, new_n7847);
not_10 g05499(new_n7847, new_n7848);
xor_4  g05500(new_n7821, new_n7791, new_n7849);
xor_4  g05501(new_n7769_1, new_n7741, new_n7850);
or_5   g05502(new_n7850, new_n7849, new_n7851);
xor_4  g05503(new_n7850, new_n7849, new_n7852);
not_10 g05504(new_n7852, new_n7853);
xor_4  g05505(new_n7819, new_n7794_1, new_n7854);
xor_4  g05506(new_n7767, new_n7744, new_n7855);
or_5   g05507(new_n7855, new_n7854, new_n7856);
xor_4  g05508(new_n7855, new_n7854, new_n7857);
not_10 g05509(new_n7857, new_n7858);
xor_4  g05510(new_n7817, new_n7797, new_n7859);
xor_4  g05511(new_n7765, new_n7747, new_n7860);
or_5   g05512(new_n7860, new_n7859, new_n7861);
xor_4  g05513(new_n7860, new_n7859, new_n7862);
not_10 g05514(new_n7862, new_n7863);
xor_4  g05515(new_n7815, new_n7800, new_n7864);
not_10 g05516(new_n7864, new_n7865);
xor_4  g05517(new_n7763, new_n7749, new_n7866);
not_10 g05518(new_n7866, new_n7867);
nand_5 g05519(new_n7867, new_n7865, new_n7868);
xor_4  g05520(new_n7867, new_n7865, new_n7869);
not_10 g05521(new_n7869, new_n7870);
xnor_4 g05522(n26882, n15271, new_n7871);
xor_4  g05523(new_n7871, new_n7813, new_n7872);
xnor_4 g05524(n16722, n6385, new_n7873);
xor_4  g05525(new_n7873, new_n7761, new_n7874);
nand_5 g05526(new_n7874, new_n7872, new_n7875);
xor_4  g05527(new_n7874, new_n7872, new_n7876_1);
not_10 g05528(new_n7876_1, new_n7877);
xnor_4 g05529(n25877, n22619, new_n7878);
xnor_4 g05530(new_n7878, new_n7810, new_n7879);
xnor_4 g05531(n20138, n11486, new_n7880);
xor_4  g05532(new_n7880, new_n7758, new_n7881);
nand_5 g05533(new_n7881, new_n7879, new_n7882);
xnor_4 g05534(n24323, n6775, new_n7883);
xnor_4 g05535(n13781, n9251, new_n7884_1);
nor_5  g05536(new_n7884_1, new_n7883, new_n7885);
not_10 g05537(new_n7885, new_n7886);
xor_4  g05538(new_n7881, new_n7879, new_n7887);
nand_5 g05539(new_n7887, new_n7886, new_n7888);
and_5  g05540(new_n7888, new_n7882, new_n7889);
or_5   g05541(new_n7889, new_n7877, new_n7890);
and_5  g05542(new_n7890, new_n7875, new_n7891);
or_5   g05543(new_n7891, new_n7870, new_n7892);
and_5  g05544(new_n7892, new_n7868, new_n7893);
or_5   g05545(new_n7893, new_n7863, new_n7894);
and_5  g05546(new_n7894, new_n7861, new_n7895);
or_5   g05547(new_n7895, new_n7858, new_n7896);
and_5  g05548(new_n7896, new_n7856, new_n7897);
or_5   g05549(new_n7897, new_n7853, new_n7898);
and_5  g05550(new_n7898, new_n7851, new_n7899);
or_5   g05551(new_n7899, new_n7848, new_n7900);
and_5  g05552(new_n7900, new_n7846, new_n7901);
or_5   g05553(new_n7901, new_n7841_1, new_n7902);
and_5  g05554(new_n7902, new_n7839, new_n7903);
or_5   g05555(new_n7903, new_n7836, new_n7904);
and_5  g05556(new_n7904, new_n7834_1, new_n7905);
xor_4  g05557(new_n7905, new_n7831, new_n7906);
not_10 g05558(new_n7906, new_n7907);
not_10 g05559(n9554, new_n7908);
not_10 g05560(n26408, new_n7909);
not_10 g05561(n18227, new_n7910);
not_10 g05562(n7377, new_n7911);
not_10 g05563(n11630, new_n7912);
not_10 g05564(n13453, new_n7913);
nor_5  g05565(n15508, n2809, new_n7914);
and_5  g05566(new_n7914, new_n6648, new_n7915);
and_5  g05567(new_n7915, new_n6634_1, new_n7916);
and_5  g05568(new_n7916, new_n7913, new_n7917_1);
and_5  g05569(new_n7917_1, new_n7912, new_n7918);
and_5  g05570(new_n7918, new_n7911, new_n7919);
and_5  g05571(new_n7919, new_n7910, new_n7920);
and_5  g05572(new_n7920, new_n7909, new_n7921);
and_5  g05573(new_n7921, new_n7908, new_n7922);
xor_4  g05574(new_n7921, new_n7908, new_n7923);
nor_5  g05575(new_n7923, n9259, new_n7924);
xor_4  g05576(new_n7920, new_n7909, new_n7925);
nor_5  g05577(new_n7925, n21489, new_n7926);
xor_4  g05578(new_n7925, n21489, new_n7927);
not_10 g05579(new_n7927, new_n7928);
xor_4  g05580(new_n7919, new_n7910, new_n7929);
or_5   g05581(new_n7929, n20213, new_n7930);
xor_4  g05582(new_n7929, n20213, new_n7931);
not_10 g05583(new_n7931, new_n7932);
xor_4  g05584(new_n7918, new_n7911, new_n7933);
or_5   g05585(new_n7933, n13912, new_n7934);
xor_4  g05586(new_n7933, n13912, new_n7935);
not_10 g05587(new_n7935, new_n7936);
xor_4  g05588(new_n7917_1, new_n7912, new_n7937_1);
or_5   g05589(new_n7937_1, n7670, new_n7938);
xor_4  g05590(new_n7937_1, new_n3588, new_n7939);
xor_4  g05591(new_n7916, new_n7913, new_n7940);
or_5   g05592(new_n7940, n9598, new_n7941);
xor_4  g05593(new_n7940, n9598, new_n7942);
not_10 g05594(new_n7942, new_n7943_1);
xor_4  g05595(new_n7915, new_n6634_1, new_n7944);
or_5   g05596(new_n7944, n22290, new_n7945);
xor_4  g05597(new_n7914, new_n6648, new_n7946);
nor_5  g05598(new_n7946, n11273, new_n7947);
xor_4  g05599(new_n7946, n11273, new_n7948);
not_10 g05600(new_n7948, new_n7949_1);
xor_4  g05601(n15508, n2809, new_n7950_1);
or_5   g05602(new_n7950_1, n25565, new_n7951);
and_5  g05603(n21993, n15508, new_n7952);
not_10 g05604(new_n7952, new_n7953);
xor_4  g05605(new_n7950_1, n25565, new_n7954);
nand_5 g05606(new_n7954, new_n7953, new_n7955);
and_5  g05607(new_n7955, new_n7951, new_n7956);
nor_5  g05608(new_n7956, new_n7949_1, new_n7957);
or_5   g05609(new_n7957, new_n7947, new_n7958);
xor_4  g05610(new_n7944, n22290, new_n7959_1);
nand_5 g05611(new_n7959_1, new_n7958, new_n7960);
and_5  g05612(new_n7960, new_n7945, new_n7961);
or_5   g05613(new_n7961, new_n7943_1, new_n7962);
and_5  g05614(new_n7962, new_n7941, new_n7963_1);
or_5   g05615(new_n7963_1, new_n7939, new_n7964);
and_5  g05616(new_n7964, new_n7938, new_n7965);
or_5   g05617(new_n7965, new_n7936, new_n7966);
and_5  g05618(new_n7966, new_n7934, new_n7967);
or_5   g05619(new_n7967, new_n7932, new_n7968_1);
and_5  g05620(new_n7968_1, new_n7930, new_n7969);
nor_5  g05621(new_n7969, new_n7928, new_n7970);
nor_5  g05622(new_n7970, new_n7926, new_n7971);
and_5  g05623(new_n7923, n9259, new_n7972);
nor_5  g05624(new_n7972, new_n7971, new_n7973);
nor_5  g05625(new_n7973, new_n7924, new_n7974);
nor_5  g05626(new_n7974, new_n7922, new_n7975);
xor_4  g05627(new_n7975, new_n7907, new_n7976);
xor_4  g05628(new_n7903, new_n7836, new_n7977);
not_10 g05629(new_n7977, new_n7978);
xor_4  g05630(new_n7923, n9259, new_n7979);
xnor_4 g05631(new_n7979, new_n7971, new_n7980);
not_10 g05632(new_n7980, new_n7981);
nor_5  g05633(new_n7981, new_n7978, new_n7982);
xor_4  g05634(new_n7981, new_n7978, new_n7983);
xor_4  g05635(new_n7901, new_n7841_1, new_n7984);
not_10 g05636(new_n7984, new_n7985);
xor_4  g05637(new_n7969, new_n7928, new_n7986);
not_10 g05638(new_n7986, new_n7987);
and_5  g05639(new_n7987, new_n7985, new_n7988);
xor_4  g05640(new_n7986, new_n7985, new_n7989);
xor_4  g05641(new_n7899, new_n7848, new_n7990);
not_10 g05642(new_n7990, new_n7991);
xor_4  g05643(new_n7967, new_n7932, new_n7992_1);
not_10 g05644(new_n7992_1, new_n7993);
nand_5 g05645(new_n7993, new_n7991, new_n7994);
xor_4  g05646(new_n7993, new_n7991, new_n7995);
xor_4  g05647(new_n7897, new_n7853, new_n7996);
not_10 g05648(new_n7996, new_n7997);
xor_4  g05649(new_n7965, new_n7936, new_n7998);
not_10 g05650(new_n7998, new_n7999_1);
or_5   g05651(new_n7999_1, new_n7997, new_n8000);
and_5  g05652(new_n7999_1, new_n7997, new_n8001);
xor_4  g05653(new_n7895, new_n7858, new_n8002);
xor_4  g05654(new_n7963_1, new_n7939, new_n8003);
nand_5 g05655(new_n8003, new_n8002, new_n8004);
not_10 g05656(new_n8002, new_n8005);
xnor_4 g05657(new_n8003, new_n8005, new_n8006_1);
xor_4  g05658(new_n7961, new_n7943_1, new_n8007);
not_10 g05659(new_n8007, new_n8008);
xor_4  g05660(new_n7893, new_n7863, new_n8009);
not_10 g05661(new_n8009, new_n8010);
or_5   g05662(new_n8010, new_n8008, new_n8011);
xor_4  g05663(new_n8010, new_n8008, new_n8012);
xor_4  g05664(new_n7891, new_n7870, new_n8013);
xor_4  g05665(new_n7959_1, new_n7958, new_n8014);
nand_5 g05666(new_n8014, new_n8013, new_n8015);
nor_5  g05667(new_n8014, new_n8013, new_n8016);
xor_4  g05668(new_n7889, new_n7877, new_n8017);
not_10 g05669(new_n8017, new_n8018);
xor_4  g05670(new_n7887, new_n7886, new_n8019);
not_10 g05671(new_n8019, new_n8020);
xor_4  g05672(new_n7954, new_n7953, new_n8021);
not_10 g05673(new_n8021, new_n8022);
or_5   g05674(new_n8022, new_n8020, new_n8023);
xor_4  g05675(n21993, n15508, new_n8024);
xor_4  g05676(new_n7884_1, new_n7883, new_n8025);
nand_5 g05677(new_n8025, new_n8024, new_n8026);
xnor_4 g05678(new_n8021, new_n8020, new_n8027_1);
nand_5 g05679(new_n8027_1, new_n8026, new_n8028);
and_5  g05680(new_n8028, new_n8023, new_n8029);
and_5  g05681(new_n8029, new_n8018, new_n8030);
xor_4  g05682(new_n7956, new_n7948, new_n8031_1);
xor_4  g05683(new_n8029, new_n8018, new_n8032);
and_5  g05684(new_n8032, new_n8031_1, new_n8033);
or_5   g05685(new_n8033, new_n8030, new_n8034);
or_5   g05686(new_n8034, new_n8016, new_n8035);
nand_5 g05687(new_n8035, new_n8015, new_n8036);
nand_5 g05688(new_n8036, new_n8012, new_n8037);
nand_5 g05689(new_n8037, new_n8011, new_n8038);
nand_5 g05690(new_n8038, new_n8006_1, new_n8039);
and_5  g05691(new_n8039, new_n8004, new_n8040);
or_5   g05692(new_n8040, new_n8001, new_n8041);
and_5  g05693(new_n8041, new_n8000, new_n8042_1);
nand_5 g05694(new_n8042_1, new_n7995, new_n8043);
and_5  g05695(new_n8043, new_n7994, new_n8044);
nor_5  g05696(new_n8044, new_n7989, new_n8045);
nor_5  g05697(new_n8045, new_n7988, new_n8046);
and_5  g05698(new_n8046, new_n7983, new_n8047);
nor_5  g05699(new_n8047, new_n7982, new_n8048);
xor_4  g05700(new_n8048, new_n7976, n829);
xnor_4 g05701(n23272, n14826, new_n8050);
or_5   g05702(n23493, n11481, new_n8051);
xor_4  g05703(n23493, n11481, new_n8052_1);
not_10 g05704(new_n8052_1, new_n8053);
or_5   g05705(n16439, n10275, new_n8054);
xor_4  g05706(n16439, n10275, new_n8055);
not_10 g05707(new_n8055, new_n8056);
or_5   g05708(n15241, n15146, new_n8057);
xor_4  g05709(n15241, n15146, new_n8058);
not_10 g05710(new_n8058, new_n8059);
or_5   g05711(n11579, n7678, new_n8060);
xor_4  g05712(n11579, n7678, new_n8061);
not_10 g05713(new_n8061, new_n8062);
or_5   g05714(n3785, n21, new_n8063);
xor_4  g05715(n3785, n21, new_n8064);
not_10 g05716(new_n8064, new_n8065);
or_5   g05717(n20250, n1682, new_n8066);
xor_4  g05718(n20250, n1682, new_n8067_1);
not_10 g05719(new_n8067_1, new_n8068);
or_5   g05720(n7963, n5822, new_n8069);
xor_4  g05721(n7963, n5822, new_n8070);
not_10 g05722(new_n8070, new_n8071);
or_5   g05723(n26443, n10017, new_n8072);
and_5  g05724(n3618, n1681, new_n8073);
not_10 g05725(new_n8073, new_n8074);
xor_4  g05726(n26443, n10017, new_n8075);
nand_5 g05727(new_n8075, new_n8074, new_n8076);
and_5  g05728(new_n8076, new_n8072, new_n8077);
or_5   g05729(new_n8077, new_n8071, new_n8078);
and_5  g05730(new_n8078, new_n8069, new_n8079);
or_5   g05731(new_n8079, new_n8068, new_n8080);
and_5  g05732(new_n8080, new_n8066, new_n8081);
or_5   g05733(new_n8081, new_n8065, new_n8082);
and_5  g05734(new_n8082, new_n8063, new_n8083);
or_5   g05735(new_n8083, new_n8062, new_n8084);
and_5  g05736(new_n8084, new_n8060, new_n8085);
or_5   g05737(new_n8085, new_n8059, new_n8086);
and_5  g05738(new_n8086, new_n8057, new_n8087);
or_5   g05739(new_n8087, new_n8056, new_n8088);
and_5  g05740(new_n8088, new_n8054, new_n8089);
or_5   g05741(new_n8089, new_n8053, new_n8090);
and_5  g05742(new_n8090, new_n8051, new_n8091);
xor_4  g05743(new_n8091, new_n8050, new_n8092);
nor_5  g05744(new_n8092, n22764, new_n8093);
xor_4  g05745(new_n8092, n22764, new_n8094);
not_10 g05746(new_n8094, new_n8095_1);
not_10 g05747(n26264, new_n8096);
xor_4  g05748(new_n8089, new_n8053, new_n8097);
not_10 g05749(new_n8097, new_n8098);
nand_5 g05750(new_n8098, new_n8096, new_n8099);
xor_4  g05751(new_n8098, new_n8096, new_n8100);
not_10 g05752(new_n8100, new_n8101);
not_10 g05753(n7841, new_n8102);
xor_4  g05754(new_n8087, new_n8056, new_n8103_1);
not_10 g05755(new_n8103_1, new_n8104);
nand_5 g05756(new_n8104, new_n8102, new_n8105);
xor_4  g05757(new_n8104, new_n8102, new_n8106);
not_10 g05758(new_n8106, new_n8107);
not_10 g05759(n16812, new_n8108);
xor_4  g05760(new_n8085, new_n8059, new_n8109_1);
not_10 g05761(new_n8109_1, new_n8110);
nand_5 g05762(new_n8110, new_n8108, new_n8111);
xor_4  g05763(new_n8110, new_n8108, new_n8112);
not_10 g05764(new_n8112, new_n8113);
not_10 g05765(n25068, new_n8114);
xor_4  g05766(new_n8083, new_n8062, new_n8115);
not_10 g05767(new_n8115, new_n8116);
nand_5 g05768(new_n8116, new_n8114, new_n8117);
xor_4  g05769(new_n8116, new_n8114, new_n8118);
not_10 g05770(new_n8118, new_n8119);
not_10 g05771(n2331, new_n8120);
xor_4  g05772(new_n8081, new_n8065, new_n8121);
not_10 g05773(new_n8121, new_n8122);
nand_5 g05774(new_n8122, new_n8120, new_n8123);
xor_4  g05775(new_n8122, new_n8120, new_n8124);
not_10 g05776(n22631, new_n8125);
xor_4  g05777(new_n8079, new_n8068, new_n8126);
not_10 g05778(new_n8126, new_n8127_1);
nand_5 g05779(new_n8127_1, new_n8125, new_n8128);
xor_4  g05780(new_n8127_1, new_n8125, new_n8129);
not_10 g05781(n16743, new_n8130_1);
xor_4  g05782(new_n8077, new_n8071, new_n8131);
not_10 g05783(new_n8131, new_n8132);
or_5   g05784(new_n8132, new_n8130_1, new_n8133);
xor_4  g05785(new_n8132, new_n8130_1, new_n8134);
not_10 g05786(n15258, new_n8135_1);
not_10 g05787(n4588, new_n8136);
and_5  g05788(new_n2546, new_n8136, new_n8137);
nand_5 g05789(new_n8137, new_n8135_1, new_n8138);
xnor_4 g05790(new_n8075, new_n8073, new_n8139_1);
not_10 g05791(new_n8139_1, new_n8140);
xor_4  g05792(new_n8137, new_n8135_1, new_n8141);
nand_5 g05793(new_n8141, new_n8140, new_n8142);
and_5  g05794(new_n8142, new_n8138, new_n8143);
nand_5 g05795(new_n8143, new_n8134, new_n8144);
and_5  g05796(new_n8144, new_n8133, new_n8145);
nand_5 g05797(new_n8145, new_n8129, new_n8146);
nand_5 g05798(new_n8146, new_n8128, new_n8147);
nand_5 g05799(new_n8147, new_n8124, new_n8148_1);
and_5  g05800(new_n8148_1, new_n8123, new_n8149_1);
or_5   g05801(new_n8149_1, new_n8119, new_n8150);
and_5  g05802(new_n8150, new_n8117, new_n8151);
or_5   g05803(new_n8151, new_n8113, new_n8152);
and_5  g05804(new_n8152, new_n8111, new_n8153);
or_5   g05805(new_n8153, new_n8107, new_n8154);
and_5  g05806(new_n8154, new_n8105, new_n8155);
or_5   g05807(new_n8155, new_n8101, new_n8156);
and_5  g05808(new_n8156, new_n8099, new_n8157);
nor_5  g05809(new_n8157, new_n8095_1, new_n8158);
or_5   g05810(new_n8158, new_n8093, new_n8159_1);
nor_5  g05811(n23272, n14826, new_n8160);
nor_5  g05812(new_n8091, new_n8050, new_n8161);
nor_5  g05813(new_n8161, new_n8160, new_n8162);
or_5   g05814(new_n8162, new_n8159_1, new_n8163);
and_5  g05815(new_n4449, n12702, new_n8164);
not_10 g05816(new_n8164, new_n8165);
xor_4  g05817(n18105, n12702, new_n8166);
or_5   g05818(new_n5592, n24196, new_n8167);
xor_4  g05819(n26797, n24196, new_n8168);
or_5   g05820(new_n5593_1, n16376, new_n8169);
xor_4  g05821(n23913, n16376, new_n8170);
or_5   g05822(n25381, new_n5594, new_n8171);
xor_4  g05823(n25381, n22554, new_n8172);
or_5   g05824(new_n5595, n12587, new_n8173);
xor_4  g05825(n20429, n12587, new_n8174);
or_5   g05826(new_n5596, n268, new_n8175);
xor_4  g05827(n3909, n268, new_n8176);
or_5   g05828(n24879, new_n5597, new_n8177);
xnor_4 g05829(n24879, n23974, new_n8178);
or_5   g05830(new_n4456, n2146, new_n8179_1);
or_5   g05831(n6785, new_n5598, new_n8180);
not_10 g05832(n22173, new_n8181);
and_5  g05833(n24032, new_n8181, new_n8182);
not_10 g05834(n22843, new_n8183);
nor_5  g05835(new_n8183, n583, new_n8184);
not_10 g05836(n24032, new_n8185);
and_5  g05837(new_n8185, n22173, new_n8186);
not_10 g05838(new_n8186, new_n8187);
and_5  g05839(new_n8187, new_n8184, new_n8188);
nor_5  g05840(new_n8188, new_n8182, new_n8189);
not_10 g05841(new_n8189, new_n8190);
nand_5 g05842(new_n8190, new_n8180, new_n8191);
and_5  g05843(new_n8191, new_n8179_1, new_n8192);
nand_5 g05844(new_n8192, new_n8178, new_n8193);
and_5  g05845(new_n8193, new_n8177, new_n8194_1);
or_5   g05846(new_n8194_1, new_n8176, new_n8195);
and_5  g05847(new_n8195, new_n8175, new_n8196);
or_5   g05848(new_n8196, new_n8174, new_n8197);
and_5  g05849(new_n8197, new_n8173, new_n8198);
or_5   g05850(new_n8198, new_n8172, new_n8199);
and_5  g05851(new_n8199, new_n8171, new_n8200);
or_5   g05852(new_n8200, new_n8170, new_n8201);
and_5  g05853(new_n8201, new_n8169, new_n8202);
or_5   g05854(new_n8202, new_n8168, new_n8203);
and_5  g05855(new_n8203, new_n8167, new_n8204);
nor_5  g05856(new_n8204, new_n8166, new_n8205);
not_10 g05857(new_n8205, new_n8206);
and_5  g05858(new_n8206, new_n8165, new_n8207);
xor_4  g05859(new_n8204, new_n8166, new_n8208);
or_5   g05860(new_n8208, n1536, new_n8209);
not_10 g05861(n1536, new_n8210);
xor_4  g05862(new_n8208, new_n8210, new_n8211);
xor_4  g05863(new_n8202, new_n8168, new_n8212);
or_5   g05864(new_n8212, n19454, new_n8213);
not_10 g05865(n19454, new_n8214);
xor_4  g05866(new_n8212, new_n8214, new_n8215_1);
xor_4  g05867(new_n8200, new_n8170, new_n8216);
or_5   g05868(new_n8216, n9445, new_n8217);
not_10 g05869(n9445, new_n8218);
xor_4  g05870(new_n8216, new_n8218, new_n8219);
xor_4  g05871(new_n8198, new_n8172, new_n8220);
or_5   g05872(new_n8220, n1279, new_n8221);
not_10 g05873(n1279, new_n8222);
xor_4  g05874(new_n8220, new_n8222, new_n8223);
xor_4  g05875(new_n8196, new_n8174, new_n8224);
or_5   g05876(new_n8224, n8324, new_n8225);
not_10 g05877(n8324, new_n8226);
xor_4  g05878(new_n8224, new_n8226, new_n8227);
xor_4  g05879(new_n8194_1, new_n8176, new_n8228);
or_5   g05880(new_n8228, n12546, new_n8229);
not_10 g05881(n12546, new_n8230);
xor_4  g05882(new_n8228, new_n8230, new_n8231);
xor_4  g05883(new_n8192, new_n8178, new_n8232);
or_5   g05884(new_n8232, n21078, new_n8233);
not_10 g05885(n21078, new_n8234);
xor_4  g05886(new_n8232, new_n8234, new_n8235);
not_10 g05887(n24485, new_n8236);
xnor_4 g05888(n6785, n2146, new_n8237);
xor_4  g05889(new_n8237, new_n8190, new_n8238);
nor_5  g05890(new_n8238, new_n8236, new_n8239);
and_5  g05891(new_n8238, new_n8236, new_n8240);
not_10 g05892(n2420, new_n8241);
xnor_4 g05893(n24032, n22173, new_n8242);
xor_4  g05894(new_n8242, new_n8184, new_n8243);
and_5  g05895(new_n8243, new_n8241, new_n8244_1);
nor_5  g05896(new_n2549, new_n2548, new_n8245);
not_10 g05897(new_n8245, new_n8246);
xor_4  g05898(new_n8243, new_n8241, new_n8247);
and_5  g05899(new_n8247, new_n8246, new_n8248);
nor_5  g05900(new_n8248, new_n8244_1, new_n8249);
not_10 g05901(new_n8249, new_n8250);
nor_5  g05902(new_n8250, new_n8240, new_n8251);
nor_5  g05903(new_n8251, new_n8239, new_n8252);
not_10 g05904(new_n8252, new_n8253);
or_5   g05905(new_n8253, new_n8235, new_n8254);
and_5  g05906(new_n8254, new_n8233, new_n8255_1);
or_5   g05907(new_n8255_1, new_n8231, new_n8256_1);
and_5  g05908(new_n8256_1, new_n8229, new_n8257);
or_5   g05909(new_n8257, new_n8227, new_n8258);
and_5  g05910(new_n8258, new_n8225, new_n8259_1);
or_5   g05911(new_n8259_1, new_n8223, new_n8260);
and_5  g05912(new_n8260, new_n8221, new_n8261);
or_5   g05913(new_n8261, new_n8219, new_n8262);
and_5  g05914(new_n8262, new_n8217, new_n8263);
or_5   g05915(new_n8263, new_n8215_1, new_n8264);
and_5  g05916(new_n8264, new_n8213, new_n8265);
or_5   g05917(new_n8265, new_n8211, new_n8266);
and_5  g05918(new_n8266, new_n8209, new_n8267_1);
and_5  g05919(new_n8267_1, new_n8207, new_n8268);
xor_4  g05920(new_n8162, new_n8159_1, new_n8269);
xor_4  g05921(new_n8267_1, new_n8207, new_n8270);
or_5   g05922(new_n8270, new_n8269, new_n8271);
xor_4  g05923(new_n8270, new_n8269, new_n8272);
not_10 g05924(new_n8272, new_n8273);
xor_4  g05925(new_n8157, new_n8095_1, new_n8274);
xor_4  g05926(new_n8265, new_n8211, new_n8275);
nand_5 g05927(new_n8275, new_n8274, new_n8276_1);
not_10 g05928(new_n8274, new_n8277);
xnor_4 g05929(new_n8275, new_n8277, new_n8278);
xor_4  g05930(new_n8155, new_n8101, new_n8279);
xor_4  g05931(new_n8263, new_n8215_1, new_n8280);
nand_5 g05932(new_n8280, new_n8279, new_n8281);
not_10 g05933(new_n8279, new_n8282);
xnor_4 g05934(new_n8280, new_n8282, new_n8283);
xor_4  g05935(new_n8153, new_n8107, new_n8284);
xor_4  g05936(new_n8261, new_n8219, new_n8285_1);
nand_5 g05937(new_n8285_1, new_n8284, new_n8286);
not_10 g05938(new_n8284, new_n8287);
xnor_4 g05939(new_n8285_1, new_n8287, new_n8288_1);
xor_4  g05940(new_n8151, new_n8113, new_n8289);
xor_4  g05941(new_n8259_1, new_n8223, new_n8290);
nand_5 g05942(new_n8290, new_n8289, new_n8291);
not_10 g05943(new_n8289, new_n8292);
xnor_4 g05944(new_n8290, new_n8292, new_n8293);
xnor_4 g05945(new_n8149_1, new_n8118, new_n8294);
xor_4  g05946(new_n8257, new_n8227, new_n8295);
nand_5 g05947(new_n8295, new_n8294, new_n8296);
not_10 g05948(new_n8294, new_n8297);
xnor_4 g05949(new_n8295, new_n8297, new_n8298);
and_5  g05950(new_n8146, new_n8128, new_n8299);
xnor_4 g05951(new_n8299, new_n8124, new_n8300);
xor_4  g05952(new_n8255_1, new_n8231, new_n8301);
nand_5 g05953(new_n8301, new_n8300, new_n8302);
not_10 g05954(new_n8300, new_n8303);
xnor_4 g05955(new_n8301, new_n8303, new_n8304);
xor_4  g05956(new_n8145, new_n8129, new_n8305_1);
xnor_4 g05957(new_n8252, new_n8235, new_n8306_1);
nand_5 g05958(new_n8306_1, new_n8305_1, new_n8307);
not_10 g05959(new_n8305_1, new_n8308);
xnor_4 g05960(new_n8306_1, new_n8308, new_n8309_1);
xor_4  g05961(new_n8143, new_n8134, new_n8310);
xor_4  g05962(new_n8238, n24485, new_n8311);
xor_4  g05963(new_n8311, new_n8250, new_n8312);
or_5   g05964(new_n8312, new_n8310, new_n8313);
xnor_4 g05965(new_n8312, new_n8310, new_n8314);
xor_4  g05966(new_n8247, new_n8246, new_n8315);
not_10 g05967(new_n8315, new_n8316);
xnor_4 g05968(new_n8141, new_n8139_1, new_n8317);
not_10 g05969(new_n8317, new_n8318);
and_5  g05970(new_n8318, new_n8316, new_n8319);
and_5  g05971(new_n2550, new_n2547_1, new_n8320_1);
xor_4  g05972(new_n8318, new_n8316, new_n8321_1);
and_5  g05973(new_n8321_1, new_n8320_1, new_n8322);
nor_5  g05974(new_n8322, new_n8319, new_n8323);
not_10 g05975(new_n8323, new_n8324_1);
or_5   g05976(new_n8324_1, new_n8314, new_n8325);
nand_5 g05977(new_n8325, new_n8313, new_n8326);
nand_5 g05978(new_n8326, new_n8309_1, new_n8327);
nand_5 g05979(new_n8327, new_n8307, new_n8328);
nand_5 g05980(new_n8328, new_n8304, new_n8329);
nand_5 g05981(new_n8329, new_n8302, new_n8330);
nand_5 g05982(new_n8330, new_n8298, new_n8331);
nand_5 g05983(new_n8331, new_n8296, new_n8332);
nand_5 g05984(new_n8332, new_n8293, new_n8333);
nand_5 g05985(new_n8333, new_n8291, new_n8334);
nand_5 g05986(new_n8334, new_n8288_1, new_n8335);
nand_5 g05987(new_n8335, new_n8286, new_n8336);
nand_5 g05988(new_n8336, new_n8283, new_n8337);
nand_5 g05989(new_n8337, new_n8281, new_n8338);
nand_5 g05990(new_n8338, new_n8278, new_n8339_1);
and_5  g05991(new_n8339_1, new_n8276_1, new_n8340);
or_5   g05992(new_n8340, new_n8273, new_n8341);
and_5  g05993(new_n8341, new_n8271, new_n8342);
xor_4  g05994(new_n8342, new_n8268, new_n8343);
xor_4  g05995(new_n8343, new_n8163, n849);
xnor_4 g05996(new_n2534, new_n2533_1, n858);
not_10 g05997(n1314, new_n8346);
not_10 g05998(n3506, new_n8347);
not_10 g05999(n14899, new_n8348);
not_10 g06000(n18444, new_n8349);
not_10 g06001(n24638, new_n8350);
not_10 g06002(n21674, new_n8351);
not_10 g06003(n17251, new_n8352);
not_10 g06004(n14790, new_n8353);
nor_5  g06005(n16994, n9246, new_n8354);
and_5  g06006(new_n8354, new_n3556, new_n8355);
and_5  g06007(new_n8355, new_n8353, new_n8356);
and_5  g06008(new_n8356, new_n8352, new_n8357);
and_5  g06009(new_n8357, new_n8351, new_n8358);
and_5  g06010(new_n8358, new_n8350, new_n8359);
and_5  g06011(new_n8359, new_n8349, new_n8360);
and_5  g06012(new_n8360, new_n8348, new_n8361);
xor_4  g06013(new_n8361, new_n8347, new_n8362);
not_10 g06014(new_n8362, new_n8363_1);
xor_4  g06015(new_n8363_1, new_n8346, new_n8364);
not_10 g06016(n3306, new_n8365);
xor_4  g06017(new_n8360, new_n8348, new_n8366);
not_10 g06018(new_n8366, new_n8367);
or_5   g06019(new_n8367, new_n8365, new_n8368);
nand_5 g06020(new_n8367, new_n8365, new_n8369);
xor_4  g06021(new_n8359, new_n8349, new_n8370);
nor_5  g06022(new_n8370, n22335, new_n8371);
not_10 g06023(n22335, new_n8372);
xor_4  g06024(new_n8370, new_n8372, new_n8373);
xor_4  g06025(new_n8358, new_n8350, new_n8374);
or_5   g06026(new_n8374, n24048, new_n8375);
not_10 g06027(n24048, new_n8376_1);
xor_4  g06028(new_n8374, new_n8376_1, new_n8377);
xor_4  g06029(new_n8357, new_n8351, new_n8378);
or_5   g06030(new_n8378, n1525, new_n8379);
xnor_4 g06031(new_n8378, n1525, new_n8380);
xor_4  g06032(new_n8356, new_n8352, new_n8381_1);
or_5   g06033(new_n8381_1, n16988, new_n8382);
xor_4  g06034(new_n8381_1, n16988, new_n8383);
not_10 g06035(new_n8383, new_n8384);
xor_4  g06036(new_n8355, new_n8353, new_n8385);
or_5   g06037(new_n8385, n21779, new_n8386);
xor_4  g06038(new_n8354, new_n3556, new_n8387);
nor_5  g06039(new_n8387, n5376, new_n8388);
xor_4  g06040(new_n8387, new_n4650, new_n8389);
xor_4  g06041(n16994, n9246, new_n8390);
or_5   g06042(new_n8390, n5128, new_n8391);
nand_5 g06043(n23120, n9246, new_n8392);
xor_4  g06044(new_n8390, n5128, new_n8393);
nand_5 g06045(new_n8393, new_n8392, new_n8394);
and_5  g06046(new_n8394, new_n8391, new_n8395);
nor_5  g06047(new_n8395, new_n8389, new_n8396);
or_5   g06048(new_n8396, new_n8388, new_n8397);
xor_4  g06049(new_n8385, n21779, new_n8398);
nand_5 g06050(new_n8398, new_n8397, new_n8399_1);
and_5  g06051(new_n8399_1, new_n8386, new_n8400);
or_5   g06052(new_n8400, new_n8384, new_n8401);
and_5  g06053(new_n8401, new_n8382, new_n8402);
or_5   g06054(new_n8402, new_n8380, new_n8403);
and_5  g06055(new_n8403, new_n8379, new_n8404);
or_5   g06056(new_n8404, new_n8377, new_n8405_1);
and_5  g06057(new_n8405_1, new_n8375, new_n8406);
nor_5  g06058(new_n8406, new_n8373, new_n8407);
nor_5  g06059(new_n8407, new_n8371, new_n8408_1);
nand_5 g06060(new_n8408_1, new_n8369, new_n8409);
and_5  g06061(new_n8409, new_n8368, new_n8410);
xor_4  g06062(new_n8410, new_n8364, new_n8411);
or_5   g06063(new_n8411, n22442, new_n8412);
xor_4  g06064(new_n8411, n22442, new_n8413);
not_10 g06065(n468, new_n8414);
and_5  g06066(new_n8369, new_n8368, new_n8415);
xor_4  g06067(new_n8415, new_n8408_1, new_n8416);
or_5   g06068(new_n8416, new_n8414, new_n8417_1);
xor_4  g06069(new_n8416, new_n8414, new_n8418);
xor_4  g06070(new_n8406, new_n8373, new_n8419);
or_5   g06071(new_n8419, n5400, new_n8420);
not_10 g06072(n5400, new_n8421);
xor_4  g06073(new_n8419, new_n8421, new_n8422);
xor_4  g06074(new_n8404, new_n8377, new_n8423);
or_5   g06075(new_n8423, n23923, new_n8424);
xor_4  g06076(new_n8423, n23923, new_n8425);
xor_4  g06077(new_n8402, new_n8380, new_n8426);
nand_5 g06078(new_n8426, n329, new_n8427);
nor_5  g06079(new_n8426, n329, new_n8428);
xor_4  g06080(new_n8398, new_n8397, new_n8429);
or_5   g06081(new_n8429, n2409, new_n8430);
not_10 g06082(n2409, new_n8431);
xor_4  g06083(new_n8429, new_n8431, new_n8432_1);
xor_4  g06084(new_n8395, new_n8389, new_n8433);
or_5   g06085(new_n8433, n8869, new_n8434);
xor_4  g06086(new_n8393, new_n8392, new_n8435);
nor_5  g06087(new_n8435, n10372, new_n8436);
not_10 g06088(n7428, new_n8437);
xor_4  g06089(n23120, n9246, new_n8438);
or_5   g06090(new_n8438, new_n8437, new_n8439_1);
xor_4  g06091(new_n8435, n10372, new_n8440);
and_5  g06092(new_n8440, new_n8439_1, new_n8441);
or_5   g06093(new_n8441, new_n8436, new_n8442);
xor_4  g06094(new_n8433, n8869, new_n8443);
nand_5 g06095(new_n8443, new_n8442, new_n8444);
and_5  g06096(new_n8444, new_n8434, new_n8445);
or_5   g06097(new_n8445, new_n8432_1, new_n8446);
and_5  g06098(new_n8446, new_n8430, new_n8447);
nor_5  g06099(new_n8447, n24170, new_n8448);
xor_4  g06100(new_n8400, new_n8383, new_n8449);
xor_4  g06101(new_n8447, n24170, new_n8450);
and_5  g06102(new_n8450, new_n8449, new_n8451);
or_5   g06103(new_n8451, new_n8448, new_n8452);
or_5   g06104(new_n8452, new_n8428, new_n8453_1);
and_5  g06105(new_n8453_1, new_n8427, new_n8454);
nand_5 g06106(new_n8454, new_n8425, new_n8455);
and_5  g06107(new_n8455, new_n8424, new_n8456);
or_5   g06108(new_n8456, new_n8422, new_n8457);
and_5  g06109(new_n8457, new_n8420, new_n8458);
nand_5 g06110(new_n8458, new_n8418, new_n8459);
and_5  g06111(new_n8459, new_n8417_1, new_n8460);
nand_5 g06112(new_n8460, new_n8413, new_n8461);
and_5  g06113(new_n8461, new_n8412, new_n8462);
and_5  g06114(new_n8363_1, new_n8346, new_n8463);
or_5   g06115(new_n8410, new_n8463, new_n8464);
nand_5 g06116(new_n8361, new_n8347, new_n8465);
or_5   g06117(new_n8363_1, new_n8346, new_n8466);
and_5  g06118(new_n8466, new_n8465, new_n8467);
and_5  g06119(new_n8467, new_n8464, new_n8468);
xor_4  g06120(new_n8468, new_n8462, new_n8469);
and_5  g06121(new_n3471, new_n3407, new_n8470);
nor_5  g06122(new_n3528_1, new_n3473, new_n8471);
nor_5  g06123(new_n8471, new_n8470, new_n8472);
nand_5 g06124(new_n3423, new_n3409, new_n8473);
nor_5  g06125(new_n3424, n25494, new_n8474);
and_5  g06126(new_n3424, n25494, new_n8475);
nor_5  g06127(new_n3470, new_n8475, new_n8476);
or_5   g06128(new_n8476, new_n8474, new_n8477);
and_5  g06129(new_n8477, new_n8473, new_n8478);
xor_4  g06130(new_n8478, new_n8472, new_n8479);
xor_4  g06131(new_n8479, new_n8469, new_n8480_1);
xor_4  g06132(new_n8460, new_n8413, new_n8481);
nor_5  g06133(new_n8481, new_n3530, new_n8482);
xor_4  g06134(new_n8481, new_n3529, new_n8483);
xor_4  g06135(new_n8458, new_n8418, new_n8484);
and_5  g06136(new_n8484, new_n3662, new_n8485);
xor_4  g06137(new_n8484, new_n3663, new_n8486);
not_10 g06138(new_n3667, new_n8487);
xor_4  g06139(new_n8456, new_n8422, new_n8488);
nor_5  g06140(new_n8488, new_n8487, new_n8489_1);
not_10 g06141(new_n8489_1, new_n8490);
xor_4  g06142(new_n8488, new_n3667, new_n8491);
not_10 g06143(new_n3672, new_n8492);
xor_4  g06144(new_n8454, new_n8425, new_n8493);
nor_5  g06145(new_n8493, new_n8492, new_n8494);
not_10 g06146(new_n3677, new_n8495);
xor_4  g06147(new_n8426, n329, new_n8496);
xor_4  g06148(new_n8496, new_n8452, new_n8497);
or_5   g06149(new_n8497, new_n8495, new_n8498);
xor_4  g06150(new_n8497, new_n3677, new_n8499);
xor_4  g06151(new_n8450, new_n8449, new_n8500);
or_5   g06152(new_n8500, new_n3685, new_n8501);
xor_4  g06153(new_n8445, new_n8432_1, new_n8502);
or_5   g06154(new_n8502, new_n3690, new_n8503);
xor_4  g06155(new_n8502, new_n3690, new_n8504);
xor_4  g06156(new_n8443, new_n8442, new_n8505_1);
or_5   g06157(new_n8505_1, new_n3693, new_n8506);
xor_4  g06158(new_n8440, new_n8439_1, new_n8507);
or_5   g06159(new_n8507, new_n3701, new_n8508);
not_10 g06160(new_n3703, new_n8509);
xor_4  g06161(new_n8438, new_n8437, new_n8510_1);
nor_5  g06162(new_n8510_1, new_n8509, new_n8511);
xor_4  g06163(new_n8507, new_n3701, new_n8512);
not_10 g06164(new_n8512, new_n8513);
or_5   g06165(new_n8513, new_n8511, new_n8514);
and_5  g06166(new_n8514, new_n8508, new_n8515);
xor_4  g06167(new_n8505_1, new_n3693, new_n8516);
not_10 g06168(new_n8516, new_n8517);
or_5   g06169(new_n8517, new_n8515, new_n8518);
nand_5 g06170(new_n8518, new_n8506, new_n8519_1);
nand_5 g06171(new_n8519_1, new_n8504, new_n8520);
and_5  g06172(new_n8520, new_n8503, new_n8521);
xor_4  g06173(new_n8500, new_n3682, new_n8522);
or_5   g06174(new_n8522, new_n8521, new_n8523);
and_5  g06175(new_n8523, new_n8501, new_n8524);
or_5   g06176(new_n8524, new_n8499, new_n8525);
and_5  g06177(new_n8525, new_n8498, new_n8526_1);
xor_4  g06178(new_n8493, new_n3672, new_n8527);
or_5   g06179(new_n8527, new_n8526_1, new_n8528);
not_10 g06180(new_n8528, new_n8529);
nor_5  g06181(new_n8529, new_n8494, new_n8530);
or_5   g06182(new_n8530, new_n8491, new_n8531);
and_5  g06183(new_n8531, new_n8490, new_n8532);
or_5   g06184(new_n8532, new_n8486, new_n8533);
not_10 g06185(new_n8533, new_n8534);
nor_5  g06186(new_n8534, new_n8485, new_n8535_1);
or_5   g06187(new_n8535_1, new_n8483, new_n8536);
not_10 g06188(new_n8536, new_n8537);
nor_5  g06189(new_n8537, new_n8482, new_n8538);
xor_4  g06190(new_n8538, new_n8480_1, n873);
xor_4  g06191(n4812, n2731, new_n8540);
or_5   g06192(new_n3189, n19911, new_n8541);
xnor_4 g06193(n24278, n19911, new_n8542);
or_5   g06194(n24618, new_n3819, new_n8543);
or_5   g06195(new_n3190, n13708, new_n8544);
and_5  g06196(n18409, new_n3241, new_n8545);
and_5  g06197(new_n3821, n3952, new_n8546);
not_10 g06198(new_n8546, new_n8547);
not_10 g06199(n12315, new_n8548);
and_5  g06200(new_n8548, n5704, new_n8549);
and_5  g06201(new_n8549, new_n8547, new_n8550_1);
nor_5  g06202(new_n8550_1, new_n8545, new_n8551);
not_10 g06203(new_n8551, new_n8552);
nand_5 g06204(new_n8552, new_n8544, new_n8553);
and_5  g06205(new_n8553, new_n8543, new_n8554);
nand_5 g06206(new_n8554, new_n8542, new_n8555);
and_5  g06207(new_n8555, new_n8541, new_n8556);
xor_4  g06208(new_n8556, new_n8540, new_n8557);
xor_4  g06209(new_n8557, new_n5207, new_n8558);
xor_4  g06210(new_n8554, new_n8542, new_n8559);
or_5   g06211(new_n8559, new_n5211_1, new_n8560);
xnor_4 g06212(n24618, n13708, new_n8561);
xor_4  g06213(new_n8561, new_n8552, new_n8562);
nor_5  g06214(new_n8562, new_n5216, new_n8563_1);
xnor_4 g06215(new_n8562, new_n5216, new_n8564);
xnor_4 g06216(n12315, n5704, new_n8565);
nor_5  g06217(new_n8565, new_n5224, new_n8566);
nand_5 g06218(new_n8566, new_n5229, new_n8567);
xnor_4 g06219(new_n8566, new_n5229, new_n8568);
xnor_4 g06220(n18409, n3952, new_n8569);
xor_4  g06221(new_n8569, new_n8549, new_n8570);
or_5   g06222(new_n8570, new_n8568, new_n8571);
and_5  g06223(new_n8571, new_n8567, new_n8572);
nor_5  g06224(new_n8572, new_n8564, new_n8573);
nor_5  g06225(new_n8573, new_n8563_1, new_n8574);
xor_4  g06226(new_n8559, new_n5211_1, new_n8575);
nand_5 g06227(new_n8575, new_n8574, new_n8576);
and_5  g06228(new_n8576, new_n8560, new_n8577);
xor_4  g06229(new_n8577, new_n8558, n879);
xor_4  g06230(new_n8127_1, n18157, new_n8579);
or_5   g06231(new_n8132, n12161, new_n8580);
and_5  g06232(new_n8140, n5026, new_n8581_1);
and_5  g06233(new_n2546, n8581, new_n8582);
xor_4  g06234(new_n8140, n5026, new_n8583);
and_5  g06235(new_n8583, new_n8582, new_n8584);
nor_5  g06236(new_n8584, new_n8581_1, new_n8585);
xor_4  g06237(new_n8132, n12161, new_n8586);
nand_5 g06238(new_n8586, new_n8585, new_n8587);
and_5  g06239(new_n8587, new_n8580, new_n8588);
xnor_4 g06240(new_n8588, new_n8579, new_n8589);
xor_4  g06241(new_n8586, new_n8585, new_n8590);
not_10 g06242(new_n8590, new_n8591);
xor_4  g06243(new_n6649, n14684, new_n8592);
not_10 g06244(n6631, new_n8593);
nand_5 g06245(new_n6653, new_n8593, new_n8594_1);
nand_5 g06246(new_n6655_1, n24732, new_n8595);
xor_4  g06247(new_n6653, new_n8593, new_n8596);
nand_5 g06248(new_n8596, new_n8595, new_n8597);
and_5  g06249(new_n8597, new_n8594_1, new_n8598);
xor_4  g06250(new_n8598, new_n8592, new_n8599);
or_5   g06251(new_n8599, new_n8591, new_n8600);
xor_4  g06252(new_n8599, new_n8591, new_n8601);
not_10 g06253(new_n8601, new_n8602);
xor_4  g06254(new_n8596, new_n8595, new_n8603);
xor_4  g06255(new_n8583, new_n8582, new_n8604);
or_5   g06256(new_n8604, new_n8603, new_n8605);
xor_4  g06257(new_n6655_1, n24732, new_n8606);
not_10 g06258(new_n8606, new_n8607);
xor_4  g06259(new_n2546, n8581, new_n8608_1);
or_5   g06260(new_n8608_1, new_n8607, new_n8609);
xor_4  g06261(new_n8604, new_n8603, new_n8610);
not_10 g06262(new_n8610, new_n8611);
or_5   g06263(new_n8611, new_n8609, new_n8612);
and_5  g06264(new_n8612, new_n8605, new_n8613);
or_5   g06265(new_n8613, new_n8602, new_n8614_1);
and_5  g06266(new_n8614_1, new_n8600, new_n8615);
xor_4  g06267(new_n8615, new_n8589, new_n8616);
xor_4  g06268(new_n6645, new_n4166, new_n8617);
nand_5 g06269(new_n6649, new_n4167, new_n8618);
or_5   g06270(new_n8598, new_n8592, new_n8619);
and_5  g06271(new_n8619, new_n8618, new_n8620_1);
xor_4  g06272(new_n8620_1, new_n8617, new_n8621);
xor_4  g06273(new_n8621, new_n8616, n887);
xor_4  g06274(new_n6084_1, new_n4931, new_n8623);
not_10 g06275(new_n8623, new_n8624);
or_5   g06276(new_n6089, new_n4935, new_n8625);
xor_4  g06277(new_n6089, new_n4935, new_n8626);
not_10 g06278(new_n8626, new_n8627);
or_5   g06279(new_n6093, new_n4939_1, new_n8628);
xor_4  g06280(new_n6093, new_n4939_1, new_n8629);
not_10 g06281(new_n8629, new_n8630);
or_5   g06282(new_n6097, new_n4943, new_n8631);
xor_4  g06283(new_n6097, new_n4943, new_n8632);
not_10 g06284(new_n8632, new_n8633);
or_5   g06285(new_n6101, new_n4946, new_n8634);
not_10 g06286(n20259, new_n8635);
and_5  g06287(new_n6104_1, new_n8635, new_n8636);
and_5  g06288(new_n5851, n3925, new_n8637_1);
not_10 g06289(new_n8637_1, new_n8638_1);
xor_4  g06290(new_n6104_1, new_n8635, new_n8639);
and_5  g06291(new_n8639, new_n8638_1, new_n8640);
nor_5  g06292(new_n8640, new_n8636, new_n8641);
xor_4  g06293(new_n6101, new_n4946, new_n8642);
nand_5 g06294(new_n8642, new_n8641, new_n8643);
and_5  g06295(new_n8643, new_n8634, new_n8644);
or_5   g06296(new_n8644, new_n8633, new_n8645);
and_5  g06297(new_n8645, new_n8631, new_n8646);
or_5   g06298(new_n8646, new_n8630, new_n8647);
and_5  g06299(new_n8647, new_n8628, new_n8648);
or_5   g06300(new_n8648, new_n8627, new_n8649);
and_5  g06301(new_n8649, new_n8625, new_n8650);
xor_4  g06302(new_n8650, new_n8624, new_n8651);
not_10 g06303(n25119, new_n8652);
xor_4  g06304(new_n2958, new_n8652, new_n8653);
not_10 g06305(n1163, new_n8654);
or_5   g06306(new_n2964, new_n8654, new_n8655);
not_10 g06307(n18537, new_n8656_1);
nand_5 g06308(new_n2970, new_n8656_1, new_n8657);
xor_4  g06309(new_n2970, new_n8656_1, new_n8658);
not_10 g06310(new_n8658, new_n8659);
not_10 g06311(n7057, new_n8660);
nand_5 g06312(new_n2976, new_n8660, new_n8661);
xor_4  g06313(new_n2976, new_n8660, new_n8662_1);
not_10 g06314(n8381, new_n8663);
or_5   g06315(new_n2981, new_n8663, new_n8664);
xor_4  g06316(new_n2981, new_n8663, new_n8665);
and_5  g06317(new_n2991, n12495, new_n8666);
or_5   g06318(new_n8666, n20235, new_n8667);
xor_4  g06319(new_n8666, n20235, new_n8668);
nand_5 g06320(new_n8668, new_n2987, new_n8669);
and_5  g06321(new_n8669, new_n8667, new_n8670);
nand_5 g06322(new_n8670, new_n8665, new_n8671);
and_5  g06323(new_n8671, new_n8664, new_n8672);
nand_5 g06324(new_n8672, new_n8662_1, new_n8673);
and_5  g06325(new_n8673, new_n8661, new_n8674);
or_5   g06326(new_n8674, new_n8659, new_n8675);
and_5  g06327(new_n8675, new_n8657, new_n8676);
xor_4  g06328(new_n2964, new_n8654, new_n8677);
nand_5 g06329(new_n8677, new_n8676, new_n8678_1);
and_5  g06330(new_n8678_1, new_n8655, new_n8679);
xor_4  g06331(new_n8679, new_n8653, new_n8680);
xor_4  g06332(new_n8680, new_n8651, new_n8681);
not_10 g06333(new_n8681, new_n8682);
xor_4  g06334(new_n8648, new_n8627, new_n8683);
not_10 g06335(new_n8683, new_n8684);
xor_4  g06336(new_n8677, new_n8676, new_n8685);
nor_5  g06337(new_n8685, new_n8684, new_n8686);
xnor_4 g06338(new_n8685, new_n8683, new_n8687_1);
not_10 g06339(new_n8687_1, new_n8688);
xor_4  g06340(new_n8674, new_n8659, new_n8689);
xor_4  g06341(new_n8646, new_n8630, new_n8690);
and_5  g06342(new_n8690, new_n8689, new_n8691);
xor_4  g06343(new_n8690, new_n8689, new_n8692);
not_10 g06344(new_n8692, new_n8693);
xor_4  g06345(new_n8672, new_n8662_1, new_n8694_1);
xor_4  g06346(new_n8644, new_n8633, new_n8695);
and_5  g06347(new_n8695, new_n8694_1, new_n8696);
xor_4  g06348(new_n8695, new_n8694_1, new_n8697);
not_10 g06349(new_n8697, new_n8698);
xor_4  g06350(new_n8670, new_n8665, new_n8699);
not_10 g06351(new_n8699, new_n8700);
xor_4  g06352(new_n8642, new_n8641, new_n8701);
and_5  g06353(new_n8701, new_n8700, new_n8702);
not_10 g06354(new_n8702, new_n8703);
not_10 g06355(new_n8701, new_n8704);
xnor_4 g06356(new_n8704, new_n8700, new_n8705);
xor_4  g06357(new_n8639, new_n8638_1, new_n8706);
not_10 g06358(new_n8706, new_n8707);
xor_4  g06359(new_n8668, new_n2987, new_n8708);
and_5  g06360(new_n8708, new_n8707, new_n8709);
not_10 g06361(new_n8709, new_n8710);
xor_4  g06362(new_n5851, n3925, new_n8711);
xor_4  g06363(new_n2991, n12495, new_n8712);
not_10 g06364(new_n8712, new_n8713);
and_5  g06365(new_n8713, new_n8711, new_n8714);
xnor_4 g06366(new_n8708, new_n8706, new_n8715);
and_5  g06367(new_n8715, new_n8714, new_n8716_1);
not_10 g06368(new_n8716_1, new_n8717);
and_5  g06369(new_n8717, new_n8710, new_n8718);
not_10 g06370(new_n8718, new_n8719);
and_5  g06371(new_n8719, new_n8705, new_n8720);
not_10 g06372(new_n8720, new_n8721_1);
and_5  g06373(new_n8721_1, new_n8703, new_n8722);
nor_5  g06374(new_n8722, new_n8698, new_n8723);
nor_5  g06375(new_n8723, new_n8696, new_n8724);
nor_5  g06376(new_n8724, new_n8693, new_n8725);
nor_5  g06377(new_n8725, new_n8691, new_n8726);
nor_5  g06378(new_n8726, new_n8688, new_n8727);
nor_5  g06379(new_n8727, new_n8686, new_n8728);
xnor_4 g06380(new_n8728, new_n8682, n904);
nor_5  g06381(n18962, n10158, new_n8730);
and_5  g06382(new_n8730, new_n7532, new_n8731);
and_5  g06383(new_n8731, new_n7528, new_n8732);
xor_4  g06384(new_n8732, new_n7525, new_n8733);
xor_4  g06385(new_n8733, n21471, new_n8734);
xor_4  g06386(new_n8731, new_n7528, new_n8735);
nand_5 g06387(new_n8735, n18737, new_n8736);
xor_4  g06388(new_n8735, new_n5247, new_n8737);
xor_4  g06389(new_n8730, new_n7532, new_n8738);
nand_5 g06390(new_n8738, n14603, new_n8739);
xor_4  g06391(new_n8738, n14603, new_n8740);
xor_4  g06392(n18962, n10158, new_n8741);
or_5   g06393(new_n8741, n20794, new_n8742);
and_5  g06394(n23333, n18962, new_n8743);
not_10 g06395(new_n8743, new_n8744_1);
xor_4  g06396(new_n8741, n20794, new_n8745_1);
nand_5 g06397(new_n8745_1, new_n8744_1, new_n8746);
and_5  g06398(new_n8746, new_n8742, new_n8747);
nand_5 g06399(new_n8747, new_n8740, new_n8748);
and_5  g06400(new_n8748, new_n8739, new_n8749);
or_5   g06401(new_n8749, new_n8737, new_n8750);
and_5  g06402(new_n8750, new_n8736, new_n8751);
xor_4  g06403(new_n8751, new_n8734, new_n8752);
not_10 g06404(new_n8752, new_n8753);
xor_4  g06405(new_n8753, n19472, new_n8754);
xor_4  g06406(new_n8749, new_n8737, new_n8755);
or_5   g06407(new_n8755, n25370, new_n8756);
xor_4  g06408(new_n8747, new_n8740, new_n8757);
nand_5 g06409(new_n8757, n24786, new_n8758);
xor_4  g06410(new_n8757, n24786, new_n8759);
not_10 g06411(new_n8759, new_n8760);
xor_4  g06412(n23333, n18962, new_n8761);
and_5  g06413(new_n8761, n23065, new_n8762);
and_5  g06414(new_n8762, new_n8745_1, new_n8763);
not_10 g06415(new_n8763, new_n8764);
xor_4  g06416(new_n8745_1, new_n8743, new_n8765);
or_5   g06417(new_n8765, new_n8762, new_n8766);
and_5  g06418(new_n8766, new_n8764, new_n8767);
nand_5 g06419(new_n8767, n27120, new_n8768);
and_5  g06420(new_n8768, new_n8764, new_n8769);
or_5   g06421(new_n8769, new_n8760, new_n8770);
and_5  g06422(new_n8770, new_n8758, new_n8771);
xor_4  g06423(new_n8755, n25370, new_n8772);
nand_5 g06424(new_n8772, new_n8771, new_n8773);
and_5  g06425(new_n8773, new_n8756, new_n8774);
xor_4  g06426(new_n8774, new_n8754, new_n8775);
xor_4  g06427(new_n8775, new_n6728, new_n8776);
xor_4  g06428(new_n8772, new_n8771, new_n8777);
nand_5 g06429(new_n8777, new_n6733, new_n8778);
xnor_4 g06430(new_n8777, new_n6731, new_n8779);
not_10 g06431(new_n8779, new_n8780);
xor_4  g06432(new_n8767, n27120, new_n8781);
or_5   g06433(new_n8781, new_n6739, new_n8782_1);
xor_4  g06434(new_n8761, n23065, new_n8783);
and_5  g06435(new_n8783, new_n6736_1, new_n8784);
xnor_4 g06436(new_n8781, new_n6739, new_n8785);
or_5   g06437(new_n8785, new_n8784, new_n8786);
and_5  g06438(new_n8786, new_n8782_1, new_n8787);
or_5   g06439(new_n8787, new_n6747, new_n8788);
xor_4  g06440(new_n8769, new_n8760, new_n8789);
not_10 g06441(new_n8789, new_n8790);
xor_4  g06442(new_n8787, new_n6747, new_n8791);
nand_5 g06443(new_n8791, new_n8790, new_n8792);
and_5  g06444(new_n8792, new_n8788, new_n8793);
or_5   g06445(new_n8793, new_n8780, new_n8794);
and_5  g06446(new_n8794, new_n8778, new_n8795);
xor_4  g06447(new_n8795, new_n8776, n948);
xor_4  g06448(n25972, n10250, new_n8797);
not_10 g06449(n21915, new_n8798);
or_5   g06450(new_n8798, n7674, new_n8799);
xnor_4 g06451(n21915, n7674, new_n8800);
not_10 g06452(new_n8800, new_n8801);
not_10 g06453(n13775, new_n8802);
or_5   g06454(new_n8802, n6397, new_n8803_1);
xnor_4 g06455(n13775, n6397, new_n8804);
not_10 g06456(new_n8804, new_n8805);
not_10 g06457(n1293, new_n8806_1);
or_5   g06458(n19196, new_n8806_1, new_n8807);
xnor_4 g06459(n19196, n1293, new_n8808);
not_10 g06460(new_n8808, new_n8809_1);
not_10 g06461(n19042, new_n8810);
or_5   g06462(n23586, new_n8810, new_n8811);
xnor_4 g06463(n23586, n19042, new_n8812);
not_10 g06464(new_n8812, new_n8813);
not_10 g06465(n19472, new_n8814);
or_5   g06466(n21226, new_n8814, new_n8815);
xnor_4 g06467(n21226, n19472, new_n8816);
not_10 g06468(new_n8816, new_n8817);
not_10 g06469(n25370, new_n8818);
or_5   g06470(new_n8818, n4426, new_n8819);
xnor_4 g06471(n25370, n4426, new_n8820);
not_10 g06472(n20036, new_n8821_1);
or_5   g06473(n24786, new_n8821_1, new_n8822);
not_10 g06474(n24786, new_n8823);
or_5   g06475(new_n8823, n20036, new_n8824_1);
nor_5  g06476(n27120, new_n4122, new_n8825);
and_5  g06477(n27120, new_n4122, new_n8826);
not_10 g06478(new_n8826, new_n8827_1);
nor_5  g06479(n23065, new_n4125, new_n8828);
and_5  g06480(new_n8828, new_n8827_1, new_n8829);
nor_5  g06481(new_n8829, new_n8825, new_n8830);
not_10 g06482(new_n8830, new_n8831);
nand_5 g06483(new_n8831, new_n8824_1, new_n8832);
and_5  g06484(new_n8832, new_n8822, new_n8833);
nand_5 g06485(new_n8833, new_n8820, new_n8834);
and_5  g06486(new_n8834, new_n8819, new_n8835);
or_5   g06487(new_n8835, new_n8817, new_n8836);
and_5  g06488(new_n8836, new_n8815, new_n8837);
or_5   g06489(new_n8837, new_n8813, new_n8838);
and_5  g06490(new_n8838, new_n8811, new_n8839);
or_5   g06491(new_n8839, new_n8809_1, new_n8840);
and_5  g06492(new_n8840, new_n8807, new_n8841);
or_5   g06493(new_n8841, new_n8805, new_n8842);
and_5  g06494(new_n8842, new_n8803_1, new_n8843);
or_5   g06495(new_n8843, new_n8801, new_n8844);
and_5  g06496(new_n8844, new_n8799, new_n8845);
xor_4  g06497(new_n8845, new_n8797, new_n8846);
xnor_4 g06498(n20040, n2978, new_n8847);
not_10 g06499(new_n8847, new_n8848);
or_5   g06500(new_n7511, n19531, new_n8849_1);
xnor_4 g06501(n23697, n19531, new_n8850);
not_10 g06502(new_n8850, new_n8851);
or_5   g06503(n18345, new_n7515, new_n8852);
xnor_4 g06504(n18345, n2289, new_n8853);
not_10 g06505(new_n8853, new_n8854);
or_5   g06506(n13190, new_n7519, new_n8855);
xnor_4 g06507(n13190, n1112, new_n8856_1);
not_10 g06508(new_n8856_1, new_n8857);
or_5   g06509(new_n7522, n3460, new_n8858);
xnor_4 g06510(n20179, n3460, new_n8859);
not_10 g06511(new_n8859, new_n8860);
or_5   g06512(new_n7525, n5226, new_n8861_1);
xnor_4 g06513(n19228, n5226, new_n8862_1);
not_10 g06514(new_n8862_1, new_n8863);
or_5   g06515(n17664, new_n7528, new_n8864);
xnor_4 g06516(n17664, n15539, new_n8865);
not_10 g06517(n23369, new_n8866);
or_5   g06518(new_n8866, n8052, new_n8867);
or_5   g06519(n23369, new_n7532, new_n8868);
and_5  g06520(new_n7534, n1136, new_n8869_1);
not_10 g06521(n1136, new_n8870);
and_5  g06522(n10158, new_n8870, new_n8871);
and_5  g06523(n19234, new_n7538, new_n8872);
not_10 g06524(new_n8872, new_n8873);
nor_5  g06525(new_n8873, new_n8871, new_n8874);
nor_5  g06526(new_n8874, new_n8869_1, new_n8875);
not_10 g06527(new_n8875, new_n8876);
nand_5 g06528(new_n8876, new_n8868, new_n8877);
and_5  g06529(new_n8877, new_n8867, new_n8878);
nand_5 g06530(new_n8878, new_n8865, new_n8879);
and_5  g06531(new_n8879, new_n8864, new_n8880);
or_5   g06532(new_n8880, new_n8863, new_n8881);
and_5  g06533(new_n8881, new_n8861_1, new_n8882);
or_5   g06534(new_n8882, new_n8860, new_n8883);
and_5  g06535(new_n8883, new_n8858, new_n8884_1);
or_5   g06536(new_n8884_1, new_n8857, new_n8885);
and_5  g06537(new_n8885, new_n8855, new_n8886);
or_5   g06538(new_n8886, new_n8854, new_n8887);
and_5  g06539(new_n8887, new_n8852, new_n8888);
or_5   g06540(new_n8888, new_n8851, new_n8889);
and_5  g06541(new_n8889, new_n8849_1, new_n8890);
xor_4  g06542(new_n8890, new_n8848, new_n8891);
not_10 g06543(new_n8891, new_n8892);
not_10 g06544(n12507, new_n8893);
not_10 g06545(n22764, new_n8894);
nor_5  g06546(n15258, n4588, new_n8895);
and_5  g06547(new_n8895, new_n8130_1, new_n8896);
and_5  g06548(new_n8896, new_n8125, new_n8897);
and_5  g06549(new_n8897, new_n8120, new_n8898);
and_5  g06550(new_n8898, new_n8114, new_n8899);
and_5  g06551(new_n8899, new_n8108, new_n8900);
and_5  g06552(new_n8900, new_n8102, new_n8901);
and_5  g06553(new_n8901, new_n8096, new_n8902);
xor_4  g06554(new_n8902, new_n8894, new_n8903);
xor_4  g06555(new_n8903, new_n8893, new_n8904);
xor_4  g06556(new_n8901, new_n8096, new_n8905);
nand_5 g06557(new_n8905, n15077, new_n8906);
nor_5  g06558(new_n8905, n15077, new_n8907);
xor_4  g06559(new_n8900, new_n8102, new_n8908);
and_5  g06560(new_n8908, n3710, new_n8909_1);
nor_5  g06561(new_n8908, n3710, new_n8910);
xor_4  g06562(new_n8899, new_n8108, new_n8911_1);
nor_5  g06563(new_n8911_1, n26318, new_n8912);
not_10 g06564(n26318, new_n8913);
xor_4  g06565(new_n8911_1, new_n8913, new_n8914);
xor_4  g06566(new_n8898, new_n8114, new_n8915);
or_5   g06567(new_n8915, n26054, new_n8916);
not_10 g06568(n26054, new_n8917);
xor_4  g06569(new_n8915, new_n8917, new_n8918);
xor_4  g06570(new_n8897, new_n8120, new_n8919);
or_5   g06571(new_n8919, n19081, new_n8920_1);
not_10 g06572(n19081, new_n8921);
xor_4  g06573(new_n8919, new_n8921, new_n8922);
xor_4  g06574(new_n8896, new_n8125, new_n8923);
or_5   g06575(new_n8923, n8309, new_n8924);
xor_4  g06576(new_n8895, new_n8130_1, new_n8925);
nor_5  g06577(new_n8925, n19144, new_n8926);
xor_4  g06578(new_n8925, n19144, new_n8927);
not_10 g06579(new_n8927, new_n8928);
xor_4  g06580(n15258, n4588, new_n8929);
or_5   g06581(new_n8929, n12593, new_n8930);
nand_5 g06582(n13714, n4588, new_n8931);
xor_4  g06583(new_n8929, n12593, new_n8932);
nand_5 g06584(new_n8932, new_n8931, new_n8933);
and_5  g06585(new_n8933, new_n8930, new_n8934);
nor_5  g06586(new_n8934, new_n8928, new_n8935);
or_5   g06587(new_n8935, new_n8926, new_n8936);
xor_4  g06588(new_n8923, n8309, new_n8937);
nand_5 g06589(new_n8937, new_n8936, new_n8938);
and_5  g06590(new_n8938, new_n8924, new_n8939);
or_5   g06591(new_n8939, new_n8922, new_n8940);
and_5  g06592(new_n8940, new_n8920_1, new_n8941);
or_5   g06593(new_n8941, new_n8918, new_n8942);
and_5  g06594(new_n8942, new_n8916, new_n8943_1);
nor_5  g06595(new_n8943_1, new_n8914, new_n8944);
nor_5  g06596(new_n8944, new_n8912, new_n8945);
not_10 g06597(new_n8945, new_n8946);
nor_5  g06598(new_n8946, new_n8910, new_n8947);
nor_5  g06599(new_n8947, new_n8909_1, new_n8948);
or_5   g06600(new_n8948, new_n8907, new_n8949);
and_5  g06601(new_n8949, new_n8906, new_n8950);
xor_4  g06602(new_n8950, new_n8904, new_n8951);
xor_4  g06603(new_n8951, new_n8892, new_n8952);
xor_4  g06604(new_n8888, new_n8851, new_n8953);
not_10 g06605(n15077, new_n8954);
xor_4  g06606(new_n8905, new_n8954, new_n8955);
xor_4  g06607(new_n8955, new_n8948, new_n8956);
nand_5 g06608(new_n8956, new_n8953, new_n8957);
not_10 g06609(new_n8953, new_n8958);
xnor_4 g06610(new_n8956, new_n8958, new_n8959);
xor_4  g06611(new_n8886, new_n8854, new_n8960);
not_10 g06612(n3710, new_n8961);
xor_4  g06613(new_n8908, new_n8961, new_n8962);
xor_4  g06614(new_n8962, new_n8946, new_n8963);
or_5   g06615(new_n8963, new_n8960, new_n8964_1);
not_10 g06616(new_n8960, new_n8965);
xor_4  g06617(new_n8963, new_n8965, new_n8966);
xor_4  g06618(new_n8884_1, new_n8857, new_n8967);
not_10 g06619(new_n8967, new_n8968);
xor_4  g06620(new_n8943_1, new_n8914, new_n8969);
nand_5 g06621(new_n8969, new_n8968, new_n8970);
xor_4  g06622(new_n8969, new_n8967, new_n8971_1);
xor_4  g06623(new_n8882, new_n8860, new_n8972);
not_10 g06624(new_n8972, new_n8973);
xor_4  g06625(new_n8941, new_n8918, new_n8974);
nand_5 g06626(new_n8974, new_n8973, new_n8975);
xor_4  g06627(new_n8974, new_n8972, new_n8976);
xor_4  g06628(new_n8880, new_n8863, new_n8977);
not_10 g06629(new_n8977, new_n8978);
xor_4  g06630(new_n8939, new_n8922, new_n8979);
nand_5 g06631(new_n8979, new_n8978, new_n8980);
xor_4  g06632(new_n8979, new_n8978, new_n8981);
not_10 g06633(new_n8981, new_n8982_1);
xor_4  g06634(new_n8878, new_n8865, new_n8983);
not_10 g06635(new_n8983, new_n8984);
xor_4  g06636(new_n8937, new_n8936, new_n8985);
nand_5 g06637(new_n8985, new_n8984, new_n8986);
xor_4  g06638(new_n8985, new_n8984, new_n8987);
xor_4  g06639(new_n8934, new_n8928, new_n8988);
xnor_4 g06640(n23369, n8052, new_n8989);
xor_4  g06641(new_n8989, new_n8876, new_n8990);
or_5   g06642(new_n8990, new_n8988, new_n8991);
xor_4  g06643(new_n8990, new_n8988, new_n8992);
not_10 g06644(new_n8992, new_n8993_1);
xor_4  g06645(new_n8932, new_n8931, new_n8994);
xnor_4 g06646(n10158, n1136, new_n8995);
xnor_4 g06647(new_n8995, new_n8873, new_n8996);
or_5   g06648(new_n8996, new_n8994, new_n8997);
xnor_4 g06649(n19234, n18962, new_n8998);
not_10 g06650(new_n8998, new_n8999);
xor_4  g06651(n13714, n4588, new_n9000);
and_5  g06652(new_n9000, new_n8999, new_n9001);
xor_4  g06653(new_n8996, new_n8994, new_n9002);
nand_5 g06654(new_n9002, new_n9001, new_n9003_1);
and_5  g06655(new_n9003_1, new_n8997, new_n9004);
or_5   g06656(new_n9004, new_n8993_1, new_n9005);
and_5  g06657(new_n9005, new_n8991, new_n9006);
nand_5 g06658(new_n9006, new_n8987, new_n9007);
and_5  g06659(new_n9007, new_n8986, new_n9008);
or_5   g06660(new_n9008, new_n8982_1, new_n9009);
and_5  g06661(new_n9009, new_n8980, new_n9010);
or_5   g06662(new_n9010, new_n8976, new_n9011);
and_5  g06663(new_n9011, new_n8975, new_n9012_1);
or_5   g06664(new_n9012_1, new_n8971_1, new_n9013);
and_5  g06665(new_n9013, new_n8970, new_n9014);
or_5   g06666(new_n9014, new_n8966, new_n9015);
and_5  g06667(new_n9015, new_n8964_1, new_n9016);
nand_5 g06668(new_n9016, new_n8959, new_n9017);
and_5  g06669(new_n9017, new_n8957, new_n9018);
xor_4  g06670(new_n9018, new_n8952, new_n9019);
xor_4  g06671(new_n9019, new_n8846, new_n9020);
xor_4  g06672(new_n8843, new_n8801, new_n9021);
xor_4  g06673(new_n9016, new_n8959, new_n9022);
or_5   g06674(new_n9022, new_n9021, new_n9023);
xor_4  g06675(new_n9022, new_n9021, new_n9024);
not_10 g06676(new_n9024, new_n9025);
xor_4  g06677(new_n8841, new_n8805, new_n9026);
not_10 g06678(new_n9026, new_n9027);
xor_4  g06679(new_n9014, new_n8966, new_n9028);
nand_5 g06680(new_n9028, new_n9027, new_n9029);
xor_4  g06681(new_n9028, new_n9027, new_n9030);
not_10 g06682(new_n9030, new_n9031);
xor_4  g06683(new_n8839, new_n8809_1, new_n9032_1);
not_10 g06684(new_n9032_1, new_n9033);
xor_4  g06685(new_n9012_1, new_n8971_1, new_n9034);
nand_5 g06686(new_n9034, new_n9033, new_n9035);
xor_4  g06687(new_n9034, new_n9033, new_n9036);
not_10 g06688(new_n9036, new_n9037);
xor_4  g06689(new_n8837, new_n8813, new_n9038);
not_10 g06690(new_n9038, new_n9039);
xor_4  g06691(new_n9010, new_n8976, new_n9040);
nand_5 g06692(new_n9040, new_n9039, new_n9041);
xor_4  g06693(new_n9040, new_n9039, new_n9042_1);
not_10 g06694(new_n9042_1, new_n9043);
xor_4  g06695(new_n8835, new_n8817, new_n9044);
not_10 g06696(new_n9044, new_n9045);
xor_4  g06697(new_n9008, new_n8982_1, new_n9046_1);
nand_5 g06698(new_n9046_1, new_n9045, new_n9047_1);
xor_4  g06699(new_n9046_1, new_n9045, new_n9048);
not_10 g06700(new_n9048, new_n9049);
xor_4  g06701(new_n9006, new_n8987, new_n9050);
not_10 g06702(new_n9050, new_n9051);
xor_4  g06703(new_n8833, new_n8820, new_n9052);
or_5   g06704(new_n9052, new_n9051, new_n9053);
xor_4  g06705(new_n9052, new_n9051, new_n9054);
xor_4  g06706(new_n9004, new_n8993_1, new_n9055);
not_10 g06707(new_n9055, new_n9056);
xnor_4 g06708(n24786, n20036, new_n9057);
xor_4  g06709(new_n9057, new_n8831, new_n9058);
nand_5 g06710(new_n9058, new_n9056, new_n9059);
xnor_4 g06711(new_n9058, new_n9055, new_n9060);
not_10 g06712(new_n9060, new_n9061);
xnor_4 g06713(n23065, n9380, new_n9062);
xnor_4 g06714(new_n9000, new_n8998, new_n9063);
not_10 g06715(new_n9063, new_n9064);
nor_5  g06716(new_n9064, new_n9062, new_n9065);
xnor_4 g06717(n27120, n11192, new_n9066);
xnor_4 g06718(new_n9066, new_n8828, new_n9067);
or_5   g06719(new_n9067, new_n9065, new_n9068);
xor_4  g06720(new_n9002, new_n9001, new_n9069);
not_10 g06721(new_n9069, new_n9070);
xor_4  g06722(new_n9067, new_n9065, new_n9071);
nand_5 g06723(new_n9071, new_n9070, new_n9072);
and_5  g06724(new_n9072, new_n9068, new_n9073);
or_5   g06725(new_n9073, new_n9061, new_n9074);
nand_5 g06726(new_n9074, new_n9059, new_n9075);
nand_5 g06727(new_n9075, new_n9054, new_n9076);
and_5  g06728(new_n9076, new_n9053, new_n9077);
or_5   g06729(new_n9077, new_n9049, new_n9078);
and_5  g06730(new_n9078, new_n9047_1, new_n9079);
or_5   g06731(new_n9079, new_n9043, new_n9080);
and_5  g06732(new_n9080, new_n9041, new_n9081);
or_5   g06733(new_n9081, new_n9037, new_n9082);
and_5  g06734(new_n9082, new_n9035, new_n9083);
or_5   g06735(new_n9083, new_n9031, new_n9084);
and_5  g06736(new_n9084, new_n9029, new_n9085);
or_5   g06737(new_n9085, new_n9025, new_n9086);
and_5  g06738(new_n9086, new_n9023, new_n9087);
xor_4  g06739(new_n9087, new_n9020, n957);
xor_4  g06740(new_n8998, n20385, new_n9089);
not_10 g06741(n21138, new_n9090_1);
xor_4  g06742(n26167, n24129, new_n9091);
xor_4  g06743(new_n9091, new_n9090_1, new_n9092);
xor_4  g06744(new_n9092, new_n9089, n980);
and_5  g06745(new_n7832, new_n4350, new_n9094);
not_10 g06746(new_n9094, new_n9095);
xor_4  g06747(new_n7832, new_n4350, new_n9096);
or_5   g06748(new_n7837, new_n4354, new_n9097);
xor_4  g06749(new_n7837, new_n4354, new_n9098);
not_10 g06750(new_n9098, new_n9099);
or_5   g06751(new_n7842, new_n4358, new_n9100);
xnor_4 g06752(new_n7843, new_n4358, new_n9101);
not_10 g06753(new_n9101, new_n9102);
or_5   g06754(new_n7849, new_n4362, new_n9103);
xor_4  g06755(new_n7849, new_n4362, new_n9104_1);
not_10 g06756(new_n9104_1, new_n9105);
or_5   g06757(new_n7854, new_n4366, new_n9106);
xor_4  g06758(new_n7854, new_n4366, new_n9107);
not_10 g06759(new_n9107, new_n9108);
or_5   g06760(new_n7859, new_n4370, new_n9109);
xor_4  g06761(new_n7859, new_n4370, new_n9110);
not_10 g06762(new_n9110, new_n9111);
or_5   g06763(new_n7864, new_n4374_1, new_n9112);
xnor_4 g06764(new_n7865, new_n4374_1, new_n9113);
not_10 g06765(new_n9113, new_n9114);
nand_5 g06766(new_n7872, new_n4379, new_n9115);
xor_4  g06767(new_n7872, new_n4379, new_n9116);
or_5   g06768(new_n7879, new_n4384, new_n9117);
nor_5  g06769(new_n7883, new_n4387, new_n9118);
xor_4  g06770(new_n7879, new_n4384, new_n9119);
nand_5 g06771(new_n9119, new_n9118, new_n9120);
and_5  g06772(new_n9120, new_n9117, new_n9121);
nand_5 g06773(new_n9121, new_n9116, new_n9122);
and_5  g06774(new_n9122, new_n9115, new_n9123);
or_5   g06775(new_n9123, new_n9114, new_n9124);
and_5  g06776(new_n9124, new_n9112, new_n9125);
or_5   g06777(new_n9125, new_n9111, new_n9126);
and_5  g06778(new_n9126, new_n9109, new_n9127);
or_5   g06779(new_n9127, new_n9108, new_n9128);
and_5  g06780(new_n9128, new_n9106, new_n9129_1);
or_5   g06781(new_n9129_1, new_n9105, new_n9130);
and_5  g06782(new_n9130, new_n9103, new_n9131);
or_5   g06783(new_n9131, new_n9102, new_n9132);
and_5  g06784(new_n9132, new_n9100, new_n9133);
or_5   g06785(new_n9133, new_n9099, new_n9134);
and_5  g06786(new_n9134, new_n9097, new_n9135);
and_5  g06787(new_n9135, new_n9096, new_n9136);
not_10 g06788(new_n9136, new_n9137);
and_5  g06789(new_n9137, new_n9095, new_n9138);
xnor_4 g06790(new_n7829, new_n4349, new_n9139);
xor_4  g06791(new_n9139, new_n9138, new_n9140);
not_10 g06792(n12650, new_n9141);
and_5  g06793(n16544, new_n9141, new_n9142);
not_10 g06794(new_n9142, new_n9143);
xnor_4 g06795(n16544, n12650, new_n9144);
not_10 g06796(new_n9144, new_n9145);
not_10 g06797(n6814, new_n9146_1);
or_5   g06798(n10201, new_n9146_1, new_n9147);
xnor_4 g06799(n10201, n6814, new_n9148);
not_10 g06800(new_n9148, new_n9149);
not_10 g06801(n19701, new_n9150);
or_5   g06802(new_n9150, n10593, new_n9151);
xnor_4 g06803(n19701, n10593, new_n9152);
not_10 g06804(new_n9152, new_n9153);
not_10 g06805(n23529, new_n9154);
or_5   g06806(new_n9154, n18290, new_n9155);
xnor_4 g06807(n23529, n18290, new_n9156);
not_10 g06808(new_n9156, new_n9157);
not_10 g06809(n24620, new_n9158);
or_5   g06810(new_n9158, n11580, new_n9159);
xnor_4 g06811(n24620, n11580, new_n9160);
not_10 g06812(new_n9160, new_n9161);
not_10 g06813(n5211, new_n9162);
or_5   g06814(n15884, new_n9162, new_n9163);
xnor_4 g06815(n15884, n5211, new_n9164_1);
not_10 g06816(new_n9164_1, new_n9165);
not_10 g06817(n12956, new_n9166_1);
or_5   g06818(new_n9166_1, n6356, new_n9167);
xnor_4 g06819(n12956, n6356, new_n9168);
not_10 g06820(n27104, new_n9169);
or_5   g06821(new_n9169, n18295, new_n9170);
not_10 g06822(n18295, new_n9171);
or_5   g06823(n27104, new_n9171, new_n9172_1);
not_10 g06824(n6502, new_n9173);
and_5  g06825(n27188, new_n9173, new_n9174);
not_10 g06826(n27188, new_n9175);
and_5  g06827(new_n9175, n6502, new_n9176);
not_10 g06828(new_n9176, new_n9177);
not_10 g06829(n15780, new_n9178);
and_5  g06830(new_n9178, n6611, new_n9179);
and_5  g06831(new_n9179, new_n9177, new_n9180);
nor_5  g06832(new_n9180, new_n9174, new_n9181);
not_10 g06833(new_n9181, new_n9182_1);
nand_5 g06834(new_n9182_1, new_n9172_1, new_n9183);
and_5  g06835(new_n9183, new_n9170, new_n9184);
nand_5 g06836(new_n9184, new_n9168, new_n9185);
and_5  g06837(new_n9185, new_n9167, new_n9186);
or_5   g06838(new_n9186, new_n9165, new_n9187);
and_5  g06839(new_n9187, new_n9163, new_n9188);
or_5   g06840(new_n9188, new_n9161, new_n9189);
and_5  g06841(new_n9189, new_n9159, new_n9190);
or_5   g06842(new_n9190, new_n9157, new_n9191_1);
and_5  g06843(new_n9191_1, new_n9155, new_n9192);
or_5   g06844(new_n9192, new_n9153, new_n9193);
and_5  g06845(new_n9193, new_n9151, new_n9194);
or_5   g06846(new_n9194, new_n9149, new_n9195);
and_5  g06847(new_n9195, new_n9147, new_n9196);
nor_5  g06848(new_n9196, new_n9145, new_n9197);
not_10 g06849(new_n9197, new_n9198);
and_5  g06850(new_n9198, new_n9143, new_n9199);
xor_4  g06851(new_n9199, new_n9140, new_n9200);
xor_4  g06852(new_n9196, new_n9145, new_n9201);
xor_4  g06853(new_n9135, new_n9096, new_n9202);
nor_5  g06854(new_n9202, new_n9201, new_n9203);
xor_4  g06855(new_n9202, new_n9201, new_n9204);
not_10 g06856(new_n9204, new_n9205);
xor_4  g06857(new_n9194, new_n9149, new_n9206);
xor_4  g06858(new_n9133, new_n9099, new_n9207);
not_10 g06859(new_n9207, new_n9208);
nor_5  g06860(new_n9208, new_n9206, new_n9209);
not_10 g06861(new_n9209, new_n9210);
xor_4  g06862(new_n9208, new_n9206, new_n9211);
xor_4  g06863(new_n9192, new_n9153, new_n9212);
xor_4  g06864(new_n9131, new_n9102, new_n9213);
not_10 g06865(new_n9213, new_n9214);
nor_5  g06866(new_n9214, new_n9212, new_n9215);
not_10 g06867(new_n9215, new_n9216);
xor_4  g06868(new_n9214, new_n9212, new_n9217_1);
xor_4  g06869(new_n9190, new_n9157, new_n9218);
xor_4  g06870(new_n9129_1, new_n9105, new_n9219);
not_10 g06871(new_n9219, new_n9220_1);
nor_5  g06872(new_n9220_1, new_n9218, new_n9221);
not_10 g06873(new_n9221, new_n9222);
xor_4  g06874(new_n9220_1, new_n9218, new_n9223);
xor_4  g06875(new_n9188, new_n9161, new_n9224);
xor_4  g06876(new_n9127, new_n9108, new_n9225);
not_10 g06877(new_n9225, new_n9226);
nor_5  g06878(new_n9226, new_n9224, new_n9227);
not_10 g06879(new_n9227, new_n9228);
xor_4  g06880(new_n9226, new_n9224, new_n9229);
xor_4  g06881(new_n9186, new_n9165, new_n9230);
xor_4  g06882(new_n9125, new_n9111, new_n9231);
not_10 g06883(new_n9231, new_n9232);
nor_5  g06884(new_n9232, new_n9230, new_n9233);
not_10 g06885(new_n9233, new_n9234);
xor_4  g06886(new_n9232, new_n9230, new_n9235);
xor_4  g06887(new_n9123, new_n9114, new_n9236);
not_10 g06888(new_n9236, new_n9237);
xor_4  g06889(new_n9184, new_n9168, new_n9238);
nor_5  g06890(new_n9238, new_n9237, new_n9239);
not_10 g06891(new_n9239, new_n9240);
xor_4  g06892(new_n9121, new_n9116, new_n9241);
xnor_4 g06893(n27104, n18295, new_n9242);
xor_4  g06894(new_n9242, new_n9182_1, new_n9243);
and_5  g06895(new_n9243, new_n9241, new_n9244);
not_10 g06896(new_n9241, new_n9245);
xnor_4 g06897(new_n9243, new_n9245, new_n9246_1);
xnor_4 g06898(n15780, n6611, new_n9247);
xor_4  g06899(new_n7883, new_n4387, new_n9248);
not_10 g06900(new_n9248, new_n9249);
nor_5  g06901(new_n9249, new_n9247, new_n9250);
xnor_4 g06902(n27188, n6502, new_n9251_1);
xnor_4 g06903(new_n9251_1, new_n9179, new_n9252);
nor_5  g06904(new_n9252, new_n9250, new_n9253);
xor_4  g06905(new_n9119, new_n9118, new_n9254);
not_10 g06906(new_n9254, new_n9255);
xor_4  g06907(new_n9252, new_n9250, new_n9256);
and_5  g06908(new_n9256, new_n9255, new_n9257);
nor_5  g06909(new_n9257, new_n9253, new_n9258);
not_10 g06910(new_n9258, new_n9259_1);
and_5  g06911(new_n9259_1, new_n9246_1, new_n9260);
nor_5  g06912(new_n9260, new_n9244, new_n9261_1);
not_10 g06913(new_n9261_1, new_n9262);
xor_4  g06914(new_n9238, new_n9237, new_n9263);
and_5  g06915(new_n9263, new_n9262, new_n9264);
not_10 g06916(new_n9264, new_n9265);
and_5  g06917(new_n9265, new_n9240, new_n9266);
not_10 g06918(new_n9266, new_n9267);
and_5  g06919(new_n9267, new_n9235, new_n9268);
not_10 g06920(new_n9268, new_n9269);
and_5  g06921(new_n9269, new_n9234, new_n9270);
not_10 g06922(new_n9270, new_n9271);
and_5  g06923(new_n9271, new_n9229, new_n9272);
not_10 g06924(new_n9272, new_n9273);
and_5  g06925(new_n9273, new_n9228, new_n9274);
not_10 g06926(new_n9274, new_n9275);
and_5  g06927(new_n9275, new_n9223, new_n9276);
not_10 g06928(new_n9276, new_n9277);
and_5  g06929(new_n9277, new_n9222, new_n9278);
not_10 g06930(new_n9278, new_n9279);
and_5  g06931(new_n9279, new_n9217_1, new_n9280);
not_10 g06932(new_n9280, new_n9281);
and_5  g06933(new_n9281, new_n9216, new_n9282);
not_10 g06934(new_n9282, new_n9283);
and_5  g06935(new_n9283, new_n9211, new_n9284);
not_10 g06936(new_n9284, new_n9285);
and_5  g06937(new_n9285, new_n9210, new_n9286);
nor_5  g06938(new_n9286, new_n9205, new_n9287_1);
nor_5  g06939(new_n9287_1, new_n9203, new_n9288);
not_10 g06940(new_n9288, new_n9289);
xnor_4 g06941(new_n9289, new_n9200, n982);
not_10 g06942(n4306, new_n9291);
not_10 g06943(n3279, new_n9292);
not_10 g06944(n13914, new_n9293);
not_10 g06945(n14702, new_n9294);
not_10 g06946(n2999, new_n9295);
not_10 g06947(n2547, new_n9296);
not_10 g06948(n2680, new_n9297);
not_10 g06949(n1667, new_n9298);
nor_5  g06950(n26808, n7339, new_n9299);
and_5  g06951(new_n9299, new_n9298, new_n9300);
and_5  g06952(new_n9300, new_n9297, new_n9301);
and_5  g06953(new_n9301, new_n9296, new_n9302);
and_5  g06954(new_n9302, new_n9295, new_n9303);
and_5  g06955(new_n9303, new_n9294, new_n9304);
and_5  g06956(new_n9304, new_n9293, new_n9305);
and_5  g06957(new_n9305, new_n9292, new_n9306);
xor_4  g06958(new_n9306, new_n9291, new_n9307);
xor_4  g06959(n23166, n18105, new_n9308_1);
not_10 g06960(n10577, new_n9309);
or_5   g06961(n24196, new_n9309, new_n9310);
xor_4  g06962(n24196, n10577, new_n9311);
not_10 g06963(n6381, new_n9312);
or_5   g06964(n16376, new_n9312, new_n9313);
xor_4  g06965(n16376, n6381, new_n9314);
not_10 g06966(n14345, new_n9315);
or_5   g06967(n25381, new_n9315, new_n9316);
xor_4  g06968(n25381, n14345, new_n9317);
not_10 g06969(n11356, new_n9318_1);
or_5   g06970(n12587, new_n9318_1, new_n9319);
xor_4  g06971(n12587, n11356, new_n9320);
not_10 g06972(n3164, new_n9321);
or_5   g06973(new_n9321, n268, new_n9322);
xor_4  g06974(n3164, n268, new_n9323_1);
not_10 g06975(n10611, new_n9324);
or_5   g06976(n24879, new_n9324, new_n9325);
xnor_4 g06977(n24879, n10611, new_n9326);
or_5   g06978(new_n4456, n2783, new_n9327);
not_10 g06979(n2783, new_n9328);
or_5   g06980(n6785, new_n9328, new_n9329);
not_10 g06981(n15490, new_n9330);
and_5  g06982(n24032, new_n9330, new_n9331);
and_5  g06983(new_n8185, n15490, new_n9332);
not_10 g06984(n18, new_n9333);
and_5  g06985(n22843, new_n9333, new_n9334);
not_10 g06986(new_n9334, new_n9335);
nor_5  g06987(new_n9335, new_n9332, new_n9336);
nor_5  g06988(new_n9336, new_n9331, new_n9337);
not_10 g06989(new_n9337, new_n9338);
nand_5 g06990(new_n9338, new_n9329, new_n9339);
and_5  g06991(new_n9339, new_n9327, new_n9340);
nand_5 g06992(new_n9340, new_n9326, new_n9341);
and_5  g06993(new_n9341, new_n9325, new_n9342);
or_5   g06994(new_n9342, new_n9323_1, new_n9343);
and_5  g06995(new_n9343, new_n9322, new_n9344_1);
or_5   g06996(new_n9344_1, new_n9320, new_n9345);
and_5  g06997(new_n9345, new_n9319, new_n9346);
or_5   g06998(new_n9346, new_n9317, new_n9347);
and_5  g06999(new_n9347, new_n9316, new_n9348);
or_5   g07000(new_n9348, new_n9314, new_n9349);
and_5  g07001(new_n9349, new_n9313, new_n9350);
or_5   g07002(new_n9350, new_n9311, new_n9351);
and_5  g07003(new_n9351, new_n9310, new_n9352);
xor_4  g07004(new_n9352, new_n9308_1, new_n9353);
xnor_4 g07005(new_n9353, new_n9307, new_n9354);
xor_4  g07006(new_n9305, new_n9292, new_n9355);
xor_4  g07007(new_n9350, new_n9311, new_n9356);
nand_5 g07008(new_n9356, new_n9355, new_n9357);
xor_4  g07009(new_n9356, new_n9355, new_n9358);
xor_4  g07010(new_n9304, new_n9293, new_n9359);
xor_4  g07011(new_n9348, new_n9314, new_n9360);
or_5   g07012(new_n9360, new_n9359, new_n9361);
xnor_4 g07013(new_n9360, new_n9359, new_n9362);
xor_4  g07014(new_n9303, new_n9294, new_n9363);
xor_4  g07015(new_n9346, new_n9317, new_n9364_1);
or_5   g07016(new_n9364_1, new_n9363, new_n9365);
xnor_4 g07017(new_n9364_1, new_n9363, new_n9366);
xor_4  g07018(new_n9302, new_n9295, new_n9367);
xor_4  g07019(new_n9344_1, new_n9320, new_n9368);
or_5   g07020(new_n9368, new_n9367, new_n9369);
xor_4  g07021(new_n9301, new_n9296, new_n9370);
xor_4  g07022(new_n9342, new_n9323_1, new_n9371_1);
nor_5  g07023(new_n9371_1, new_n9370, new_n9372_1);
xnor_4 g07024(new_n9371_1, new_n9370, new_n9373);
xor_4  g07025(new_n9300, new_n9297, new_n9374);
xor_4  g07026(new_n9340, new_n9326, new_n9375);
or_5   g07027(new_n9375, new_n9374, new_n9376);
xor_4  g07028(new_n9299, n1667, new_n9377);
xnor_4 g07029(n6785, n2783, new_n9378);
xor_4  g07030(new_n9378, new_n9338, new_n9379);
and_5  g07031(new_n9379, new_n9377, new_n9380_1);
xor_4  g07032(new_n9379, new_n9377, new_n9381);
xnor_4 g07033(n26808, n7339, new_n9382_1);
xnor_4 g07034(n24032, n15490, new_n9383);
xnor_4 g07035(new_n9383, new_n9335, new_n9384);
or_5   g07036(new_n9384, new_n9382_1, new_n9385);
not_10 g07037(n26808, new_n9386);
xnor_4 g07038(n22843, n18, new_n9387);
nor_5  g07039(new_n9387, new_n9386, new_n9388);
xor_4  g07040(new_n9384, new_n9382_1, new_n9389);
nand_5 g07041(new_n9389, new_n9388, new_n9390);
and_5  g07042(new_n9390, new_n9385, new_n9391);
and_5  g07043(new_n9391, new_n9381, new_n9392);
or_5   g07044(new_n9392, new_n9380_1, new_n9393);
xor_4  g07045(new_n9375, new_n9374, new_n9394);
nand_5 g07046(new_n9394, new_n9393, new_n9395);
and_5  g07047(new_n9395, new_n9376, new_n9396_1);
nor_5  g07048(new_n9396_1, new_n9373, new_n9397);
or_5   g07049(new_n9397, new_n9372_1, new_n9398);
xor_4  g07050(new_n9368, new_n9367, new_n9399_1);
nand_5 g07051(new_n9399_1, new_n9398, new_n9400);
and_5  g07052(new_n9400, new_n9369, new_n9401);
or_5   g07053(new_n9401, new_n9366, new_n9402);
and_5  g07054(new_n9402, new_n9365, new_n9403_1);
or_5   g07055(new_n9403_1, new_n9362, new_n9404);
and_5  g07056(new_n9404, new_n9361, new_n9405);
nand_5 g07057(new_n9405, new_n9358, new_n9406);
and_5  g07058(new_n9406, new_n9357, new_n9407);
xor_4  g07059(new_n9407, new_n9354, new_n9408);
xor_4  g07060(new_n9408, new_n4538, new_n9409);
xor_4  g07061(new_n9405, new_n9358, new_n9410);
nor_5  g07062(new_n9410, new_n4543, new_n9411);
not_10 g07063(new_n9411, new_n9412);
xor_4  g07064(new_n9410, new_n4543, new_n9413);
xor_4  g07065(new_n9403_1, new_n9362, new_n9414);
and_5  g07066(new_n9414, new_n4548, new_n9415);
xor_4  g07067(new_n9414, new_n4548, new_n9416);
not_10 g07068(new_n9416, new_n9417);
xor_4  g07069(new_n9401, new_n9366, new_n9418);
and_5  g07070(new_n9418, new_n4553, new_n9419_1);
xor_4  g07071(new_n9418, new_n4553, new_n9420);
not_10 g07072(new_n9420, new_n9421);
xor_4  g07073(new_n9399_1, new_n9398, new_n9422);
and_5  g07074(new_n9422, new_n4558, new_n9423_1);
xor_4  g07075(new_n9422, new_n4558, new_n9424);
not_10 g07076(new_n9424, new_n9425);
xor_4  g07077(new_n9396_1, new_n9373, new_n9426);
and_5  g07078(new_n9426, new_n4562, new_n9427);
xor_4  g07079(new_n9426, new_n4562, new_n9428);
not_10 g07080(new_n9428, new_n9429);
xor_4  g07081(new_n9394, new_n9393, new_n9430_1);
and_5  g07082(new_n9430_1, new_n4568, new_n9431);
not_10 g07083(new_n9431, new_n9432);
xor_4  g07084(new_n9430_1, new_n4568, new_n9433);
xor_4  g07085(new_n9391, new_n9381, new_n9434);
nor_5  g07086(new_n9434, new_n4586, new_n9435_1);
xnor_4 g07087(new_n9434, new_n4586, new_n9436);
xor_4  g07088(new_n9389, new_n9388, new_n9437);
nand_5 g07089(new_n9437, new_n4582, new_n9438);
xor_4  g07090(new_n9387, new_n9386, new_n9439);
and_5  g07091(new_n9439, new_n4580, new_n9440);
xor_4  g07092(new_n9437, new_n4582, new_n9441);
nand_5 g07093(new_n9441, new_n9440, new_n9442);
and_5  g07094(new_n9442, new_n9438, new_n9443);
nor_5  g07095(new_n9443, new_n9436, new_n9444);
nor_5  g07096(new_n9444, new_n9435_1, new_n9445_1);
and_5  g07097(new_n9445_1, new_n9433, new_n9446);
not_10 g07098(new_n9446, new_n9447);
and_5  g07099(new_n9447, new_n9432, new_n9448);
nor_5  g07100(new_n9448, new_n9429, new_n9449);
nor_5  g07101(new_n9449, new_n9427, new_n9450);
nor_5  g07102(new_n9450, new_n9425, new_n9451_1);
nor_5  g07103(new_n9451_1, new_n9423_1, new_n9452);
nor_5  g07104(new_n9452, new_n9421, new_n9453);
nor_5  g07105(new_n9453, new_n9419_1, new_n9454);
nor_5  g07106(new_n9454, new_n9417, new_n9455);
nor_5  g07107(new_n9455, new_n9415, new_n9456);
not_10 g07108(new_n9456, new_n9457);
and_5  g07109(new_n9457, new_n9413, new_n9458_1);
not_10 g07110(new_n9458_1, new_n9459_1);
and_5  g07111(new_n9459_1, new_n9412, new_n9460_1);
xor_4  g07112(new_n9460_1, new_n9409, n984);
xnor_4 g07113(new_n9452, new_n9421, n1005);
xnor_4 g07114(new_n3388, new_n3337, n1016);
xor_4  g07115(new_n4104, new_n4089_1, n1020);
xor_4  g07116(n18290, n12875, new_n9465);
not_10 g07117(new_n9465, new_n9466);
or_5   g07118(n11580, n2035, new_n9467);
xor_4  g07119(n11580, n2035, new_n9468);
not_10 g07120(new_n9468, new_n9469);
or_5   g07121(n15884, n5213, new_n9470);
xor_4  g07122(n15884, n5213, new_n9471);
not_10 g07123(new_n9471, new_n9472);
or_5   g07124(n6356, n4665, new_n9473);
xor_4  g07125(n6356, n4665, new_n9474);
not_10 g07126(new_n9474, new_n9475);
or_5   g07127(n27104, n19005, new_n9476);
xor_4  g07128(n27104, n19005, new_n9477);
not_10 g07129(new_n9477, new_n9478);
or_5   g07130(n27188, n4326, new_n9479);
and_5  g07131(n6611, n5438, new_n9480);
not_10 g07132(new_n9480, new_n9481);
xor_4  g07133(n27188, n4326, new_n9482);
nand_5 g07134(new_n9482, new_n9481, new_n9483);
and_5  g07135(new_n9483, new_n9479, new_n9484);
or_5   g07136(new_n9484, new_n9478, new_n9485);
and_5  g07137(new_n9485, new_n9476, new_n9486);
or_5   g07138(new_n9486, new_n9475, new_n9487);
and_5  g07139(new_n9487, new_n9473, new_n9488);
or_5   g07140(new_n9488, new_n9472, new_n9489);
and_5  g07141(new_n9489, new_n9470, new_n9490);
or_5   g07142(new_n9490, new_n9469, new_n9491);
and_5  g07143(new_n9491, new_n9467, new_n9492);
xor_4  g07144(new_n9492, new_n9466, new_n9493_1);
not_10 g07145(new_n9493_1, new_n9494);
xor_4  g07146(new_n9494, n23529, new_n9495);
not_10 g07147(new_n9495, new_n9496);
xor_4  g07148(new_n9490, new_n9469, new_n9497);
not_10 g07149(new_n9497, new_n9498);
or_5   g07150(new_n9498, n24620, new_n9499);
xor_4  g07151(new_n9498, n24620, new_n9500);
not_10 g07152(new_n9500, new_n9501);
xor_4  g07153(new_n9488, new_n9472, new_n9502);
not_10 g07154(new_n9502, new_n9503);
or_5   g07155(new_n9503, n5211, new_n9504);
xor_4  g07156(new_n9503, n5211, new_n9505);
not_10 g07157(new_n9505, new_n9506);
xor_4  g07158(new_n9486, new_n9475, new_n9507_1);
not_10 g07159(new_n9507_1, new_n9508_1);
or_5   g07160(new_n9508_1, n12956, new_n9509);
xor_4  g07161(new_n9508_1, n12956, new_n9510);
xor_4  g07162(new_n9484, new_n9478, new_n9511);
not_10 g07163(new_n9511, new_n9512_1);
or_5   g07164(new_n9512_1, n18295, new_n9513);
xnor_4 g07165(new_n9482, new_n9480, new_n9514);
not_10 g07166(new_n9514, new_n9515);
and_5  g07167(new_n9515, n6502, new_n9516);
xor_4  g07168(n6611, n5438, new_n9517);
and_5  g07169(new_n9517, n15780, new_n9518);
xor_4  g07170(new_n9515, n6502, new_n9519);
and_5  g07171(new_n9519, new_n9518, new_n9520);
nor_5  g07172(new_n9520, new_n9516, new_n9521);
xor_4  g07173(new_n9512_1, n18295, new_n9522);
nand_5 g07174(new_n9522, new_n9521, new_n9523);
nand_5 g07175(new_n9523, new_n9513, new_n9524);
nand_5 g07176(new_n9524, new_n9510, new_n9525);
and_5  g07177(new_n9525, new_n9509, new_n9526);
or_5   g07178(new_n9526, new_n9506, new_n9527);
and_5  g07179(new_n9527, new_n9504, new_n9528);
or_5   g07180(new_n9528, new_n9501, new_n9529);
and_5  g07181(new_n9529, new_n9499, new_n9530);
xor_4  g07182(new_n9530, new_n9496, new_n9531);
xnor_4 g07183(n17250, n4409, new_n9532);
or_5   g07184(n23160, n3570, new_n9533);
xnor_4 g07185(n23160, n3570, new_n9534);
or_5   g07186(n16524, n13668, new_n9535);
xnor_4 g07187(n16524, n13668, new_n9536);
or_5   g07188(n21276, n11056, new_n9537);
xnor_4 g07189(n21276, n11056, new_n9538);
or_5   g07190(n26748, n15271, new_n9539);
xnor_4 g07191(n26748, n15271, new_n9540);
or_5   g07192(n25877, n10057, new_n9541);
and_5  g07193(n24323, n8920, new_n9542);
not_10 g07194(new_n9542, new_n9543);
xor_4  g07195(n25877, n10057, new_n9544);
nand_5 g07196(new_n9544, new_n9543, new_n9545);
and_5  g07197(new_n9545, new_n9541, new_n9546);
or_5   g07198(new_n9546, new_n9540, new_n9547);
and_5  g07199(new_n9547, new_n9539, new_n9548);
or_5   g07200(new_n9548, new_n9538, new_n9549);
and_5  g07201(new_n9549, new_n9537, new_n9550);
or_5   g07202(new_n9550, new_n9536, new_n9551);
and_5  g07203(new_n9551, new_n9535, new_n9552_1);
or_5   g07204(new_n9552_1, new_n9534, new_n9553);
and_5  g07205(new_n9553, new_n9533, new_n9554_1);
xor_4  g07206(new_n9554_1, new_n9532, new_n9555);
xor_4  g07207(new_n9555, new_n7789, new_n9556_1);
not_10 g07208(new_n9556_1, new_n9557_1);
xor_4  g07209(new_n9552_1, new_n9534, new_n9558_1);
or_5   g07210(new_n9558_1, new_n7792, new_n9559);
xor_4  g07211(new_n9558_1, new_n7792, new_n9560);
not_10 g07212(new_n9560, new_n9561);
xor_4  g07213(new_n9550, new_n9536, new_n9562);
or_5   g07214(new_n9562, new_n7795, new_n9563);
xor_4  g07215(new_n9562, new_n7795, new_n9564);
not_10 g07216(new_n9564, new_n9565);
xor_4  g07217(new_n9548, new_n9538, new_n9566);
or_5   g07218(new_n9566, new_n7798, new_n9567);
xor_4  g07219(new_n9566, new_n7798, new_n9568);
not_10 g07220(new_n9568, new_n9569);
xor_4  g07221(new_n9546, new_n9540, new_n9570);
or_5   g07222(new_n9570, new_n7803, new_n9571);
xnor_4 g07223(new_n9544, new_n9542, new_n9572);
and_5  g07224(new_n9572, new_n7805, new_n9573);
xor_4  g07225(n24323, n8920, new_n9574);
and_5  g07226(new_n9574, n6775, new_n9575);
not_10 g07227(new_n9575, new_n9576);
xor_4  g07228(new_n9572, new_n7805, new_n9577);
and_5  g07229(new_n9577, new_n9576, new_n9578);
nor_5  g07230(new_n9578, new_n9573, new_n9579);
xor_4  g07231(new_n9570, new_n7803, new_n9580);
nand_5 g07232(new_n9580, new_n9579, new_n9581);
and_5  g07233(new_n9581, new_n9571, new_n9582);
or_5   g07234(new_n9582, new_n9569, new_n9583);
and_5  g07235(new_n9583, new_n9567, new_n9584);
or_5   g07236(new_n9584, new_n9565, new_n9585);
and_5  g07237(new_n9585, new_n9563, new_n9586);
or_5   g07238(new_n9586, new_n9561, new_n9587);
and_5  g07239(new_n9587, new_n9559, new_n9588);
xor_4  g07240(new_n9588, new_n9557_1, new_n9589);
xor_4  g07241(new_n9589, new_n9531, new_n9590);
not_10 g07242(new_n9590, new_n9591);
xor_4  g07243(new_n9528, new_n9501, new_n9592);
xor_4  g07244(new_n9586, new_n9561, new_n9593);
and_5  g07245(new_n9593, new_n9592, new_n9594);
xor_4  g07246(new_n9593, new_n9592, new_n9595);
not_10 g07247(new_n9595, new_n9596);
xnor_4 g07248(new_n9526, new_n9505, new_n9597);
xor_4  g07249(new_n9584, new_n9565, new_n9598_1);
and_5  g07250(new_n9598_1, new_n9597, new_n9599);
xor_4  g07251(new_n9598_1, new_n9597, new_n9600);
not_10 g07252(new_n9600, new_n9601);
xor_4  g07253(new_n9524, new_n9510, new_n9602);
xor_4  g07254(new_n9582, new_n9569, new_n9603);
and_5  g07255(new_n9603, new_n9602, new_n9604);
xor_4  g07256(new_n9603, new_n9602, new_n9605);
not_10 g07257(new_n9605, new_n9606);
xor_4  g07258(new_n9522, new_n9521, new_n9607);
xor_4  g07259(new_n9580, new_n9579, new_n9608);
and_5  g07260(new_n9608, new_n9607, new_n9609);
not_10 g07261(new_n9608, new_n9610);
xnor_4 g07262(new_n9610, new_n9607, new_n9611);
xor_4  g07263(new_n9577, new_n9576, new_n9612);
xor_4  g07264(new_n9519, new_n9518, new_n9613);
nor_5  g07265(new_n9613, new_n9612, new_n9614);
xor_4  g07266(new_n9574, n6775, new_n9615);
not_10 g07267(new_n9615, new_n9616_1);
xor_4  g07268(new_n9517, n15780, new_n9617);
nor_5  g07269(new_n9617, new_n9616_1, new_n9618);
not_10 g07270(new_n9612, new_n9619);
xnor_4 g07271(new_n9613, new_n9619, new_n9620);
and_5  g07272(new_n9620, new_n9618, new_n9621);
nor_5  g07273(new_n9621, new_n9614, new_n9622_1);
not_10 g07274(new_n9622_1, new_n9623);
and_5  g07275(new_n9623, new_n9611, new_n9624);
nor_5  g07276(new_n9624, new_n9609, new_n9625);
nor_5  g07277(new_n9625, new_n9606, new_n9626_1);
nor_5  g07278(new_n9626_1, new_n9604, new_n9627);
nor_5  g07279(new_n9627, new_n9601, new_n9628);
nor_5  g07280(new_n9628, new_n9599, new_n9629);
nor_5  g07281(new_n9629, new_n9596, new_n9630);
nor_5  g07282(new_n9630, new_n9594, new_n9631);
xnor_4 g07283(new_n9631, new_n9591, n1044);
nor_5  g07284(n22619, n6775, new_n9633_1);
and_5  g07285(new_n9633_1, new_n7803, new_n9634);
xor_4  g07286(new_n9634, new_n7798, new_n9635_1);
xor_4  g07287(new_n9635_1, n7305, new_n9636);
not_10 g07288(new_n9636, new_n9637);
xor_4  g07289(new_n9633_1, new_n7803, new_n9638);
nand_5 g07290(new_n9638, n25872, new_n9639);
xor_4  g07291(new_n9638, new_n4946, new_n9640);
xor_4  g07292(n22619, n6775, new_n9641);
nand_5 g07293(new_n9641, n20259, new_n9642);
and_5  g07294(n6775, n3925, new_n9643);
xor_4  g07295(new_n9641, n20259, new_n9644);
nand_5 g07296(new_n9644, new_n9643, new_n9645);
and_5  g07297(new_n9645, new_n9642, new_n9646_1);
or_5   g07298(new_n9646_1, new_n9640, new_n9647);
and_5  g07299(new_n9647, new_n9639, new_n9648_1);
xor_4  g07300(new_n9648_1, new_n9637, new_n9649);
not_10 g07301(new_n9649, new_n9650);
nor_5  g07302(n9399, n2088, new_n9651);
and_5  g07303(new_n9651, new_n4322, new_n9652);
xor_4  g07304(new_n9652, new_n4319_1, new_n9653);
xor_4  g07305(new_n9653, n3480, new_n9654);
not_10 g07306(new_n9654, new_n9655_1);
xor_4  g07307(new_n9651, new_n4322, new_n9656);
nand_5 g07308(new_n9656, n16722, new_n9657);
xor_4  g07309(new_n9656, n16722, new_n9658);
not_10 g07310(new_n5841_1, new_n9659);
nand_5 g07311(new_n5846, new_n9659, new_n9660);
and_5  g07312(new_n9660, new_n5843, new_n9661);
nand_5 g07313(new_n9661, new_n9658, new_n9662);
and_5  g07314(new_n9662, new_n9657, new_n9663);
xor_4  g07315(new_n9663, new_n9655_1, new_n9664);
not_10 g07316(new_n9664, new_n9665);
xor_4  g07317(new_n9665, new_n9650, new_n9666);
xor_4  g07318(new_n9661, new_n9658, new_n9667);
xor_4  g07319(new_n9646_1, new_n9640, new_n9668);
nand_5 g07320(new_n9668, new_n9667, new_n9669);
not_10 g07321(new_n9667, new_n9670);
xnor_4 g07322(new_n9668, new_n9670, new_n9671);
xor_4  g07323(new_n9644, new_n9643, new_n9672);
not_10 g07324(new_n9672, new_n9673);
or_5   g07325(new_n9673, new_n5847, new_n9674);
xor_4  g07326(n6775, n3925, new_n9675);
and_5  g07327(new_n9675, new_n5830, new_n9676);
xnor_4 g07328(new_n9672, new_n5847, new_n9677);
nand_5 g07329(new_n9677, new_n9676, new_n9678);
nand_5 g07330(new_n9678, new_n9674, new_n9679);
nand_5 g07331(new_n9679, new_n9671, new_n9680);
and_5  g07332(new_n9680, new_n9669, new_n9681);
xnor_4 g07333(new_n9681, new_n9666, new_n9682);
not_10 g07334(new_n9682, new_n9683);
xor_4  g07335(n12956, n7057, new_n9684);
or_5   g07336(new_n9171, n8381, new_n9685);
or_5   g07337(n18295, new_n8663, new_n9686);
and_5  g07338(new_n5061, n6502, new_n9687);
and_5  g07339(n20235, new_n9173, new_n9688);
not_10 g07340(new_n9688, new_n9689_1);
and_5  g07341(n15780, new_n5062_1, new_n9690);
and_5  g07342(new_n9690, new_n9689_1, new_n9691);
nor_5  g07343(new_n9691, new_n9687, new_n9692);
not_10 g07344(new_n9692, new_n9693);
nand_5 g07345(new_n9693, new_n9686, new_n9694);
and_5  g07346(new_n9694, new_n9685, new_n9695_1);
xor_4  g07347(new_n9695_1, new_n9684, new_n9696);
xor_4  g07348(new_n9696, new_n9683, new_n9697);
and_5  g07349(new_n9678, new_n9674, new_n9698);
xnor_4 g07350(new_n9698, new_n9671, new_n9699_1);
not_10 g07351(new_n9699_1, new_n9700);
xnor_4 g07352(n18295, n8381, new_n9701);
xor_4  g07353(new_n9701, new_n9693, new_n9702);
nand_5 g07354(new_n9702, new_n9700, new_n9703);
xor_4  g07355(new_n9702, new_n9700, new_n9704);
xor_4  g07356(n15780, n12495, new_n9705);
xor_4  g07357(new_n9675, new_n5830, new_n9706);
nand_5 g07358(new_n9706, new_n9705, new_n9707);
xnor_4 g07359(n20235, n6502, new_n9708);
xor_4  g07360(new_n9708, new_n9690, new_n9709);
and_5  g07361(new_n9709, new_n9707, new_n9710);
xor_4  g07362(new_n9677, new_n9676, new_n9711);
not_10 g07363(new_n9711, new_n9712);
xor_4  g07364(new_n9709, new_n9707, new_n9713);
and_5  g07365(new_n9713, new_n9712, new_n9714);
or_5   g07366(new_n9714, new_n9710, new_n9715);
nand_5 g07367(new_n9715, new_n9704, new_n9716);
and_5  g07368(new_n9716, new_n9703, new_n9717);
xor_4  g07369(new_n9717, new_n9697, n1060);
xnor_4 g07370(new_n3386, new_n3342, n1069);
xor_4  g07371(n9832, n3959, new_n9720);
not_10 g07372(new_n9720, new_n9721);
or_5   g07373(n11566, n1558, new_n9722);
xnor_4 g07374(n11566, n1558, new_n9723);
or_5   g07375(n26744, n21749, new_n9724);
xor_4  g07376(n26744, n21749, new_n9725);
not_10 g07377(new_n9725, new_n9726_1);
or_5   g07378(n26625, n7769, new_n9727);
and_5  g07379(n21138, n14230, new_n9728);
xnor_4 g07380(n26625, n7769, new_n9729);
or_5   g07381(new_n9729, new_n9728, new_n9730);
and_5  g07382(new_n9730, new_n9727, new_n9731);
or_5   g07383(new_n9731, new_n9726_1, new_n9732);
and_5  g07384(new_n9732, new_n9724, new_n9733);
or_5   g07385(new_n9733, new_n9723, new_n9734);
and_5  g07386(new_n9734, new_n9722, new_n9735);
xor_4  g07387(new_n9735, new_n9721, new_n9736);
not_10 g07388(new_n9736, new_n9737);
not_10 g07389(n19575, new_n9738);
not_10 g07390(n15378, new_n9739);
not_10 g07391(n17095, new_n9740);
nor_5  g07392(n26167, n22591, new_n9741);
and_5  g07393(new_n9741, new_n9740, new_n9742);
and_5  g07394(new_n9742, new_n9739, new_n9743);
xor_4  g07395(new_n9743, new_n9738, new_n9744);
xor_4  g07396(new_n6816, n5226, new_n9745);
not_10 g07397(n17664, new_n9746);
or_5   g07398(new_n6820, new_n9746, new_n9747);
xor_4  g07399(new_n6820, new_n9746, new_n9748);
not_10 g07400(new_n9748, new_n9749);
or_5   g07401(new_n6824, new_n8866, new_n9750);
xor_4  g07402(new_n6824, new_n8866, new_n9751);
nand_5 g07403(new_n6830, new_n8870, new_n9752);
and_5  g07404(new_n6827, n19234, new_n9753_1);
not_10 g07405(new_n9753_1, new_n9754);
xor_4  g07406(new_n6830, new_n8870, new_n9755);
nand_5 g07407(new_n9755, new_n9754, new_n9756);
and_5  g07408(new_n9756, new_n9752, new_n9757);
nand_5 g07409(new_n9757, new_n9751, new_n9758);
and_5  g07410(new_n9758, new_n9750, new_n9759);
or_5   g07411(new_n9759, new_n9749, new_n9760);
and_5  g07412(new_n9760, new_n9747, new_n9761_1);
xor_4  g07413(new_n9761_1, new_n9745, new_n9762);
xnor_4 g07414(new_n9762, new_n9744, new_n9763_1);
xor_4  g07415(new_n9759, new_n9749, new_n9764);
xor_4  g07416(new_n9742, new_n9739, new_n9765);
or_5   g07417(new_n9765, new_n9764, new_n9766);
xor_4  g07418(new_n9765, new_n9764, new_n9767_1);
not_10 g07419(new_n9767_1, new_n9768);
xor_4  g07420(new_n9757, new_n9751, new_n9769);
xor_4  g07421(new_n9741, new_n9740, new_n9770);
or_5   g07422(new_n9770, new_n9769, new_n9771_1);
xor_4  g07423(new_n9770, new_n9769, new_n9772);
xor_4  g07424(new_n9755, new_n9754, new_n9773);
not_10 g07425(new_n9773, new_n9774);
and_5  g07426(new_n7247, n26167, new_n9775);
xor_4  g07427(new_n9775, n22591, new_n9776);
nand_5 g07428(new_n9776, new_n9774, new_n9777);
nand_5 g07429(new_n7246, n26167, new_n9778_1);
or_5   g07430(new_n9778_1, n22591, new_n9779);
and_5  g07431(new_n9779, new_n9777, new_n9780);
nand_5 g07432(new_n9780, new_n9772, new_n9781);
and_5  g07433(new_n9781, new_n9771_1, new_n9782);
or_5   g07434(new_n9782, new_n9768, new_n9783_1);
and_5  g07435(new_n9783_1, new_n9766, new_n9784);
xor_4  g07436(new_n9784, new_n9763_1, new_n9785);
xor_4  g07437(new_n9785, new_n9737, new_n9786);
xor_4  g07438(new_n9782, new_n9768, new_n9787);
xor_4  g07439(new_n9733, new_n9723, new_n9788);
not_10 g07440(new_n9788, new_n9789);
nand_5 g07441(new_n9789, new_n9787, new_n9790);
xor_4  g07442(new_n9789, new_n9787, new_n9791);
xnor_4 g07443(new_n9780, new_n9772, new_n9792);
xor_4  g07444(new_n9731, new_n9726_1, new_n9793);
and_5  g07445(new_n9793, new_n9792, new_n9794);
not_10 g07446(new_n9794, new_n9795);
xor_4  g07447(new_n9793, new_n9792, new_n9796);
xor_4  g07448(new_n9776, new_n9774, new_n9797);
xor_4  g07449(n26625, n7769, new_n9798);
xnor_4 g07450(new_n9798, new_n9728, new_n9799);
or_5   g07451(new_n9799, new_n9797, new_n9800);
and_5  g07452(new_n7248, new_n7244, new_n9801);
xor_4  g07453(new_n9799, new_n9797, new_n9802);
nand_5 g07454(new_n9802, new_n9801, new_n9803_1);
and_5  g07455(new_n9803_1, new_n9800, new_n9804);
and_5  g07456(new_n9804, new_n9796, new_n9805);
not_10 g07457(new_n9805, new_n9806);
and_5  g07458(new_n9806, new_n9795, new_n9807);
nand_5 g07459(new_n9807, new_n9791, new_n9808);
and_5  g07460(new_n9808, new_n9790, new_n9809);
xor_4  g07461(new_n9809, new_n9786, n1111);
not_10 g07462(n25475, new_n9811);
xor_4  g07463(new_n2596, new_n9811, new_n9812);
not_10 g07464(new_n9812, new_n9813);
not_10 g07465(n23849, new_n9814);
or_5   g07466(new_n2601, new_n9814, new_n9815);
xor_4  g07467(new_n2601, new_n9814, new_n9816);
not_10 g07468(new_n9816, new_n9817);
or_5   g07469(new_n2606, new_n4436, new_n9818);
not_10 g07470(n11011, new_n9819);
and_5  g07471(new_n2609, new_n9819, new_n9820);
xor_4  g07472(new_n2609, new_n9819, new_n9821);
not_10 g07473(new_n9821, new_n9822);
not_10 g07474(n16029, new_n9823);
nand_5 g07475(new_n2614, new_n9823, new_n9824);
xor_4  g07476(new_n2614, new_n9823, new_n9825);
not_10 g07477(n16476, new_n9826);
or_5   g07478(new_n2618, new_n9826, new_n9827);
xor_4  g07479(new_n2618, new_n9826, new_n9828);
not_10 g07480(new_n9828, new_n9829);
or_5   g07481(new_n2623, new_n5564_1, new_n9830);
not_10 g07482(n22433, new_n9831);
and_5  g07483(new_n2626, new_n9831, new_n9832_1);
and_5  g07484(new_n2628, n14090, new_n9833_1);
not_10 g07485(new_n9833_1, new_n9834);
xor_4  g07486(new_n2626, new_n9831, new_n9835);
and_5  g07487(new_n9835, new_n9834, new_n9836);
nor_5  g07488(new_n9836, new_n9832_1, new_n9837);
xor_4  g07489(new_n2623, new_n5564_1, new_n9838_1);
nand_5 g07490(new_n9838_1, new_n9837, new_n9839);
and_5  g07491(new_n9839, new_n9830, new_n9840);
or_5   g07492(new_n9840, new_n9829, new_n9841);
and_5  g07493(new_n9841, new_n9827, new_n9842);
nand_5 g07494(new_n9842, new_n9825, new_n9843);
and_5  g07495(new_n9843, new_n9824, new_n9844);
nor_5  g07496(new_n9844, new_n9822, new_n9845);
nor_5  g07497(new_n9845, new_n9820, new_n9846);
xor_4  g07498(new_n2606, new_n4436, new_n9847);
nand_5 g07499(new_n9847, new_n9846, new_n9848);
and_5  g07500(new_n9848, new_n9818, new_n9849);
or_5   g07501(new_n9849, new_n9817, new_n9850);
and_5  g07502(new_n9850, new_n9815, new_n9851);
xor_4  g07503(new_n9851, new_n9813, new_n9852);
and_5  g07504(new_n9652, new_n4319_1, new_n9853);
and_5  g07505(new_n9853, new_n4316, new_n9854);
and_5  g07506(new_n9854, new_n4313, new_n9855);
and_5  g07507(new_n9855, new_n4310, new_n9856);
and_5  g07508(new_n9856, new_n4307, new_n9857);
xor_4  g07509(new_n9857, new_n4304, new_n9858);
xor_4  g07510(new_n9858, new_n2715, new_n9859);
xor_4  g07511(new_n9856, new_n4307, new_n9860);
nand_5 g07512(new_n9860, new_n2718, new_n9861);
xnor_4 g07513(new_n9860, new_n2720, new_n9862);
xor_4  g07514(new_n9855, new_n4310, new_n9863);
or_5   g07515(new_n9863, new_n2723, new_n9864);
xor_4  g07516(new_n9863, new_n2725, new_n9865);
xor_4  g07517(new_n9854, new_n4313, new_n9866);
or_5   g07518(new_n9866, new_n2728, new_n9867_1);
xor_4  g07519(new_n9866, new_n2730, new_n9868);
xor_4  g07520(new_n9853, new_n4316, new_n9869);
or_5   g07521(new_n9869, new_n2733, new_n9870);
nor_5  g07522(new_n9653, new_n2737, new_n9871);
xnor_4 g07523(new_n9653, new_n2738, new_n9872_1);
or_5   g07524(new_n9656, new_n2743_1, new_n9873);
xnor_4 g07525(new_n9656, new_n2744, new_n9874);
nand_5 g07526(new_n9659, new_n2754, new_n9875);
and_5  g07527(new_n2752, new_n4329, new_n9876);
xor_4  g07528(new_n9659, new_n2754, new_n9877);
nand_5 g07529(new_n9877, new_n9876, new_n9878);
nand_5 g07530(new_n9878, new_n9875, new_n9879);
nand_5 g07531(new_n9879, new_n9874, new_n9880);
nand_5 g07532(new_n9880, new_n9873, new_n9881);
and_5  g07533(new_n9881, new_n9872_1, new_n9882);
or_5   g07534(new_n9882, new_n9871, new_n9883);
xnor_4 g07535(new_n9869, new_n2762, new_n9884);
nand_5 g07536(new_n9884, new_n9883, new_n9885);
and_5  g07537(new_n9885, new_n9870, new_n9886);
or_5   g07538(new_n9886, new_n9868, new_n9887);
and_5  g07539(new_n9887, new_n9867_1, new_n9888);
or_5   g07540(new_n9888, new_n9865, new_n9889);
and_5  g07541(new_n9889, new_n9864, new_n9890_1);
nand_5 g07542(new_n9890_1, new_n9862, new_n9891);
and_5  g07543(new_n9891, new_n9861, new_n9892);
xor_4  g07544(new_n9892, new_n9859, new_n9893);
xor_4  g07545(new_n9893, new_n9852, new_n9894);
xor_4  g07546(new_n9849, new_n9817, new_n9895);
xor_4  g07547(new_n9890_1, new_n9862, new_n9896);
and_5  g07548(new_n9896, new_n9895, new_n9897);
xor_4  g07549(new_n9896, new_n9895, new_n9898);
xor_4  g07550(new_n9847, new_n9846, new_n9899);
not_10 g07551(new_n9899, new_n9900);
xor_4  g07552(new_n9888, new_n9865, new_n9901);
nand_5 g07553(new_n9901, new_n9900, new_n9902);
xor_4  g07554(new_n9901, new_n9900, new_n9903);
xor_4  g07555(new_n9844, new_n9822, new_n9904);
xor_4  g07556(new_n9886, new_n9868, new_n9905);
nor_5  g07557(new_n9905, new_n9904, new_n9906);
xnor_4 g07558(new_n9905, new_n9904, new_n9907);
xor_4  g07559(new_n9842, new_n9825, new_n9908);
xor_4  g07560(new_n9884, new_n9883, new_n9909);
or_5   g07561(new_n9909, new_n9908, new_n9910);
not_10 g07562(new_n9908, new_n9911);
xor_4  g07563(new_n9909, new_n9911, new_n9912);
xor_4  g07564(new_n9881, new_n9872_1, new_n9913);
xor_4  g07565(new_n9840, new_n9829, new_n9914);
not_10 g07566(new_n9914, new_n9915);
or_5   g07567(new_n9915, new_n9913, new_n9916);
xor_4  g07568(new_n9914, new_n9913, new_n9917_1);
xnor_4 g07569(new_n9879, new_n9874, new_n9918);
xor_4  g07570(new_n9838_1, new_n9837, new_n9919_1);
nand_5 g07571(new_n9919_1, new_n9918, new_n9920);
not_10 g07572(new_n9919_1, new_n9921);
xnor_4 g07573(new_n9921, new_n9918, new_n9922);
xor_4  g07574(new_n9877, new_n9876, new_n9923);
xor_4  g07575(new_n9835, new_n9834, new_n9924);
nand_5 g07576(new_n9924, new_n9923, new_n9925);
xor_4  g07577(new_n2628, n14090, new_n9926_1);
not_10 g07578(new_n9926_1, new_n9927);
xor_4  g07579(new_n2752, new_n4329, new_n9928);
or_5   g07580(new_n9928, new_n9927, new_n9929);
not_10 g07581(new_n9924, new_n9930);
xnor_4 g07582(new_n9930, new_n9923, new_n9931);
nand_5 g07583(new_n9931, new_n9929, new_n9932);
and_5  g07584(new_n9932, new_n9925, new_n9933);
nand_5 g07585(new_n9933, new_n9922, new_n9934_1);
and_5  g07586(new_n9934_1, new_n9920, new_n9935);
or_5   g07587(new_n9935, new_n9917_1, new_n9936);
and_5  g07588(new_n9936, new_n9916, new_n9937);
or_5   g07589(new_n9937, new_n9912, new_n9938_1);
and_5  g07590(new_n9938_1, new_n9910, new_n9939);
nor_5  g07591(new_n9939, new_n9907, new_n9940);
nor_5  g07592(new_n9940, new_n9906, new_n9941);
nand_5 g07593(new_n9941, new_n9903, new_n9942_1);
and_5  g07594(new_n9942_1, new_n9902, new_n9943);
and_5  g07595(new_n9943, new_n9898, new_n9944);
nor_5  g07596(new_n9944, new_n9897, new_n9945);
xnor_4 g07597(new_n9945, new_n9894, n1119);
not_10 g07598(new_n8013, new_n9947);
xnor_4 g07599(new_n8014, new_n9947, new_n9948);
xor_4  g07600(new_n9948, new_n8034, n1120);
xor_4  g07601(n9246, n3925, new_n9950);
xnor_4 g07602(new_n9950, new_n7884_1, new_n9951);
not_10 g07603(new_n9951, new_n9952);
xnor_4 g07604(n12495, n7428, new_n9953);
xor_4  g07605(new_n9953, new_n9952, n1196);
xor_4  g07606(n16223, n15636, new_n9955);
or_5   g07607(new_n5567, n19494, new_n9956);
or_5   g07608(n20077, new_n2365, new_n9957);
and_5  g07609(n6794, new_n2370, new_n9958);
nand_5 g07610(new_n9958, new_n9957, new_n9959);
and_5  g07611(new_n9959, new_n9956, new_n9960);
xor_4  g07612(new_n9960, new_n9955, new_n9961);
xnor_4 g07613(new_n9961, new_n8018, new_n9962);
not_10 g07614(new_n8025, new_n9963);
xnor_4 g07615(n6794, n2387, new_n9964);
or_5   g07616(new_n9964, new_n9963, new_n9965);
xnor_4 g07617(n20077, n19494, new_n9966);
xor_4  g07618(new_n9966, new_n9958, new_n9967_1);
nand_5 g07619(new_n9967_1, new_n9965, new_n9968_1);
xor_4  g07620(new_n9967_1, new_n9965, new_n9969);
nand_5 g07621(new_n9969, new_n8019, new_n9970);
nand_5 g07622(new_n9970, new_n9968_1, new_n9971);
xnor_4 g07623(new_n9971, new_n9962, n1237);
not_10 g07624(new_n5743, new_n9973);
xnor_4 g07625(new_n9973, new_n5536, new_n9974);
xor_4  g07626(new_n9974, new_n5825, n1239);
not_10 g07627(n2416, new_n9976);
xnor_4 g07628(n22764, n1536, new_n9977);
or_5   g07629(n26264, n19454, new_n9978);
xnor_4 g07630(n26264, n19454, new_n9979);
or_5   g07631(n9445, n7841, new_n9980);
xnor_4 g07632(n9445, n7841, new_n9981);
or_5   g07633(n16812, n1279, new_n9982);
xnor_4 g07634(n16812, n1279, new_n9983);
or_5   g07635(n25068, n8324, new_n9984);
xnor_4 g07636(n25068, n8324, new_n9985);
or_5   g07637(n12546, n2331, new_n9986);
xnor_4 g07638(n12546, n2331, new_n9987);
or_5   g07639(n22631, n21078, new_n9988);
xnor_4 g07640(n22631, n21078, new_n9989);
or_5   g07641(n24485, n16743, new_n9990);
xnor_4 g07642(n24485, n16743, new_n9991);
or_5   g07643(n15258, n2420, new_n9992);
nand_5 g07644(n22201, n4588, new_n9993);
xor_4  g07645(n15258, n2420, new_n9994);
nand_5 g07646(new_n9994, new_n9993, new_n9995);
and_5  g07647(new_n9995, new_n9992, new_n9996);
or_5   g07648(new_n9996, new_n9991, new_n9997);
and_5  g07649(new_n9997, new_n9990, new_n9998);
or_5   g07650(new_n9998, new_n9989, new_n9999);
and_5  g07651(new_n9999, new_n9988, new_n10000);
or_5   g07652(new_n10000, new_n9987, new_n10001);
and_5  g07653(new_n10001, new_n9986, new_n10002);
or_5   g07654(new_n10002, new_n9985, new_n10003);
and_5  g07655(new_n10003, new_n9984, new_n10004);
or_5   g07656(new_n10004, new_n9983, new_n10005);
and_5  g07657(new_n10005, new_n9982, new_n10006);
or_5   g07658(new_n10006, new_n9981, new_n10007);
and_5  g07659(new_n10007, new_n9980, new_n10008);
or_5   g07660(new_n10008, new_n9979, new_n10009_1);
and_5  g07661(new_n10009_1, new_n9978, new_n10010_1);
xor_4  g07662(new_n10010_1, new_n9977, new_n10011);
and_5  g07663(new_n10011, new_n9976, new_n10012);
xor_4  g07664(new_n10011, new_n9976, new_n10013);
not_10 g07665(new_n10013, new_n10014);
not_10 g07666(n21905, new_n10015);
xor_4  g07667(new_n10008, new_n9979, new_n10016);
nand_5 g07668(new_n10016, new_n10015, new_n10017_1);
xor_4  g07669(new_n10016, new_n10015, new_n10018_1);
not_10 g07670(new_n10018_1, new_n10019_1);
not_10 g07671(n22918, new_n10020);
xor_4  g07672(new_n10006, new_n9981, new_n10021_1);
nand_5 g07673(new_n10021_1, new_n10020, new_n10022);
xor_4  g07674(new_n10021_1, new_n10020, new_n10023);
not_10 g07675(new_n10023, new_n10024);
not_10 g07676(n25923, new_n10025);
xor_4  g07677(new_n10004, new_n9983, new_n10026);
nand_5 g07678(new_n10026, new_n10025, new_n10027);
xor_4  g07679(new_n10026, new_n10025, new_n10028);
not_10 g07680(new_n10028, new_n10029);
not_10 g07681(n6790, new_n10030);
xor_4  g07682(new_n10002, new_n9985, new_n10031);
nand_5 g07683(new_n10031, new_n10030, new_n10032);
xor_4  g07684(new_n10031, new_n10030, new_n10033);
not_10 g07685(new_n10033, new_n10034);
not_10 g07686(n22879, new_n10035);
xor_4  g07687(new_n10000, new_n9987, new_n10036);
nand_5 g07688(new_n10036, new_n10035, new_n10037);
xor_4  g07689(new_n10036, new_n10035, new_n10038);
not_10 g07690(new_n10038, new_n10039);
not_10 g07691(n2117, new_n10040);
xor_4  g07692(new_n9998, new_n9989, new_n10041);
nand_5 g07693(new_n10041, new_n10040, new_n10042);
xor_4  g07694(new_n10041, new_n10040, new_n10043);
not_10 g07695(new_n10043, new_n10044);
not_10 g07696(n5882, new_n10045);
xor_4  g07697(new_n9996, new_n9991, new_n10046);
nand_5 g07698(new_n10046, new_n10045, new_n10047);
not_10 g07699(n11775, new_n10048);
xor_4  g07700(new_n9994, new_n9993, new_n10049);
and_5  g07701(new_n10049, new_n10048, new_n10050);
not_10 g07702(new_n10050, new_n10051);
xor_4  g07703(n22201, n4588, new_n10052);
and_5  g07704(new_n10052, n27134, new_n10053_1);
not_10 g07705(new_n10053_1, new_n10054);
xor_4  g07706(new_n10049, new_n10048, new_n10055_1);
and_5  g07707(new_n10055_1, new_n10054, new_n10056);
not_10 g07708(new_n10056, new_n10057_1);
and_5  g07709(new_n10057_1, new_n10051, new_n10058);
xor_4  g07710(new_n10046, n5882, new_n10059);
or_5   g07711(new_n10059, new_n10058, new_n10060);
and_5  g07712(new_n10060, new_n10047, new_n10061);
or_5   g07713(new_n10061, new_n10044, new_n10062);
and_5  g07714(new_n10062, new_n10042, new_n10063);
or_5   g07715(new_n10063, new_n10039, new_n10064);
and_5  g07716(new_n10064, new_n10037, new_n10065);
or_5   g07717(new_n10065, new_n10034, new_n10066);
and_5  g07718(new_n10066, new_n10032, new_n10067);
or_5   g07719(new_n10067, new_n10029, new_n10068);
and_5  g07720(new_n10068, new_n10027, new_n10069);
or_5   g07721(new_n10069, new_n10024, new_n10070);
and_5  g07722(new_n10070, new_n10022, new_n10071);
or_5   g07723(new_n10071, new_n10019_1, new_n10072);
and_5  g07724(new_n10072, new_n10017_1, new_n10073);
nor_5  g07725(new_n10073, new_n10014, new_n10074);
nor_5  g07726(new_n10074, new_n10012, new_n10075);
nor_5  g07727(n22764, n1536, new_n10076);
nor_5  g07728(new_n10010_1, new_n9977, new_n10077);
nor_5  g07729(new_n10077, new_n10076, new_n10078);
nand_5 g07730(new_n10078, new_n10075, new_n10079);
or_5   g07731(n23493, n8405, new_n10080);
or_5   g07732(n22359, n10275, new_n10081);
or_5   g07733(n15146, n5532, new_n10082);
or_5   g07734(n11579, n3962, new_n10083);
or_5   g07735(n23513, n21, new_n10084);
xnor_4 g07736(n23513, n21, new_n10085);
or_5   g07737(n6427, n1682, new_n10086);
nand_5 g07738(n6427, n1682, new_n10087);
nor_5  g07739(n7963, n6590, new_n10088);
nor_5  g07740(n20349, n10017, new_n10089);
and_5  g07741(n15936, n3618, new_n10090);
and_5  g07742(n20349, n10017, new_n10091);
nor_5  g07743(new_n10091, new_n10090, new_n10092);
nor_5  g07744(new_n10092, new_n10089, new_n10093);
and_5  g07745(n7963, n6590, new_n10094);
nor_5  g07746(new_n10094, new_n10093, new_n10095);
nor_5  g07747(new_n10095, new_n10088, new_n10096_1);
not_10 g07748(new_n10096_1, new_n10097);
nand_5 g07749(new_n10097, new_n10087, new_n10098);
and_5  g07750(new_n10098, new_n10086, new_n10099);
or_5   g07751(new_n10099, new_n10085, new_n10100);
and_5  g07752(new_n10100, new_n10084, new_n10101_1);
xnor_4 g07753(n11579, n3962, new_n10102);
or_5   g07754(new_n10102, new_n10101_1, new_n10103);
and_5  g07755(new_n10103, new_n10083, new_n10104);
xnor_4 g07756(n15146, n5532, new_n10105);
or_5   g07757(new_n10105, new_n10104, new_n10106);
and_5  g07758(new_n10106, new_n10082, new_n10107);
xnor_4 g07759(n22359, n10275, new_n10108);
or_5   g07760(new_n10108, new_n10107, new_n10109);
and_5  g07761(new_n10109, new_n10081, new_n10110);
xnor_4 g07762(n23493, n8405, new_n10111_1);
or_5   g07763(new_n10111_1, new_n10110, new_n10112);
and_5  g07764(new_n10112, new_n10080, new_n10113);
xnor_4 g07765(n14826, n13549, new_n10114);
xor_4  g07766(new_n10114, new_n10113, new_n10115);
and_5  g07767(new_n10115, new_n4449, new_n10116);
xor_4  g07768(new_n10115, n18105, new_n10117_1);
xor_4  g07769(new_n10111_1, new_n10110, new_n10118);
nand_5 g07770(new_n10118, new_n4450, new_n10119);
xor_4  g07771(new_n10118, new_n4450, new_n10120);
not_10 g07772(new_n10120, new_n10121);
xor_4  g07773(new_n10108, new_n10107, new_n10122);
nand_5 g07774(new_n10122, new_n4451_1, new_n10123);
xor_4  g07775(new_n10122, n16376, new_n10124);
xor_4  g07776(new_n10105, new_n10104, new_n10125_1);
nand_5 g07777(new_n10125_1, new_n4452, new_n10126);
xor_4  g07778(new_n10125_1, n25381, new_n10127);
xor_4  g07779(new_n10102, new_n10101_1, new_n10128);
nand_5 g07780(new_n10128, new_n4453, new_n10129);
xor_4  g07781(new_n10128, n12587, new_n10130);
xor_4  g07782(new_n10099, new_n10085, new_n10131);
nand_5 g07783(new_n10131, new_n4454, new_n10132);
xor_4  g07784(new_n10131, n268, new_n10133);
xor_4  g07785(n6427, n1682, new_n10134);
xor_4  g07786(new_n10134, new_n10097, new_n10135);
nand_5 g07787(new_n10135, new_n4455, new_n10136);
xor_4  g07788(new_n10135, n24879, new_n10137);
xnor_4 g07789(n7963, n6590, new_n10138);
xnor_4 g07790(new_n10138, new_n10093, new_n10139);
or_5   g07791(new_n10139, n6785, new_n10140);
xnor_4 g07792(n20349, n10017, new_n10141);
xnor_4 g07793(new_n10141, new_n10090, new_n10142);
nor_5  g07794(new_n10142, n24032, new_n10143);
xnor_4 g07795(n15936, n3618, new_n10144);
or_5   g07796(new_n10144, new_n8183, new_n10145);
xor_4  g07797(new_n10142, n24032, new_n10146);
and_5  g07798(new_n10146, new_n10145, new_n10147);
or_5   g07799(new_n10147, new_n10143, new_n10148);
xor_4  g07800(new_n10139, n6785, new_n10149);
nand_5 g07801(new_n10149, new_n10148, new_n10150);
and_5  g07802(new_n10150, new_n10140, new_n10151);
or_5   g07803(new_n10151, new_n10137, new_n10152);
and_5  g07804(new_n10152, new_n10136, new_n10153);
or_5   g07805(new_n10153, new_n10133, new_n10154);
and_5  g07806(new_n10154, new_n10132, new_n10155);
or_5   g07807(new_n10155, new_n10130, new_n10156);
and_5  g07808(new_n10156, new_n10129, new_n10157);
or_5   g07809(new_n10157, new_n10127, new_n10158_1);
and_5  g07810(new_n10158_1, new_n10126, new_n10159);
or_5   g07811(new_n10159, new_n10124, new_n10160);
and_5  g07812(new_n10160, new_n10123, new_n10161);
or_5   g07813(new_n10161, new_n10121, new_n10162);
and_5  g07814(new_n10162, new_n10119, new_n10163);
nor_5  g07815(new_n10163, new_n10117_1, new_n10164);
nor_5  g07816(new_n10164, new_n10116, new_n10165_1);
or_5   g07817(new_n10114, new_n10113, new_n10166);
or_5   g07818(n14826, n13549, new_n10167);
and_5  g07819(new_n10167, new_n10166, new_n10168);
and_5  g07820(new_n10168, new_n10165_1, new_n10169);
not_10 g07821(new_n10169, new_n10170);
xor_4  g07822(new_n10170, new_n10079, new_n10171);
xor_4  g07823(new_n10078, new_n10075, new_n10172);
not_10 g07824(new_n10172, new_n10173);
xor_4  g07825(new_n10168, new_n10165_1, new_n10174);
and_5  g07826(new_n10174, new_n10173, new_n10175);
not_10 g07827(new_n10174, new_n10176);
xnor_4 g07828(new_n10176, new_n10173, new_n10177);
xor_4  g07829(new_n10073, new_n10014, new_n10178);
xnor_4 g07830(new_n10163, new_n10117_1, new_n10179);
and_5  g07831(new_n10179, new_n10178, new_n10180);
xor_4  g07832(new_n10163, new_n10117_1, new_n10181);
xnor_4 g07833(new_n10181, new_n10178, new_n10182);
not_10 g07834(new_n10182, new_n10183);
xor_4  g07835(new_n10071, new_n10019_1, new_n10184);
xor_4  g07836(new_n10161, new_n10121, new_n10185);
not_10 g07837(new_n10185, new_n10186);
and_5  g07838(new_n10186, new_n10184, new_n10187);
not_10 g07839(new_n10187, new_n10188);
xor_4  g07840(new_n10186, new_n10184, new_n10189);
xor_4  g07841(new_n10069, new_n10024, new_n10190);
xnor_4 g07842(new_n10159, new_n10124, new_n10191);
and_5  g07843(new_n10191, new_n10190, new_n10192);
xor_4  g07844(new_n10159, new_n10124, new_n10193);
xnor_4 g07845(new_n10193, new_n10190, new_n10194);
not_10 g07846(new_n10194, new_n10195);
xor_4  g07847(new_n10067, new_n10029, new_n10196);
xnor_4 g07848(new_n10157, new_n10127, new_n10197);
and_5  g07849(new_n10197, new_n10196, new_n10198);
xor_4  g07850(new_n10157, new_n10127, new_n10199);
xnor_4 g07851(new_n10199, new_n10196, new_n10200);
not_10 g07852(new_n10200, new_n10201_1);
xor_4  g07853(new_n10065, new_n10034, new_n10202);
xnor_4 g07854(new_n10155, new_n10130, new_n10203);
and_5  g07855(new_n10203, new_n10202, new_n10204);
xor_4  g07856(new_n10155, new_n10130, new_n10205);
xnor_4 g07857(new_n10205, new_n10202, new_n10206);
not_10 g07858(new_n10206, new_n10207);
xor_4  g07859(new_n10063, new_n10039, new_n10208);
xnor_4 g07860(new_n10153, new_n10133, new_n10209);
and_5  g07861(new_n10209, new_n10208, new_n10210);
xor_4  g07862(new_n10153, new_n10133, new_n10211);
xnor_4 g07863(new_n10211, new_n10208, new_n10212);
not_10 g07864(new_n10212, new_n10213);
xor_4  g07865(new_n10061, new_n10044, new_n10214);
xnor_4 g07866(new_n10151, new_n10137, new_n10215);
and_5  g07867(new_n10215, new_n10214, new_n10216);
xor_4  g07868(new_n10151, new_n10137, new_n10217);
xnor_4 g07869(new_n10217, new_n10214, new_n10218);
not_10 g07870(new_n10218, new_n10219);
xor_4  g07871(new_n10059, new_n10058, new_n10220);
not_10 g07872(new_n10220, new_n10221);
xor_4  g07873(new_n10149, new_n10148, new_n10222);
nor_5  g07874(new_n10222, new_n10221, new_n10223);
not_10 g07875(new_n10223, new_n10224);
xor_4  g07876(new_n10222, new_n10221, new_n10225);
xor_4  g07877(new_n10055_1, new_n10054, new_n10226);
not_10 g07878(new_n10226, new_n10227);
xor_4  g07879(new_n10146, new_n10145, new_n10228);
nor_5  g07880(new_n10228, new_n10227, new_n10229);
not_10 g07881(new_n10229, new_n10230);
xor_4  g07882(new_n10052, n27134, new_n10231);
not_10 g07883(new_n10231, new_n10232);
xor_4  g07884(new_n10144, new_n8183, new_n10233);
and_5  g07885(new_n10233, new_n10232, new_n10234);
xor_4  g07886(new_n10228, new_n10227, new_n10235);
and_5  g07887(new_n10235, new_n10234, new_n10236_1);
not_10 g07888(new_n10236_1, new_n10237);
and_5  g07889(new_n10237, new_n10230, new_n10238);
not_10 g07890(new_n10238, new_n10239_1);
and_5  g07891(new_n10239_1, new_n10225, new_n10240);
not_10 g07892(new_n10240, new_n10241);
and_5  g07893(new_n10241, new_n10224, new_n10242);
nor_5  g07894(new_n10242, new_n10219, new_n10243);
nor_5  g07895(new_n10243, new_n10216, new_n10244_1);
nor_5  g07896(new_n10244_1, new_n10213, new_n10245);
nor_5  g07897(new_n10245, new_n10210, new_n10246);
nor_5  g07898(new_n10246, new_n10207, new_n10247);
nor_5  g07899(new_n10247, new_n10204, new_n10248);
nor_5  g07900(new_n10248, new_n10201_1, new_n10249);
nor_5  g07901(new_n10249, new_n10198, new_n10250_1);
nor_5  g07902(new_n10250_1, new_n10195, new_n10251);
nor_5  g07903(new_n10251, new_n10192, new_n10252);
not_10 g07904(new_n10252, new_n10253);
and_5  g07905(new_n10253, new_n10189, new_n10254);
not_10 g07906(new_n10254, new_n10255);
and_5  g07907(new_n10255, new_n10188, new_n10256);
nor_5  g07908(new_n10256, new_n10183, new_n10257);
nor_5  g07909(new_n10257, new_n10180, new_n10258);
not_10 g07910(new_n10258, new_n10259);
and_5  g07911(new_n10259, new_n10177, new_n10260);
nor_5  g07912(new_n10260, new_n10175, new_n10261_1);
xnor_4 g07913(new_n10261_1, new_n10171, n1302);
and_5  g07914(new_n2650, n12507, new_n10263);
not_10 g07915(new_n10263, new_n10264);
xnor_4 g07916(n13951, n12507, new_n10265);
not_10 g07917(new_n10265, new_n10266);
or_5   g07918(n22793, new_n8954, new_n10267);
xnor_4 g07919(n22793, n15077, new_n10268);
not_10 g07920(new_n10268, new_n10269);
or_5   g07921(n8439, new_n8961, new_n10270);
xnor_4 g07922(n8439, n3710, new_n10271);
not_10 g07923(new_n10271, new_n10272);
or_5   g07924(new_n8913, n25523, new_n10273);
xnor_4 g07925(n26318, n25523, new_n10274);
not_10 g07926(new_n10274, new_n10275_1);
or_5   g07927(new_n8917, n5579, new_n10276);
xnor_4 g07928(n26054, n5579, new_n10277);
not_10 g07929(new_n10277, new_n10278);
or_5   g07930(n23430, new_n8921, new_n10279);
xnor_4 g07931(n23430, n19081, new_n10280);
not_10 g07932(new_n10280, new_n10281);
not_10 g07933(n8309, new_n10282);
or_5   g07934(n10411, new_n10282, new_n10283);
xnor_4 g07935(n10411, n8309, new_n10284);
or_5   g07936(n19144, new_n2657, new_n10285);
not_10 g07937(n19144, new_n10286);
or_5   g07938(new_n10286, n16971, new_n10287_1);
not_10 g07939(n12593, new_n10288);
and_5  g07940(new_n10288, n11503, new_n10289);
not_10 g07941(n11503, new_n10290);
and_5  g07942(n12593, new_n10290, new_n10291);
not_10 g07943(new_n10291, new_n10292);
not_10 g07944(n13714, new_n10293);
and_5  g07945(n18151, new_n10293, new_n10294);
and_5  g07946(new_n10294, new_n10292, new_n10295_1);
nor_5  g07947(new_n10295_1, new_n10289, new_n10296);
not_10 g07948(new_n10296, new_n10297);
nand_5 g07949(new_n10297, new_n10287_1, new_n10298);
and_5  g07950(new_n10298, new_n10285, new_n10299);
nand_5 g07951(new_n10299, new_n10284, new_n10300);
and_5  g07952(new_n10300, new_n10283, new_n10301);
or_5   g07953(new_n10301, new_n10281, new_n10302);
and_5  g07954(new_n10302, new_n10279, new_n10303);
or_5   g07955(new_n10303, new_n10278, new_n10304);
and_5  g07956(new_n10304, new_n10276, new_n10305);
or_5   g07957(new_n10305, new_n10275_1, new_n10306);
and_5  g07958(new_n10306, new_n10273, new_n10307);
or_5   g07959(new_n10307, new_n10272, new_n10308);
and_5  g07960(new_n10308, new_n10270, new_n10309);
or_5   g07961(new_n10309, new_n10269, new_n10310);
and_5  g07962(new_n10310, new_n10267, new_n10311);
nor_5  g07963(new_n10311, new_n10266, new_n10312);
not_10 g07964(new_n10312, new_n10313);
and_5  g07965(new_n10313, new_n10264, new_n10314);
not_10 g07966(new_n10314, new_n10315);
nor_5  g07967(n12650, n11220, new_n10316);
not_10 g07968(new_n10316, new_n10317);
xor_4  g07969(n12650, n11220, new_n10318);
not_10 g07970(new_n10318, new_n10319);
or_5   g07971(n22379, n10201, new_n10320);
xor_4  g07972(n22379, n10201, new_n10321_1);
not_10 g07973(new_n10321_1, new_n10322);
or_5   g07974(n10593, n1662, new_n10323);
xor_4  g07975(n10593, n1662, new_n10324);
not_10 g07976(new_n10324, new_n10325);
or_5   g07977(n18290, n12875, new_n10326_1);
or_5   g07978(new_n9492, new_n9466, new_n10327_1);
and_5  g07979(new_n10327_1, new_n10326_1, new_n10328);
or_5   g07980(new_n10328, new_n10325, new_n10329);
and_5  g07981(new_n10329, new_n10323, new_n10330_1);
or_5   g07982(new_n10330_1, new_n10322, new_n10331);
and_5  g07983(new_n10331, new_n10320, new_n10332);
nor_5  g07984(new_n10332, new_n10319, new_n10333);
not_10 g07985(new_n10333, new_n10334);
and_5  g07986(new_n10334, new_n10317, new_n10335);
or_5   g07987(n22270, n2944, new_n10336);
or_5   g07988(new_n2708, new_n2668, new_n10337);
and_5  g07989(new_n10337, new_n10336, new_n10338);
xor_4  g07990(new_n10338, new_n10335, new_n10339);
xor_4  g07991(new_n10332, new_n10319, new_n10340_1);
not_10 g07992(new_n10340_1, new_n10341);
nand_5 g07993(new_n10341, new_n2709, new_n10342);
xor_4  g07994(new_n10330_1, new_n10322, new_n10343);
not_10 g07995(new_n10343, new_n10344);
or_5   g07996(new_n10344, new_n2713, new_n10345_1);
xnor_4 g07997(new_n10344, new_n2715, new_n10346);
not_10 g07998(new_n10346, new_n10347);
xor_4  g07999(new_n10328, new_n10325, new_n10348);
not_10 g08000(new_n10348, new_n10349);
or_5   g08001(new_n10349, new_n2718, new_n10350);
xnor_4 g08002(new_n10349, new_n2720, new_n10351);
not_10 g08003(new_n10351, new_n10352);
or_5   g08004(new_n9494, new_n2723, new_n10353);
nor_5  g08005(new_n9498, new_n2728, new_n10354);
not_10 g08006(new_n10354, new_n10355);
xnor_4 g08007(new_n9498, new_n2730, new_n10356_1);
nand_5 g08008(new_n9503, new_n2733, new_n10357);
or_5   g08009(new_n9508_1, new_n2737, new_n10358);
xnor_4 g08010(new_n9508_1, new_n2738, new_n10359);
not_10 g08011(new_n10359, new_n10360);
or_5   g08012(new_n9512_1, new_n2743_1, new_n10361);
xnor_4 g08013(new_n9512_1, new_n2744, new_n10362);
nand_5 g08014(new_n9514, new_n2754, new_n10363);
not_10 g08015(new_n9517, new_n10364);
and_5  g08016(new_n10364, new_n2752, new_n10365);
xnor_4 g08017(new_n9515, new_n2754, new_n10366);
nand_5 g08018(new_n10366, new_n10365, new_n10367);
nand_5 g08019(new_n10367, new_n10363, new_n10368);
nand_5 g08020(new_n10368, new_n10362, new_n10369);
and_5  g08021(new_n10369, new_n10361, new_n10370);
or_5   g08022(new_n10370, new_n10360, new_n10371);
and_5  g08023(new_n10371, new_n10358, new_n10372_1);
xnor_4 g08024(new_n9503, new_n2762, new_n10373);
nand_5 g08025(new_n10373, new_n10372_1, new_n10374);
and_5  g08026(new_n10374, new_n10357, new_n10375);
and_5  g08027(new_n10375, new_n10356_1, new_n10376);
not_10 g08028(new_n10376, new_n10377);
and_5  g08029(new_n10377, new_n10355, new_n10378);
xor_4  g08030(new_n9494, new_n2725, new_n10379);
or_5   g08031(new_n10379, new_n10378, new_n10380);
and_5  g08032(new_n10380, new_n10353, new_n10381);
or_5   g08033(new_n10381, new_n10352, new_n10382);
and_5  g08034(new_n10382, new_n10350, new_n10383);
or_5   g08035(new_n10383, new_n10347, new_n10384);
and_5  g08036(new_n10384, new_n10345_1, new_n10385_1);
xnor_4 g08037(new_n10341, new_n2710, new_n10386);
nand_5 g08038(new_n10386, new_n10385_1, new_n10387_1);
and_5  g08039(new_n10387_1, new_n10342, new_n10388_1);
xor_4  g08040(new_n10388_1, new_n10339, new_n10389);
xnor_4 g08041(new_n10389, new_n10315, new_n10390_1);
not_10 g08042(new_n10390_1, new_n10391);
xor_4  g08043(new_n10311, new_n10266, new_n10392);
xor_4  g08044(new_n10386, new_n10385_1, new_n10393);
nor_5  g08045(new_n10393, new_n10392, new_n10394);
xor_4  g08046(new_n10393, new_n10392, new_n10395);
not_10 g08047(new_n10395, new_n10396);
xor_4  g08048(new_n10309, new_n10269, new_n10397);
xor_4  g08049(new_n10383, new_n10347, new_n10398);
not_10 g08050(new_n10398, new_n10399);
nor_5  g08051(new_n10399, new_n10397, new_n10400);
xor_4  g08052(new_n10399, new_n10397, new_n10401);
xor_4  g08053(new_n10307, new_n10272, new_n10402);
xnor_4 g08054(new_n10381, new_n10351, new_n10403);
not_10 g08055(new_n10403, new_n10404_1);
nor_5  g08056(new_n10404_1, new_n10402, new_n10405_1);
xnor_4 g08057(new_n10403, new_n10402, new_n10406);
xor_4  g08058(new_n10305, new_n10275_1, new_n10407);
not_10 g08059(new_n10407, new_n10408);
xnor_4 g08060(new_n9494, new_n2725, new_n10409_1);
xnor_4 g08061(new_n10409_1, new_n10378, new_n10410);
and_5  g08062(new_n10410, new_n10408, new_n10411_1);
xor_4  g08063(new_n10410, new_n10408, new_n10412);
xor_4  g08064(new_n10303, new_n10278, new_n10413);
xor_4  g08065(new_n10375, new_n10356_1, new_n10414);
not_10 g08066(new_n10414, new_n10415);
nor_5  g08067(new_n10415, new_n10413, new_n10416);
xor_4  g08068(new_n10301, new_n10281, new_n10417);
xor_4  g08069(new_n10373, new_n10372_1, new_n10418);
nor_5  g08070(new_n10418, new_n10417, new_n10419);
xor_4  g08071(new_n10418, new_n10417, new_n10420_1);
not_10 g08072(new_n10420_1, new_n10421);
xnor_4 g08073(new_n10370, new_n10359, new_n10422);
not_10 g08074(new_n10422, new_n10423);
xor_4  g08075(new_n10299, new_n10284, new_n10424);
nor_5  g08076(new_n10424, new_n10423, new_n10425);
xor_4  g08077(new_n10368, new_n10362, new_n10426);
xnor_4 g08078(n19144, n16971, new_n10427);
xor_4  g08079(new_n10427, new_n10297, new_n10428);
and_5  g08080(new_n10428, new_n10426, new_n10429);
not_10 g08081(new_n10429, new_n10430);
xor_4  g08082(new_n10428, new_n10426, new_n10431);
xnor_4 g08083(new_n9517, new_n2752, new_n10432_1);
xnor_4 g08084(n18151, n13714, new_n10433);
or_5   g08085(new_n10433, new_n10432_1, new_n10434);
xnor_4 g08086(n12593, n11503, new_n10435);
xor_4  g08087(new_n10435, new_n10294, new_n10436);
nor_5  g08088(new_n10436, new_n10434, new_n10437);
xnor_4 g08089(new_n10366, new_n10365, new_n10438);
xor_4  g08090(new_n10436, new_n10434, new_n10439);
and_5  g08091(new_n10439, new_n10438, new_n10440);
nor_5  g08092(new_n10440, new_n10437, new_n10441);
and_5  g08093(new_n10441, new_n10431, new_n10442);
not_10 g08094(new_n10442, new_n10443);
and_5  g08095(new_n10443, new_n10430, new_n10444);
xnor_4 g08096(new_n10424, new_n10422, new_n10445);
not_10 g08097(new_n10445, new_n10446);
nor_5  g08098(new_n10446, new_n10444, new_n10447);
nor_5  g08099(new_n10447, new_n10425, new_n10448);
nor_5  g08100(new_n10448, new_n10421, new_n10449);
nor_5  g08101(new_n10449, new_n10419, new_n10450);
not_10 g08102(new_n10450, new_n10451);
xor_4  g08103(new_n10415, new_n10413, new_n10452);
and_5  g08104(new_n10452, new_n10451, new_n10453);
nor_5  g08105(new_n10453, new_n10416, new_n10454);
not_10 g08106(new_n10454, new_n10455);
and_5  g08107(new_n10455, new_n10412, new_n10456);
nor_5  g08108(new_n10456, new_n10411_1, new_n10457);
not_10 g08109(new_n10457, new_n10458);
and_5  g08110(new_n10458, new_n10406, new_n10459);
nor_5  g08111(new_n10459, new_n10405_1, new_n10460);
not_10 g08112(new_n10460, new_n10461);
and_5  g08113(new_n10461, new_n10401, new_n10462);
nor_5  g08114(new_n10462, new_n10400, new_n10463);
nor_5  g08115(new_n10463, new_n10396, new_n10464);
nor_5  g08116(new_n10464, new_n10394, new_n10465);
xnor_4 g08117(new_n10465, new_n10391, n1332);
or_5   g08118(new_n5591, n14692, new_n10467);
xor_4  g08119(new_n5591, n14692, new_n10468);
not_10 g08120(new_n10468, new_n10469);
not_10 g08121(n4100, new_n10470);
nand_5 g08122(new_n5662, new_n10470, new_n10471);
xor_4  g08123(new_n5662, n4100, new_n10472);
not_10 g08124(n21957, new_n10473);
nand_5 g08125(new_n5668, new_n10473, new_n10474);
xor_4  g08126(new_n5668, n21957, new_n10475);
not_10 g08127(n15761, new_n10476);
nand_5 g08128(new_n5673, new_n10476, new_n10477);
xor_4  g08129(new_n5673, n15761, new_n10478);
not_10 g08130(n11201, new_n10479);
nand_5 g08131(new_n5678, new_n10479, new_n10480);
xor_4  g08132(new_n5678, n11201, new_n10481);
not_10 g08133(n18690, new_n10482);
nand_5 g08134(new_n5684, new_n10482, new_n10483);
xor_4  g08135(new_n5684, n18690, new_n10484_1);
not_10 g08136(n12153, new_n10485);
nand_5 g08137(new_n5689, new_n10485, new_n10486);
xor_4  g08138(new_n5689, new_n10485, new_n10487);
nand_5 g08139(new_n5697, n13044, new_n10488);
or_5   g08140(new_n5697, n13044, new_n10489_1);
nor_5  g08141(new_n5863, n18745, new_n10490);
and_5  g08142(new_n5864, new_n5862, new_n10491);
nor_5  g08143(new_n10491, new_n10490, new_n10492);
nand_5 g08144(new_n10492, new_n10489_1, new_n10493);
and_5  g08145(new_n10493, new_n10488, new_n10494);
nand_5 g08146(new_n10494, new_n10487, new_n10495);
and_5  g08147(new_n10495, new_n10486, new_n10496);
or_5   g08148(new_n10496, new_n10484_1, new_n10497);
and_5  g08149(new_n10497, new_n10483, new_n10498);
or_5   g08150(new_n10498, new_n10481, new_n10499);
and_5  g08151(new_n10499, new_n10480, new_n10500);
or_5   g08152(new_n10500, new_n10478, new_n10501);
and_5  g08153(new_n10501, new_n10477, new_n10502);
or_5   g08154(new_n10502, new_n10475, new_n10503);
and_5  g08155(new_n10503, new_n10474, new_n10504);
or_5   g08156(new_n10504, new_n10472, new_n10505);
and_5  g08157(new_n10505, new_n10471, new_n10506);
or_5   g08158(new_n10506, new_n10469, new_n10507);
and_5  g08159(new_n10507, new_n10467, new_n10508);
and_5  g08160(new_n10508, new_n5590, new_n10509);
not_10 g08161(new_n10509, new_n10510);
not_10 g08162(n15182, new_n10511);
not_10 g08163(n27037, new_n10512);
not_10 g08164(n10405, new_n10513);
and_5  g08165(new_n5874, new_n5507, new_n10514_1);
and_5  g08166(new_n10514_1, new_n10513, new_n10515);
and_5  g08167(new_n10515, new_n4041, new_n10516);
and_5  g08168(new_n10516, new_n4009, new_n10517);
and_5  g08169(new_n10517, new_n6259, new_n10518);
and_5  g08170(new_n10518, new_n10512, new_n10519);
and_5  g08171(new_n10519, new_n10511, new_n10520);
and_5  g08172(new_n10520, new_n5480, new_n10521);
not_10 g08173(n15766, new_n10522);
not_10 g08174(n25629, new_n10523);
not_10 g08175(n7692, new_n10524);
not_10 g08176(n23039, new_n10525_1);
not_10 g08177(n13677, new_n10526);
not_10 g08178(n18926, new_n10527);
not_10 g08179(n5330, new_n10528);
nor_5  g08180(n25926, n7657, new_n10529);
and_5  g08181(new_n10529, new_n10528, new_n10530);
and_5  g08182(new_n10530, new_n3978, new_n10531);
and_5  g08183(new_n10531, new_n10527, new_n10532);
and_5  g08184(new_n10532, new_n10526, new_n10533);
and_5  g08185(new_n10533, new_n10525_1, new_n10534);
and_5  g08186(new_n10534, new_n10524, new_n10535);
and_5  g08187(new_n10535, new_n10523, new_n10536);
and_5  g08188(new_n10536, new_n10522, new_n10537);
not_10 g08189(n23895, new_n10538);
xor_4  g08190(new_n10536, new_n10522, new_n10539);
not_10 g08191(new_n10539, new_n10540_1);
and_5  g08192(new_n10540_1, new_n10538, new_n10541);
xor_4  g08193(new_n10535, new_n10523, new_n10542);
nor_5  g08194(new_n10542, n17351, new_n10543);
xor_4  g08195(new_n10542, new_n5484, new_n10544);
xor_4  g08196(new_n10534, new_n10524, new_n10545);
or_5   g08197(new_n10545, n11736, new_n10546);
xor_4  g08198(new_n10545, new_n5488, new_n10547);
xor_4  g08199(new_n10533, new_n10525_1, new_n10548);
or_5   g08200(new_n10548, n23200, new_n10549);
xor_4  g08201(new_n10548, new_n5492, new_n10550);
xor_4  g08202(new_n10532, new_n10526, new_n10551);
or_5   g08203(new_n10551, n17959, new_n10552);
xor_4  g08204(new_n10531, new_n10527, new_n10553);
nor_5  g08205(new_n10553, n7566, new_n10554);
xor_4  g08206(new_n10553, n7566, new_n10555);
xor_4  g08207(new_n10530, new_n3978, new_n10556);
nand_5 g08208(new_n10556, n7731, new_n10557);
nor_5  g08209(new_n10556, n7731, new_n10558);
xor_4  g08210(new_n10529, new_n10528, new_n10559);
and_5  g08211(new_n10559, n12341, new_n10560);
xor_4  g08212(new_n10559, n12341, new_n10561_1);
not_10 g08213(new_n10561_1, new_n10562);
nand_5 g08214(new_n5868, n20986, new_n10563);
nand_5 g08215(new_n5869, new_n5867, new_n10564_1);
and_5  g08216(new_n10564_1, new_n10563, new_n10565);
nor_5  g08217(new_n10565, new_n10562, new_n10566);
nor_5  g08218(new_n10566, new_n10560, new_n10567);
or_5   g08219(new_n10567, new_n10558, new_n10568);
and_5  g08220(new_n10568, new_n10557, new_n10569);
and_5  g08221(new_n10569, new_n10555, new_n10570);
or_5   g08222(new_n10570, new_n10554, new_n10571);
xor_4  g08223(new_n10551, n17959, new_n10572);
nand_5 g08224(new_n10572, new_n10571, new_n10573);
and_5  g08225(new_n10573, new_n10552, new_n10574);
or_5   g08226(new_n10574, new_n10550, new_n10575);
and_5  g08227(new_n10575, new_n10549, new_n10576);
or_5   g08228(new_n10576, new_n10547, new_n10577_1);
and_5  g08229(new_n10577_1, new_n10546, new_n10578);
nor_5  g08230(new_n10578, new_n10544, new_n10579);
nor_5  g08231(new_n10579, new_n10543, new_n10580);
nor_5  g08232(new_n10540_1, new_n10538, new_n10581);
nor_5  g08233(new_n10581, new_n10580, new_n10582);
nor_5  g08234(new_n10582, new_n10541, new_n10583);
nor_5  g08235(new_n10583, new_n10537, new_n10584);
nor_5  g08236(new_n10584, new_n10521, new_n10585);
xor_4  g08237(new_n10520, n8614, new_n10586);
or_5   g08238(new_n10581, new_n10541, new_n10587);
xor_4  g08239(new_n10587, new_n10580, new_n10588_1);
nor_5  g08240(new_n10588_1, new_n10586, new_n10589);
xor_4  g08241(new_n10519, new_n10511, new_n10590);
not_10 g08242(new_n10590, new_n10591);
xor_4  g08243(new_n10578, new_n10544, new_n10592);
nand_5 g08244(new_n10592, new_n10591, new_n10593_1);
xor_4  g08245(new_n10592, new_n10590, new_n10594);
xor_4  g08246(new_n10518, new_n10512, new_n10595_1);
not_10 g08247(new_n10595_1, new_n10596);
xor_4  g08248(new_n10576, new_n10547, new_n10597);
nand_5 g08249(new_n10597, new_n10596, new_n10598);
xor_4  g08250(new_n10597, new_n10596, new_n10599);
not_10 g08251(new_n10599, new_n10600);
xor_4  g08252(new_n10517, new_n6259, new_n10601);
not_10 g08253(new_n10601, new_n10602);
xor_4  g08254(new_n10574, new_n10550, new_n10603);
nand_5 g08255(new_n10603, new_n10602, new_n10604);
xor_4  g08256(new_n10603, new_n10601, new_n10605);
xor_4  g08257(new_n10516, new_n4009, new_n10606);
not_10 g08258(new_n10606, new_n10607);
xor_4  g08259(new_n10572, new_n10571, new_n10608);
nand_5 g08260(new_n10608, new_n10607, new_n10609);
xor_4  g08261(new_n10608, new_n10607, new_n10610);
not_10 g08262(new_n10610, new_n10611_1);
xor_4  g08263(new_n10515, new_n4041, new_n10612);
not_10 g08264(new_n10612, new_n10613);
xor_4  g08265(new_n10569, new_n10555, new_n10614_1);
nand_5 g08266(new_n10614_1, new_n10613, new_n10615);
xor_4  g08267(new_n10614_1, new_n10612, new_n10616);
xor_4  g08268(new_n10514_1, new_n10513, new_n10617_1);
xor_4  g08269(new_n10556, n7731, new_n10618);
xnor_4 g08270(new_n10618, new_n10567, new_n10619);
or_5   g08271(new_n10619, new_n10617_1, new_n10620);
not_10 g08272(new_n10619, new_n10621);
xnor_4 g08273(new_n10621, new_n10617_1, new_n10622);
not_10 g08274(new_n10622, new_n10623);
xor_4  g08275(new_n10565, new_n10562, new_n10624);
xor_4  g08276(new_n5874, new_n5507, new_n10625);
or_5   g08277(new_n10625, new_n10624, new_n10626);
not_10 g08278(new_n10624, new_n10627);
xnor_4 g08279(new_n10625, new_n10627, new_n10628_1);
nand_5 g08280(new_n5878, new_n5871, new_n10629);
nand_5 g08281(new_n10629, new_n5877, new_n10630);
nand_5 g08282(new_n10630, new_n10628_1, new_n10631);
and_5  g08283(new_n10631, new_n10626, new_n10632);
or_5   g08284(new_n10632, new_n10623, new_n10633);
and_5  g08285(new_n10633, new_n10620, new_n10634);
or_5   g08286(new_n10634, new_n10616, new_n10635);
and_5  g08287(new_n10635, new_n10615, new_n10636);
or_5   g08288(new_n10636, new_n10611_1, new_n10637);
and_5  g08289(new_n10637, new_n10609, new_n10638);
or_5   g08290(new_n10638, new_n10605, new_n10639);
and_5  g08291(new_n10639, new_n10604, new_n10640);
or_5   g08292(new_n10640, new_n10600, new_n10641);
and_5  g08293(new_n10641, new_n10598, new_n10642);
or_5   g08294(new_n10642, new_n10594, new_n10643);
and_5  g08295(new_n10643, new_n10593_1, new_n10644);
xor_4  g08296(new_n10588_1, new_n10586, new_n10645);
and_5  g08297(new_n10645, new_n10644, new_n10646);
nor_5  g08298(new_n10646, new_n10589, new_n10647_1);
and_5  g08299(new_n10647_1, new_n10585, new_n10648);
xor_4  g08300(new_n10648, new_n10510, new_n10649);
xor_4  g08301(new_n10508, new_n5590, new_n10650_1);
xor_4  g08302(new_n10584, new_n10521, new_n10651);
xor_4  g08303(new_n10651, new_n10647_1, new_n10652);
nor_5  g08304(new_n10652, new_n10650_1, new_n10653_1);
xor_4  g08305(new_n10652, new_n10650_1, new_n10654);
xnor_4 g08306(new_n10506, new_n10469, new_n10655);
xor_4  g08307(new_n10645, new_n10644, new_n10656);
and_5  g08308(new_n10656, new_n10655, new_n10657);
not_10 g08309(new_n10655, new_n10658);
xor_4  g08310(new_n10656, new_n10658, new_n10659);
xor_4  g08311(new_n10642, new_n10594, new_n10660);
xor_4  g08312(new_n10504, new_n10472, new_n10661);
or_5   g08313(new_n10661, new_n10660, new_n10662);
xor_4  g08314(new_n10640, new_n10600, new_n10663);
not_10 g08315(new_n10663, new_n10664);
xor_4  g08316(new_n10502, new_n10475, new_n10665);
not_10 g08317(new_n10665, new_n10666);
or_5   g08318(new_n10666, new_n10664, new_n10667);
xor_4  g08319(new_n10666, new_n10664, new_n10668);
xor_4  g08320(new_n10638, new_n10605, new_n10669);
xor_4  g08321(new_n10500, new_n10478, new_n10670);
nor_5  g08322(new_n10670, new_n10669, new_n10671);
xor_4  g08323(new_n10636, new_n10611_1, new_n10672);
not_10 g08324(new_n10672, new_n10673);
xor_4  g08325(new_n10498, new_n10481, new_n10674);
not_10 g08326(new_n10674, new_n10675);
or_5   g08327(new_n10675, new_n10673, new_n10676);
xor_4  g08328(new_n10675, new_n10673, new_n10677);
xor_4  g08329(new_n10634, new_n10616, new_n10678);
xor_4  g08330(new_n10496, new_n10484_1, new_n10679);
nor_5  g08331(new_n10679, new_n10678, new_n10680);
xor_4  g08332(new_n10679, new_n10678, new_n10681);
xnor_4 g08333(new_n10632, new_n10622, new_n10682);
not_10 g08334(new_n10682, new_n10683);
xor_4  g08335(new_n10494, new_n10487, new_n10684);
not_10 g08336(new_n10684, new_n10685);
or_5   g08337(new_n10685, new_n10683, new_n10686);
xor_4  g08338(new_n10685, new_n10683, new_n10687);
xor_4  g08339(new_n10630, new_n10628_1, new_n10688);
not_10 g08340(new_n10688, new_n10689);
and_5  g08341(new_n10489_1, new_n10488, new_n10690);
xor_4  g08342(new_n10690, new_n10492, new_n10691);
or_5   g08343(new_n10691, new_n10689, new_n10692_1);
nand_5 g08344(new_n5879, new_n5865, new_n10693);
not_10 g08345(new_n5860, new_n10694_1);
nand_5 g08346(new_n5880, new_n10694_1, new_n10695);
nand_5 g08347(new_n10695, new_n10693, new_n10696);
xor_4  g08348(new_n10691, new_n10689, new_n10697);
nand_5 g08349(new_n10697, new_n10696, new_n10698);
nand_5 g08350(new_n10698, new_n10692_1, new_n10699);
nand_5 g08351(new_n10699, new_n10687, new_n10700);
and_5  g08352(new_n10700, new_n10686, new_n10701_1);
and_5  g08353(new_n10701_1, new_n10681, new_n10702);
nor_5  g08354(new_n10702, new_n10680, new_n10703);
nand_5 g08355(new_n10703, new_n10677, new_n10704);
and_5  g08356(new_n10704, new_n10676, new_n10705);
xor_4  g08357(new_n10670, new_n10669, new_n10706);
and_5  g08358(new_n10706, new_n10705, new_n10707);
nor_5  g08359(new_n10707, new_n10671, new_n10708);
nand_5 g08360(new_n10708, new_n10668, new_n10709);
and_5  g08361(new_n10709, new_n10667, new_n10710_1);
xor_4  g08362(new_n10661, new_n10660, new_n10711);
nand_5 g08363(new_n10711, new_n10710_1, new_n10712_1);
and_5  g08364(new_n10712_1, new_n10662, new_n10713);
nor_5  g08365(new_n10713, new_n10659, new_n10714);
nor_5  g08366(new_n10714, new_n10657, new_n10715);
and_5  g08367(new_n10715, new_n10654, new_n10716);
nor_5  g08368(new_n10716, new_n10653_1, new_n10717);
not_10 g08369(new_n10717, new_n10718);
xor_4  g08370(new_n10718, new_n10649, n1357);
xor_4  g08371(new_n8104, n25240, new_n10720);
not_10 g08372(new_n10720, new_n10721);
or_5   g08373(new_n8110, n10125, new_n10722);
xor_4  g08374(new_n8110, n10125, new_n10723);
not_10 g08375(new_n10723, new_n10724);
or_5   g08376(new_n8116, n8067, new_n10725);
xor_4  g08377(new_n8116, n8067, new_n10726);
not_10 g08378(new_n10726, new_n10727);
or_5   g08379(new_n8122, n20923, new_n10728);
xor_4  g08380(new_n8122, n20923, new_n10729);
not_10 g08381(new_n10729, new_n10730);
or_5   g08382(new_n8127_1, n18157, new_n10731);
nand_5 g08383(new_n8587, new_n8580, new_n10732);
nand_5 g08384(new_n10732, new_n8579, new_n10733);
and_5  g08385(new_n10733, new_n10731, new_n10734);
or_5   g08386(new_n10734, new_n10730, new_n10735);
and_5  g08387(new_n10735, new_n10728, new_n10736);
or_5   g08388(new_n10736, new_n10727, new_n10737);
and_5  g08389(new_n10737, new_n10725, new_n10738);
or_5   g08390(new_n10738, new_n10724, new_n10739_1);
and_5  g08391(new_n10739_1, new_n10722, new_n10740);
xor_4  g08392(new_n10740, new_n10721, new_n10741);
not_10 g08393(new_n10741, new_n10742);
not_10 g08394(n5077, new_n10743);
xnor_4 g08395(n6381, n1099, new_n10744);
or_5   g08396(n14345, n2113, new_n10745);
xnor_4 g08397(n14345, n2113, new_n10746);
or_5   g08398(n21134, n11356, new_n10747);
xor_4  g08399(n21134, n11356, new_n10748);
nand_5 g08400(n6369, n3164, new_n10749);
or_5   g08401(n6369, n3164, new_n10750);
nor_5  g08402(n25797, n10611, new_n10751);
nor_5  g08403(new_n6644, new_n6635, new_n10752);
nor_5  g08404(new_n10752, new_n10751, new_n10753);
nand_5 g08405(new_n10753, new_n10750, new_n10754);
and_5  g08406(new_n10754, new_n10749, new_n10755);
nand_5 g08407(new_n10755, new_n10748, new_n10756_1);
and_5  g08408(new_n10756_1, new_n10747, new_n10757);
or_5   g08409(new_n10757, new_n10746, new_n10758);
and_5  g08410(new_n10758, new_n10745, new_n10759);
xor_4  g08411(new_n10759, new_n10744, new_n10760);
xor_4  g08412(new_n10760, new_n10743, new_n10761);
not_10 g08413(n15546, new_n10762);
xor_4  g08414(new_n10757, new_n10746, new_n10763_1);
or_5   g08415(new_n10763_1, new_n10762, new_n10764);
xor_4  g08416(new_n10763_1, new_n10762, new_n10765);
not_10 g08417(n26452, new_n10766);
xor_4  g08418(new_n10755, new_n10748, new_n10767);
nand_5 g08419(new_n10767, new_n10766, new_n10768);
xor_4  g08420(n6369, n3164, new_n10769);
xor_4  g08421(new_n10769, new_n10753, new_n10770);
nand_5 g08422(new_n10770, n19905, new_n10771);
xor_4  g08423(new_n10770, new_n4165_1, new_n10772);
or_5   g08424(new_n6645, new_n4166, new_n10773);
nand_5 g08425(new_n8620_1, new_n8617, new_n10774);
and_5  g08426(new_n10774, new_n10773, new_n10775_1);
or_5   g08427(new_n10775_1, new_n10772, new_n10776);
and_5  g08428(new_n10776, new_n10771, new_n10777);
xor_4  g08429(new_n10767, new_n10766, new_n10778);
nand_5 g08430(new_n10778, new_n10777, new_n10779);
and_5  g08431(new_n10779, new_n10768, new_n10780_1);
nand_5 g08432(new_n10780_1, new_n10765, new_n10781);
and_5  g08433(new_n10781, new_n10764, new_n10782);
xor_4  g08434(new_n10782, new_n10761, new_n10783);
xor_4  g08435(new_n10783, new_n10742, new_n10784);
xor_4  g08436(new_n10738, new_n10724, new_n10785);
xor_4  g08437(new_n10780_1, new_n10765, new_n10786);
nand_5 g08438(new_n10786, new_n10785, new_n10787);
xor_4  g08439(new_n10786, new_n10785, new_n10788);
not_10 g08440(new_n10788, new_n10789);
xor_4  g08441(new_n10736, new_n10727, new_n10790);
not_10 g08442(new_n10790, new_n10791);
xor_4  g08443(new_n10778, new_n10777, new_n10792_1);
or_5   g08444(new_n10792_1, new_n10791, new_n10793);
xor_4  g08445(new_n10792_1, new_n10791, new_n10794);
xnor_4 g08446(new_n10734, new_n10729, new_n10795);
xor_4  g08447(new_n10775_1, new_n10772, new_n10796);
nand_5 g08448(new_n10796, new_n10795, new_n10797);
xor_4  g08449(new_n10796, new_n10795, new_n10798);
not_10 g08450(new_n8589, new_n10799);
and_5  g08451(new_n8615, new_n10799, new_n10800);
nor_5  g08452(new_n8621, new_n8616, new_n10801);
nor_5  g08453(new_n10801, new_n10800, new_n10802);
nand_5 g08454(new_n10802, new_n10798, new_n10803);
nand_5 g08455(new_n10803, new_n10797, new_n10804);
nand_5 g08456(new_n10804, new_n10794, new_n10805);
and_5  g08457(new_n10805, new_n10793, new_n10806);
or_5   g08458(new_n10806, new_n10789, new_n10807);
nand_5 g08459(new_n10807, new_n10787, new_n10808);
xnor_4 g08460(new_n10808, new_n10784, n1371);
xnor_4 g08461(n17250, n15241, new_n10810);
not_10 g08462(new_n10810, new_n10811);
nand_5 g08463(n23160, new_n4368, new_n10812);
not_10 g08464(n3785, new_n10813);
and_5  g08465(n16524, new_n10813, new_n10814);
xnor_4 g08466(n16524, n3785, new_n10815);
or_5   g08467(new_n6664, n11056, new_n10816);
and_5  g08468(new_n7801, n5822, new_n10817_1);
xor_4  g08469(n15271, n5822, new_n10818);
or_5   g08470(new_n4382, n25877, new_n10819);
nand_5 g08471(new_n5837, new_n5836, new_n10820);
and_5  g08472(new_n10820, new_n10819, new_n10821);
nor_5  g08473(new_n10821, new_n10818, new_n10822);
or_5   g08474(new_n10822, new_n10817_1, new_n10823);
xnor_4 g08475(n20250, n11056, new_n10824);
nand_5 g08476(new_n10824, new_n10823, new_n10825);
and_5  g08477(new_n10825, new_n10816, new_n10826);
and_5  g08478(new_n10826, new_n10815, new_n10827);
or_5   g08479(new_n10827, new_n10814, new_n10828);
xnor_4 g08480(n23160, n7678, new_n10829);
nand_5 g08481(new_n10829, new_n10828, new_n10830);
and_5  g08482(new_n10830, new_n10812, new_n10831);
xor_4  g08483(new_n10831, new_n10811, new_n10832);
not_10 g08484(new_n10832, new_n10833);
not_10 g08485(n13783, new_n10834_1);
xor_4  g08486(new_n9863, new_n10834_1, new_n10835);
or_5   g08487(new_n9866, n26660, new_n10836);
xor_4  g08488(new_n9866, n26660, new_n10837);
nand_5 g08489(new_n9869, n3018, new_n10838);
nor_5  g08490(new_n9869, n3018, new_n10839);
and_5  g08491(new_n9653, n3480, new_n10840);
nor_5  g08492(new_n9663, new_n9655_1, new_n10841);
nor_5  g08493(new_n10841, new_n10840, new_n10842);
or_5   g08494(new_n10842, new_n10839, new_n10843);
and_5  g08495(new_n10843, new_n10838, new_n10844);
nand_5 g08496(new_n10844, new_n10837, new_n10845);
and_5  g08497(new_n10845, new_n10836, new_n10846);
xor_4  g08498(new_n10846, new_n10835, new_n10847);
xnor_4 g08499(new_n10847, new_n10833, new_n10848);
xor_4  g08500(new_n10844, new_n10837, new_n10849);
not_10 g08501(new_n10849, new_n10850);
xor_4  g08502(new_n10829, new_n10828, new_n10851_1);
nand_5 g08503(new_n10851_1, new_n10850, new_n10852);
xor_4  g08504(new_n10851_1, new_n10850, new_n10853);
xor_4  g08505(new_n10826, new_n10815, new_n10854);
not_10 g08506(n3018, new_n10855);
xor_4  g08507(new_n9869, new_n10855, new_n10856);
xor_4  g08508(new_n10856, new_n10842, new_n10857);
or_5   g08509(new_n10857, new_n10854, new_n10858);
not_10 g08510(new_n10854, new_n10859);
xor_4  g08511(new_n10857, new_n10859, new_n10860);
xor_4  g08512(new_n10824, new_n10823, new_n10861);
nand_5 g08513(new_n10861, new_n9665, new_n10862);
xor_4  g08514(new_n10861, new_n9665, new_n10863);
xor_4  g08515(new_n10821, new_n10818, new_n10864);
or_5   g08516(new_n10864, new_n9670, new_n10865);
xnor_4 g08517(new_n10864, new_n9670, new_n10866);
nand_5 g08518(new_n5839, new_n5835, new_n10867);
xor_4  g08519(new_n5846, new_n5841_1, new_n10868);
nand_5 g08520(new_n10868, new_n5840_1, new_n10869);
and_5  g08521(new_n10869, new_n10867, new_n10870);
or_5   g08522(new_n10870, new_n10866, new_n10871);
and_5  g08523(new_n10871, new_n10865, new_n10872);
nand_5 g08524(new_n10872, new_n10863, new_n10873);
and_5  g08525(new_n10873, new_n10862, new_n10874_1);
or_5   g08526(new_n10874_1, new_n10860, new_n10875);
and_5  g08527(new_n10875, new_n10858, new_n10876);
nand_5 g08528(new_n10876, new_n10853, new_n10877);
and_5  g08529(new_n10877, new_n10852, new_n10878);
xor_4  g08530(new_n10878, new_n10848, new_n10879);
xor_4  g08531(new_n10879, new_n5672, new_n10880);
xor_4  g08532(new_n10876, new_n10853, new_n10881);
not_10 g08533(new_n10881, new_n10882);
nand_5 g08534(new_n10882, new_n5678, new_n10883);
xor_4  g08535(new_n10882, new_n5678, new_n10884);
xor_4  g08536(new_n10874_1, new_n10860, new_n10885);
nor_5  g08537(new_n10885, new_n5684, new_n10886);
xor_4  g08538(new_n10872, new_n10863, new_n10887);
nand_5 g08539(new_n10887, new_n5689, new_n10888);
xnor_4 g08540(new_n10887, new_n5688, new_n10889);
xor_4  g08541(new_n10870, new_n10866, new_n10890);
and_5  g08542(new_n10890, new_n5697, new_n10891);
and_5  g08543(new_n5832, new_n5863, new_n10892);
and_5  g08544(new_n5848, new_n5833_1, new_n10893);
or_5   g08545(new_n10893, new_n10892, new_n10894);
xnor_4 g08546(new_n10890, new_n5696_1, new_n10895);
and_5  g08547(new_n10895, new_n10894, new_n10896);
nor_5  g08548(new_n10896, new_n10891, new_n10897);
nand_5 g08549(new_n10897, new_n10889, new_n10898);
and_5  g08550(new_n10898, new_n10888, new_n10899);
xnor_4 g08551(new_n10885, new_n5683, new_n10900);
and_5  g08552(new_n10900, new_n10899, new_n10901);
nor_5  g08553(new_n10901, new_n10886, new_n10902);
nand_5 g08554(new_n10902, new_n10884, new_n10903);
and_5  g08555(new_n10903, new_n10883, new_n10904);
xor_4  g08556(new_n10904, new_n10880, n1385);
xor_4  g08557(n26808, n24732, new_n10906);
and_5  g08558(n26808, n24732, new_n10907);
xor_4  g08559(n7339, n6631, new_n10908);
xnor_4 g08560(new_n10908, new_n10907, new_n10909);
not_10 g08561(new_n10909, new_n10910);
nor_5  g08562(new_n10910, new_n10906, new_n10911);
xnor_4 g08563(n14684, n1667, new_n10912);
or_5   g08564(n7339, n6631, new_n10913);
not_10 g08565(new_n10907, new_n10914);
nand_5 g08566(new_n10908, new_n10914, new_n10915);
and_5  g08567(new_n10915, new_n10913, new_n10916);
xor_4  g08568(new_n10916, new_n10912, new_n10917);
and_5  g08569(new_n10917, new_n10911, new_n10918);
xnor_4 g08570(n17035, n2680, new_n10919);
or_5   g08571(n14684, n1667, new_n10920);
or_5   g08572(new_n10916, new_n10912, new_n10921);
and_5  g08573(new_n10921, new_n10920, new_n10922);
xor_4  g08574(new_n10922, new_n10919, new_n10923);
and_5  g08575(new_n10923, new_n10918, new_n10924_1);
xnor_4 g08576(n19905, n2547, new_n10925);
or_5   g08577(n17035, n2680, new_n10926);
or_5   g08578(new_n10922, new_n10919, new_n10927);
and_5  g08579(new_n10927, new_n10926, new_n10928);
xor_4  g08580(new_n10928, new_n10925, new_n10929);
and_5  g08581(new_n10929, new_n10924_1, new_n10930);
xor_4  g08582(n26452, n2999, new_n10931);
not_10 g08583(new_n10931, new_n10932);
or_5   g08584(n19905, n2547, new_n10933);
or_5   g08585(new_n10928, new_n10925, new_n10934);
and_5  g08586(new_n10934, new_n10933, new_n10935);
xor_4  g08587(new_n10935, new_n10932, new_n10936);
and_5  g08588(new_n10936, new_n10930, new_n10937);
xor_4  g08589(n15546, n14702, new_n10938);
not_10 g08590(new_n10938, new_n10939);
or_5   g08591(n26452, n2999, new_n10940);
or_5   g08592(new_n10935, new_n10932, new_n10941);
and_5  g08593(new_n10941, new_n10940, new_n10942);
xor_4  g08594(new_n10942, new_n10939, new_n10943_1);
and_5  g08595(new_n10943_1, new_n10937, new_n10944);
xor_4  g08596(n13914, n5077, new_n10945);
not_10 g08597(new_n10945, new_n10946);
or_5   g08598(n15546, n14702, new_n10947);
or_5   g08599(new_n10942, new_n10939, new_n10948);
and_5  g08600(new_n10948, new_n10947, new_n10949);
xor_4  g08601(new_n10949, new_n10946, new_n10950);
and_5  g08602(new_n10950, new_n10944, new_n10951);
xor_4  g08603(n18035, n3279, new_n10952);
not_10 g08604(new_n10952, new_n10953);
or_5   g08605(n13914, n5077, new_n10954);
or_5   g08606(new_n10949, new_n10946, new_n10955);
and_5  g08607(new_n10955, new_n10954, new_n10956);
xor_4  g08608(new_n10956, new_n10953, new_n10957);
and_5  g08609(new_n10957, new_n10951, new_n10958);
xor_4  g08610(n8827, n4306, new_n10959);
not_10 g08611(new_n10959, new_n10960);
or_5   g08612(n18035, n3279, new_n10961_1);
or_5   g08613(new_n10956, new_n10953, new_n10962);
and_5  g08614(new_n10962, new_n10961_1, new_n10963);
xor_4  g08615(new_n10963, new_n10960, new_n10964);
xor_4  g08616(new_n10964, new_n10958, new_n10965);
not_10 g08617(new_n10965, new_n10966);
xnor_4 g08618(new_n10966, new_n8092, new_n10967);
xor_4  g08619(new_n10957, new_n10951, new_n10968);
nor_5  g08620(new_n10968, new_n8098, new_n10969);
xor_4  g08621(new_n10968, new_n8097, new_n10970);
not_10 g08622(new_n10950, new_n10971);
xnor_4 g08623(new_n10971, new_n10944, new_n10972);
or_5   g08624(new_n10972, new_n8104, new_n10973);
xor_4  g08625(new_n10972, new_n8103_1, new_n10974);
not_10 g08626(new_n10943_1, new_n10975);
xnor_4 g08627(new_n10975, new_n10937, new_n10976);
or_5   g08628(new_n10976, new_n8110, new_n10977);
xor_4  g08629(new_n10976, new_n8109_1, new_n10978);
not_10 g08630(new_n10936, new_n10979);
xnor_4 g08631(new_n10979, new_n10930, new_n10980);
or_5   g08632(new_n10980, new_n8116, new_n10981);
xor_4  g08633(new_n10980, new_n8115, new_n10982);
xor_4  g08634(new_n10929, new_n10924_1, new_n10983);
or_5   g08635(new_n10983, new_n8122, new_n10984);
xor_4  g08636(new_n10983, new_n8121, new_n10985);
xor_4  g08637(new_n10923, new_n10918, new_n10986);
or_5   g08638(new_n10986, new_n8127_1, new_n10987);
xor_4  g08639(new_n10986, new_n8126, new_n10988);
xor_4  g08640(new_n10917, new_n10911, new_n10989);
or_5   g08641(new_n10989, new_n8132, new_n10990);
xor_4  g08642(new_n10989, new_n8131, new_n10991);
and_5  g08643(new_n10906, new_n2546, new_n10992);
or_5   g08644(new_n10992, new_n8140, new_n10993);
and_5  g08645(new_n10908, new_n10906, new_n10994);
nor_5  g08646(new_n10994, new_n10911, new_n10995);
not_10 g08647(new_n10995, new_n10996);
nand_5 g08648(new_n10992, new_n8075, new_n10997);
and_5  g08649(new_n10997, new_n10993, new_n10998);
nand_5 g08650(new_n10998, new_n10996, new_n10999);
and_5  g08651(new_n10999, new_n10993, new_n11000);
or_5   g08652(new_n11000, new_n10991, new_n11001);
and_5  g08653(new_n11001, new_n10990, new_n11002);
or_5   g08654(new_n11002, new_n10988, new_n11003);
and_5  g08655(new_n11003, new_n10987, new_n11004);
or_5   g08656(new_n11004, new_n10985, new_n11005_1);
and_5  g08657(new_n11005_1, new_n10984, new_n11006);
or_5   g08658(new_n11006, new_n10982, new_n11007);
and_5  g08659(new_n11007, new_n10981, new_n11008);
or_5   g08660(new_n11008, new_n10978, new_n11009);
and_5  g08661(new_n11009, new_n10977, new_n11010);
or_5   g08662(new_n11010, new_n10974, new_n11011_1);
and_5  g08663(new_n11011_1, new_n10973, new_n11012);
nor_5  g08664(new_n11012, new_n10970, new_n11013);
nor_5  g08665(new_n11013, new_n10969, new_n11014);
xor_4  g08666(new_n11014, new_n10967, new_n11015);
xor_4  g08667(new_n11015, new_n9353, new_n11016);
not_10 g08668(new_n11016, new_n11017);
xor_4  g08669(new_n11012, new_n10970, new_n11018);
and_5  g08670(new_n11018, new_n9356, new_n11019);
xor_4  g08671(new_n11018, new_n9356, new_n11020);
not_10 g08672(new_n11020, new_n11021);
xor_4  g08673(new_n11010, new_n10974, new_n11022);
and_5  g08674(new_n11022, new_n9360, new_n11023_1);
xor_4  g08675(new_n11022, new_n9360, new_n11024);
not_10 g08676(new_n11024, new_n11025_1);
xor_4  g08677(new_n11008, new_n10978, new_n11026);
and_5  g08678(new_n11026, new_n9364_1, new_n11027);
xor_4  g08679(new_n11026, new_n9364_1, new_n11028);
not_10 g08680(new_n11028, new_n11029);
xor_4  g08681(new_n11006, new_n10982, new_n11030);
and_5  g08682(new_n11030, new_n9368, new_n11031);
xor_4  g08683(new_n11030, new_n9368, new_n11032);
not_10 g08684(new_n11032, new_n11033);
xor_4  g08685(new_n11004, new_n10985, new_n11034);
and_5  g08686(new_n11034, new_n9371_1, new_n11035);
xor_4  g08687(new_n11034, new_n9371_1, new_n11036);
not_10 g08688(new_n11036, new_n11037);
xor_4  g08689(new_n11002, new_n10988, new_n11038);
and_5  g08690(new_n11038, new_n9375, new_n11039);
not_10 g08691(new_n9379, new_n11040);
xor_4  g08692(new_n11000, new_n10991, new_n11041);
and_5  g08693(new_n11041, new_n11040, new_n11042);
xnor_4 g08694(new_n11041, new_n9379, new_n11043);
not_10 g08695(new_n11043, new_n11044_1);
xor_4  g08696(new_n10906, new_n2546, new_n11045);
nor_5  g08697(new_n11045, new_n9387, new_n11046);
not_10 g08698(new_n11046, new_n11047);
nor_5  g08699(new_n11047, new_n9384, new_n11048);
not_10 g08700(new_n11048, new_n11049);
xor_4  g08701(new_n11047, new_n9384, new_n11050);
xor_4  g08702(new_n10998, new_n10996, new_n11051);
and_5  g08703(new_n11051, new_n11050, new_n11052);
not_10 g08704(new_n11052, new_n11053);
and_5  g08705(new_n11053, new_n11049, new_n11054);
nor_5  g08706(new_n11054, new_n11044_1, new_n11055);
nor_5  g08707(new_n11055, new_n11042, new_n11056_1);
xor_4  g08708(new_n11038, new_n9375, new_n11057);
not_10 g08709(new_n11057, new_n11058);
nor_5  g08710(new_n11058, new_n11056_1, new_n11059);
nor_5  g08711(new_n11059, new_n11039, new_n11060);
nor_5  g08712(new_n11060, new_n11037, new_n11061);
nor_5  g08713(new_n11061, new_n11035, new_n11062);
nor_5  g08714(new_n11062, new_n11033, new_n11063_1);
nor_5  g08715(new_n11063_1, new_n11031, new_n11064);
nor_5  g08716(new_n11064, new_n11029, new_n11065);
nor_5  g08717(new_n11065, new_n11027, new_n11066);
nor_5  g08718(new_n11066, new_n11025_1, new_n11067);
nor_5  g08719(new_n11067, new_n11023_1, new_n11068);
nor_5  g08720(new_n11068, new_n11021, new_n11069);
nor_5  g08721(new_n11069, new_n11019, new_n11070);
xnor_4 g08722(new_n11070, new_n11017, n1498);
xor_4  g08723(n20658, n9090, new_n11072);
xor_4  g08724(new_n11072, new_n6009, new_n11073);
xor_4  g08725(new_n11073, new_n5024_1, n1501);
not_10 g08726(n752, new_n11075);
not_10 g08727(n1611, new_n11076);
not_10 g08728(n25094, new_n11077);
not_10 g08729(n21538, new_n11078_1);
not_10 g08730(n5131, new_n11079);
nor_5  g08731(n15506, n11473, new_n11080_1);
and_5  g08732(new_n11080_1, new_n11079, new_n11081);
and_5  g08733(new_n11081, new_n11078_1, new_n11082);
and_5  g08734(new_n11082, new_n11077, new_n11083);
and_5  g08735(new_n11083, new_n11076, new_n11084);
xor_4  g08736(new_n11084, new_n11075, new_n11085);
xnor_4 g08737(new_n11085, new_n9900, new_n11086);
xor_4  g08738(new_n11083, n1611, new_n11087);
nand_5 g08739(new_n11087, new_n9904, new_n11088);
xor_4  g08740(new_n11083, new_n11076, new_n11089);
xnor_4 g08741(new_n11089, new_n9904, new_n11090);
not_10 g08742(new_n11090, new_n11091);
xor_4  g08743(new_n11082, new_n11077, new_n11092);
or_5   g08744(new_n11092, new_n9911, new_n11093);
xor_4  g08745(new_n11092, new_n9911, new_n11094_1);
xor_4  g08746(new_n11081, new_n11078_1, new_n11095);
nand_5 g08747(new_n11095, new_n9914, new_n11096);
xor_4  g08748(new_n11080_1, new_n11079, new_n11097);
or_5   g08749(new_n11097, new_n9919_1, new_n11098);
xor_4  g08750(new_n11097, new_n9921, new_n11099);
not_10 g08751(n15506, new_n11100);
nor_5  g08752(new_n9927, new_n11100, new_n11101_1);
xor_4  g08753(n15506, n11473, new_n11102);
or_5   g08754(new_n11102, new_n11101_1, new_n11103_1);
not_10 g08755(n11473, new_n11104);
nand_5 g08756(new_n11101_1, new_n11104, new_n11105);
and_5  g08757(new_n11105, new_n11103_1, new_n11106);
nand_5 g08758(new_n11106, new_n9924, new_n11107);
and_5  g08759(new_n11107, new_n11103_1, new_n11108);
or_5   g08760(new_n11108, new_n11099, new_n11109);
and_5  g08761(new_n11109, new_n11098, new_n11110);
xor_4  g08762(new_n11095, new_n9914, new_n11111);
nand_5 g08763(new_n11111, new_n11110, new_n11112);
and_5  g08764(new_n11112, new_n11096, new_n11113);
nand_5 g08765(new_n11113, new_n11094_1, new_n11114);
and_5  g08766(new_n11114, new_n11093, new_n11115);
or_5   g08767(new_n11115, new_n11091, new_n11116);
and_5  g08768(new_n11116, new_n11088, new_n11117);
xor_4  g08769(new_n11117, new_n11086, new_n11118);
not_10 g08770(new_n11118, new_n11119);
xor_4  g08771(n20470, n3366, new_n11120_1);
nand_5 g08772(n26565, n21222, new_n11121_1);
or_5   g08773(n26565, n21222, new_n11122);
nor_5  g08774(n9832, n3959, new_n11123);
nor_5  g08775(new_n9735, new_n9721, new_n11124);
nor_5  g08776(new_n11124, new_n11123, new_n11125);
nand_5 g08777(new_n11125, new_n11122, new_n11126);
and_5  g08778(new_n11126, new_n11121_1, new_n11127_1);
xor_4  g08779(new_n11127_1, new_n11120_1, new_n11128);
not_10 g08780(new_n11128, new_n11129);
xor_4  g08781(new_n11129, new_n11119, new_n11130);
xor_4  g08782(new_n11115, new_n11091, new_n11131);
xor_4  g08783(n26565, n21222, new_n11132_1);
xor_4  g08784(new_n11132_1, new_n11125, new_n11133);
and_5  g08785(new_n11133, new_n11131, new_n11134_1);
xor_4  g08786(new_n11133, new_n11131, new_n11135);
not_10 g08787(new_n11135, new_n11136);
xor_4  g08788(new_n11113, new_n11094_1, new_n11137);
and_5  g08789(new_n11137, new_n9737, new_n11138_1);
xor_4  g08790(new_n11137, new_n9737, new_n11139);
not_10 g08791(new_n11139, new_n11140);
xor_4  g08792(new_n11111, new_n11110, new_n11141);
nor_5  g08793(new_n11141, new_n9788, new_n11142);
not_10 g08794(new_n11142, new_n11143);
xor_4  g08795(new_n11141, new_n9788, new_n11144);
not_10 g08796(new_n9793, new_n11145);
xor_4  g08797(new_n11108, new_n11099, new_n11146);
nor_5  g08798(new_n11146, new_n11145, new_n11147);
not_10 g08799(new_n9799, new_n11148);
xor_4  g08800(new_n11106, new_n9924, new_n11149);
nand_5 g08801(new_n11149, new_n11148, new_n11150);
xor_4  g08802(new_n9927, new_n11100, new_n11151);
nor_5  g08803(new_n11151, new_n7245, new_n11152);
xnor_4 g08804(new_n11149, new_n9799, new_n11153);
nand_5 g08805(new_n11153, new_n11152, new_n11154);
and_5  g08806(new_n11154, new_n11150, new_n11155);
xnor_4 g08807(new_n11146, new_n9793, new_n11156);
and_5  g08808(new_n11156, new_n11155, new_n11157);
nor_5  g08809(new_n11157, new_n11147, new_n11158);
and_5  g08810(new_n11158, new_n11144, new_n11159);
not_10 g08811(new_n11159, new_n11160);
and_5  g08812(new_n11160, new_n11143, new_n11161);
nor_5  g08813(new_n11161, new_n11140, new_n11162);
nor_5  g08814(new_n11162, new_n11138_1, new_n11163);
nor_5  g08815(new_n11163, new_n11136, new_n11164);
nor_5  g08816(new_n11164, new_n11134_1, new_n11165);
xor_4  g08817(new_n11165, new_n11130, n1518);
not_10 g08818(n14826, new_n11167);
and_5  g08819(n17458, new_n11167, new_n11168);
not_10 g08820(new_n11168, new_n11169);
xor_4  g08821(n17458, n14826, new_n11170);
not_10 g08822(n1222, new_n11171);
or_5   g08823(n23493, new_n11171, new_n11172);
xnor_4 g08824(n23493, n1222, new_n11173);
not_10 g08825(new_n11173, new_n11174);
not_10 g08826(n25240, new_n11175);
or_5   g08827(new_n11175, n10275, new_n11176);
xnor_4 g08828(n25240, n10275, new_n11177);
not_10 g08829(new_n11177, new_n11178);
not_10 g08830(n10125, new_n11179);
or_5   g08831(n15146, new_n11179, new_n11180);
xnor_4 g08832(n15146, n10125, new_n11181);
not_10 g08833(new_n11181, new_n11182_1);
not_10 g08834(n8067, new_n11183);
or_5   g08835(n11579, new_n11183, new_n11184_1);
xnor_4 g08836(n11579, n8067, new_n11185);
not_10 g08837(new_n11185, new_n11186);
not_10 g08838(n20923, new_n11187);
or_5   g08839(new_n11187, n21, new_n11188);
xor_4  g08840(n20923, n21, new_n11189);
not_10 g08841(n18157, new_n11190);
or_5   g08842(new_n11190, n1682, new_n11191);
xnor_4 g08843(n18157, n1682, new_n11192_1);
and_5  g08844(new_n7268_1, n7963, new_n11193);
or_5   g08845(new_n7268_1, n7963, new_n11194);
and_5  g08846(n10017, new_n7272, new_n11195);
nor_5  g08847(n10017, new_n7272, new_n11196);
and_5  g08848(new_n7274, n3618, new_n11197);
not_10 g08849(new_n11197, new_n11198);
nor_5  g08850(new_n11198, new_n11196, new_n11199);
nor_5  g08851(new_n11199, new_n11195, new_n11200);
not_10 g08852(new_n11200, new_n11201_1);
and_5  g08853(new_n11201_1, new_n11194, new_n11202);
nor_5  g08854(new_n11202, new_n11193, new_n11203);
nand_5 g08855(new_n11203, new_n11192_1, new_n11204);
and_5  g08856(new_n11204, new_n11191, new_n11205);
or_5   g08857(new_n11205, new_n11189, new_n11206);
and_5  g08858(new_n11206, new_n11188, new_n11207);
or_5   g08859(new_n11207, new_n11186, new_n11208);
and_5  g08860(new_n11208, new_n11184_1, new_n11209);
or_5   g08861(new_n11209, new_n11182_1, new_n11210);
and_5  g08862(new_n11210, new_n11180, new_n11211);
or_5   g08863(new_n11211, new_n11178, new_n11212);
and_5  g08864(new_n11212, new_n11176, new_n11213);
or_5   g08865(new_n11213, new_n11174, new_n11214);
and_5  g08866(new_n11214, new_n11172, new_n11215);
nor_5  g08867(new_n11215, new_n11170, new_n11216);
not_10 g08868(new_n11216, new_n11217);
and_5  g08869(new_n11217, new_n11169, new_n11218);
not_10 g08870(n2944, new_n11219);
not_10 g08871(n767, new_n11220_1);
not_10 g08872(n7330, new_n11221);
not_10 g08873(n22492, new_n11222);
not_10 g08874(n12821, new_n11223_1);
and_5  g08875(new_n4196, new_n4192, new_n11224);
and_5  g08876(new_n11224, new_n11223_1, new_n11225);
and_5  g08877(new_n11225, new_n11222, new_n11226);
and_5  g08878(new_n11226, new_n11221, new_n11227);
and_5  g08879(new_n11227, new_n11220_1, new_n11228);
xor_4  g08880(new_n11228, new_n11219, new_n11229);
nand_5 g08881(new_n11229, n19282, new_n11230);
nand_5 g08882(new_n11228, new_n11219, new_n11231);
xor_4  g08883(new_n11227, new_n11220_1, new_n11232);
nor_5  g08884(new_n11232, n12657, new_n11233);
xor_4  g08885(new_n11232, n12657, new_n11234_1);
xor_4  g08886(new_n11226, new_n11221, new_n11235);
nand_5 g08887(new_n11235, n17077, new_n11236);
xor_4  g08888(new_n11235, n17077, new_n11237);
not_10 g08889(new_n11237, new_n11238);
xor_4  g08890(new_n11225, new_n11222, new_n11239);
nand_5 g08891(new_n11239, n26510, new_n11240);
xnor_4 g08892(new_n11239, n26510, new_n11241);
xor_4  g08893(new_n11224, new_n11223_1, new_n11242);
nand_5 g08894(new_n11242, n23068, new_n11243);
nor_5  g08895(new_n11242, n23068, new_n11244);
and_5  g08896(new_n4197, n19514, new_n11245_1);
nor_5  g08897(new_n4217, new_n4199, new_n11246);
nor_5  g08898(new_n11246, new_n11245_1, new_n11247);
or_5   g08899(new_n11247, new_n11244, new_n11248);
and_5  g08900(new_n11248, new_n11243, new_n11249);
or_5   g08901(new_n11249, new_n11241, new_n11250);
and_5  g08902(new_n11250, new_n11240, new_n11251);
or_5   g08903(new_n11251, new_n11238, new_n11252);
and_5  g08904(new_n11252, new_n11236, new_n11253);
and_5  g08905(new_n11253, new_n11234_1, new_n11254);
nor_5  g08906(new_n11254, new_n11233, new_n11255);
or_5   g08907(new_n11229, n19282, new_n11256);
nand_5 g08908(new_n11256, new_n11255, new_n11257);
and_5  g08909(new_n11257, new_n11231, new_n11258);
and_5  g08910(new_n11258, new_n11230, new_n11259);
or_5   g08911(new_n11259, new_n11218, new_n11260);
xor_4  g08912(new_n11215, new_n11170, new_n11261_1);
xor_4  g08913(new_n11229, n19282, new_n11262);
xnor_4 g08914(new_n11262, new_n11255, new_n11263);
not_10 g08915(new_n11263, new_n11264);
or_5   g08916(new_n11264, new_n11261_1, new_n11265);
xnor_4 g08917(new_n11264, new_n11261_1, new_n11266_1);
xor_4  g08918(new_n11213, new_n11174, new_n11267);
xor_4  g08919(new_n11253, new_n11234_1, new_n11268);
not_10 g08920(new_n11268, new_n11269);
or_5   g08921(new_n11269, new_n11267, new_n11270);
xnor_4 g08922(new_n11269, new_n11267, new_n11271);
xor_4  g08923(new_n11211, new_n11178, new_n11272);
not_10 g08924(new_n11272, new_n11273_1);
xor_4  g08925(new_n11251, new_n11238, new_n11274);
not_10 g08926(new_n11274, new_n11275_1);
nand_5 g08927(new_n11275_1, new_n11273_1, new_n11276);
xnor_4 g08928(new_n11275_1, new_n11273_1, new_n11277);
xor_4  g08929(new_n11209, new_n11182_1, new_n11278);
xor_4  g08930(new_n11249, new_n11241, new_n11279);
or_5   g08931(new_n11279, new_n11278, new_n11280);
not_10 g08932(new_n11278, new_n11281);
xor_4  g08933(new_n11279, new_n11281, new_n11282);
xor_4  g08934(new_n11207, new_n11186, new_n11283);
xor_4  g08935(new_n11242, n23068, new_n11284);
xnor_4 g08936(new_n11284, new_n11247, new_n11285);
or_5   g08937(new_n11285, new_n11283, new_n11286);
not_10 g08938(new_n11283, new_n11287);
xor_4  g08939(new_n11285, new_n11287, new_n11288);
xor_4  g08940(new_n11205, new_n11189, new_n11289);
or_5   g08941(new_n11289, new_n4218, new_n11290_1);
xor_4  g08942(new_n11203, new_n11192_1, new_n11291);
nor_5  g08943(new_n11291, new_n4249, new_n11292);
xor_4  g08944(new_n11291, new_n4250, new_n11293);
not_10 g08945(new_n4268, new_n11294);
xnor_4 g08946(n12161, n7963, new_n11295);
xor_4  g08947(new_n11295, new_n11201_1, new_n11296);
nand_5 g08948(new_n11296, new_n11294, new_n11297);
xnor_4 g08949(new_n11296, new_n11294, new_n11298);
xnor_4 g08950(n8581, n3618, new_n11299);
not_10 g08951(new_n11299, new_n11300);
and_5  g08952(new_n11300, new_n4262, new_n11301);
not_10 g08953(new_n11301, new_n11302_1);
xnor_4 g08954(n10017, n5026, new_n11303);
xnor_4 g08955(new_n11303, new_n11198, new_n11304);
nand_5 g08956(new_n11304, new_n11302_1, new_n11305);
xor_4  g08957(new_n11304, new_n11302_1, new_n11306);
nand_5 g08958(new_n11306, new_n4258, new_n11307);
and_5  g08959(new_n11307, new_n11305, new_n11308);
or_5   g08960(new_n11308, new_n11298, new_n11309);
and_5  g08961(new_n11309, new_n11297, new_n11310);
nor_5  g08962(new_n11310, new_n11293, new_n11311);
or_5   g08963(new_n11311, new_n11292, new_n11312);
xnor_4 g08964(new_n11289, new_n4219, new_n11313_1);
nand_5 g08965(new_n11313_1, new_n11312, new_n11314);
and_5  g08966(new_n11314, new_n11290_1, new_n11315);
or_5   g08967(new_n11315, new_n11288, new_n11316);
and_5  g08968(new_n11316, new_n11286, new_n11317);
or_5   g08969(new_n11317, new_n11282, new_n11318);
and_5  g08970(new_n11318, new_n11280, new_n11319);
or_5   g08971(new_n11319, new_n11277, new_n11320);
and_5  g08972(new_n11320, new_n11276, new_n11321);
or_5   g08973(new_n11321, new_n11271, new_n11322);
and_5  g08974(new_n11322, new_n11270, new_n11323);
or_5   g08975(new_n11323, new_n11266_1, new_n11324);
and_5  g08976(new_n11324, new_n11265, new_n11325_1);
xor_4  g08977(new_n11259, new_n11218, new_n11326_1);
nand_5 g08978(new_n11326_1, new_n11325_1, new_n11327);
and_5  g08979(new_n11327, new_n11260, new_n11328);
not_10 g08980(n20040, new_n11329);
and_5  g08981(new_n11329, n2978, new_n11330_1);
not_10 g08982(new_n11330_1, new_n11331);
nor_5  g08983(new_n8890, new_n8848, new_n11332);
not_10 g08984(new_n11332, new_n11333);
and_5  g08985(new_n11333, new_n11331, new_n11334);
xor_4  g08986(new_n11334, new_n11328, new_n11335);
xor_4  g08987(new_n11326_1, new_n11325_1, new_n11336);
nor_5  g08988(new_n11336, new_n11334, new_n11337);
xor_4  g08989(new_n11323, new_n11266_1, new_n11338);
and_5  g08990(new_n11338, new_n8892, new_n11339);
xor_4  g08991(new_n11338, new_n8892, new_n11340);
not_10 g08992(new_n11340, new_n11341);
xor_4  g08993(new_n11321, new_n11271, new_n11342);
and_5  g08994(new_n11342, new_n8958, new_n11343);
xor_4  g08995(new_n11342, new_n8958, new_n11344);
not_10 g08996(new_n11344, new_n11345);
xor_4  g08997(new_n11319, new_n11277, new_n11346);
and_5  g08998(new_n11346, new_n8965, new_n11347_1);
xor_4  g08999(new_n11346, new_n8965, new_n11348_1);
not_10 g09000(new_n11348_1, new_n11349);
xor_4  g09001(new_n11317, new_n11282, new_n11350);
and_5  g09002(new_n11350, new_n8968, new_n11351);
xor_4  g09003(new_n11350, new_n8968, new_n11352_1);
not_10 g09004(new_n11352_1, new_n11353);
xor_4  g09005(new_n11315, new_n11288, new_n11354);
and_5  g09006(new_n11354, new_n8973, new_n11355);
not_10 g09007(new_n11355, new_n11356_1);
xor_4  g09008(new_n11354, new_n8973, new_n11357);
xor_4  g09009(new_n11313_1, new_n11312, new_n11358);
nor_5  g09010(new_n11358, new_n8978, new_n11359);
xor_4  g09011(new_n11310, new_n11293, new_n11360);
nand_5 g09012(new_n11360, new_n8984, new_n11361);
xor_4  g09013(new_n11360, new_n8984, new_n11362);
not_10 g09014(new_n11362, new_n11363);
xor_4  g09015(new_n11308, new_n11298, new_n11364);
nand_5 g09016(new_n11364, new_n8990, new_n11365);
not_10 g09017(new_n8996, new_n11366);
xnor_4 g09018(new_n11299, new_n4262, new_n11367);
and_5  g09019(new_n11367, new_n8999, new_n11368);
and_5  g09020(new_n11368, new_n11366, new_n11369);
xor_4  g09021(new_n11306, new_n4258, new_n11370);
xor_4  g09022(new_n11368, new_n8996, new_n11371);
nor_5  g09023(new_n11371, new_n11370, new_n11372);
or_5   g09024(new_n11372, new_n11369, new_n11373);
xor_4  g09025(new_n11364, new_n8990, new_n11374);
not_10 g09026(new_n11374, new_n11375_1);
or_5   g09027(new_n11375_1, new_n11373, new_n11376);
and_5  g09028(new_n11376, new_n11365, new_n11377);
or_5   g09029(new_n11377, new_n11363, new_n11378);
and_5  g09030(new_n11378, new_n11361, new_n11379_1);
xor_4  g09031(new_n11358, new_n8978, new_n11380);
and_5  g09032(new_n11380, new_n11379_1, new_n11381);
nor_5  g09033(new_n11381, new_n11359, new_n11382);
and_5  g09034(new_n11382, new_n11357, new_n11383);
not_10 g09035(new_n11383, new_n11384);
and_5  g09036(new_n11384, new_n11356_1, new_n11385);
nor_5  g09037(new_n11385, new_n11353, new_n11386_1);
nor_5  g09038(new_n11386_1, new_n11351, new_n11387);
nor_5  g09039(new_n11387, new_n11349, new_n11388);
nor_5  g09040(new_n11388, new_n11347_1, new_n11389);
nor_5  g09041(new_n11389, new_n11345, new_n11390);
nor_5  g09042(new_n11390, new_n11343, new_n11391_1);
nor_5  g09043(new_n11391_1, new_n11341, new_n11392);
nor_5  g09044(new_n11392, new_n11339, new_n11393);
xor_4  g09045(new_n11336, new_n11334, new_n11394);
not_10 g09046(new_n11394, new_n11395);
nor_5  g09047(new_n11395, new_n11393, new_n11396);
nor_5  g09048(new_n11396, new_n11337, new_n11397);
xor_4  g09049(new_n11397, new_n11335, n1527);
xor_4  g09050(n25345, n23463, new_n11399);
not_10 g09051(n13074, new_n11400);
or_5   g09052(new_n11400, n9655, new_n11401);
xor_4  g09053(n13074, n9655, new_n11402);
not_10 g09054(n10739, new_n11403_1);
or_5   g09055(n13490, new_n11403_1, new_n11404);
xor_4  g09056(n13490, n10739, new_n11405);
or_5   g09057(n22660, new_n2350, new_n11406);
xor_4  g09058(n22660, n21753, new_n11407);
or_5   g09059(new_n2354, n1777, new_n11408);
xor_4  g09060(n21832, n1777, new_n11409);
or_5   g09061(new_n2358, n8745, new_n11410);
or_5   g09062(n16223, new_n6823, new_n11411);
or_5   g09063(new_n9960, new_n9955, new_n11412);
and_5  g09064(new_n11412, new_n11411, new_n11413);
xnor_4 g09065(n26913, n8745, new_n11414);
nand_5 g09066(new_n11414, new_n11413, new_n11415);
and_5  g09067(new_n11415, new_n11410, new_n11416);
or_5   g09068(new_n11416, new_n11409, new_n11417);
and_5  g09069(new_n11417, new_n11408, new_n11418);
or_5   g09070(new_n11418, new_n11407, new_n11419_1);
and_5  g09071(new_n11419_1, new_n11406, new_n11420);
or_5   g09072(new_n11420, new_n11405, new_n11421);
and_5  g09073(new_n11421, new_n11404, new_n11422);
or_5   g09074(new_n11422, new_n11402, new_n11423);
and_5  g09075(new_n11423, new_n11401, new_n11424_1);
xor_4  g09076(new_n11424_1, new_n11399, new_n11425);
xor_4  g09077(new_n11425, new_n7985, new_n11426);
xor_4  g09078(new_n11422, new_n11402, new_n11427);
or_5   g09079(new_n11427, new_n7991, new_n11428);
xor_4  g09080(new_n11427, new_n7991, new_n11429);
xor_4  g09081(new_n11420, new_n11405, new_n11430);
or_5   g09082(new_n11430, new_n7997, new_n11431);
xor_4  g09083(new_n11430, new_n7997, new_n11432);
xor_4  g09084(new_n11418, new_n11407, new_n11433);
or_5   g09085(new_n11433, new_n8005, new_n11434);
xor_4  g09086(new_n11433, new_n8005, new_n11435);
xor_4  g09087(new_n11416, new_n11409, new_n11436);
or_5   g09088(new_n11436, new_n8010, new_n11437);
xor_4  g09089(new_n11436, new_n8010, new_n11438);
xor_4  g09090(new_n11414, new_n11413, new_n11439_1);
or_5   g09091(new_n11439_1, new_n9947, new_n11440);
nand_5 g09092(new_n9961, new_n8017, new_n11441);
nand_5 g09093(new_n9971, new_n9962, new_n11442);
nand_5 g09094(new_n11442, new_n11441, new_n11443);
xor_4  g09095(new_n11439_1, new_n9947, new_n11444);
nand_5 g09096(new_n11444, new_n11443, new_n11445);
nand_5 g09097(new_n11445, new_n11440, new_n11446);
nand_5 g09098(new_n11446, new_n11438, new_n11447);
nand_5 g09099(new_n11447, new_n11437, new_n11448);
nand_5 g09100(new_n11448, new_n11435, new_n11449);
nand_5 g09101(new_n11449, new_n11434, new_n11450);
nand_5 g09102(new_n11450, new_n11432, new_n11451);
nand_5 g09103(new_n11451, new_n11431, new_n11452);
nand_5 g09104(new_n11452, new_n11429, new_n11453);
and_5  g09105(new_n11453, new_n11428, new_n11454);
xor_4  g09106(new_n11454, new_n11426, n1580);
xnor_4 g09107(n18962, n12315, new_n11456);
or_5   g09108(new_n11456, new_n7467, new_n11457);
and_5  g09109(n18962, new_n8548, new_n11458);
xnor_4 g09110(n10158, n3952, new_n11459);
xor_4  g09111(new_n11459, new_n11458, new_n11460);
xor_4  g09112(new_n11460, new_n11457, new_n11461);
xnor_4 g09113(new_n11461, new_n7473, n1586);
xnor_4 g09114(n19539, n1483, new_n11463);
not_10 g09115(new_n11463, new_n11464);
not_10 g09116(n8194, new_n11465);
or_5   g09117(n24093, new_n11465, new_n11466);
xnor_4 g09118(n24093, n8194, new_n11467);
not_10 g09119(new_n11467, new_n11468);
not_10 g09120(n23657, new_n11469);
or_5   g09121(new_n11469, n23035, new_n11470_1);
xnor_4 g09122(n23657, n23035, new_n11471);
not_10 g09123(new_n11471, new_n11472_1);
not_10 g09124(n16911, new_n11473_1);
or_5   g09125(new_n11473_1, n7773, new_n11474);
or_5   g09126(new_n6496, new_n6465_1, new_n11475);
and_5  g09127(new_n11475, new_n11474, new_n11476);
or_5   g09128(new_n11476, new_n11472_1, new_n11477);
and_5  g09129(new_n11477, new_n11470_1, new_n11478);
or_5   g09130(new_n11478, new_n11468, new_n11479_1);
and_5  g09131(new_n11479_1, new_n11466, new_n11480);
xor_4  g09132(new_n11480, new_n11464, new_n11481_1);
xnor_4 g09133(n25494, n1314, new_n11482);
not_10 g09134(new_n11482, new_n11483);
or_5   g09135(n10117, new_n8365, new_n11484);
xnor_4 g09136(n10117, n3306, new_n11485);
not_10 g09137(new_n11485, new_n11486_1);
or_5   g09138(new_n8372, n13460, new_n11487);
xnor_4 g09139(n22335, n13460, new_n11488);
not_10 g09140(new_n11488, new_n11489);
or_5   g09141(new_n8376_1, n6104, new_n11490);
and_5  g09142(new_n3437, n1525, new_n11491);
nor_5  g09143(new_n4666, new_n4640, new_n11492);
or_5   g09144(new_n11492, new_n11491, new_n11493);
xnor_4 g09145(n24048, n6104, new_n11494);
nand_5 g09146(new_n11494, new_n11493, new_n11495);
and_5  g09147(new_n11495, new_n11490, new_n11496_1);
or_5   g09148(new_n11496_1, new_n11489, new_n11497);
and_5  g09149(new_n11497, new_n11487, new_n11498);
or_5   g09150(new_n11498, new_n11486_1, new_n11499);
and_5  g09151(new_n11499, new_n11484, new_n11500);
xor_4  g09152(new_n11500, new_n11483, new_n11501);
not_10 g09153(new_n11501, new_n11502);
xnor_4 g09154(n25296, n23717, new_n11503_1);
not_10 g09155(new_n11503_1, new_n11504);
not_10 g09156(n7788, new_n11505);
or_5   g09157(n20013, new_n11505, new_n11506_1);
xnor_4 g09158(n20013, n7788, new_n11507);
not_10 g09159(new_n11507, new_n11508);
not_10 g09160(n5443, new_n11509);
or_5   g09161(new_n11509, n1320, new_n11510);
xor_4  g09162(n5443, n1320, new_n11511);
not_10 g09163(n18584, new_n11512);
or_5   g09164(n19803, new_n11512, new_n11513);
or_5   g09165(new_n6462, new_n6458, new_n11514);
and_5  g09166(new_n11514, new_n11513, new_n11515_1);
or_5   g09167(new_n11515_1, new_n11511, new_n11516);
and_5  g09168(new_n11516, new_n11510, new_n11517);
or_5   g09169(new_n11517, new_n11508, new_n11518);
and_5  g09170(new_n11518, new_n11506_1, new_n11519);
xor_4  g09171(new_n11519, new_n11504, new_n11520);
not_10 g09172(new_n11520, new_n11521);
xnor_4 g09173(new_n11521, new_n11502, new_n11522);
xor_4  g09174(new_n11498, new_n11486_1, new_n11523);
not_10 g09175(new_n11523, new_n11524);
xor_4  g09176(new_n11517, new_n11508, new_n11525);
not_10 g09177(new_n11525, new_n11526);
or_5   g09178(new_n11526, new_n11524, new_n11527);
xor_4  g09179(new_n11526, new_n11524, new_n11528);
xor_4  g09180(new_n11496_1, new_n11489, new_n11529);
xor_4  g09181(new_n11515_1, new_n11511, new_n11530);
or_5   g09182(new_n11530, new_n11529, new_n11531);
xor_4  g09183(new_n11530, new_n11529, new_n11532);
xor_4  g09184(new_n11494, new_n11493, new_n11533);
nand_5 g09185(new_n11533, new_n6463, new_n11534);
xnor_4 g09186(new_n11533, new_n6463, new_n11535);
nand_5 g09187(new_n4695, new_n4667, new_n11536);
or_5   g09188(new_n4730, new_n4696, new_n11537);
and_5  g09189(new_n11537, new_n11536, new_n11538_1);
or_5   g09190(new_n11538_1, new_n11535, new_n11539);
and_5  g09191(new_n11539, new_n11534, new_n11540);
nand_5 g09192(new_n11540, new_n11532, new_n11541);
and_5  g09193(new_n11541, new_n11531, new_n11542);
nand_5 g09194(new_n11542, new_n11528, new_n11543);
and_5  g09195(new_n11543, new_n11527, new_n11544);
xor_4  g09196(new_n11544, new_n11522, new_n11545);
xor_4  g09197(new_n11545, new_n11481_1, new_n11546);
xor_4  g09198(new_n11478, new_n11468, new_n11547);
xor_4  g09199(new_n11542, new_n11528, new_n11548_1);
or_5   g09200(new_n11548_1, new_n11547, new_n11549);
xor_4  g09201(new_n11548_1, new_n11547, new_n11550);
not_10 g09202(new_n11550, new_n11551);
xor_4  g09203(new_n11476, new_n11472_1, new_n11552);
xor_4  g09204(new_n11540, new_n11532, new_n11553);
not_10 g09205(new_n11553, new_n11554);
or_5   g09206(new_n11554, new_n11552, new_n11555);
xor_4  g09207(new_n11554, new_n11552, new_n11556);
xor_4  g09208(new_n11538_1, new_n11535, new_n11557);
or_5   g09209(new_n11557, new_n6497, new_n11558);
xor_4  g09210(new_n11557, new_n6497, new_n11559);
not_10 g09211(new_n11559, new_n11560);
or_5   g09212(new_n6553, new_n4731_1, new_n11561);
or_5   g09213(new_n6558_1, new_n4734, new_n11562);
xor_4  g09214(new_n6558_1, new_n4734, new_n11563);
not_10 g09215(new_n11563, new_n11564_1);
nand_5 g09216(new_n6564, new_n4738, new_n11565);
nand_5 g09217(new_n6569, new_n4741, new_n11566_1);
xnor_4 g09218(new_n6569, new_n4745_1, new_n11567);
nor_5  g09219(new_n6574, new_n4749, new_n11568);
not_10 g09220(new_n11568, new_n11569);
nand_5 g09221(new_n11569, new_n6578, new_n11570);
xnor_4 g09222(new_n11568, new_n6578, new_n11571);
not_10 g09223(new_n11571, new_n11572);
or_5   g09224(new_n11572, new_n4754, new_n11573);
nand_5 g09225(new_n11573, new_n11570, new_n11574);
nand_5 g09226(new_n11574, new_n11567, new_n11575);
and_5  g09227(new_n11575, new_n11566_1, new_n11576);
xor_4  g09228(new_n6564, new_n4738, new_n11577);
not_10 g09229(new_n11577, new_n11578);
or_5   g09230(new_n11578, new_n11576, new_n11579_1);
and_5  g09231(new_n11579_1, new_n11565, new_n11580_1);
or_5   g09232(new_n11580_1, new_n11564_1, new_n11581);
and_5  g09233(new_n11581, new_n11562, new_n11582);
xor_4  g09234(new_n6553, new_n4731_1, new_n11583);
not_10 g09235(new_n11583, new_n11584);
or_5   g09236(new_n11584, new_n11582, new_n11585);
and_5  g09237(new_n11585, new_n11561, new_n11586);
or_5   g09238(new_n11586, new_n11560, new_n11587);
nand_5 g09239(new_n11587, new_n11558, new_n11588);
nand_5 g09240(new_n11588, new_n11556, new_n11589);
and_5  g09241(new_n11589, new_n11555, new_n11590);
or_5   g09242(new_n11590, new_n11551, new_n11591_1);
and_5  g09243(new_n11591_1, new_n11549, new_n11592);
xor_4  g09244(new_n11592, new_n11546, n1590);
xor_4  g09245(new_n7703, new_n7684, n1602);
xor_4  g09246(new_n2831, new_n2779_1, n1634);
xnor_4 g09247(new_n11590, new_n11551, n1636);
nor_5  g09248(n10514, n4514, new_n11597);
not_10 g09249(new_n11597, new_n11598);
xor_4  g09250(n10514, n4514, new_n11599);
not_10 g09251(new_n11599, new_n11600);
or_5   g09252(n18649, n3984, new_n11601);
xor_4  g09253(n18649, n3984, new_n11602);
nand_5 g09254(n19652, n6218, new_n11603);
nor_5  g09255(n19652, n6218, new_n11604);
nor_5  g09256(n20470, n3366, new_n11605);
and_5  g09257(new_n11127_1, new_n11120_1, new_n11606);
or_5   g09258(new_n11606, new_n11605, new_n11607_1);
or_5   g09259(new_n11607_1, new_n11604, new_n11608);
and_5  g09260(new_n11608, new_n11603, new_n11609);
nand_5 g09261(new_n11609, new_n11602, new_n11610);
and_5  g09262(new_n11610, new_n11601, new_n11611);
nor_5  g09263(new_n11611, new_n11600, new_n11612);
not_10 g09264(new_n11612, new_n11613);
and_5  g09265(new_n11613, new_n11598, new_n11614);
xnor_4 g09266(n18880, n2978, new_n11615_1);
or_5   g09267(n25475, n23697, new_n11616);
or_5   g09268(new_n6804, new_n6775_1, new_n11617);
and_5  g09269(new_n11617, new_n11616, new_n11618);
xor_4  g09270(new_n11618, new_n11615_1, new_n11619);
nor_5  g09271(new_n11619, new_n11329, new_n11620);
xor_4  g09272(new_n11619, new_n11329, new_n11621);
not_10 g09273(new_n11621, new_n11622);
not_10 g09274(n19531, new_n11623);
or_5   g09275(new_n6805, new_n11623, new_n11624);
xor_4  g09276(new_n6805, new_n11623, new_n11625);
not_10 g09277(n18345, new_n11626);
nand_5 g09278(new_n6808, new_n11626, new_n11627);
xor_4  g09279(new_n6808, new_n11626, new_n11628);
not_10 g09280(new_n11628, new_n11629);
not_10 g09281(n13190, new_n11630_1);
nand_5 g09282(new_n6811, new_n11630_1, new_n11631);
xor_4  g09283(new_n6811, new_n11630_1, new_n11632);
not_10 g09284(n3460, new_n11633);
or_5   g09285(new_n6814_1, new_n11633, new_n11634);
not_10 g09286(n5226, new_n11635);
nor_5  g09287(new_n6816, new_n11635, new_n11636);
not_10 g09288(new_n11636, new_n11637);
nor_5  g09289(new_n9761_1, new_n9745, new_n11638);
not_10 g09290(new_n11638, new_n11639);
and_5  g09291(new_n11639, new_n11637, new_n11640);
xor_4  g09292(new_n6814_1, n3460, new_n11641);
or_5   g09293(new_n11641, new_n11640, new_n11642);
and_5  g09294(new_n11642, new_n11634, new_n11643);
nand_5 g09295(new_n11643, new_n11632, new_n11644);
and_5  g09296(new_n11644, new_n11631, new_n11645);
or_5   g09297(new_n11645, new_n11629, new_n11646);
and_5  g09298(new_n11646, new_n11627, new_n11647_1);
nand_5 g09299(new_n11647_1, new_n11625, new_n11648);
and_5  g09300(new_n11648, new_n11624, new_n11649);
nor_5  g09301(new_n11649, new_n11622, new_n11650);
nor_5  g09302(new_n11650, new_n11620, new_n11651);
not_10 g09303(new_n11651, new_n11652);
nor_5  g09304(n18880, n2978, new_n11653);
not_10 g09305(new_n11653, new_n11654);
nor_5  g09306(new_n11618, new_n11615_1, new_n11655);
not_10 g09307(new_n11655, new_n11656);
and_5  g09308(new_n11656, new_n11654, new_n11657);
xor_4  g09309(new_n11657, new_n11652, new_n11658);
not_10 g09310(n7569, new_n11659);
not_10 g09311(n17037, new_n11660);
not_10 g09312(n5386, new_n11661);
not_10 g09313(n26191, new_n11662);
not_10 g09314(n26512, new_n11663);
and_5  g09315(new_n9743, new_n9738, new_n11664);
and_5  g09316(new_n11664, new_n11663, new_n11665);
and_5  g09317(new_n11665, new_n11662, new_n11666);
and_5  g09318(new_n11666, new_n11661, new_n11667_1);
and_5  g09319(new_n11667_1, new_n11660, new_n11668);
and_5  g09320(new_n11668, new_n11659, new_n11669);
not_10 g09321(new_n11669, new_n11670);
xor_4  g09322(new_n11670, new_n11658, new_n11671);
xor_4  g09323(new_n11649, new_n11622, new_n11672);
xor_4  g09324(new_n11668, new_n11659, new_n11673);
nor_5  g09325(new_n11673, new_n11672, new_n11674_1);
xor_4  g09326(new_n11673, new_n11672, new_n11675);
not_10 g09327(new_n11675, new_n11676);
xor_4  g09328(new_n11647_1, new_n11625, new_n11677);
xor_4  g09329(new_n11667_1, new_n11660, new_n11678);
or_5   g09330(new_n11678, new_n11677, new_n11679);
not_10 g09331(new_n11677, new_n11680);
xnor_4 g09332(new_n11678, new_n11680, new_n11681);
xor_4  g09333(new_n11645, new_n11629, new_n11682_1);
xor_4  g09334(new_n11666, n5386, new_n11683);
nand_5 g09335(new_n11683, new_n11682_1, new_n11684);
xor_4  g09336(new_n11683, new_n11682_1, new_n11685);
not_10 g09337(new_n11685, new_n11686);
xor_4  g09338(new_n11643, new_n11632, new_n11687);
not_10 g09339(new_n11687, new_n11688);
xor_4  g09340(new_n11665, new_n11662, new_n11689);
or_5   g09341(new_n11689, new_n11688, new_n11690);
xor_4  g09342(new_n11664, new_n11663, new_n11691);
xor_4  g09343(new_n6814_1, new_n11633, new_n11692);
xnor_4 g09344(new_n11692, new_n11640, new_n11693);
nand_5 g09345(new_n11693, new_n11691, new_n11694);
not_10 g09346(new_n11693, new_n11695);
xnor_4 g09347(new_n11695, new_n11691, new_n11696);
or_5   g09348(new_n9762, new_n9744, new_n11697);
or_5   g09349(new_n9784, new_n9763_1, new_n11698);
and_5  g09350(new_n11698, new_n11697, new_n11699);
nand_5 g09351(new_n11699, new_n11696, new_n11700);
and_5  g09352(new_n11700, new_n11694, new_n11701);
xor_4  g09353(new_n11689, new_n11688, new_n11702);
nand_5 g09354(new_n11702, new_n11701, new_n11703);
and_5  g09355(new_n11703, new_n11690, new_n11704);
or_5   g09356(new_n11704, new_n11686, new_n11705);
nand_5 g09357(new_n11705, new_n11684, new_n11706);
nand_5 g09358(new_n11706, new_n11681, new_n11707);
and_5  g09359(new_n11707, new_n11679, new_n11708);
nor_5  g09360(new_n11708, new_n11676, new_n11709);
nor_5  g09361(new_n11709, new_n11674_1, new_n11710_1);
xor_4  g09362(new_n11710_1, new_n11671, new_n11711);
xnor_4 g09363(new_n11711, new_n11614, new_n11712_1);
not_10 g09364(new_n11712_1, new_n11713);
xor_4  g09365(new_n11708, new_n11676, new_n11714);
xor_4  g09366(new_n11611, new_n11600, new_n11715);
not_10 g09367(new_n11715, new_n11716);
and_5  g09368(new_n11716, new_n11714, new_n11717);
xor_4  g09369(new_n11716, new_n11714, new_n11718);
not_10 g09370(new_n11718, new_n11719);
xor_4  g09371(new_n11706, new_n11681, new_n11720);
not_10 g09372(new_n11720, new_n11721);
xor_4  g09373(new_n11609, new_n11602, new_n11722);
nor_5  g09374(new_n11722, new_n11721, new_n11723);
xor_4  g09375(new_n11722, new_n11721, new_n11724_1);
xor_4  g09376(new_n11704, new_n11686, new_n11725);
xor_4  g09377(n19652, n6218, new_n11726);
xnor_4 g09378(new_n11726, new_n11607_1, new_n11727);
and_5  g09379(new_n11727, new_n11725, new_n11728);
xor_4  g09380(new_n11726, new_n11607_1, new_n11729);
xnor_4 g09381(new_n11729, new_n11725, new_n11730);
not_10 g09382(new_n11730, new_n11731);
xor_4  g09383(new_n11702, new_n11701, new_n11732);
and_5  g09384(new_n11732, new_n11129, new_n11733);
not_10 g09385(new_n11733, new_n11734);
xnor_4 g09386(new_n11732, new_n11128, new_n11735);
not_10 g09387(new_n11133, new_n11736_1);
xor_4  g09388(new_n11699, new_n11696, new_n11737);
and_5  g09389(new_n11737, new_n11736_1, new_n11738);
nor_5  g09390(new_n11737, new_n11736_1, new_n11739);
nor_5  g09391(new_n9785, new_n9737, new_n11740);
and_5  g09392(new_n9809, new_n9786, new_n11741_1);
nor_5  g09393(new_n11741_1, new_n11740, new_n11742);
nor_5  g09394(new_n11742, new_n11739, new_n11743);
nor_5  g09395(new_n11743, new_n11738, new_n11744);
and_5  g09396(new_n11744, new_n11735, new_n11745);
not_10 g09397(new_n11745, new_n11746);
and_5  g09398(new_n11746, new_n11734, new_n11747);
nor_5  g09399(new_n11747, new_n11731, new_n11748);
nor_5  g09400(new_n11748, new_n11728, new_n11749_1);
not_10 g09401(new_n11749_1, new_n11750);
and_5  g09402(new_n11750, new_n11724_1, new_n11751);
nor_5  g09403(new_n11751, new_n11723, new_n11752);
nor_5  g09404(new_n11752, new_n11719, new_n11753);
nor_5  g09405(new_n11753, new_n11717, new_n11754);
xnor_4 g09406(new_n11754, new_n11713, n1684);
not_10 g09407(n3984, new_n11756);
xor_4  g09408(new_n6250, new_n11756, new_n11757);
or_5   g09409(new_n6254, n19652, new_n11758);
not_10 g09410(n19652, new_n11759);
xor_4  g09411(new_n6254, new_n11759, new_n11760);
or_5   g09412(new_n6257, n3366, new_n11761);
not_10 g09413(n3366, new_n11762);
xor_4  g09414(new_n6257, new_n11762, new_n11763);
or_5   g09415(new_n4018, n26565, new_n11764);
not_10 g09416(n26565, new_n11765);
xor_4  g09417(new_n4018, new_n11765, new_n11766);
or_5   g09418(new_n4020, n3959, new_n11767);
not_10 g09419(n3959, new_n11768);
xor_4  g09420(new_n4020, new_n11768, new_n11769);
or_5   g09421(new_n4022, n11566, new_n11770_1);
not_10 g09422(n11566, new_n11771_1);
xor_4  g09423(new_n4022, new_n11771_1, new_n11772);
or_5   g09424(new_n4026, n26744, new_n11773);
not_10 g09425(n26744, new_n11774);
xor_4  g09426(new_n4026, new_n11774, new_n11775_1);
or_5   g09427(new_n4030, n26625, new_n11776);
nand_5 g09428(n19922, n14230, new_n11777);
xor_4  g09429(new_n4030, n26625, new_n11778);
nand_5 g09430(new_n11778, new_n11777, new_n11779);
and_5  g09431(new_n11779, new_n11776, new_n11780);
or_5   g09432(new_n11780, new_n11775_1, new_n11781);
and_5  g09433(new_n11781, new_n11773, new_n11782);
or_5   g09434(new_n11782, new_n11772, new_n11783);
and_5  g09435(new_n11783, new_n11770_1, new_n11784);
or_5   g09436(new_n11784, new_n11769, new_n11785);
and_5  g09437(new_n11785, new_n11767, new_n11786);
or_5   g09438(new_n11786, new_n11766, new_n11787);
and_5  g09439(new_n11787, new_n11764, new_n11788);
or_5   g09440(new_n11788, new_n11763, new_n11789);
and_5  g09441(new_n11789, new_n11761, new_n11790);
or_5   g09442(new_n11790, new_n11760, new_n11791);
and_5  g09443(new_n11791, new_n11758, new_n11792);
xor_4  g09444(new_n11792, new_n11757, new_n11793);
or_5   g09445(new_n11793, n13026, new_n11794);
not_10 g09446(n13026, new_n11795);
xor_4  g09447(new_n11793, new_n11795, new_n11796);
xor_4  g09448(new_n11790, new_n11760, new_n11797);
or_5   g09449(new_n11797, n2175, new_n11798);
not_10 g09450(n2175, new_n11799);
xor_4  g09451(new_n11797, new_n11799, new_n11800);
xor_4  g09452(new_n11788, new_n11763, new_n11801);
or_5   g09453(new_n11801, n752, new_n11802);
xor_4  g09454(new_n11801, new_n11075, new_n11803);
xor_4  g09455(new_n11786, new_n11766, new_n11804);
or_5   g09456(new_n11804, n1611, new_n11805);
xor_4  g09457(new_n11784, new_n11769, new_n11806);
nor_5  g09458(new_n11806, n25094, new_n11807);
xor_4  g09459(new_n11806, new_n11077, new_n11808);
xor_4  g09460(new_n11782, new_n11772, new_n11809);
or_5   g09461(new_n11809, n21538, new_n11810);
xor_4  g09462(new_n11809, new_n11078_1, new_n11811);
xor_4  g09463(new_n11780, new_n11775_1, new_n11812);
or_5   g09464(new_n11812, n5131, new_n11813);
xor_4  g09465(new_n11778, new_n11777, new_n11814);
nor_5  g09466(new_n11814, n11473, new_n11815);
xor_4  g09467(n19922, n14230, new_n11816);
or_5   g09468(new_n11816, new_n11100, new_n11817);
xor_4  g09469(new_n11814, n11473, new_n11818_1);
and_5  g09470(new_n11818_1, new_n11817, new_n11819);
or_5   g09471(new_n11819, new_n11815, new_n11820);
xor_4  g09472(new_n11812, n5131, new_n11821);
nand_5 g09473(new_n11821, new_n11820, new_n11822);
and_5  g09474(new_n11822, new_n11813, new_n11823);
or_5   g09475(new_n11823, new_n11811, new_n11824);
and_5  g09476(new_n11824, new_n11810, new_n11825);
nor_5  g09477(new_n11825, new_n11808, new_n11826);
or_5   g09478(new_n11826, new_n11807, new_n11827);
xor_4  g09479(new_n11804, n1611, new_n11828);
nand_5 g09480(new_n11828, new_n11827, new_n11829);
and_5  g09481(new_n11829, new_n11805, new_n11830);
or_5   g09482(new_n11830, new_n11803, new_n11831);
and_5  g09483(new_n11831, new_n11802, new_n11832);
or_5   g09484(new_n11832, new_n11800, new_n11833);
and_5  g09485(new_n11833, new_n11798, new_n11834);
or_5   g09486(new_n11834, new_n11796, new_n11835);
and_5  g09487(new_n11835, new_n11794, new_n11836);
and_5  g09488(new_n11836, n23912, new_n11837_1);
not_10 g09489(n23912, new_n11838);
xor_4  g09490(new_n11836, new_n11838, new_n11839);
nor_5  g09491(new_n6250, n3984, new_n11840);
nor_5  g09492(new_n11792, new_n11757, new_n11841_1);
nor_5  g09493(new_n11841_1, new_n11840, new_n11842_1);
not_10 g09494(n4514, new_n11843_1);
nand_5 g09495(new_n6245_1, new_n11843_1, new_n11844);
or_5   g09496(new_n6245_1, new_n11843_1, new_n11845);
and_5  g09497(new_n11845, new_n11844, new_n11846);
xor_4  g09498(new_n11846, new_n11842_1, new_n11847);
nor_5  g09499(new_n11847, new_n11839, new_n11848);
or_5   g09500(new_n11848, new_n11837_1, new_n11849);
not_10 g09501(new_n6248_1, new_n11850);
nand_5 g09502(new_n11844, new_n11842_1, new_n11851);
and_5  g09503(new_n11851, new_n11850, new_n11852);
and_5  g09504(new_n11852, new_n11845, new_n11853);
or_5   g09505(new_n11853, new_n11849, new_n11854);
or_5   g09506(new_n4468, n15766, new_n11855);
xor_4  g09507(new_n4468, n15766, new_n11856);
not_10 g09508(new_n11856, new_n11857);
or_5   g09509(new_n4474, n25629, new_n11858);
xor_4  g09510(new_n4474, n25629, new_n11859);
not_10 g09511(new_n11859, new_n11860);
nand_5 g09512(new_n4479, new_n10524, new_n11861);
xor_4  g09513(new_n4479, new_n10524, new_n11862);
not_10 g09514(new_n11862, new_n11863);
nand_5 g09515(new_n4486, new_n10525_1, new_n11864);
xor_4  g09516(new_n4486, new_n10525_1, new_n11865);
not_10 g09517(new_n11865, new_n11866);
or_5   g09518(new_n3971_1, n13677, new_n11867);
nand_5 g09519(new_n3997, new_n3972, new_n11868);
and_5  g09520(new_n11868, new_n11867, new_n11869);
or_5   g09521(new_n11869, new_n11866, new_n11870);
and_5  g09522(new_n11870, new_n11864, new_n11871);
or_5   g09523(new_n11871, new_n11863, new_n11872);
and_5  g09524(new_n11872, new_n11861, new_n11873);
or_5   g09525(new_n11873, new_n11860, new_n11874);
and_5  g09526(new_n11874, new_n11858, new_n11875);
or_5   g09527(new_n11875, new_n11857, new_n11876);
and_5  g09528(new_n11876, new_n11855, new_n11877);
and_5  g09529(new_n11877, new_n4447, new_n11878);
xor_4  g09530(new_n11877, new_n4447, new_n11879);
xor_4  g09531(new_n11853, new_n11849, new_n11880);
nor_5  g09532(new_n11880, new_n11879, new_n11881);
xor_4  g09533(new_n11880, new_n11879, new_n11882);
not_10 g09534(new_n11882, new_n11883);
xor_4  g09535(new_n11875, new_n11857, new_n11884);
xor_4  g09536(new_n11847, new_n11839, new_n11885);
and_5  g09537(new_n11885, new_n11884, new_n11886);
xor_4  g09538(new_n11873, new_n11860, new_n11887);
not_10 g09539(new_n11887, new_n11888);
xor_4  g09540(new_n11834, new_n11796, new_n11889);
nor_5  g09541(new_n11889, new_n11888, new_n11890);
not_10 g09542(new_n11890, new_n11891);
xor_4  g09543(new_n11889, new_n11888, new_n11892);
not_10 g09544(new_n11892, new_n11893);
xnor_4 g09545(new_n11871, new_n11862, new_n11894);
not_10 g09546(new_n11894, new_n11895);
xor_4  g09547(new_n11832, new_n11800, new_n11896);
nor_5  g09548(new_n11896, new_n11895, new_n11897);
not_10 g09549(new_n11897, new_n11898_1);
xor_4  g09550(new_n11896, new_n11895, new_n11899);
not_10 g09551(new_n11899, new_n11900);
xor_4  g09552(new_n11869, new_n11866, new_n11901);
not_10 g09553(new_n11901, new_n11902);
xor_4  g09554(new_n11830, new_n11803, new_n11903);
nor_5  g09555(new_n11903, new_n11902, new_n11904);
not_10 g09556(new_n11904, new_n11905_1);
xor_4  g09557(new_n11903, new_n11902, new_n11906);
xor_4  g09558(new_n11828, new_n11827, new_n11907);
nor_5  g09559(new_n11907, new_n3999, new_n11908);
not_10 g09560(new_n11908, new_n11909);
xor_4  g09561(new_n11907, new_n3999, new_n11910);
xor_4  g09562(new_n11825, new_n11808, new_n11911);
nor_5  g09563(new_n11911, new_n4082, new_n11912);
xor_4  g09564(new_n11823, new_n11811, new_n11913);
nor_5  g09565(new_n11913, new_n4086, new_n11914);
xor_4  g09566(new_n11913, new_n4086, new_n11915);
not_10 g09567(new_n11915, new_n11916);
xor_4  g09568(new_n11821, new_n11820, new_n11917);
nor_5  g09569(new_n11917, new_n4090, new_n11918);
xor_4  g09570(new_n11818_1, new_n11817, new_n11919);
nor_5  g09571(new_n11919, new_n4096, new_n11920);
not_10 g09572(new_n2555_1, new_n11921);
xor_4  g09573(new_n11816, new_n11100, new_n11922);
nor_5  g09574(new_n11922, new_n11921, new_n11923);
xor_4  g09575(new_n11919, new_n4096, new_n11924);
not_10 g09576(new_n11924, new_n11925);
nor_5  g09577(new_n11925, new_n11923, new_n11926_1);
nor_5  g09578(new_n11926_1, new_n11920, new_n11927);
xor_4  g09579(new_n11917, new_n4090, new_n11928);
not_10 g09580(new_n11928, new_n11929);
nor_5  g09581(new_n11929, new_n11927, new_n11930);
nor_5  g09582(new_n11930, new_n11918, new_n11931);
nor_5  g09583(new_n11931, new_n11916, new_n11932);
nor_5  g09584(new_n11932, new_n11914, new_n11933);
xnor_4 g09585(new_n11911, new_n4079, new_n11934);
not_10 g09586(new_n11934, new_n11935);
nor_5  g09587(new_n11935, new_n11933, new_n11936);
nor_5  g09588(new_n11936, new_n11912, new_n11937);
not_10 g09589(new_n11937, new_n11938);
and_5  g09590(new_n11938, new_n11910, new_n11939);
not_10 g09591(new_n11939, new_n11940);
and_5  g09592(new_n11940, new_n11909, new_n11941);
not_10 g09593(new_n11941, new_n11942);
and_5  g09594(new_n11942, new_n11906, new_n11943);
not_10 g09595(new_n11943, new_n11944);
and_5  g09596(new_n11944, new_n11905_1, new_n11945);
nor_5  g09597(new_n11945, new_n11900, new_n11946);
not_10 g09598(new_n11946, new_n11947);
and_5  g09599(new_n11947, new_n11898_1, new_n11948);
nor_5  g09600(new_n11948, new_n11893, new_n11949);
not_10 g09601(new_n11949, new_n11950);
and_5  g09602(new_n11950, new_n11891, new_n11951);
xor_4  g09603(new_n11885, new_n11884, new_n11952);
not_10 g09604(new_n11952, new_n11953);
nor_5  g09605(new_n11953, new_n11951, new_n11954);
nor_5  g09606(new_n11954, new_n11886, new_n11955);
nor_5  g09607(new_n11955, new_n11883, new_n11956);
nor_5  g09608(new_n11956, new_n11881, new_n11957);
xor_4  g09609(new_n11957, new_n11878, new_n11958);
xor_4  g09610(new_n11958, new_n11854, n1701);
xnor_4 g09611(new_n3932_1, new_n3901, n1703);
xor_4  g09612(new_n4600, new_n4546, n1721);
not_10 g09613(new_n9199, new_n11962);
nor_5  g09614(new_n7829, new_n4349, new_n11963);
nor_5  g09615(new_n9139, new_n9138, new_n11964);
nor_5  g09616(new_n11964, new_n11963, new_n11965_1);
nor_5  g09617(new_n11965_1, new_n11962, new_n11966);
nor_5  g09618(new_n9199, new_n9140, new_n11967);
and_5  g09619(new_n9289, new_n9200, new_n11968);
nor_5  g09620(new_n11968, new_n11967, new_n11969);
or_5   g09621(new_n11969, new_n11966, new_n11970);
and_5  g09622(new_n11965_1, new_n11962, new_n11971);
or_5   g09623(new_n11971, new_n11968, new_n11972);
and_5  g09624(new_n11972, new_n11970, n1760);
xnor_4 g09625(new_n4102, new_n4094, n1791);
xor_4  g09626(new_n3368, new_n3367, n1808);
and_5  g09627(new_n7829, new_n7778, new_n11976);
nor_5  g09628(new_n7905, new_n7831, new_n11977);
nor_5  g09629(new_n11977, new_n11976, new_n11978);
not_10 g09630(n13494, new_n11979);
and_5  g09631(new_n11979, n4319, new_n11980_1);
xor_4  g09632(n13494, n4319, new_n11981);
not_10 g09633(n23463, new_n11982);
or_5   g09634(n25345, new_n11982, new_n11983);
or_5   g09635(new_n11424_1, new_n11399, new_n11984);
and_5  g09636(new_n11984, new_n11983, new_n11985);
nor_5  g09637(new_n11985, new_n11981, new_n11986);
nor_5  g09638(new_n11986, new_n11980_1, new_n11987);
and_5  g09639(new_n11987, new_n11978, new_n11988);
nor_5  g09640(new_n11987, new_n7907, new_n11989);
xor_4  g09641(new_n11987, new_n7907, new_n11990);
xor_4  g09642(new_n11985, new_n11981, new_n11991);
and_5  g09643(new_n11991, new_n7978, new_n11992);
xnor_4 g09644(new_n11991, new_n7978, new_n11993);
nand_5 g09645(new_n11425, new_n7985, new_n11994);
nand_5 g09646(new_n11454, new_n11426, new_n11995);
and_5  g09647(new_n11995, new_n11994, new_n11996);
nor_5  g09648(new_n11996, new_n11993, new_n11997);
nor_5  g09649(new_n11997, new_n11992, new_n11998);
and_5  g09650(new_n11998, new_n11990, new_n11999);
nor_5  g09651(new_n11999, new_n11989, new_n12000_1);
or_5   g09652(new_n12000_1, new_n11988, new_n12001);
nor_5  g09653(new_n11987, new_n11978, new_n12002);
or_5   g09654(new_n12002, new_n11999, new_n12003_1);
and_5  g09655(new_n12003_1, new_n12001, n1821);
xor_4  g09656(new_n6968, new_n6966, n1832);
xnor_4 g09657(n9934, n2272, new_n12006);
or_5   g09658(n25331, n18496, new_n12007);
xnor_4 g09659(n25331, n18496, new_n12008);
or_5   g09660(n26224, n18483, new_n12009);
xnor_4 g09661(n26224, n18483, new_n12010);
or_5   g09662(n21934, n19327, new_n12011_1);
xnor_4 g09663(n21934, n19327, new_n12012);
or_5   g09664(n22597, n18901, new_n12013);
xnor_4 g09665(n22597, n18901, new_n12014);
or_5   g09666(n26107, n4376, new_n12015);
xnor_4 g09667(n26107, n4376, new_n12016);
or_5   g09668(n14570, n342, new_n12017);
xnor_4 g09669(n14570, n342, new_n12018);
or_5   g09670(n26553, n23775, new_n12019);
xnor_4 g09671(n26553, n23775, new_n12020);
or_5   g09672(n8259, n4964, new_n12021);
and_5  g09673(n11479, n7876, new_n12022);
xnor_4 g09674(n8259, n4964, new_n12023);
or_5   g09675(new_n12023, new_n12022, new_n12024);
and_5  g09676(new_n12024, new_n12021, new_n12025);
or_5   g09677(new_n12025, new_n12020, new_n12026);
and_5  g09678(new_n12026, new_n12019, new_n12027);
or_5   g09679(new_n12027, new_n12018, new_n12028);
and_5  g09680(new_n12028, new_n12017, new_n12029);
or_5   g09681(new_n12029, new_n12016, new_n12030);
and_5  g09682(new_n12030, new_n12015, new_n12031);
or_5   g09683(new_n12031, new_n12014, new_n12032);
and_5  g09684(new_n12032, new_n12013, new_n12033);
or_5   g09685(new_n12033, new_n12012, new_n12034);
and_5  g09686(new_n12034, new_n12011_1, new_n12035);
or_5   g09687(new_n12035, new_n12010, new_n12036);
and_5  g09688(new_n12036, new_n12009, new_n12037);
or_5   g09689(new_n12037, new_n12008, new_n12038);
and_5  g09690(new_n12038, new_n12007, new_n12039);
xor_4  g09691(new_n12039, new_n12006, new_n12040);
xor_4  g09692(new_n12040, n2160, new_n12041);
not_10 g09693(new_n12041, new_n12042);
xor_4  g09694(new_n12037, new_n12008, new_n12043);
or_5   g09695(new_n12043, n10763, new_n12044);
xor_4  g09696(new_n12043, n10763, new_n12045);
xor_4  g09697(new_n12035, new_n12010, new_n12046);
nand_5 g09698(new_n12046, n7437, new_n12047);
xor_4  g09699(new_n12046, n7437, new_n12048);
not_10 g09700(new_n12048, new_n12049);
xor_4  g09701(new_n12033, new_n12012, new_n12050);
nand_5 g09702(new_n12050, n20700, new_n12051);
not_10 g09703(n20700, new_n12052);
xor_4  g09704(new_n12050, new_n12052, new_n12053);
xor_4  g09705(new_n12031, new_n12014, new_n12054);
nand_5 g09706(new_n12054, n7099, new_n12055);
not_10 g09707(n7099, new_n12056);
xor_4  g09708(new_n12054, new_n12056, new_n12057);
xor_4  g09709(new_n12029, new_n12016, new_n12058);
nand_5 g09710(new_n12058, n12811, new_n12059);
not_10 g09711(n12811, new_n12060);
xor_4  g09712(new_n12058, new_n12060, new_n12061);
xor_4  g09713(new_n12027, new_n12018, new_n12062);
nand_5 g09714(new_n12062, n1118, new_n12063);
not_10 g09715(n1118, new_n12064);
xor_4  g09716(new_n12062, new_n12064, new_n12065);
xor_4  g09717(new_n12025, new_n12020, new_n12066);
nand_5 g09718(new_n12066, n25974, new_n12067);
xor_4  g09719(new_n12066, n25974, new_n12068);
not_10 g09720(n1451, new_n12069);
xor_4  g09721(n11479, n7876, new_n12070);
nor_5  g09722(new_n12070, new_n12069, new_n12071);
or_5   g09723(new_n12071, n1630, new_n12072_1);
xnor_4 g09724(new_n12023, new_n12022, new_n12073);
xor_4  g09725(new_n12071, n1630, new_n12074);
nand_5 g09726(new_n12074, new_n12073, new_n12075);
and_5  g09727(new_n12075, new_n12072_1, new_n12076);
nand_5 g09728(new_n12076, new_n12068, new_n12077);
and_5  g09729(new_n12077, new_n12067, new_n12078);
or_5   g09730(new_n12078, new_n12065, new_n12079);
and_5  g09731(new_n12079, new_n12063, new_n12080);
or_5   g09732(new_n12080, new_n12061, new_n12081);
and_5  g09733(new_n12081, new_n12059, new_n12082);
or_5   g09734(new_n12082, new_n12057, new_n12083);
and_5  g09735(new_n12083, new_n12055, new_n12084);
or_5   g09736(new_n12084, new_n12053, new_n12085);
and_5  g09737(new_n12085, new_n12051, new_n12086);
or_5   g09738(new_n12086, new_n12049, new_n12087);
and_5  g09739(new_n12087, new_n12047, new_n12088);
nand_5 g09740(new_n12088, new_n12045, new_n12089);
and_5  g09741(new_n12089, new_n12044, new_n12090);
xor_4  g09742(new_n12090, new_n12042, new_n12091);
not_10 g09743(n21784, new_n12092);
not_10 g09744(n5521, new_n12093);
not_10 g09745(n11926, new_n12094);
and_5  g09746(new_n3850_1, new_n3841, new_n12095);
and_5  g09747(new_n12095, new_n12094, new_n12096);
and_5  g09748(new_n12096, new_n12093, new_n12097);
xor_4  g09749(new_n12097, new_n12092, new_n12098);
xor_4  g09750(new_n12098, new_n7313_1, new_n12099);
not_10 g09751(new_n12099, new_n12100);
xor_4  g09752(new_n12096, new_n12093, new_n12101);
or_5   g09753(new_n12101, new_n7317, new_n12102);
xor_4  g09754(new_n12101, new_n7317, new_n12103);
not_10 g09755(new_n12103, new_n12104);
xor_4  g09756(new_n12095, new_n12094, new_n12105);
or_5   g09757(new_n12105, new_n7322, new_n12106);
xor_4  g09758(new_n12105, new_n7322, new_n12107);
not_10 g09759(new_n12107, new_n12108);
or_5   g09760(new_n3851, new_n3839, new_n12109);
or_5   g09761(new_n3894, new_n3853, new_n12110);
and_5  g09762(new_n12110, new_n12109, new_n12111);
or_5   g09763(new_n12111, new_n12108, new_n12112);
and_5  g09764(new_n12112, new_n12106, new_n12113_1);
or_5   g09765(new_n12113_1, new_n12104, new_n12114);
and_5  g09766(new_n12114, new_n12102, new_n12115);
xor_4  g09767(new_n12115, new_n12100, new_n12116);
not_10 g09768(new_n12116, new_n12117);
xor_4  g09769(new_n12117, new_n12091, new_n12118);
xor_4  g09770(new_n12088, new_n12045, new_n12119);
xor_4  g09771(new_n12113_1, new_n12104, new_n12120);
not_10 g09772(new_n12120, new_n12121_1);
nor_5  g09773(new_n12121_1, new_n12119, new_n12122);
not_10 g09774(new_n12122, new_n12123);
xor_4  g09775(new_n12121_1, new_n12119, new_n12124);
xor_4  g09776(new_n12086, new_n12049, new_n12125);
not_10 g09777(new_n12125, new_n12126);
xor_4  g09778(new_n12111, new_n12108, new_n12127);
not_10 g09779(new_n12127, new_n12128);
nor_5  g09780(new_n12128, new_n12126, new_n12129);
not_10 g09781(new_n12129, new_n12130);
xor_4  g09782(new_n12128, new_n12126, new_n12131_1);
xor_4  g09783(new_n12084, new_n12053, new_n12132);
and_5  g09784(new_n12132, new_n3895, new_n12133);
not_10 g09785(new_n12133, new_n12134);
not_10 g09786(new_n3895, new_n12135);
xnor_4 g09787(new_n12132, new_n12135, new_n12136);
xor_4  g09788(new_n12082, new_n12057, new_n12137);
and_5  g09789(new_n12137, new_n3897, new_n12138);
not_10 g09790(new_n12138, new_n12139);
xnor_4 g09791(new_n12137, new_n3898, new_n12140);
xor_4  g09792(new_n12080, new_n12061, new_n12141);
and_5  g09793(new_n12141, new_n3902, new_n12142);
not_10 g09794(new_n12142, new_n12143);
xnor_4 g09795(new_n12141, new_n3903, new_n12144);
xor_4  g09796(new_n12078, new_n12065, new_n12145);
and_5  g09797(new_n12145, new_n3907, new_n12146_1);
not_10 g09798(new_n12146_1, new_n12147);
xnor_4 g09799(new_n12145, new_n3908, new_n12148);
xor_4  g09800(new_n12076, new_n12068, new_n12149);
and_5  g09801(new_n12149, new_n3912, new_n12150);
xnor_4 g09802(new_n12149, new_n3913, new_n12151);
xor_4  g09803(new_n12070, new_n12069, new_n12152_1);
not_10 g09804(new_n12152_1, new_n12153_1);
and_5  g09805(new_n12153_1, new_n3921, new_n12154);
xor_4  g09806(new_n12074, new_n12073, new_n12155);
and_5  g09807(new_n12155, new_n12154, new_n12156);
xor_4  g09808(new_n12155, new_n12154, new_n12157_1);
and_5  g09809(new_n12157_1, new_n3917, new_n12158_1);
nor_5  g09810(new_n12158_1, new_n12156, new_n12159);
and_5  g09811(new_n12159, new_n12151, new_n12160);
nor_5  g09812(new_n12160, new_n12150, new_n12161_1);
not_10 g09813(new_n12161_1, new_n12162);
and_5  g09814(new_n12162, new_n12148, new_n12163);
not_10 g09815(new_n12163, new_n12164);
and_5  g09816(new_n12164, new_n12147, new_n12165);
not_10 g09817(new_n12165, new_n12166);
and_5  g09818(new_n12166, new_n12144, new_n12167);
not_10 g09819(new_n12167, new_n12168);
and_5  g09820(new_n12168, new_n12143, new_n12169);
not_10 g09821(new_n12169, new_n12170);
and_5  g09822(new_n12170, new_n12140, new_n12171);
not_10 g09823(new_n12171, new_n12172);
and_5  g09824(new_n12172, new_n12139, new_n12173);
not_10 g09825(new_n12173, new_n12174);
and_5  g09826(new_n12174, new_n12136, new_n12175);
not_10 g09827(new_n12175, new_n12176);
and_5  g09828(new_n12176, new_n12134, new_n12177);
not_10 g09829(new_n12177, new_n12178);
and_5  g09830(new_n12178, new_n12131_1, new_n12179_1);
not_10 g09831(new_n12179_1, new_n12180);
and_5  g09832(new_n12180, new_n12130, new_n12181);
not_10 g09833(new_n12181, new_n12182);
and_5  g09834(new_n12182, new_n12124, new_n12183);
not_10 g09835(new_n12183, new_n12184);
and_5  g09836(new_n12184, new_n12123, new_n12185);
xor_4  g09837(new_n12185, new_n12118, n1859);
xnor_4 g09838(new_n5238, new_n5209, n1860);
and_5  g09839(new_n11657, new_n11652, new_n12188);
not_10 g09840(n10250, new_n12189);
nor_5  g09841(n21915, n15182, new_n12190);
nor_5  g09842(new_n6875, new_n6849, new_n12191);
nor_5  g09843(new_n12191, new_n12190, new_n12192_1);
xor_4  g09844(n25972, n8614, new_n12193);
xor_4  g09845(new_n12193, new_n12192_1, new_n12194);
not_10 g09846(new_n12194, new_n12195);
or_5   g09847(new_n12195, new_n12189, new_n12196);
xor_4  g09848(new_n12195, n10250, new_n12197);
nand_5 g09849(new_n6877, n7674, new_n12198);
not_10 g09850(n7674, new_n12199);
xor_4  g09851(new_n6877, new_n12199, new_n12200);
nand_5 g09852(new_n6880, n6397, new_n12201);
not_10 g09853(n6397, new_n12202);
xor_4  g09854(new_n6880, new_n12202, new_n12203);
nand_5 g09855(new_n6885, n19196, new_n12204);
not_10 g09856(n19196, new_n12205);
xor_4  g09857(new_n6885, new_n12205, new_n12206);
nand_5 g09858(new_n6890, n23586, new_n12207);
or_5   g09859(new_n6895, n21226, new_n12208);
xor_4  g09860(new_n6895, n21226, new_n12209_1);
not_10 g09861(n4426, new_n12210);
or_5   g09862(new_n6900, new_n12210, new_n12211);
xor_4  g09863(new_n6900, new_n12210, new_n12212);
nand_5 g09864(new_n4120, new_n8821_1, new_n12213);
or_5   g09865(new_n4131, new_n4122, new_n12214);
and_5  g09866(new_n4135, n9380, new_n12215);
xor_4  g09867(new_n4131, new_n4122, new_n12216);
nand_5 g09868(new_n12216, new_n12215, new_n12217);
and_5  g09869(new_n12217, new_n12214, new_n12218);
xor_4  g09870(new_n4120, new_n8821_1, new_n12219);
nand_5 g09871(new_n12219, new_n12218, new_n12220);
and_5  g09872(new_n12220, new_n12213, new_n12221);
nand_5 g09873(new_n12221, new_n12212, new_n12222);
and_5  g09874(new_n12222, new_n12211, new_n12223_1);
nand_5 g09875(new_n12223_1, new_n12209_1, new_n12224);
and_5  g09876(new_n12224, new_n12208, new_n12225_1);
xor_4  g09877(new_n6890, n23586, new_n12226);
nand_5 g09878(new_n12226, new_n12225_1, new_n12227);
and_5  g09879(new_n12227, new_n12207, new_n12228_1);
or_5   g09880(new_n12228_1, new_n12206, new_n12229);
and_5  g09881(new_n12229, new_n12204, new_n12230);
or_5   g09882(new_n12230, new_n12203, new_n12231);
and_5  g09883(new_n12231, new_n12201, new_n12232);
or_5   g09884(new_n12232, new_n12200, new_n12233);
and_5  g09885(new_n12233, new_n12198, new_n12234);
or_5   g09886(new_n12234, new_n12197, new_n12235_1);
and_5  g09887(new_n12235_1, new_n12196, new_n12236);
and_5  g09888(n25972, n8614, new_n12237);
not_10 g09889(new_n12192_1, new_n12238);
nor_5  g09890(n25972, n8614, new_n12239);
nor_5  g09891(new_n12239, new_n12238, new_n12240);
nor_5  g09892(new_n12240, new_n12237, new_n12241);
nor_5  g09893(new_n12241, new_n12236, new_n12242);
not_10 g09894(new_n12242, new_n12243);
and_5  g09895(new_n12243, new_n12188, new_n12244);
xnor_4 g09896(new_n12243, new_n12188, new_n12245);
not_10 g09897(new_n12241, new_n12246);
xor_4  g09898(new_n12246, new_n12236, new_n12247);
and_5  g09899(new_n12247, new_n11658, new_n12248);
xor_4  g09900(new_n12247, new_n11658, new_n12249);
not_10 g09901(new_n12249, new_n12250);
not_10 g09902(new_n11672, new_n12251);
xor_4  g09903(new_n12234, new_n12197, new_n12252);
nor_5  g09904(new_n12252, new_n12251, new_n12253);
xnor_4 g09905(new_n12252, new_n11672, new_n12254);
not_10 g09906(new_n12254, new_n12255);
xor_4  g09907(new_n12232, new_n12200, new_n12256);
nor_5  g09908(new_n12256, new_n11680, new_n12257);
not_10 g09909(new_n12257, new_n12258);
xor_4  g09910(new_n12256, new_n11680, new_n12259);
xor_4  g09911(new_n12230, new_n12203, new_n12260);
nor_5  g09912(new_n12260, new_n11682_1, new_n12261);
xor_4  g09913(new_n12260, new_n11682_1, new_n12262);
not_10 g09914(new_n12262, new_n12263);
xor_4  g09915(new_n12228_1, new_n12206, new_n12264);
nor_5  g09916(new_n12264, new_n11687, new_n12265);
not_10 g09917(new_n12265, new_n12266);
xnor_4 g09918(new_n12264, new_n11688, new_n12267);
xor_4  g09919(new_n12226, new_n12225_1, new_n12268);
nor_5  g09920(new_n12268, new_n11695, new_n12269);
xnor_4 g09921(new_n12268, new_n11693, new_n12270);
not_10 g09922(new_n12270, new_n12271);
xor_4  g09923(new_n12223_1, new_n12209_1, new_n12272);
and_5  g09924(new_n12272, new_n9762, new_n12273);
xor_4  g09925(new_n12272, new_n9762, new_n12274);
not_10 g09926(new_n12274, new_n12275);
not_10 g09927(new_n9764, new_n12276);
xor_4  g09928(new_n12221, new_n12212, new_n12277);
nor_5  g09929(new_n12277, new_n12276, new_n12278);
xnor_4 g09930(new_n12277, new_n9764, new_n12279);
not_10 g09931(new_n12279, new_n12280);
xor_4  g09932(new_n12219, new_n12218, new_n12281);
and_5  g09933(new_n12281, new_n9769, new_n12282);
xor_4  g09934(new_n12281, new_n9769, new_n12283);
not_10 g09935(new_n12283, new_n12284);
xor_4  g09936(new_n12216, new_n12215, new_n12285);
nor_5  g09937(new_n12285, new_n9773, new_n12286);
not_10 g09938(new_n12286, new_n12287);
xor_4  g09939(new_n4135, n9380, new_n12288);
nor_5  g09940(new_n12288, new_n7247, new_n12289);
xor_4  g09941(new_n12285, new_n9773, new_n12290);
and_5  g09942(new_n12290, new_n12289, new_n12291);
not_10 g09943(new_n12291, new_n12292);
and_5  g09944(new_n12292, new_n12287, new_n12293);
nor_5  g09945(new_n12293, new_n12284, new_n12294);
nor_5  g09946(new_n12294, new_n12282, new_n12295);
nor_5  g09947(new_n12295, new_n12280, new_n12296);
nor_5  g09948(new_n12296, new_n12278, new_n12297);
nor_5  g09949(new_n12297, new_n12275, new_n12298);
nor_5  g09950(new_n12298, new_n12273, new_n12299);
nor_5  g09951(new_n12299, new_n12271, new_n12300);
nor_5  g09952(new_n12300, new_n12269, new_n12301);
not_10 g09953(new_n12301, new_n12302_1);
and_5  g09954(new_n12302_1, new_n12267, new_n12303);
not_10 g09955(new_n12303, new_n12304_1);
and_5  g09956(new_n12304_1, new_n12266, new_n12305);
nor_5  g09957(new_n12305, new_n12263, new_n12306);
nor_5  g09958(new_n12306, new_n12261, new_n12307);
not_10 g09959(new_n12307, new_n12308);
and_5  g09960(new_n12308, new_n12259, new_n12309);
not_10 g09961(new_n12309, new_n12310);
and_5  g09962(new_n12310, new_n12258, new_n12311);
nor_5  g09963(new_n12311, new_n12255, new_n12312);
nor_5  g09964(new_n12312, new_n12253, new_n12313);
nor_5  g09965(new_n12313, new_n12250, new_n12314);
nor_5  g09966(new_n12314, new_n12248, new_n12315_1);
nor_5  g09967(new_n12315_1, new_n12245, new_n12316);
or_5   g09968(new_n12316, new_n12244, n1861);
nor_5  g09969(n13714, n12593, new_n12318);
and_5  g09970(new_n12318, new_n10286, new_n12319);
and_5  g09971(new_n12319, new_n10282, new_n12320);
and_5  g09972(new_n12320, new_n8921, new_n12321);
and_5  g09973(new_n12321, new_n8917, new_n12322);
xor_4  g09974(new_n12322, new_n8913, new_n12323);
xor_4  g09975(new_n12323, new_n5382, new_n12324_1);
xor_4  g09976(new_n12321, new_n8917, new_n12325_1);
or_5   g09977(new_n12325_1, new_n5418, new_n12326);
not_10 g09978(new_n5415, new_n12327);
xor_4  g09979(new_n12320, new_n8921, new_n12328);
nor_5  g09980(new_n12328, new_n12327, new_n12329_1);
xor_4  g09981(new_n12328, new_n12327, new_n12330_1);
xor_4  g09982(new_n12319, new_n10282, new_n12331);
or_5   g09983(new_n12331, new_n5390, new_n12332);
xor_4  g09984(new_n12318, new_n10286, new_n12333);
nor_5  g09985(new_n12333, new_n5406, new_n12334);
not_10 g09986(new_n12334, new_n12335);
xor_4  g09987(new_n12333, new_n5406, new_n12336);
nor_5  g09988(new_n5400_1, new_n10293, new_n12337);
xor_4  g09989(new_n12337, n12593, new_n12338);
nand_5 g09990(new_n12338, new_n5397, new_n12339);
nand_5 g09991(new_n5400_1, n13714, new_n12340);
or_5   g09992(new_n12340, n12593, new_n12341_1);
and_5  g09993(new_n12341_1, new_n12339, new_n12342);
and_5  g09994(new_n12342, new_n12336, new_n12343);
not_10 g09995(new_n12343, new_n12344);
and_5  g09996(new_n12344, new_n12335, new_n12345);
xnor_4 g09997(new_n12331, new_n5390, new_n12346_1);
or_5   g09998(new_n12346_1, new_n12345, new_n12347);
nand_5 g09999(new_n12347, new_n12332, new_n12348);
and_5  g10000(new_n12348, new_n12330_1, new_n12349_1);
or_5   g10001(new_n12349_1, new_n12329_1, new_n12350);
xor_4  g10002(new_n12325_1, new_n5418, new_n12351);
nand_5 g10003(new_n12351, new_n12350, new_n12352);
and_5  g10004(new_n12352, new_n12326, new_n12353);
xnor_4 g10005(new_n12353, new_n12324_1, new_n12354);
not_10 g10006(new_n12354, new_n12355);
and_5  g10007(new_n8732, new_n7525, new_n12356);
and_5  g10008(new_n12356, new_n7522, new_n12357);
xor_4  g10009(new_n12357, new_n7519, new_n12358);
xnor_4 g10010(new_n12358, new_n7326, new_n12359);
xor_4  g10011(new_n12356, new_n7522, new_n12360);
nand_5 g10012(new_n12360, new_n7330_1, new_n12361);
xor_4  g10013(new_n12360, new_n7330_1, new_n12362);
or_5   g10014(new_n8733, new_n7334, new_n12363);
xnor_4 g10015(new_n8733, new_n7334, new_n12364_1);
or_5   g10016(new_n8735, new_n7338, new_n12365);
not_10 g10017(new_n7338, new_n12366);
xnor_4 g10018(new_n8735, new_n12366, new_n12367);
nand_5 g10019(new_n8738, new_n7343, new_n12368);
or_5   g10020(new_n8738, new_n7343, new_n12369);
not_10 g10021(new_n7348, new_n12370);
nor_5  g10022(new_n8741, new_n12370, new_n12371);
nor_5  g10023(new_n7350, new_n7538, new_n12372);
not_10 g10024(new_n12372, new_n12373);
xor_4  g10025(new_n8741, new_n12370, new_n12374);
and_5  g10026(new_n12374, new_n12373, new_n12375);
nor_5  g10027(new_n12375, new_n12371, new_n12376);
nand_5 g10028(new_n12376, new_n12369, new_n12377);
and_5  g10029(new_n12377, new_n12368, new_n12378);
nand_5 g10030(new_n12378, new_n12367, new_n12379);
and_5  g10031(new_n12379, new_n12365, new_n12380_1);
or_5   g10032(new_n12380_1, new_n12364_1, new_n12381);
and_5  g10033(new_n12381, new_n12363, new_n12382);
nand_5 g10034(new_n12382, new_n12362, new_n12383_1);
and_5  g10035(new_n12383_1, new_n12361, new_n12384_1);
xor_4  g10036(new_n12384_1, new_n12359, new_n12385);
xor_4  g10037(new_n12385, new_n12355, new_n12386);
not_10 g10038(new_n12386, new_n12387);
xor_4  g10039(new_n12382, new_n12362, new_n12388);
not_10 g10040(new_n12388, new_n12389);
xor_4  g10041(new_n12351, new_n12350, new_n12390);
and_5  g10042(new_n12390, new_n12389, new_n12391);
xor_4  g10043(new_n12390, new_n12389, new_n12392);
xor_4  g10044(new_n12348, new_n12330_1, new_n12393);
xor_4  g10045(new_n12380_1, new_n12364_1, new_n12394);
and_5  g10046(new_n12394, new_n12393, new_n12395);
xor_4  g10047(new_n12394, new_n12393, new_n12396);
not_10 g10048(new_n12396, new_n12397_1);
xor_4  g10049(new_n12331, new_n5390, new_n12398_1);
xnor_4 g10050(new_n12398_1, new_n12345, new_n12399);
xor_4  g10051(new_n12378, new_n12367, new_n12400);
and_5  g10052(new_n12400, new_n12399, new_n12401);
xor_4  g10053(new_n12400, new_n12399, new_n12402);
not_10 g10054(new_n12402, new_n12403);
xor_4  g10055(new_n12342, new_n12336, new_n12404);
not_10 g10056(new_n12404, new_n12405);
xor_4  g10057(new_n8738, new_n7343, new_n12406);
xor_4  g10058(new_n12406, new_n12376, new_n12407);
nor_5  g10059(new_n12407, new_n12405, new_n12408_1);
xnor_4 g10060(new_n12407, new_n12404, new_n12409);
not_10 g10061(new_n12409, new_n12410);
xor_4  g10062(new_n12374, new_n12373, new_n12411);
xor_4  g10063(new_n12338, new_n5397, new_n12412);
not_10 g10064(new_n12412, new_n12413);
and_5  g10065(new_n12413, new_n12411, new_n12414);
xor_4  g10066(new_n7350, n18962, new_n12415);
xor_4  g10067(new_n5400_1, new_n10293, new_n12416);
nor_5  g10068(new_n12416, new_n12415, new_n12417);
not_10 g10069(new_n12417, new_n12418);
xor_4  g10070(new_n12413, new_n12411, new_n12419);
and_5  g10071(new_n12419, new_n12418, new_n12420);
nor_5  g10072(new_n12420, new_n12414, new_n12421);
nor_5  g10073(new_n12421, new_n12410, new_n12422);
nor_5  g10074(new_n12422, new_n12408_1, new_n12423);
nor_5  g10075(new_n12423, new_n12403, new_n12424);
nor_5  g10076(new_n12424, new_n12401, new_n12425);
nor_5  g10077(new_n12425, new_n12397_1, new_n12426);
nor_5  g10078(new_n12426, new_n12395, new_n12427);
not_10 g10079(new_n12427, new_n12428);
and_5  g10080(new_n12428, new_n12392, new_n12429);
nor_5  g10081(new_n12429, new_n12391, new_n12430);
xnor_4 g10082(new_n12430, new_n12387, n1891);
xor_4  g10083(n20169, n1949, new_n12432);
or_5   g10084(new_n4013, n8285, new_n12433);
or_5   g10085(n9323, new_n4003, new_n12434);
not_10 g10086(n6729, new_n12435);
and_5  g10087(n10792, new_n12435, new_n12436);
nor_5  g10088(n10792, new_n12435, new_n12437);
not_10 g10089(new_n12437, new_n12438);
not_10 g10090(n21687, new_n12439);
and_5  g10091(new_n12439, n19922, new_n12440);
and_5  g10092(new_n12440, new_n12438, new_n12441);
nor_5  g10093(new_n12441, new_n12436, new_n12442);
not_10 g10094(new_n12442, new_n12443);
nand_5 g10095(new_n12443, new_n12434, new_n12444);
and_5  g10096(new_n12444, new_n12433, new_n12445);
xor_4  g10097(new_n12445, new_n12432, new_n12446_1);
xor_4  g10098(new_n12446_1, new_n6605, new_n12447);
xnor_4 g10099(n9323, n8285, new_n12448);
xor_4  g10100(new_n12448, new_n12443, new_n12449_1);
and_5  g10101(new_n12449_1, new_n6607, new_n12450);
xor_4  g10102(new_n12449_1, new_n6607, new_n12451);
not_10 g10103(new_n12451, new_n12452);
xnor_4 g10104(n21687, n19922, new_n12453);
nor_5  g10105(new_n12453, new_n6612_1, new_n12454);
xnor_4 g10106(n10792, n6729, new_n12455);
xnor_4 g10107(new_n12455, new_n12440, new_n12456);
nor_5  g10108(new_n12456, new_n12454, new_n12457);
not_10 g10109(new_n12457, new_n12458);
xor_4  g10110(new_n12456, new_n12454, new_n12459);
and_5  g10111(new_n12459, new_n6616, new_n12460);
not_10 g10112(new_n12460, new_n12461_1);
and_5  g10113(new_n12461_1, new_n12458, new_n12462_1);
nor_5  g10114(new_n12462_1, new_n12452, new_n12463);
nor_5  g10115(new_n12463, new_n12450, new_n12464);
xor_4  g10116(new_n12464, new_n12447, n1925);
xor_4  g10117(new_n7710, new_n7674_1, n1942);
xnor_4 g10118(new_n6451, new_n6388, n1972);
not_10 g10119(new_n11218, new_n12468);
and_5  g10120(new_n8951, new_n8891, new_n12469_1);
not_10 g10121(new_n12469_1, new_n12470);
nor_5  g10122(new_n9018, new_n8952, new_n12471);
not_10 g10123(new_n12471, new_n12472);
and_5  g10124(new_n12472, new_n12470, new_n12473);
not_10 g10125(new_n11334, new_n12474);
nand_5 g10126(new_n8902, new_n8894, new_n12475);
nand_5 g10127(new_n8903, n12507, new_n12476);
nor_5  g10128(new_n8903, n12507, new_n12477);
or_5   g10129(new_n8950, new_n12477, new_n12478);
and_5  g10130(new_n12478, new_n12476, new_n12479);
and_5  g10131(new_n12479, new_n12475, new_n12480);
and_5  g10132(new_n12480, new_n12474, new_n12481);
and_5  g10133(new_n12481, new_n12473, new_n12482);
nor_5  g10134(new_n12480, new_n12474, new_n12483);
not_10 g10135(new_n12483, new_n12484);
nor_5  g10136(new_n12484, new_n12473, new_n12485);
nor_5  g10137(new_n12485, new_n12482, new_n12486);
nand_5 g10138(new_n12486, new_n12468, new_n12487);
xor_4  g10139(new_n12486, new_n12468, new_n12488);
xnor_4 g10140(new_n12480, new_n11334, new_n12489);
xor_4  g10141(new_n12489, new_n12473, new_n12490);
nor_5  g10142(new_n12490, new_n11218, new_n12491);
xor_4  g10143(new_n12490, new_n11218, new_n12492);
nor_5  g10144(new_n11261_1, new_n9019, new_n12493);
nor_5  g10145(new_n11267, new_n9022, new_n12494);
xor_4  g10146(new_n11267, new_n9022, new_n12495_1);
not_10 g10147(new_n12495_1, new_n12496);
and_5  g10148(new_n11273_1, new_n9028, new_n12497);
xnor_4 g10149(new_n11272, new_n9028, new_n12498);
not_10 g10150(new_n12498, new_n12499);
and_5  g10151(new_n11281, new_n9034, new_n12500);
xnor_4 g10152(new_n11278, new_n9034, new_n12501);
not_10 g10153(new_n12501, new_n12502);
and_5  g10154(new_n11287, new_n9040, new_n12503);
xnor_4 g10155(new_n11283, new_n9040, new_n12504);
not_10 g10156(new_n12504, new_n12505);
xnor_4 g10157(new_n11205, new_n11189, new_n12506);
and_5  g10158(new_n12506, new_n9046_1, new_n12507_1);
xnor_4 g10159(new_n11289, new_n9046_1, new_n12508);
not_10 g10160(new_n12508, new_n12509);
nor_5  g10161(new_n11291, new_n9051, new_n12510);
xor_4  g10162(new_n11291, new_n9051, new_n12511);
and_5  g10163(new_n11296, new_n9056, new_n12512);
xnor_4 g10164(new_n11296, new_n9055, new_n12513);
not_10 g10165(new_n12513, new_n12514);
nor_5  g10166(new_n11299, new_n9064, new_n12515_1);
not_10 g10167(new_n12515_1, new_n12516_1);
and_5  g10168(new_n12516_1, new_n11304, new_n12517);
xnor_4 g10169(new_n12515_1, new_n11304, new_n12518);
and_5  g10170(new_n12518, new_n9070, new_n12519);
nor_5  g10171(new_n12519, new_n12517, new_n12520);
nor_5  g10172(new_n12520, new_n12514, new_n12521);
nor_5  g10173(new_n12521, new_n12512, new_n12522);
not_10 g10174(new_n12522, new_n12523);
and_5  g10175(new_n12523, new_n12511, new_n12524);
nor_5  g10176(new_n12524, new_n12510, new_n12525);
nor_5  g10177(new_n12525, new_n12509, new_n12526);
nor_5  g10178(new_n12526, new_n12507_1, new_n12527);
nor_5  g10179(new_n12527, new_n12505, new_n12528);
nor_5  g10180(new_n12528, new_n12503, new_n12529);
nor_5  g10181(new_n12529, new_n12502, new_n12530);
nor_5  g10182(new_n12530, new_n12500, new_n12531);
nor_5  g10183(new_n12531, new_n12499, new_n12532);
nor_5  g10184(new_n12532, new_n12497, new_n12533);
nor_5  g10185(new_n12533, new_n12496, new_n12534);
nor_5  g10186(new_n12534, new_n12494, new_n12535);
xor_4  g10187(new_n11261_1, new_n9019, new_n12536);
not_10 g10188(new_n12536, new_n12537);
nor_5  g10189(new_n12537, new_n12535, new_n12538);
nor_5  g10190(new_n12538, new_n12493, new_n12539);
not_10 g10191(new_n12539, new_n12540_1);
and_5  g10192(new_n12540_1, new_n12492, new_n12541);
nor_5  g10193(new_n12541, new_n12491, new_n12542);
nand_5 g10194(new_n12542, new_n12488, new_n12543);
and_5  g10195(new_n12543, new_n12487, n1981);
xnor_4 g10196(new_n12537, new_n12535, n2004);
not_10 g10197(n6105, new_n12546_1);
and_5  g10198(new_n12546_1, n5140, new_n12547);
not_10 g10199(new_n12547, new_n12548);
xnor_4 g10200(n6105, n5140, new_n12549);
not_10 g10201(new_n12549, new_n12550);
not_10 g10202(n6204, new_n12551);
or_5   g10203(new_n12551, n3795, new_n12552_1);
xnor_4 g10204(n6204, n3795, new_n12553);
not_10 g10205(new_n12553, new_n12554);
not_10 g10206(n3349, new_n12555);
or_5   g10207(n25464, new_n12555, new_n12556);
xnor_4 g10208(n25464, n3349, new_n12557);
not_10 g10209(new_n12557, new_n12558);
or_5   g10210(n4590, new_n6499, new_n12559);
xnor_4 g10211(n4590, n1742, new_n12560);
not_10 g10212(new_n12560, new_n12561);
or_5   g10213(n26752, new_n6515, new_n12562_1);
xnor_4 g10214(n26752, n4858, new_n12563);
not_10 g10215(new_n12563, new_n12564);
or_5   g10216(new_n6520, n6513, new_n12565);
xnor_4 g10217(n8244, n6513, new_n12566_1);
not_10 g10218(new_n12566_1, new_n12567);
or_5   g10219(new_n6525, n3918, new_n12568);
xnor_4 g10220(n9493, n3918, new_n12569_1);
not_10 g10221(n919, new_n12570);
or_5   g10222(n15167, new_n12570, new_n12571);
or_5   g10223(new_n6529, n919, new_n12572);
not_10 g10224(n21095, new_n12573);
and_5  g10225(n25316, new_n12573, new_n12574);
nor_5  g10226(n25316, new_n12573, new_n12575);
not_10 g10227(new_n12575, new_n12576);
not_10 g10228(n8656, new_n12577);
and_5  g10229(n20385, new_n12577, new_n12578);
and_5  g10230(new_n12578, new_n12576, new_n12579);
nor_5  g10231(new_n12579, new_n12574, new_n12580);
not_10 g10232(new_n12580, new_n12581);
nand_5 g10233(new_n12581, new_n12572, new_n12582);
and_5  g10234(new_n12582, new_n12571, new_n12583);
nand_5 g10235(new_n12583, new_n12569_1, new_n12584);
and_5  g10236(new_n12584, new_n12568, new_n12585);
or_5   g10237(new_n12585, new_n12567, new_n12586);
and_5  g10238(new_n12586, new_n12565, new_n12587_1);
or_5   g10239(new_n12587_1, new_n12564, new_n12588);
and_5  g10240(new_n12588, new_n12562_1, new_n12589);
or_5   g10241(new_n12589, new_n12561, new_n12590);
and_5  g10242(new_n12590, new_n12559, new_n12591);
or_5   g10243(new_n12591, new_n12558, new_n12592);
and_5  g10244(new_n12592, new_n12556, new_n12593_1);
or_5   g10245(new_n12593_1, new_n12554, new_n12594);
and_5  g10246(new_n12594, new_n12552_1, new_n12595);
nor_5  g10247(new_n12595, new_n12550, new_n12596);
not_10 g10248(new_n12596, new_n12597);
and_5  g10249(new_n12597, new_n12548, new_n12598);
or_5   g10250(new_n6245_1, n10018, new_n12599);
and_5  g10251(new_n6245_1, n10018, new_n12600);
not_10 g10252(n2184, new_n12601);
and_5  g10253(new_n6250, new_n12601, new_n12602);
xor_4  g10254(new_n6250, n2184, new_n12603);
not_10 g10255(n3541, new_n12604);
nand_5 g10256(new_n6254, new_n12604, new_n12605);
xor_4  g10257(new_n6254, n3541, new_n12606);
nand_5 g10258(new_n6257, new_n6500, new_n12607_1);
xor_4  g10259(new_n6257, n16818, new_n12608);
nand_5 g10260(new_n4018, new_n6501, new_n12609);
xor_4  g10261(new_n4018, n1269, new_n12610);
nand_5 g10262(new_n4020, new_n6502_1, new_n12611);
xor_4  g10263(new_n4020, new_n6502_1, new_n12612);
or_5   g10264(new_n4022, new_n6503, new_n12613);
xor_4  g10265(new_n4022, new_n6503, new_n12614);
nand_5 g10266(new_n4026, new_n6504, new_n12615);
not_10 g10267(n15652, new_n12616);
or_5   g10268(new_n4030, new_n12616, new_n12617);
not_10 g10269(n4939, new_n12618);
nor_5  g10270(n19922, new_n12618, new_n12619);
xor_4  g10271(new_n4030, new_n12616, new_n12620_1);
nand_5 g10272(new_n12620_1, new_n12619, new_n12621_1);
and_5  g10273(new_n12621_1, new_n12617, new_n12622);
xor_4  g10274(new_n4026, new_n6504, new_n12623);
nand_5 g10275(new_n12623, new_n12622, new_n12624);
and_5  g10276(new_n12624, new_n12615, new_n12625);
nand_5 g10277(new_n12625, new_n12614, new_n12626_1);
and_5  g10278(new_n12626_1, new_n12613, new_n12627);
nand_5 g10279(new_n12627, new_n12612, new_n12628);
and_5  g10280(new_n12628, new_n12611, new_n12629);
or_5   g10281(new_n12629, new_n12610, new_n12630);
and_5  g10282(new_n12630, new_n12609, new_n12631);
or_5   g10283(new_n12631, new_n12608, new_n12632);
and_5  g10284(new_n12632, new_n12607_1, new_n12633);
or_5   g10285(new_n12633, new_n12606, new_n12634);
and_5  g10286(new_n12634, new_n12605, new_n12635);
nor_5  g10287(new_n12635, new_n12603, new_n12636);
nor_5  g10288(new_n12636, new_n12602, new_n12637);
nor_5  g10289(new_n12637, new_n12600, new_n12638);
xor_4  g10290(new_n12638, new_n11850, new_n12639);
and_5  g10291(new_n12639, new_n12599, new_n12640);
xor_4  g10292(new_n12640, new_n6235, new_n12641);
xor_4  g10293(new_n6245_1, n10018, new_n12642);
xor_4  g10294(new_n12642, new_n12637, new_n12643);
and_5  g10295(new_n12643, new_n6277, new_n12644);
xnor_4 g10296(new_n12643, new_n6277, new_n12645);
xor_4  g10297(new_n12635, new_n12603, new_n12646);
or_5   g10298(new_n12646, new_n6285, new_n12647);
xor_4  g10299(new_n12646, new_n6284, new_n12648);
xor_4  g10300(new_n12633, new_n12606, new_n12649);
or_5   g10301(new_n12649, new_n6292, new_n12650_1);
xor_4  g10302(new_n12649, new_n6291, new_n12651);
xor_4  g10303(new_n12631, new_n12608, new_n12652);
or_5   g10304(new_n12652, new_n6296, new_n12653);
xor_4  g10305(new_n12629, new_n12610, new_n12654_1);
nor_5  g10306(new_n12654_1, new_n6300, new_n12655);
xor_4  g10307(new_n12654_1, new_n6299, new_n12656);
xor_4  g10308(new_n12627, new_n12612, new_n12657_1);
or_5   g10309(new_n12657_1, new_n6305, new_n12658);
xor_4  g10310(new_n12657_1, new_n6304, new_n12659);
xor_4  g10311(new_n12625, new_n12614, new_n12660);
nand_5 g10312(new_n12660, new_n6306, new_n12661);
xor_4  g10313(new_n12623, new_n12622, new_n12662);
nand_5 g10314(new_n12662, new_n6309, new_n12663);
xnor_4 g10315(new_n12662, new_n6308_1, new_n12664);
not_10 g10316(new_n12664, new_n12665_1);
xor_4  g10317(new_n12620_1, new_n12619, new_n12666);
or_5   g10318(new_n12666, new_n6312, new_n12667);
xor_4  g10319(n19922, n4939, new_n12668);
and_5  g10320(new_n12668, new_n6314, new_n12669);
xor_4  g10321(new_n12666, new_n6312, new_n12670_1);
nand_5 g10322(new_n12670_1, new_n12669, new_n12671);
and_5  g10323(new_n12671, new_n12667, new_n12672);
or_5   g10324(new_n12672, new_n12665_1, new_n12673);
and_5  g10325(new_n12673, new_n12663, new_n12674);
xor_4  g10326(new_n12660, new_n6306, new_n12675);
nand_5 g10327(new_n12675, new_n12674, new_n12676);
and_5  g10328(new_n12676, new_n12661, new_n12677);
or_5   g10329(new_n12677, new_n12659, new_n12678);
and_5  g10330(new_n12678, new_n12658, new_n12679);
nor_5  g10331(new_n12679, new_n12656, new_n12680);
or_5   g10332(new_n12680, new_n12655, new_n12681);
xnor_4 g10333(new_n12652, new_n6295, new_n12682);
nand_5 g10334(new_n12682, new_n12681, new_n12683);
and_5  g10335(new_n12683, new_n12653, new_n12684);
or_5   g10336(new_n12684, new_n12651, new_n12685);
and_5  g10337(new_n12685, new_n12650_1, new_n12686);
or_5   g10338(new_n12686, new_n12648, new_n12687);
and_5  g10339(new_n12687, new_n12647, new_n12688);
nor_5  g10340(new_n12688, new_n12645, new_n12689);
nor_5  g10341(new_n12689, new_n12644, new_n12690);
xor_4  g10342(new_n12690, new_n12641, new_n12691);
nor_5  g10343(new_n12691, new_n12598, new_n12692);
xor_4  g10344(new_n12691, new_n12598, new_n12693);
not_10 g10345(new_n12693, new_n12694);
xor_4  g10346(new_n12595, new_n12550, new_n12695);
not_10 g10347(new_n12695, new_n12696);
xor_4  g10348(new_n12688, new_n12645, new_n12697);
and_5  g10349(new_n12697, new_n12696, new_n12698);
xnor_4 g10350(new_n12697, new_n12695, new_n12699);
not_10 g10351(new_n12699, new_n12700);
xor_4  g10352(new_n12593_1, new_n12554, new_n12701);
not_10 g10353(new_n12701, new_n12702_1);
xor_4  g10354(new_n12686, new_n12648, new_n12703);
and_5  g10355(new_n12703, new_n12702_1, new_n12704);
xnor_4 g10356(new_n12703, new_n12701, new_n12705);
not_10 g10357(new_n12705, new_n12706);
xor_4  g10358(new_n12591, new_n12558, new_n12707_1);
not_10 g10359(new_n12707_1, new_n12708);
xor_4  g10360(new_n12684, new_n12651, new_n12709);
nand_5 g10361(new_n12709, new_n12708, new_n12710);
xnor_4 g10362(new_n12709, new_n12707_1, new_n12711);
not_10 g10363(new_n12711, new_n12712);
xor_4  g10364(new_n12589, new_n12561, new_n12713);
not_10 g10365(new_n12713, new_n12714);
xor_4  g10366(new_n12682, new_n12681, new_n12715);
nand_5 g10367(new_n12715, new_n12714, new_n12716);
xnor_4 g10368(new_n12715, new_n12713, new_n12717);
not_10 g10369(new_n12717, new_n12718);
xor_4  g10370(new_n12587_1, new_n12564, new_n12719);
not_10 g10371(new_n12719, new_n12720);
xor_4  g10372(new_n12679, new_n12656, new_n12721);
nand_5 g10373(new_n12721, new_n12720, new_n12722);
xnor_4 g10374(new_n12721, new_n12719, new_n12723);
not_10 g10375(new_n12723, new_n12724);
xor_4  g10376(new_n12585, new_n12567, new_n12725_1);
not_10 g10377(new_n12725_1, new_n12726);
xor_4  g10378(new_n12677, new_n12659, new_n12727_1);
nand_5 g10379(new_n12727_1, new_n12726, new_n12728);
xnor_4 g10380(new_n12727_1, new_n12725_1, new_n12729);
not_10 g10381(new_n12729, new_n12730);
xor_4  g10382(new_n12583, new_n12569_1, new_n12731);
not_10 g10383(new_n12731, new_n12732);
xor_4  g10384(new_n12675, new_n12674, new_n12733);
nand_5 g10385(new_n12733, new_n12732, new_n12734);
xnor_4 g10386(new_n12733, new_n12731, new_n12735);
not_10 g10387(new_n12735, new_n12736);
xor_4  g10388(new_n12672, new_n12665_1, new_n12737);
xnor_4 g10389(n15167, n919, new_n12738);
xnor_4 g10390(new_n12738, new_n12581, new_n12739);
or_5   g10391(new_n12739, new_n12737, new_n12740_1);
xor_4  g10392(new_n12738, new_n12581, new_n12741);
xnor_4 g10393(new_n12741, new_n12737, new_n12742_1);
not_10 g10394(new_n12742_1, new_n12743);
xnor_4 g10395(new_n12668, new_n6314, new_n12744);
xnor_4 g10396(n20385, n8656, new_n12745);
nor_5  g10397(new_n12745, new_n12744, new_n12746_1);
not_10 g10398(new_n12746_1, new_n12747);
xnor_4 g10399(n25316, n21095, new_n12748);
xor_4  g10400(new_n12748, new_n12578, new_n12749);
nand_5 g10401(new_n12749, new_n12747, new_n12750);
xor_4  g10402(new_n12670_1, new_n12669, new_n12751);
xor_4  g10403(new_n12749, new_n12747, new_n12752);
not_10 g10404(new_n12752, new_n12753);
or_5   g10405(new_n12753, new_n12751, new_n12754);
and_5  g10406(new_n12754, new_n12750, new_n12755);
or_5   g10407(new_n12755, new_n12743, new_n12756_1);
and_5  g10408(new_n12756_1, new_n12740_1, new_n12757);
or_5   g10409(new_n12757, new_n12736, new_n12758);
and_5  g10410(new_n12758, new_n12734, new_n12759);
or_5   g10411(new_n12759, new_n12730, new_n12760);
and_5  g10412(new_n12760, new_n12728, new_n12761);
or_5   g10413(new_n12761, new_n12724, new_n12762);
and_5  g10414(new_n12762, new_n12722, new_n12763);
or_5   g10415(new_n12763, new_n12718, new_n12764);
and_5  g10416(new_n12764, new_n12716, new_n12765);
or_5   g10417(new_n12765, new_n12712, new_n12766);
and_5  g10418(new_n12766, new_n12710, new_n12767);
nor_5  g10419(new_n12767, new_n12706, new_n12768);
nor_5  g10420(new_n12768, new_n12704, new_n12769);
nor_5  g10421(new_n12769, new_n12700, new_n12770);
nor_5  g10422(new_n12770, new_n12698, new_n12771);
nor_5  g10423(new_n12771, new_n12694, new_n12772);
nor_5  g10424(new_n12772, new_n12692, new_n12773);
or_5   g10425(new_n12640, new_n6235, new_n12774);
nand_5 g10426(new_n12638, new_n6248_1, new_n12775);
nand_5 g10427(new_n12640, new_n6235, new_n12776);
nand_5 g10428(new_n12690, new_n12776, new_n12777);
and_5  g10429(new_n12777, new_n12775, new_n12778);
nand_5 g10430(new_n12778, new_n12774, new_n12779);
nor_5  g10431(new_n12779, new_n12773, n2007);
xnor_4 g10432(new_n9073, new_n9061, n2061);
xnor_4 g10433(new_n11523, new_n7154, new_n12782);
not_10 g10434(new_n12782, new_n12783_1);
not_10 g10435(new_n11529, new_n12784);
and_5  g10436(new_n12784, new_n7160, new_n12785);
xnor_4 g10437(new_n11529, new_n7160, new_n12786);
not_10 g10438(new_n12786, new_n12787);
nor_5  g10439(new_n11533, new_n7166, new_n12788);
and_5  g10440(new_n7171, new_n4668, new_n12789);
xor_4  g10441(new_n7171, new_n4668, new_n12790);
not_10 g10442(new_n12790, new_n12791);
and_5  g10443(new_n7177, new_n4698, new_n12792);
xor_4  g10444(new_n7177, new_n4698, new_n12793);
not_10 g10445(new_n12793, new_n12794);
nor_5  g10446(new_n7182, new_n4703, new_n12795);
not_10 g10447(new_n12795, new_n12796);
and_5  g10448(new_n7186, new_n4709, new_n12797);
not_10 g10449(new_n12797, new_n12798);
xor_4  g10450(new_n7186, new_n4709, new_n12799);
or_5   g10451(new_n7192, new_n4719, new_n12800);
nor_5  g10452(new_n12800, new_n4715, new_n12801_1);
xor_4  g10453(new_n12800, new_n4715, new_n12802);
and_5  g10454(new_n12802, new_n7198, new_n12803);
nor_5  g10455(new_n12803, new_n12801_1, new_n12804);
and_5  g10456(new_n12804, new_n12799, new_n12805);
not_10 g10457(new_n12805, new_n12806);
and_5  g10458(new_n12806, new_n12798, new_n12807);
not_10 g10459(new_n12807, new_n12808);
xor_4  g10460(new_n7182, new_n4703, new_n12809);
and_5  g10461(new_n12809, new_n12808, new_n12810);
not_10 g10462(new_n12810, new_n12811_1);
and_5  g10463(new_n12811_1, new_n12796, new_n12812_1);
nor_5  g10464(new_n12812_1, new_n12794, new_n12813);
nor_5  g10465(new_n12813, new_n12792, new_n12814);
nor_5  g10466(new_n12814, new_n12791, new_n12815);
nor_5  g10467(new_n12815, new_n12789, new_n12816_1);
not_10 g10468(new_n12816_1, new_n12817);
xor_4  g10469(new_n11533, new_n7166, new_n12818);
and_5  g10470(new_n12818, new_n12817, new_n12819);
nor_5  g10471(new_n12819, new_n12788, new_n12820);
nor_5  g10472(new_n12820, new_n12787, new_n12821_1);
nor_5  g10473(new_n12821_1, new_n12785, new_n12822);
xnor_4 g10474(new_n12822, new_n12783_1, n2092);
xnor_4 g10475(n22253, n10650, new_n12824);
or_5   g10476(n12900, n1255, new_n12825);
xnor_4 g10477(n12900, n1255, new_n12826);
or_5   g10478(n20411, n9512, new_n12827);
xnor_4 g10479(n20411, n9512, new_n12828);
or_5   g10480(n17069, n16608, new_n12829);
xnor_4 g10481(n17069, n16608, new_n12830);
or_5   g10482(n21735, n15918, new_n12831);
xnor_4 g10483(n21735, n15918, new_n12832);
or_5   g10484(n24085, n17784, new_n12833);
xnor_4 g10485(n24085, n17784, new_n12834);
or_5   g10486(n14323, n14071, new_n12835);
xnor_4 g10487(n14323, n14071, new_n12836);
or_5   g10488(n2886, n1738, new_n12837);
xnor_4 g10489(n2886, n1738, new_n12838);
or_5   g10490(n12152, n1040, new_n12839);
and_5  g10491(n19107, n9090, new_n12840);
xnor_4 g10492(n12152, n1040, new_n12841);
or_5   g10493(new_n12841, new_n12840, new_n12842);
and_5  g10494(new_n12842, new_n12839, new_n12843_1);
or_5   g10495(new_n12843_1, new_n12838, new_n12844);
and_5  g10496(new_n12844, new_n12837, new_n12845);
or_5   g10497(new_n12845, new_n12836, new_n12846);
and_5  g10498(new_n12846, new_n12835, new_n12847);
or_5   g10499(new_n12847, new_n12834, new_n12848);
and_5  g10500(new_n12848, new_n12833, new_n12849);
or_5   g10501(new_n12849, new_n12832, new_n12850);
and_5  g10502(new_n12850, new_n12831, new_n12851);
or_5   g10503(new_n12851, new_n12830, new_n12852);
and_5  g10504(new_n12852, new_n12829, new_n12853);
or_5   g10505(new_n12853, new_n12828, new_n12854);
and_5  g10506(new_n12854, new_n12827, new_n12855);
or_5   g10507(new_n12855, new_n12826, new_n12856);
and_5  g10508(new_n12856, new_n12825, new_n12857);
xor_4  g10509(new_n12857, new_n12824, new_n12858);
and_5  g10510(new_n12858, n2272, new_n12859);
xor_4  g10511(new_n12858, n2272, new_n12860);
not_10 g10512(new_n12860, new_n12861_1);
xor_4  g10513(new_n12855, new_n12826, new_n12862);
nand_5 g10514(new_n12862, n25331, new_n12863);
xor_4  g10515(new_n12862, n25331, new_n12864_1);
not_10 g10516(new_n12864_1, new_n12865_1);
xor_4  g10517(new_n12853, new_n12828, new_n12866);
nand_5 g10518(new_n12866, n18483, new_n12867);
xor_4  g10519(new_n12866, n18483, new_n12868);
not_10 g10520(new_n12868, new_n12869);
xor_4  g10521(new_n12851, new_n12830, new_n12870_1);
nand_5 g10522(new_n12870_1, n21934, new_n12871_1);
xor_4  g10523(new_n12870_1, n21934, new_n12872);
not_10 g10524(new_n12872, new_n12873_1);
xor_4  g10525(new_n12849, new_n12832, new_n12874);
nand_5 g10526(new_n12874, n18901, new_n12875_1);
xor_4  g10527(new_n12874, n18901, new_n12876);
not_10 g10528(new_n12876, new_n12877);
xor_4  g10529(new_n12847, new_n12834, new_n12878);
nand_5 g10530(new_n12878, n4376, new_n12879);
xor_4  g10531(new_n12878, n4376, new_n12880);
not_10 g10532(new_n12880, new_n12881);
xor_4  g10533(new_n12845, new_n12836, new_n12882);
nand_5 g10534(new_n12882, n14570, new_n12883);
xor_4  g10535(new_n12882, n14570, new_n12884);
not_10 g10536(new_n12884, new_n12885);
xor_4  g10537(new_n12843_1, new_n12838, new_n12886);
nand_5 g10538(new_n12886, n23775, new_n12887);
xor_4  g10539(new_n12886, n23775, new_n12888);
xor_4  g10540(n19107, n9090, new_n12889);
nor_5  g10541(new_n12889, new_n7022, new_n12890);
or_5   g10542(new_n12890, n8259, new_n12891);
xnor_4 g10543(new_n12841, new_n12840, new_n12892_1);
xor_4  g10544(new_n12890, n8259, new_n12893);
nand_5 g10545(new_n12893, new_n12892_1, new_n12894);
and_5  g10546(new_n12894, new_n12891, new_n12895);
nand_5 g10547(new_n12895, new_n12888, new_n12896);
and_5  g10548(new_n12896, new_n12887, new_n12897);
or_5   g10549(new_n12897, new_n12885, new_n12898);
and_5  g10550(new_n12898, new_n12883, new_n12899);
or_5   g10551(new_n12899, new_n12881, new_n12900_1);
and_5  g10552(new_n12900_1, new_n12879, new_n12901);
or_5   g10553(new_n12901, new_n12877, new_n12902);
and_5  g10554(new_n12902, new_n12875_1, new_n12903);
or_5   g10555(new_n12903, new_n12873_1, new_n12904_1);
and_5  g10556(new_n12904_1, new_n12871_1, new_n12905);
or_5   g10557(new_n12905, new_n12869, new_n12906);
and_5  g10558(new_n12906, new_n12867, new_n12907);
or_5   g10559(new_n12907, new_n12865_1, new_n12908);
and_5  g10560(new_n12908, new_n12863, new_n12909);
nor_5  g10561(new_n12909, new_n12861_1, new_n12910);
nor_5  g10562(new_n12910, new_n12859, new_n12911);
or_5   g10563(n22253, n10650, new_n12912);
or_5   g10564(new_n12857, new_n12824, new_n12913);
and_5  g10565(new_n12913, new_n12912, new_n12914);
nor_5  g10566(new_n12914, new_n12911, new_n12915);
not_10 g10567(n9934, new_n12916);
not_10 g10568(n18496, new_n12917_1);
not_10 g10569(n26224, new_n12918);
not_10 g10570(n26107, new_n12919);
not_10 g10571(n342, new_n12920);
not_10 g10572(n26553, new_n12921);
nor_5  g10573(n7876, n4964, new_n12922);
and_5  g10574(new_n12922, new_n12921, new_n12923);
and_5  g10575(new_n12923, new_n12920, new_n12924);
and_5  g10576(new_n12924, new_n12919, new_n12925);
and_5  g10577(new_n12925, new_n3739, new_n12926);
and_5  g10578(new_n12926, new_n3724, new_n12927);
and_5  g10579(new_n12927, new_n12918, new_n12928);
and_5  g10580(new_n12928, new_n12917_1, new_n12929);
and_5  g10581(new_n12929, new_n12916, new_n12930);
not_10 g10582(new_n12930, new_n12931);
xor_4  g10583(new_n12929, new_n12916, new_n12932);
nor_5  g10584(n18409, n5704, new_n12933);
and_5  g10585(new_n12933, new_n3819, new_n12934);
and_5  g10586(new_n12934, new_n3814, new_n12935);
and_5  g10587(new_n12935, new_n3810, new_n12936);
and_5  g10588(new_n12936, new_n3806, new_n12937);
and_5  g10589(new_n12937, new_n7005, new_n12938);
and_5  g10590(new_n12938, new_n7001, new_n12939);
xor_4  g10591(new_n12939, new_n6997, new_n12940);
nor_5  g10592(new_n12940, n12861, new_n12941_1);
xor_4  g10593(new_n12940, n12861, new_n12942_1);
not_10 g10594(new_n12942_1, new_n12943);
xor_4  g10595(new_n12938, new_n7001, new_n12944);
or_5   g10596(new_n12944, n13333, new_n12945);
xnor_4 g10597(new_n12944, n13333, new_n12946);
xor_4  g10598(new_n12937, new_n7005, new_n12947);
or_5   g10599(new_n12947, n2210, new_n12948);
xor_4  g10600(new_n12947, n2210, new_n12949);
not_10 g10601(new_n12949, new_n12950);
xor_4  g10602(new_n12936, new_n3806, new_n12951);
or_5   g10603(new_n12951, n20604, new_n12952);
not_10 g10604(n20604, new_n12953);
xor_4  g10605(new_n12951, new_n12953, new_n12954);
xor_4  g10606(new_n12935, new_n3810, new_n12955);
or_5   g10607(new_n12955, n16158, new_n12956_1);
xor_4  g10608(new_n12955, new_n4613, new_n12957);
xor_4  g10609(new_n12934, new_n3814, new_n12958);
or_5   g10610(new_n12958, n5752, new_n12959);
xor_4  g10611(new_n12933, new_n3819, new_n12960);
nor_5  g10612(new_n12960, n18171, new_n12961);
xor_4  g10613(new_n12960, n18171, new_n12962);
not_10 g10614(new_n12962, new_n12963);
xor_4  g10615(n18409, n5704, new_n12964);
or_5   g10616(new_n12964, n25073, new_n12965);
nand_5 g10617(n22309, n5704, new_n12966);
xor_4  g10618(new_n12964, n25073, new_n12967);
nand_5 g10619(new_n12967, new_n12966, new_n12968);
and_5  g10620(new_n12968, new_n12965, new_n12969);
nor_5  g10621(new_n12969, new_n12963, new_n12970);
or_5   g10622(new_n12970, new_n12961, new_n12971);
xor_4  g10623(new_n12958, n5752, new_n12972);
nand_5 g10624(new_n12972, new_n12971, new_n12973);
and_5  g10625(new_n12973, new_n12959, new_n12974);
or_5   g10626(new_n12974, new_n12957, new_n12975);
and_5  g10627(new_n12975, new_n12956_1, new_n12976);
or_5   g10628(new_n12976, new_n12954, new_n12977);
and_5  g10629(new_n12977, new_n12952, new_n12978_1);
or_5   g10630(new_n12978_1, new_n12950, new_n12979);
and_5  g10631(new_n12979, new_n12948, new_n12980_1);
or_5   g10632(new_n12980_1, new_n12946, new_n12981);
and_5  g10633(new_n12981, new_n12945, new_n12982);
nor_5  g10634(new_n12982, new_n12943, new_n12983);
nor_5  g10635(new_n12983, new_n12941_1, new_n12984);
and_5  g10636(new_n12939, new_n6997, new_n12985_1);
xor_4  g10637(new_n12985_1, new_n7223, new_n12986);
xor_4  g10638(new_n12986, n8305, new_n12987_1);
xnor_4 g10639(new_n12987_1, new_n12984, new_n12988);
not_10 g10640(new_n12988, new_n12989);
and_5  g10641(new_n12989, new_n12932, new_n12990);
xor_4  g10642(new_n12989, new_n12932, new_n12991);
not_10 g10643(new_n12991, new_n12992_1);
xor_4  g10644(new_n12928, new_n12917_1, new_n12993);
xor_4  g10645(new_n12982, new_n12943, new_n12994);
not_10 g10646(new_n12994, new_n12995);
nand_5 g10647(new_n12995, new_n12993, new_n12996);
xor_4  g10648(new_n12995, new_n12993, new_n12997);
not_10 g10649(new_n12997, new_n12998);
xor_4  g10650(new_n12927, new_n12918, new_n12999);
not_10 g10651(new_n12999, new_n13000);
xor_4  g10652(new_n12980_1, new_n12946, new_n13001);
or_5   g10653(new_n13001, new_n13000, new_n13002);
xor_4  g10654(new_n13001, new_n13000, new_n13003);
not_10 g10655(new_n13003, new_n13004);
xor_4  g10656(new_n12926, new_n3724, new_n13005_1);
xor_4  g10657(new_n12978_1, new_n12950, new_n13006);
not_10 g10658(new_n13006, new_n13007);
nand_5 g10659(new_n13007, new_n13005_1, new_n13008);
xor_4  g10660(new_n13007, new_n13005_1, new_n13009);
not_10 g10661(new_n13009, new_n13010);
xor_4  g10662(new_n12925, new_n3739, new_n13011);
not_10 g10663(new_n13011, new_n13012);
xor_4  g10664(new_n12976, new_n12954, new_n13013);
or_5   g10665(new_n13013, new_n13012, new_n13014);
xor_4  g10666(new_n13013, new_n13011, new_n13015);
xor_4  g10667(new_n12924, new_n12919, new_n13016);
not_10 g10668(new_n13016, new_n13017);
xor_4  g10669(new_n12974, new_n12957, new_n13018);
or_5   g10670(new_n13018, new_n13017, new_n13019);
xor_4  g10671(new_n13018, new_n13016, new_n13020);
xor_4  g10672(new_n12923, new_n12920, new_n13021);
not_10 g10673(new_n13021, new_n13022);
xor_4  g10674(new_n12972, new_n12971, new_n13023);
or_5   g10675(new_n13023, new_n13022, new_n13024);
xor_4  g10676(new_n13023, new_n13021, new_n13025);
xor_4  g10677(new_n12969, new_n12963, new_n13026_1);
not_10 g10678(new_n13026_1, new_n13027);
xor_4  g10679(new_n12922, new_n12921, new_n13028);
nand_5 g10680(new_n13028, new_n13027, new_n13029);
xor_4  g10681(new_n13028, new_n13027, new_n13030);
xnor_4 g10682(n7876, n4964, new_n13031);
xor_4  g10683(new_n12967, new_n12966, new_n13032);
or_5   g10684(new_n13032, new_n13031, new_n13033);
xor_4  g10685(n22309, n5704, new_n13034);
and_5  g10686(new_n13034, n7876, new_n13035);
xor_4  g10687(new_n13032, new_n13031, new_n13036);
nand_5 g10688(new_n13036, new_n13035, new_n13037);
nand_5 g10689(new_n13037, new_n13033, new_n13038);
nand_5 g10690(new_n13038, new_n13030, new_n13039);
and_5  g10691(new_n13039, new_n13029, new_n13040);
or_5   g10692(new_n13040, new_n13025, new_n13041);
and_5  g10693(new_n13041, new_n13024, new_n13042);
or_5   g10694(new_n13042, new_n13020, new_n13043_1);
and_5  g10695(new_n13043_1, new_n13019, new_n13044_1);
or_5   g10696(new_n13044_1, new_n13015, new_n13045);
and_5  g10697(new_n13045, new_n13014, new_n13046);
or_5   g10698(new_n13046, new_n13010, new_n13047);
and_5  g10699(new_n13047, new_n13008, new_n13048_1);
or_5   g10700(new_n13048_1, new_n13004, new_n13049);
and_5  g10701(new_n13049, new_n13002, new_n13050);
or_5   g10702(new_n13050, new_n12998, new_n13051);
and_5  g10703(new_n13051, new_n12996, new_n13052);
nor_5  g10704(new_n13052, new_n12992_1, new_n13053);
nor_5  g10705(new_n13053, new_n12990, new_n13054_1);
and_5  g10706(new_n13054_1, new_n12931, new_n13055);
not_10 g10707(new_n13055, new_n13056);
nand_5 g10708(new_n12985_1, new_n7223, new_n13057);
nor_5  g10709(new_n12986, n8305, new_n13058);
and_5  g10710(new_n12986, n8305, new_n13059);
nor_5  g10711(new_n13059, new_n12984, new_n13060);
or_5   g10712(new_n13060, new_n13058, new_n13061);
and_5  g10713(new_n13061, new_n13057, new_n13062);
nor_5  g10714(new_n13062, new_n13056, new_n13063);
xor_4  g10715(new_n13063, new_n12915, new_n13064);
xnor_4 g10716(new_n12914, new_n12911, new_n13065);
xor_4  g10717(new_n13062, new_n13056, new_n13066);
not_10 g10718(new_n13066, new_n13067);
nor_5  g10719(new_n13067, new_n13065, new_n13068);
xnor_4 g10720(new_n13066, new_n13065, new_n13069);
xor_4  g10721(new_n12909, new_n12861_1, new_n13070);
xor_4  g10722(new_n13052, new_n12992_1, new_n13071);
not_10 g10723(new_n13071, new_n13072);
and_5  g10724(new_n13072, new_n13070, new_n13073);
xor_4  g10725(new_n13072, new_n13070, new_n13074_1);
xor_4  g10726(new_n12907, new_n12865_1, new_n13075);
xor_4  g10727(new_n13050, new_n12998, new_n13076);
not_10 g10728(new_n13076, new_n13077);
and_5  g10729(new_n13077, new_n13075, new_n13078);
xor_4  g10730(new_n13077, new_n13075, new_n13079);
xor_4  g10731(new_n12905, new_n12869, new_n13080);
not_10 g10732(new_n13080, new_n13081);
xor_4  g10733(new_n13048_1, new_n13004, new_n13082_1);
nor_5  g10734(new_n13082_1, new_n13081, new_n13083);
xor_4  g10735(new_n13082_1, new_n13081, new_n13084);
not_10 g10736(new_n13084, new_n13085);
xor_4  g10737(new_n12903, new_n12873_1, new_n13086);
xnor_4 g10738(new_n13046, new_n13009, new_n13087);
not_10 g10739(new_n13087, new_n13088);
and_5  g10740(new_n13088, new_n13086, new_n13089);
xor_4  g10741(new_n13088, new_n13086, new_n13090);
xor_4  g10742(new_n12901, new_n12877, new_n13091);
not_10 g10743(new_n13091, new_n13092);
xor_4  g10744(new_n13044_1, new_n13015, new_n13093);
nor_5  g10745(new_n13093, new_n13092, new_n13094);
xor_4  g10746(new_n13093, new_n13092, new_n13095);
not_10 g10747(new_n13095, new_n13096_1);
xor_4  g10748(new_n12899, new_n12881, new_n13097);
not_10 g10749(new_n13097, new_n13098);
xor_4  g10750(new_n13042, new_n13020, new_n13099);
nor_5  g10751(new_n13099, new_n13098, new_n13100);
xor_4  g10752(new_n13099, new_n13098, new_n13101);
not_10 g10753(new_n13101, new_n13102);
xor_4  g10754(new_n12897, new_n12885, new_n13103);
not_10 g10755(new_n13103, new_n13104);
xor_4  g10756(new_n13040, new_n13025, new_n13105);
nor_5  g10757(new_n13105, new_n13104, new_n13106);
xor_4  g10758(new_n13105, new_n13104, new_n13107);
not_10 g10759(new_n13107, new_n13108);
xor_4  g10760(new_n12895, new_n12888, new_n13109);
and_5  g10761(new_n13037, new_n13033, new_n13110_1);
xnor_4 g10762(new_n13110_1, new_n13030, new_n13111);
not_10 g10763(new_n13111, new_n13112);
and_5  g10764(new_n13112, new_n13109, new_n13113);
not_10 g10765(new_n13113, new_n13114);
xor_4  g10766(new_n13112, new_n13109, new_n13115);
xor_4  g10767(new_n13036, new_n13035, new_n13116_1);
xor_4  g10768(new_n12893, new_n12892_1, new_n13117);
and_5  g10769(new_n13117, new_n13116_1, new_n13118);
xor_4  g10770(new_n12889, n11479, new_n13119);
xor_4  g10771(new_n13034, n7876, new_n13120);
and_5  g10772(new_n13120, new_n13119, new_n13121);
not_10 g10773(new_n13116_1, new_n13122_1);
xnor_4 g10774(new_n13117, new_n13122_1, new_n13123);
and_5  g10775(new_n13123, new_n13121, new_n13124);
nor_5  g10776(new_n13124, new_n13118, new_n13125);
and_5  g10777(new_n13125, new_n13115, new_n13126);
not_10 g10778(new_n13126, new_n13127);
and_5  g10779(new_n13127, new_n13114, new_n13128);
nor_5  g10780(new_n13128, new_n13108, new_n13129);
nor_5  g10781(new_n13129, new_n13106, new_n13130);
nor_5  g10782(new_n13130, new_n13102, new_n13131);
nor_5  g10783(new_n13131, new_n13100, new_n13132);
nor_5  g10784(new_n13132, new_n13096_1, new_n13133);
nor_5  g10785(new_n13133, new_n13094, new_n13134);
not_10 g10786(new_n13134, new_n13135);
and_5  g10787(new_n13135, new_n13090, new_n13136);
nor_5  g10788(new_n13136, new_n13089, new_n13137_1);
nor_5  g10789(new_n13137_1, new_n13085, new_n13138);
nor_5  g10790(new_n13138, new_n13083, new_n13139);
not_10 g10791(new_n13139, new_n13140);
and_5  g10792(new_n13140, new_n13079, new_n13141_1);
nor_5  g10793(new_n13141_1, new_n13078, new_n13142);
not_10 g10794(new_n13142, new_n13143);
and_5  g10795(new_n13143, new_n13074_1, new_n13144_1);
nor_5  g10796(new_n13144_1, new_n13073, new_n13145);
not_10 g10797(new_n13145, new_n13146);
and_5  g10798(new_n13146, new_n13069, new_n13147);
nor_5  g10799(new_n13147, new_n13068, new_n13148);
xor_4  g10800(new_n13148, new_n13064, n2095);
xnor_4 g10801(new_n11584, new_n11582, n2105);
xor_4  g10802(n23166, n11898, new_n13151);
nand_5 g10803(n19941, n10577, new_n13152);
or_5   g10804(n19941, n10577, new_n13153);
nor_5  g10805(n6381, n1099, new_n13154);
nor_5  g10806(new_n10759, new_n10744, new_n13155);
nor_5  g10807(new_n13155, new_n13154, new_n13156);
nand_5 g10808(new_n13156, new_n13153, new_n13157);
and_5  g10809(new_n13157, new_n13152, new_n13158);
xor_4  g10810(new_n13158, new_n13151, new_n13159);
xor_4  g10811(new_n13159, n8827, new_n13160);
xor_4  g10812(n19941, n10577, new_n13161);
xor_4  g10813(new_n13161, new_n13156, new_n13162);
nand_5 g10814(new_n13162, n18035, new_n13163);
xor_4  g10815(new_n13162, n18035, new_n13164);
nand_5 g10816(new_n10760, new_n10743, new_n13165);
nand_5 g10817(new_n10782, new_n10761, new_n13166);
and_5  g10818(new_n13166, new_n13165, new_n13167);
nand_5 g10819(new_n13167, new_n13164, new_n13168_1);
and_5  g10820(new_n13168_1, new_n13163, new_n13169);
xor_4  g10821(new_n13169, new_n13160, new_n13170);
xnor_4 g10822(new_n13170, new_n6126, new_n13171);
not_10 g10823(new_n13171, new_n13172);
not_10 g10824(new_n6128, new_n13173);
xor_4  g10825(new_n13167, new_n13164, new_n13174);
and_5  g10826(new_n13174, new_n13173, new_n13175);
xnor_4 g10827(new_n13174, new_n6128, new_n13176);
not_10 g10828(new_n13176, new_n13177);
nor_5  g10829(new_n10783, new_n6135, new_n13178);
xor_4  g10830(new_n10783, new_n6135, new_n13179);
not_10 g10831(new_n13179, new_n13180);
not_10 g10832(new_n6140, new_n13181);
and_5  g10833(new_n10786, new_n13181, new_n13182);
xnor_4 g10834(new_n10786, new_n6140, new_n13183);
not_10 g10835(new_n13183, new_n13184);
nor_5  g10836(new_n10792_1, new_n6145, new_n13185);
xor_4  g10837(new_n10792_1, new_n6145, new_n13186);
not_10 g10838(new_n13186, new_n13187);
xnor_4 g10839(new_n10775_1, new_n10772, new_n13188);
nor_5  g10840(new_n13188, new_n6150, new_n13189);
xnor_4 g10841(new_n10796, new_n6150, new_n13190_1);
not_10 g10842(new_n13190_1, new_n13191);
xnor_4 g10843(new_n8620_1, new_n8617, new_n13192);
nor_5  g10844(new_n13192, new_n6155, new_n13193);
xnor_4 g10845(new_n8621, new_n6155, new_n13194);
not_10 g10846(new_n13194, new_n13195);
nor_5  g10847(new_n8599, new_n6160_1, new_n13196);
xor_4  g10848(new_n8599, new_n6160_1, new_n13197);
not_10 g10849(new_n13197, new_n13198_1);
not_10 g10850(new_n6164, new_n13199_1);
nor_5  g10851(new_n8603, new_n13199_1, new_n13200);
not_10 g10852(new_n13200, new_n13201);
and_5  g10853(new_n8606, new_n6167, new_n13202);
xor_4  g10854(new_n8603, new_n13199_1, new_n13203);
and_5  g10855(new_n13203, new_n13202, new_n13204_1);
not_10 g10856(new_n13204_1, new_n13205);
and_5  g10857(new_n13205, new_n13201, new_n13206);
nor_5  g10858(new_n13206, new_n13198_1, new_n13207);
nor_5  g10859(new_n13207, new_n13196, new_n13208);
nor_5  g10860(new_n13208, new_n13195, new_n13209_1);
nor_5  g10861(new_n13209_1, new_n13193, new_n13210);
nor_5  g10862(new_n13210, new_n13191, new_n13211);
nor_5  g10863(new_n13211, new_n13189, new_n13212);
nor_5  g10864(new_n13212, new_n13187, new_n13213);
nor_5  g10865(new_n13213, new_n13185, new_n13214);
nor_5  g10866(new_n13214, new_n13184, new_n13215);
nor_5  g10867(new_n13215, new_n13182, new_n13216);
nor_5  g10868(new_n13216, new_n13180, new_n13217);
nor_5  g10869(new_n13217, new_n13178, new_n13218);
nor_5  g10870(new_n13218, new_n13177, new_n13219);
nor_5  g10871(new_n13219, new_n13175, new_n13220);
xnor_4 g10872(new_n13220, new_n13172, n2122);
xor_4  g10873(new_n2823, new_n2799, n2147);
xnor_4 g10874(new_n10708, new_n10668, n2209);
xnor_4 g10875(new_n5831, new_n5704_1, n2214);
xor_4  g10876(new_n11358, new_n4190, new_n13225);
nand_5 g10877(new_n11360, new_n4279, new_n13226);
xor_4  g10878(new_n11360, new_n4279, new_n13227);
nor_5  g10879(new_n11364, new_n4283, new_n13228);
xor_4  g10880(new_n11364, new_n4283, new_n13229);
nand_5 g10881(new_n11370, new_n4289, new_n13230);
and_5  g10882(new_n11367, new_n4291, new_n13231);
xor_4  g10883(new_n11370, new_n4289, new_n13232);
not_10 g10884(new_n13232, new_n13233);
or_5   g10885(new_n13233, new_n13231, new_n13234);
and_5  g10886(new_n13234, new_n13230, new_n13235);
and_5  g10887(new_n13235, new_n13229, new_n13236);
nor_5  g10888(new_n13236, new_n13228, new_n13237);
nand_5 g10889(new_n13237, new_n13227, new_n13238);
and_5  g10890(new_n13238, new_n13226, new_n13239);
xor_4  g10891(new_n13239, new_n13225, n2238);
xor_4  g10892(new_n11380, new_n11379_1, n2327);
xnor_4 g10893(new_n5815, new_n5776_1, n2343);
xor_4  g10894(new_n10770, new_n7913, new_n13243);
or_5   g10895(new_n6645, new_n6634_1, new_n13244);
or_5   g10896(new_n6662, new_n6647, new_n13245);
and_5  g10897(new_n13245, new_n13244, new_n13246);
xor_4  g10898(new_n13246, new_n13243, new_n13247);
xnor_4 g10899(n20923, n16524, new_n13248);
or_5   g10900(n18157, n11056, new_n13249);
or_5   g10901(new_n6674_1, new_n6665, new_n13250);
and_5  g10902(new_n13250, new_n13249, new_n13251);
xor_4  g10903(new_n13251, new_n13248, new_n13252);
xor_4  g10904(new_n13252, new_n10813, new_n13253);
not_10 g10905(new_n13253, new_n13254);
nand_5 g10906(new_n6675, new_n6664, new_n13255);
or_5   g10907(new_n6689, new_n6677, new_n13256);
and_5  g10908(new_n13256, new_n13255, new_n13257);
xor_4  g10909(new_n13257, new_n13254, new_n13258);
xor_4  g10910(new_n13258, new_n13247, new_n13259);
not_10 g10911(new_n13259, new_n13260);
and_5  g10912(new_n6690, new_n6663, new_n13261);
not_10 g10913(new_n13261, new_n13262);
and_5  g10914(new_n6708, new_n6691_1, new_n13263_1);
not_10 g10915(new_n13263_1, new_n13264);
and_5  g10916(new_n13264, new_n13262, new_n13265);
xnor_4 g10917(new_n13265, new_n13260, n2361);
xor_4  g10918(new_n3704, new_n3703, n2363);
xnor_4 g10919(new_n4594, new_n4561, n2374);
xnor_4 g10920(n7305, n1204, new_n13269);
or_5   g10921(n25872, n19618, new_n13270_1);
or_5   g10922(new_n5887, new_n5882_1, new_n13271);
and_5  g10923(new_n13271, new_n13270_1, new_n13272);
xor_4  g10924(new_n13272, new_n13269, new_n13273_1);
and_5  g10925(new_n13273_1, new_n4880, new_n13274);
xor_4  g10926(new_n13273_1, new_n4880, new_n13275);
or_5   g10927(new_n5888, new_n4884, new_n13276);
or_5   g10928(new_n5896, new_n5889, new_n13277);
and_5  g10929(new_n13277, new_n13276, new_n13278);
and_5  g10930(new_n13278, new_n13275, new_n13279);
or_5   g10931(new_n13279, new_n13274, new_n13280);
xnor_4 g10932(n20826, n626, new_n13281);
or_5   g10933(n7305, n1204, new_n13282);
or_5   g10934(new_n13272, new_n13269, new_n13283);
and_5  g10935(new_n13283, new_n13282, new_n13284);
xor_4  g10936(new_n13284, new_n13281, new_n13285_1);
xor_4  g10937(new_n13285_1, new_n13280, new_n13286);
xor_4  g10938(new_n13286, new_n4876, new_n13287);
xor_4  g10939(new_n13287, new_n3773, new_n13288);
xor_4  g10940(new_n13278, new_n13275, new_n13289);
or_5   g10941(new_n13289, new_n3779, new_n13290);
and_5  g10942(new_n5897, new_n3783, new_n13291);
and_5  g10943(new_n5906, new_n5898, new_n13292);
or_5   g10944(new_n13292, new_n13291, new_n13293);
xor_4  g10945(new_n13289, new_n3779, new_n13294);
nand_5 g10946(new_n13294, new_n13293, new_n13295);
and_5  g10947(new_n13295, new_n13290, new_n13296);
xor_4  g10948(new_n13296, new_n13288, n2388);
xor_4  g10949(n7335, n2160, new_n13298);
not_10 g10950(new_n13298, new_n13299);
or_5   g10951(n10763, n5696, new_n13300);
or_5   g10952(new_n5372, new_n5338, new_n13301);
and_5  g10953(new_n13301, new_n13300, new_n13302);
xor_4  g10954(new_n13302, new_n13299, new_n13303);
xor_4  g10955(n11220, n3425, new_n13304);
not_10 g10956(new_n13304, new_n13305);
or_5   g10957(n22379, n9967, new_n13306);
or_5   g10958(new_n5335, new_n5300_1, new_n13307);
and_5  g10959(new_n13307, new_n13306, new_n13308);
xor_4  g10960(new_n13308, new_n13305, new_n13309);
not_10 g10961(new_n13309, new_n13310);
xor_4  g10962(new_n13310, new_n13303, new_n13311);
not_10 g10963(new_n13311, new_n13312);
or_5   g10964(new_n5373, new_n5337_1, new_n13313);
or_5   g10965(new_n5425, new_n5374, new_n13314);
and_5  g10966(new_n13314, new_n13313, new_n13315);
xor_4  g10967(new_n13315, new_n13312, new_n13316);
not_10 g10968(new_n13316, new_n13317);
not_10 g10969(n7593, new_n13318);
and_5  g10970(new_n5255_1, new_n5242, new_n13319_1);
xor_4  g10971(new_n13319_1, new_n13318, new_n13320);
xor_4  g10972(new_n13320, new_n3075, new_n13321);
nor_5  g10973(new_n5256_1, n6485, new_n13322);
not_10 g10974(new_n5257, new_n13323);
nor_5  g10975(new_n5297, new_n13323, new_n13324);
nor_5  g10976(new_n13324, new_n13322, new_n13325);
xor_4  g10977(new_n13325, new_n13321, new_n13326);
xnor_4 g10978(new_n13326, new_n13317, new_n13327);
nand_5 g10979(new_n5426, new_n5298, new_n13328);
nand_5 g10980(new_n5478, new_n5427, new_n13329);
and_5  g10981(new_n13329, new_n13328, new_n13330);
xor_4  g10982(new_n13330, new_n13327, n2440);
xnor_4 g10983(new_n11747, new_n11731, n2444);
xnor_4 g10984(new_n5101_1, new_n3242, n2513);
xor_4  g10985(new_n5998, n14323, new_n13334);
not_10 g10986(new_n13334, new_n13335);
nand_5 g10987(new_n6003, n2886, new_n13336);
xnor_4 g10988(new_n6003, n2886, new_n13337);
nand_5 g10989(new_n6014, n1040, new_n13338_1);
and_5  g10990(n20658, n9090, new_n13339);
xor_4  g10991(new_n6014, n1040, new_n13340);
nand_5 g10992(new_n13340, new_n13339, new_n13341);
and_5  g10993(new_n13341, new_n13338_1, new_n13342);
or_5   g10994(new_n13342, new_n13337, new_n13343);
and_5  g10995(new_n13343, new_n13336, new_n13344);
xor_4  g10996(new_n13344, new_n13335, new_n13345);
not_10 g10997(new_n13345, new_n13346);
xnor_4 g10998(new_n13346, n12562, new_n13347);
xor_4  g10999(new_n13342, new_n13337, new_n13348);
or_5   g11000(new_n13348, n7949, new_n13349);
not_10 g11001(n7949, new_n13350);
xor_4  g11002(new_n13348, new_n13350, new_n13351);
and_5  g11003(new_n11072, n14575, new_n13352);
or_5   g11004(new_n13352, n24374, new_n13353);
xor_4  g11005(new_n13340, new_n13339, new_n13354);
not_10 g11006(new_n13354, new_n13355);
xor_4  g11007(new_n13352, n24374, new_n13356);
nand_5 g11008(new_n13356, new_n13355, new_n13357);
and_5  g11009(new_n13357, new_n13353, new_n13358);
or_5   g11010(new_n13358, new_n13351, new_n13359);
and_5  g11011(new_n13359, new_n13349, new_n13360);
xor_4  g11012(new_n13360, new_n13347, new_n13361);
xor_4  g11013(new_n13361, new_n13105, new_n13362);
not_10 g11014(new_n13362, new_n13363);
xor_4  g11015(new_n13358, new_n13351, new_n13364);
nand_5 g11016(new_n13364, new_n13112, new_n13365);
xnor_4 g11017(new_n13364, new_n13111, new_n13366);
not_10 g11018(new_n13366, new_n13367_1);
xor_4  g11019(new_n13356, new_n13355, new_n13368);
nand_5 g11020(new_n13368, new_n13122_1, new_n13369);
xor_4  g11021(new_n11072, n14575, new_n13370);
nand_5 g11022(new_n13370, new_n13120, new_n13371);
xor_4  g11023(new_n13368, new_n13122_1, new_n13372);
nand_5 g11024(new_n13372, new_n13371, new_n13373);
and_5  g11025(new_n13373, new_n13369, new_n13374);
or_5   g11026(new_n13374, new_n13367_1, new_n13375);
and_5  g11027(new_n13375, new_n13365, new_n13376);
xnor_4 g11028(new_n13376, new_n13363, n2515);
xnor_4 g11029(new_n11064, new_n11029, n2533);
and_5  g11030(new_n7223, n3425, new_n13379);
not_10 g11031(new_n13379, new_n13380);
xnor_4 g11032(n26986, n3425, new_n13381);
not_10 g11033(new_n13381, new_n13382);
or_5   g11034(n21287, new_n3184, new_n13383);
xnor_4 g11035(n21287, n9967, new_n13384);
not_10 g11036(new_n13384, new_n13385);
or_5   g11037(new_n3185, n4256, new_n13386);
xnor_4 g11038(n20946, n4256, new_n13387);
not_10 g11039(new_n13387, new_n13388);
or_5   g11040(n22332, new_n3186, new_n13389);
xnor_4 g11041(n22332, n7751, new_n13390);
not_10 g11042(new_n13390, new_n13391);
or_5   g11043(new_n3187, n18907, new_n13392);
xor_4  g11044(n26823, n18907, new_n13393);
or_5   g11045(new_n3188, n2731, new_n13394);
or_5   g11046(new_n8556, new_n8540, new_n13395);
and_5  g11047(new_n13395, new_n13394, new_n13396);
or_5   g11048(new_n13396, new_n13393, new_n13397);
and_5  g11049(new_n13397, new_n13392, new_n13398);
or_5   g11050(new_n13398, new_n13391, new_n13399);
and_5  g11051(new_n13399, new_n13389, new_n13400);
or_5   g11052(new_n13400, new_n13388, new_n13401);
and_5  g11053(new_n13401, new_n13386, new_n13402);
or_5   g11054(new_n13402, new_n13385, new_n13403);
and_5  g11055(new_n13403, new_n13383, new_n13404);
nor_5  g11056(new_n13404, new_n13382, new_n13405);
not_10 g11057(new_n13405, new_n13406);
and_5  g11058(new_n13406, new_n13380, new_n13407_1);
and_5  g11059(new_n5140_1, new_n5134, new_n13408);
and_5  g11060(new_n7098, new_n13408, new_n13409_1);
and_5  g11061(new_n13409_1, new_n7095, new_n13410);
and_5  g11062(new_n13410, new_n7090, new_n13411);
and_5  g11063(new_n13411, new_n7146, new_n13412);
not_10 g11064(new_n13412, new_n13413);
nor_5  g11065(new_n13413, new_n7234, new_n13414);
and_5  g11066(new_n13413, new_n7236_1, new_n13415);
nor_5  g11067(new_n13415, new_n13414, new_n13416);
nor_5  g11068(new_n13416, new_n3180, new_n13417);
xor_4  g11069(new_n13411, new_n7146, new_n13418);
nor_5  g11070(new_n13418, new_n3119, new_n13419_1);
xnor_4 g11071(new_n13418, new_n3118, new_n13420);
not_10 g11072(new_n13420, new_n13421);
xor_4  g11073(new_n13410, new_n7090, new_n13422);
or_5   g11074(new_n13422, new_n3124, new_n13423);
xnor_4 g11075(new_n13422, new_n3122, new_n13424_1);
not_10 g11076(new_n13424_1, new_n13425);
xor_4  g11077(new_n13409_1, new_n7095, new_n13426);
or_5   g11078(new_n13426, new_n3128, new_n13427);
xnor_4 g11079(new_n13426, new_n3126_1, new_n13428);
not_10 g11080(new_n13428, new_n13429);
xnor_4 g11081(new_n7099_1, new_n13408, new_n13430);
or_5   g11082(new_n13430, new_n3132, new_n13431);
xnor_4 g11083(new_n13430, new_n3130, new_n13432);
not_10 g11084(new_n13432, new_n13433);
or_5   g11085(new_n5142, new_n3136_1, new_n13434);
or_5   g11086(new_n5175, new_n5144, new_n13435);
and_5  g11087(new_n13435, new_n13434, new_n13436);
or_5   g11088(new_n13436, new_n13433, new_n13437);
and_5  g11089(new_n13437, new_n13431, new_n13438);
or_5   g11090(new_n13438, new_n13429, new_n13439);
and_5  g11091(new_n13439, new_n13427, new_n13440);
or_5   g11092(new_n13440, new_n13425, new_n13441);
and_5  g11093(new_n13441, new_n13423, new_n13442);
nor_5  g11094(new_n13442, new_n13421, new_n13443);
nor_5  g11095(new_n13443, new_n13419_1, new_n13444);
and_5  g11096(new_n13416, new_n3180, new_n13445);
nor_5  g11097(new_n13445, new_n13444, new_n13446);
nor_5  g11098(new_n13446, new_n13417, new_n13447);
nor_5  g11099(new_n13447, new_n13414, new_n13448);
xor_4  g11100(new_n13448, new_n13407_1, new_n13449);
xnor_4 g11101(new_n13416, new_n3180, new_n13450);
xor_4  g11102(new_n13450, new_n13444, new_n13451);
not_10 g11103(new_n13451, new_n13452);
nor_5  g11104(new_n13452, new_n13407_1, new_n13453_1);
xor_4  g11105(new_n13452, new_n13407_1, new_n13454);
xor_4  g11106(new_n13404, new_n13382, new_n13455);
not_10 g11107(new_n13455, new_n13456_1);
xor_4  g11108(new_n13442, new_n13421, new_n13457_1);
and_5  g11109(new_n13457_1, new_n13456_1, new_n13458);
xor_4  g11110(new_n13457_1, new_n13456_1, new_n13459);
not_10 g11111(new_n13459, new_n13460_1);
xor_4  g11112(new_n13402, new_n13385, new_n13461);
not_10 g11113(new_n13461, new_n13462);
xor_4  g11114(new_n13440, new_n13425, new_n13463);
and_5  g11115(new_n13463, new_n13462, new_n13464);
xor_4  g11116(new_n13463, new_n13462, new_n13465);
not_10 g11117(new_n13465, new_n13466);
xor_4  g11118(new_n13400, new_n13388, new_n13467);
not_10 g11119(new_n13467, new_n13468);
xor_4  g11120(new_n13438, new_n13429, new_n13469);
and_5  g11121(new_n13469, new_n13468, new_n13470);
xor_4  g11122(new_n13469, new_n13468, new_n13471);
not_10 g11123(new_n13471, new_n13472);
xor_4  g11124(new_n13398, new_n13391, new_n13473);
xor_4  g11125(new_n13436, new_n13433, new_n13474);
not_10 g11126(new_n13474, new_n13475);
nor_5  g11127(new_n13475, new_n13473, new_n13476);
not_10 g11128(new_n13476, new_n13477_1);
xor_4  g11129(new_n13475, new_n13473, new_n13478);
xor_4  g11130(new_n13396, new_n13393, new_n13479);
and_5  g11131(new_n13479, new_n5177, new_n13480);
xnor_4 g11132(new_n13479, new_n5177, new_n13481);
nand_5 g11133(new_n8557, new_n5207, new_n13482);
nand_5 g11134(new_n8577, new_n8558, new_n13483);
and_5  g11135(new_n13483, new_n13482, new_n13484_1);
nor_5  g11136(new_n13484_1, new_n13481, new_n13485);
nor_5  g11137(new_n13485, new_n13480, new_n13486_1);
and_5  g11138(new_n13486_1, new_n13478, new_n13487_1);
not_10 g11139(new_n13487_1, new_n13488);
and_5  g11140(new_n13488, new_n13477_1, new_n13489);
nor_5  g11141(new_n13489, new_n13472, new_n13490_1);
nor_5  g11142(new_n13490_1, new_n13470, new_n13491);
nor_5  g11143(new_n13491, new_n13466, new_n13492);
nor_5  g11144(new_n13492, new_n13464, new_n13493);
nor_5  g11145(new_n13493, new_n13460_1, new_n13494_1);
nor_5  g11146(new_n13494_1, new_n13458, new_n13495);
not_10 g11147(new_n13495, new_n13496);
and_5  g11148(new_n13496, new_n13454, new_n13497);
nor_5  g11149(new_n13497, new_n13453_1, new_n13498);
xor_4  g11150(new_n13498, new_n13449, n2535);
nor_5  g11151(n20259, n3925, new_n13500_1);
and_5  g11152(new_n13500_1, new_n4946, new_n13501_1);
and_5  g11153(new_n13501_1, new_n4943, new_n13502);
and_5  g11154(new_n13502, new_n4939_1, new_n13503);
xor_4  g11155(new_n13503, new_n4935, new_n13504);
xor_4  g11156(new_n13504, new_n8351, new_n13505);
xor_4  g11157(new_n13502, new_n4939_1, new_n13506_1);
or_5   g11158(new_n13506_1, n17251, new_n13507);
xor_4  g11159(new_n13506_1, new_n8352, new_n13508);
xor_4  g11160(new_n13501_1, new_n4943, new_n13509);
or_5   g11161(new_n13509, n14790, new_n13510);
xor_4  g11162(new_n13500_1, new_n4946, new_n13511);
nor_5  g11163(new_n13511, n10096, new_n13512);
xor_4  g11164(new_n13511, new_n3556, new_n13513);
xor_4  g11165(n20259, n3925, new_n13514);
or_5   g11166(new_n13514, n16994, new_n13515);
nand_5 g11167(n9246, n3925, new_n13516);
xor_4  g11168(new_n13514, n16994, new_n13517);
nand_5 g11169(new_n13517, new_n13516, new_n13518);
and_5  g11170(new_n13518, new_n13515, new_n13519);
nor_5  g11171(new_n13519, new_n13513, new_n13520);
or_5   g11172(new_n13520, new_n13512, new_n13521);
xor_4  g11173(new_n13509, n14790, new_n13522);
nand_5 g11174(new_n13522, new_n13521, new_n13523);
and_5  g11175(new_n13523, new_n13510, new_n13524);
or_5   g11176(new_n13524, new_n13508, new_n13525);
and_5  g11177(new_n13525, new_n13507, new_n13526);
xor_4  g11178(new_n13526, new_n13505, new_n13527);
xnor_4 g11179(new_n13527, new_n7855, new_n13528);
not_10 g11180(new_n13528, new_n13529);
not_10 g11181(new_n7860, new_n13530);
xor_4  g11182(new_n13524, new_n13508, new_n13531);
nand_5 g11183(new_n13531, new_n13530, new_n13532);
xor_4  g11184(new_n13531, new_n7860, new_n13533);
xor_4  g11185(new_n13522, new_n13521, new_n13534);
nand_5 g11186(new_n13534, new_n7867, new_n13535);
xnor_4 g11187(new_n13534, new_n7866, new_n13536);
xor_4  g11188(new_n13519, new_n13513, new_n13537);
or_5   g11189(new_n13537, new_n7874, new_n13538);
xor_4  g11190(new_n13537, new_n7874, new_n13539);
not_10 g11191(new_n13539, new_n13540);
xor_4  g11192(new_n13517, new_n13516, new_n13541);
or_5   g11193(new_n13541, new_n7881, new_n13542);
not_10 g11194(new_n9950, new_n13543);
nor_5  g11195(new_n13543, new_n7884_1, new_n13544);
xor_4  g11196(new_n13541, new_n7881, new_n13545);
nand_5 g11197(new_n13545, new_n13544, new_n13546);
and_5  g11198(new_n13546, new_n13542, new_n13547);
or_5   g11199(new_n13547, new_n13540, new_n13548_1);
and_5  g11200(new_n13548_1, new_n13538, new_n13549_1);
nand_5 g11201(new_n13549_1, new_n13536, new_n13550);
and_5  g11202(new_n13550, new_n13535, new_n13551_1);
or_5   g11203(new_n13551_1, new_n13533, new_n13552);
and_5  g11204(new_n13552, new_n13532, new_n13553);
xor_4  g11205(new_n13553, new_n13529, new_n13554);
xor_4  g11206(n1163, n329, new_n13555);
not_10 g11207(n24170, new_n13556);
or_5   g11208(new_n13556, n18537, new_n13557);
xnor_4 g11209(n24170, n18537, new_n13558);
not_10 g11210(new_n13558, new_n13559);
or_5   g11211(n7057, new_n8431, new_n13560);
xnor_4 g11212(n7057, n2409, new_n13561);
or_5   g11213(n8869, new_n8663, new_n13562);
nand_5 g11214(n8869, new_n8663, new_n13563);
nor_5  g11215(new_n5061, n10372, new_n13564);
and_5  g11216(n12495, new_n8437, new_n13565);
and_5  g11217(new_n5061, n10372, new_n13566);
not_10 g11218(new_n13566, new_n13567);
and_5  g11219(new_n13567, new_n13565, new_n13568);
nor_5  g11220(new_n13568, new_n13564, new_n13569);
not_10 g11221(new_n13569, new_n13570);
nand_5 g11222(new_n13570, new_n13563, new_n13571);
and_5  g11223(new_n13571, new_n13562, new_n13572);
nand_5 g11224(new_n13572, new_n13561, new_n13573);
and_5  g11225(new_n13573, new_n13560, new_n13574);
or_5   g11226(new_n13574, new_n13559, new_n13575);
and_5  g11227(new_n13575, new_n13557, new_n13576);
xor_4  g11228(new_n13576, new_n13555, new_n13577);
xnor_4 g11229(new_n13577, new_n13554, new_n13578);
not_10 g11230(new_n13578, new_n13579);
xor_4  g11231(new_n13574, new_n13559, new_n13580);
not_10 g11232(new_n13580, new_n13581);
xor_4  g11233(new_n13551_1, new_n13533, new_n13582);
nand_5 g11234(new_n13582, new_n13581, new_n13583);
xor_4  g11235(new_n13582, new_n13581, new_n13584);
not_10 g11236(new_n13584, new_n13585);
xor_4  g11237(new_n13549_1, new_n13536, new_n13586);
not_10 g11238(new_n13586, new_n13587);
xor_4  g11239(new_n13572, new_n13561, new_n13588);
or_5   g11240(new_n13588, new_n13587, new_n13589);
xor_4  g11241(new_n13588, new_n13587, new_n13590);
xor_4  g11242(new_n13547, new_n13540, new_n13591);
xnor_4 g11243(n8869, n8381, new_n13592);
xor_4  g11244(new_n13592, new_n13570, new_n13593);
not_10 g11245(new_n13593, new_n13594);
or_5   g11246(new_n13594, new_n13591, new_n13595);
xnor_4 g11247(new_n13593, new_n13591, new_n13596);
not_10 g11248(new_n13596, new_n13597);
nor_5  g11249(new_n9953, new_n9952, new_n13598);
xnor_4 g11250(n20235, n10372, new_n13599);
xnor_4 g11251(new_n13599, new_n13565, new_n13600);
or_5   g11252(new_n13600, new_n13598, new_n13601);
xor_4  g11253(new_n13545, new_n13544, new_n13602_1);
xor_4  g11254(new_n13599, new_n13565, new_n13603);
xnor_4 g11255(new_n13603, new_n13598, new_n13604);
not_10 g11256(new_n13604, new_n13605);
or_5   g11257(new_n13605, new_n13602_1, new_n13606);
and_5  g11258(new_n13606, new_n13601, new_n13607);
or_5   g11259(new_n13607, new_n13597, new_n13608);
nand_5 g11260(new_n13608, new_n13595, new_n13609);
nand_5 g11261(new_n13609, new_n13590, new_n13610);
and_5  g11262(new_n13610, new_n13589, new_n13611);
or_5   g11263(new_n13611, new_n13585, new_n13612);
and_5  g11264(new_n13612, new_n13583, new_n13613);
xnor_4 g11265(new_n13613, new_n13579, n2537);
xor_4  g11266(new_n11242, new_n2966, new_n13615);
nand_5 g11267(new_n4197, new_n2971_1, new_n13616);
xnor_4 g11268(new_n4197, new_n2972, new_n13617);
or_5   g11269(new_n4200, new_n2977, new_n13618);
xnor_4 g11270(new_n4200, new_n2978_1, new_n13619);
nand_5 g11271(new_n4204_1, new_n2982, new_n13620);
xnor_4 g11272(new_n4204_1, new_n2983, new_n13621);
or_5   g11273(new_n4208, new_n2989, new_n13622);
not_10 g11274(n1152, new_n13623);
and_5  g11275(new_n3047, new_n13623, new_n13624);
xor_4  g11276(new_n4208, new_n2989, new_n13625);
nand_5 g11277(new_n13625, new_n13624, new_n13626_1);
and_5  g11278(new_n13626_1, new_n13622, new_n13627);
nand_5 g11279(new_n13627, new_n13621, new_n13628);
and_5  g11280(new_n13628, new_n13620, new_n13629);
nand_5 g11281(new_n13629, new_n13619, new_n13630);
and_5  g11282(new_n13630, new_n13618, new_n13631);
nand_5 g11283(new_n13631, new_n13617, new_n13632);
and_5  g11284(new_n13632, new_n13616, new_n13633);
xor_4  g11285(new_n13633, new_n13615, new_n13634);
xor_4  g11286(new_n13634, new_n11693, new_n13635);
not_10 g11287(new_n13635, new_n13636);
xor_4  g11288(new_n13631, new_n13617, new_n13637);
nor_5  g11289(new_n13637, new_n9762, new_n13638);
xor_4  g11290(new_n13637, new_n9762, new_n13639);
not_10 g11291(new_n13639, new_n13640);
xor_4  g11292(new_n13629, new_n13619, new_n13641);
and_5  g11293(new_n13641, new_n12276, new_n13642);
not_10 g11294(new_n13642, new_n13643);
xnor_4 g11295(new_n13641, new_n9764, new_n13644);
xor_4  g11296(new_n13627, new_n13621, new_n13645);
and_5  g11297(new_n13645, new_n9769, new_n13646);
xor_4  g11298(new_n13645, new_n9769, new_n13647);
xor_4  g11299(new_n13625, new_n13624, new_n13648);
nand_5 g11300(new_n13648, new_n9773, new_n13649);
xor_4  g11301(new_n3047, new_n13623, new_n13650);
nor_5  g11302(new_n13650, new_n7247, new_n13651);
xor_4  g11303(new_n13648, new_n9773, new_n13652);
not_10 g11304(new_n13652, new_n13653);
or_5   g11305(new_n13653, new_n13651, new_n13654);
and_5  g11306(new_n13654, new_n13649, new_n13655);
and_5  g11307(new_n13655, new_n13647, new_n13656);
nor_5  g11308(new_n13656, new_n13646, new_n13657);
and_5  g11309(new_n13657, new_n13644, new_n13658);
not_10 g11310(new_n13658, new_n13659);
and_5  g11311(new_n13659, new_n13643, new_n13660);
nor_5  g11312(new_n13660, new_n13640, new_n13661);
nor_5  g11313(new_n13661, new_n13638, new_n13662);
xnor_4 g11314(new_n13662, new_n13636, n2553);
xor_4  g11315(new_n12165, new_n12144, n2555);
xor_4  g11316(new_n10906, n12892, new_n13665);
not_10 g11317(new_n13665, new_n13666);
or_5   g11318(new_n13666, new_n10233, new_n13667);
and_5  g11319(new_n10906, n12892, new_n13668_1);
not_10 g11320(new_n13668_1, new_n13669);
xor_4  g11321(new_n10910, n12209, new_n13670);
xor_4  g11322(new_n13670, new_n13669, new_n13671);
xnor_4 g11323(new_n13671, new_n10228, new_n13672);
not_10 g11324(new_n13672, new_n13673);
xnor_4 g11325(new_n13673, new_n13667, n2560);
nor_5  g11326(n26180, n10650, new_n13675);
not_10 g11327(new_n13675, new_n13676);
xnor_4 g11328(n26180, n10650, new_n13677_1);
or_5   g11329(n24004, n12900, new_n13678);
xnor_4 g11330(n24004, n12900, new_n13679);
or_5   g11331(n20411, n12871, new_n13680);
xnor_4 g11332(n20411, n12871, new_n13681);
or_5   g11333(n23304, n17069, new_n13682);
xnor_4 g11334(n23304, n17069, new_n13683_1);
or_5   g11335(n19361, n15918, new_n13684);
xnor_4 g11336(n19361, n15918, new_n13685);
or_5   g11337(n17784, n1437, new_n13686);
xnor_4 g11338(n17784, n1437, new_n13687);
or_5   g11339(n14323, n4722, new_n13688);
xnor_4 g11340(n14323, n4722, new_n13689);
or_5   g11341(n14633, n2886, new_n13690);
xnor_4 g11342(n14633, n2886, new_n13691);
or_5   g11343(n8721, n1040, new_n13692);
and_5  g11344(n18578, n9090, new_n13693);
xnor_4 g11345(n8721, n1040, new_n13694);
or_5   g11346(new_n13694, new_n13693, new_n13695);
and_5  g11347(new_n13695, new_n13692, new_n13696);
or_5   g11348(new_n13696, new_n13691, new_n13697);
and_5  g11349(new_n13697, new_n13690, new_n13698);
or_5   g11350(new_n13698, new_n13689, new_n13699);
and_5  g11351(new_n13699, new_n13688, new_n13700);
or_5   g11352(new_n13700, new_n13687, new_n13701);
and_5  g11353(new_n13701, new_n13686, new_n13702);
or_5   g11354(new_n13702, new_n13685, new_n13703);
and_5  g11355(new_n13703, new_n13684, new_n13704);
or_5   g11356(new_n13704, new_n13683_1, new_n13705);
and_5  g11357(new_n13705, new_n13682, new_n13706);
or_5   g11358(new_n13706, new_n13681, new_n13707);
and_5  g11359(new_n13707, new_n13680, new_n13708_1);
or_5   g11360(new_n13708_1, new_n13679, new_n13709);
and_5  g11361(new_n13709, new_n13678, new_n13710_1);
nor_5  g11362(new_n13710_1, new_n13677_1, new_n13711);
not_10 g11363(new_n13711, new_n13712);
and_5  g11364(new_n13712, new_n13676, new_n13713);
nor_5  g11365(n9259, n6456, new_n13714_1);
nor_5  g11366(new_n5964_1, new_n5924, new_n13715);
nor_5  g11367(new_n13715, new_n13714_1, new_n13716);
not_10 g11368(new_n13716, new_n13717);
nor_5  g11369(new_n13717, new_n13713, new_n13718);
xor_4  g11370(new_n13717, new_n13713, new_n13719_1);
not_10 g11371(new_n13719_1, new_n13720);
xor_4  g11372(new_n13710_1, new_n13677_1, new_n13721);
nand_5 g11373(new_n13721, new_n5966, new_n13722_1);
xnor_4 g11374(new_n13721, new_n5966, new_n13723);
xor_4  g11375(new_n13708_1, new_n13679, new_n13724);
nand_5 g11376(new_n13724, new_n5972, new_n13725);
xnor_4 g11377(new_n13724, new_n5972, new_n13726);
xor_4  g11378(new_n13706, new_n13681, new_n13727);
nand_5 g11379(new_n13727, new_n5977, new_n13728);
xnor_4 g11380(new_n13727, new_n5977, new_n13729);
xor_4  g11381(new_n13704, new_n13683_1, new_n13730);
nand_5 g11382(new_n13730, new_n5983, new_n13731);
xnor_4 g11383(new_n13730, new_n5983, new_n13732);
xor_4  g11384(new_n13702, new_n13685, new_n13733);
nand_5 g11385(new_n13733, new_n5989, new_n13734);
xor_4  g11386(new_n13733, new_n5989, new_n13735);
xor_4  g11387(new_n13700, new_n13687, new_n13736);
or_5   g11388(new_n13736, new_n5995, new_n13737);
xnor_4 g11389(new_n13736, new_n5995, new_n13738);
xor_4  g11390(new_n13698, new_n13689, new_n13739);
or_5   g11391(new_n13739, new_n6001, new_n13740);
xnor_4 g11392(new_n13739, new_n6001, new_n13741);
xor_4  g11393(new_n13696, new_n13691, new_n13742);
or_5   g11394(new_n13742, new_n6006, new_n13743);
xnor_4 g11395(new_n13742, new_n6006, new_n13744);
xnor_4 g11396(n18578, n9090, new_n13745);
and_5  g11397(new_n13745, new_n6009, new_n13746);
or_5   g11398(new_n13746, new_n6013, new_n13747);
xnor_4 g11399(new_n13694, new_n13693, new_n13748);
nand_5 g11400(new_n13746, new_n5948, new_n13749);
and_5  g11401(new_n13749, new_n13747, new_n13750);
nand_5 g11402(new_n13750, new_n13748, new_n13751);
and_5  g11403(new_n13751, new_n13747, new_n13752);
or_5   g11404(new_n13752, new_n13744, new_n13753);
and_5  g11405(new_n13753, new_n13743, new_n13754_1);
or_5   g11406(new_n13754_1, new_n13741, new_n13755);
and_5  g11407(new_n13755, new_n13740, new_n13756);
or_5   g11408(new_n13756, new_n13738, new_n13757);
and_5  g11409(new_n13757, new_n13737, new_n13758);
nand_5 g11410(new_n13758, new_n13735, new_n13759);
and_5  g11411(new_n13759, new_n13734, new_n13760);
or_5   g11412(new_n13760, new_n13732, new_n13761);
and_5  g11413(new_n13761, new_n13731, new_n13762);
or_5   g11414(new_n13762, new_n13729, new_n13763);
and_5  g11415(new_n13763, new_n13728, new_n13764_1);
or_5   g11416(new_n13764_1, new_n13726, new_n13765);
and_5  g11417(new_n13765, new_n13725, new_n13766);
or_5   g11418(new_n13766, new_n13723, new_n13767);
and_5  g11419(new_n13767, new_n13722_1, new_n13768);
nor_5  g11420(new_n13768, new_n13720, new_n13769);
nor_5  g11421(new_n13769, new_n13718, new_n13770);
xor_4  g11422(new_n13768, new_n13720, new_n13771);
not_10 g11423(new_n13771, new_n13772);
and_5  g11424(new_n8347, n2743, new_n13773);
not_10 g11425(new_n13773, new_n13774);
nor_5  g11426(new_n3582_1, new_n3532, new_n13775_1);
not_10 g11427(new_n13775_1, new_n13776);
and_5  g11428(new_n13776, new_n13774, new_n13777);
not_10 g11429(new_n13777, new_n13778);
nor_5  g11430(new_n13778, new_n13772, new_n13779);
xor_4  g11431(new_n13778, new_n13772, new_n13780);
xor_4  g11432(new_n13766, new_n13723, new_n13781_1);
and_5  g11433(new_n13781_1, new_n3583, new_n13782);
xor_4  g11434(new_n13781_1, new_n3583, new_n13783_1);
xor_4  g11435(new_n13764_1, new_n13726, new_n13784);
and_5  g11436(new_n13784, new_n3602, new_n13785);
xor_4  g11437(new_n13784, new_n3602, new_n13786);
xor_4  g11438(new_n13762, new_n13729, new_n13787);
and_5  g11439(new_n13787, new_n3606, new_n13788);
xor_4  g11440(new_n13787, new_n3606, new_n13789);
xor_4  g11441(new_n13760, new_n13732, new_n13790);
and_5  g11442(new_n13790, new_n3610, new_n13791);
xor_4  g11443(new_n13790, new_n3610, new_n13792);
xor_4  g11444(new_n13758, new_n13735, new_n13793);
and_5  g11445(new_n13793, new_n3614, new_n13794);
xor_4  g11446(new_n13793, new_n3614, new_n13795);
xor_4  g11447(new_n13756, new_n13738, new_n13796);
nor_5  g11448(new_n13796, new_n3621, new_n13797);
xnor_4 g11449(new_n13796, new_n3619, new_n13798_1);
not_10 g11450(new_n13798_1, new_n13799);
xor_4  g11451(new_n13754_1, new_n13741, new_n13800);
or_5   g11452(new_n13800, new_n3646, new_n13801);
xnor_4 g11453(new_n13800, new_n3624, new_n13802);
not_10 g11454(new_n13802, new_n13803);
xor_4  g11455(new_n13752, new_n13744, new_n13804);
or_5   g11456(new_n13804, new_n3629, new_n13805);
xor_4  g11457(new_n13804, new_n3629, new_n13806);
not_10 g11458(new_n13806, new_n13807);
xor_4  g11459(new_n13750, new_n13748, new_n13808);
or_5   g11460(new_n13808, new_n3635, new_n13809);
xor_4  g11461(new_n13745, new_n6009, new_n13810);
not_10 g11462(new_n13810, new_n13811);
nor_5  g11463(new_n13811, new_n3638, new_n13812);
xor_4  g11464(new_n13808, new_n3635, new_n13813);
nand_5 g11465(new_n13813, new_n13812, new_n13814);
and_5  g11466(new_n13814, new_n13809, new_n13815);
or_5   g11467(new_n13815, new_n13807, new_n13816);
and_5  g11468(new_n13816, new_n13805, new_n13817);
or_5   g11469(new_n13817, new_n13803, new_n13818);
and_5  g11470(new_n13818, new_n13801, new_n13819);
nor_5  g11471(new_n13819, new_n13799, new_n13820);
nor_5  g11472(new_n13820, new_n13797, new_n13821);
not_10 g11473(new_n13821, new_n13822);
and_5  g11474(new_n13822, new_n13795, new_n13823);
nor_5  g11475(new_n13823, new_n13794, new_n13824);
not_10 g11476(new_n13824, new_n13825);
and_5  g11477(new_n13825, new_n13792, new_n13826);
nor_5  g11478(new_n13826, new_n13791, new_n13827);
not_10 g11479(new_n13827, new_n13828);
and_5  g11480(new_n13828, new_n13789, new_n13829);
nor_5  g11481(new_n13829, new_n13788, new_n13830);
not_10 g11482(new_n13830, new_n13831);
and_5  g11483(new_n13831, new_n13786, new_n13832);
nor_5  g11484(new_n13832, new_n13785, new_n13833);
not_10 g11485(new_n13833, new_n13834);
and_5  g11486(new_n13834, new_n13783_1, new_n13835_1);
nor_5  g11487(new_n13835_1, new_n13782, new_n13836);
not_10 g11488(new_n13836, new_n13837);
and_5  g11489(new_n13837, new_n13780, new_n13838);
nor_5  g11490(new_n13838, new_n13779, new_n13839);
xor_4  g11491(new_n13839, new_n13770, n2561);
xor_4  g11492(new_n8570, new_n8568, n2573);
xor_4  g11493(n18558, n10411, new_n13842);
or_5   g11494(new_n2657, n7149, new_n13843);
or_5   g11495(n16971, new_n2856, new_n13844);
and_5  g11496(new_n2862, n11503, new_n13845);
and_5  g11497(n14148, new_n10290, new_n13846);
not_10 g11498(new_n13846, new_n13847);
and_5  g11499(n18151, new_n13623, new_n13848);
and_5  g11500(new_n13848, new_n13847, new_n13849);
nor_5  g11501(new_n13849, new_n13845, new_n13850_1);
not_10 g11502(new_n13850_1, new_n13851_1);
nand_5 g11503(new_n13851_1, new_n13844, new_n13852);
and_5  g11504(new_n13852, new_n13843, new_n13853);
xor_4  g11505(new_n13853, new_n13842, new_n13854);
not_10 g11506(n6590, new_n13855);
or_5   g11507(n7963, new_n13855, new_n13856);
and_5  g11508(n7963, new_n13855, new_n13857);
not_10 g11509(n20349, new_n13858);
or_5   g11510(new_n13858, n10017, new_n13859);
and_5  g11511(new_n13858, n10017, new_n13860);
not_10 g11512(n3618, new_n13861);
and_5  g11513(n15936, new_n13861, new_n13862);
not_10 g11514(new_n13862, new_n13863);
or_5   g11515(new_n13863, new_n13860, new_n13864);
and_5  g11516(new_n13864, new_n13859, new_n13865);
or_5   g11517(new_n13865, new_n13857, new_n13866);
and_5  g11518(new_n13866, new_n13856, new_n13867);
xnor_4 g11519(new_n13867, new_n10134, new_n13868);
not_10 g11520(new_n13868, new_n13869);
xor_4  g11521(new_n13869, new_n13854, new_n13870);
xnor_4 g11522(n16971, n7149, new_n13871);
xor_4  g11523(new_n13871, new_n13851_1, new_n13872);
xor_4  g11524(new_n13865, new_n10138, new_n13873);
not_10 g11525(new_n13873, new_n13874);
or_5   g11526(new_n13874, new_n13872, new_n13875);
xor_4  g11527(new_n13874, new_n13872, new_n13876);
xnor_4 g11528(n18151, n1152, new_n13877);
nor_5  g11529(new_n13877, new_n10144, new_n13878);
not_10 g11530(new_n13878, new_n13879);
xnor_4 g11531(n14148, n11503, new_n13880);
xor_4  g11532(new_n13880, new_n13848, new_n13881);
nand_5 g11533(new_n13881, new_n13879, new_n13882);
xor_4  g11534(new_n13881, new_n13879, new_n13883);
not_10 g11535(new_n13883, new_n13884);
xor_4  g11536(new_n13863, new_n10141, new_n13885);
or_5   g11537(new_n13885, new_n13884, new_n13886);
and_5  g11538(new_n13886, new_n13882, new_n13887);
nand_5 g11539(new_n13887, new_n13876, new_n13888);
nand_5 g11540(new_n13888, new_n13875, new_n13889);
xor_4  g11541(new_n13889, new_n13870, new_n13890);
xnor_4 g11542(n19515, n17035, new_n13891);
not_10 g11543(new_n13891, new_n13892);
not_10 g11544(n22588, new_n13893);
or_5   g11545(new_n13893, n14684, new_n13894);
or_5   g11546(n22588, new_n4167, new_n13895);
and_5  g11547(n12209, new_n8593, new_n13896);
nor_5  g11548(n12209, new_n8593, new_n13897);
not_10 g11549(n24732, new_n13898);
and_5  g11550(new_n13898, n12892, new_n13899);
not_10 g11551(new_n13899, new_n13900);
nor_5  g11552(new_n13900, new_n13897, new_n13901);
nor_5  g11553(new_n13901, new_n13896, new_n13902);
not_10 g11554(new_n13902, new_n13903);
nand_5 g11555(new_n13903, new_n13895, new_n13904);
and_5  g11556(new_n13904, new_n13894, new_n13905);
xor_4  g11557(new_n13905, new_n13892, new_n13906);
not_10 g11558(new_n13906, new_n13907);
xor_4  g11559(new_n13907, new_n13890, new_n13908);
not_10 g11560(new_n13908, new_n13909);
xor_4  g11561(new_n13887, new_n13876, new_n13910);
xnor_4 g11562(n22588, n14684, new_n13911);
xor_4  g11563(new_n13911, new_n13903, new_n13912_1);
not_10 g11564(new_n13912_1, new_n13913);
or_5   g11565(new_n13913, new_n13910, new_n13914_1);
xor_4  g11566(n24732, n12892, new_n13915);
xor_4  g11567(new_n13877, new_n10144, new_n13916);
and_5  g11568(new_n13916, new_n13915, new_n13917);
xnor_4 g11569(n12209, n6631, new_n13918);
xnor_4 g11570(new_n13918, new_n13900, new_n13919);
not_10 g11571(new_n13919, new_n13920);
or_5   g11572(new_n13920, new_n13917, new_n13921);
xnor_4 g11573(new_n13919, new_n13917, new_n13922_1);
xor_4  g11574(new_n13885, new_n13884, new_n13923_1);
nand_5 g11575(new_n13923_1, new_n13922_1, new_n13924);
and_5  g11576(new_n13924, new_n13921, new_n13925);
xor_4  g11577(new_n13913, new_n13910, new_n13926);
not_10 g11578(new_n13926, new_n13927);
or_5   g11579(new_n13927, new_n13925, new_n13928);
and_5  g11580(new_n13928, new_n13914_1, new_n13929);
xnor_4 g11581(new_n13929, new_n13909, n2578);
not_10 g11582(new_n7975, new_n13931);
nand_5 g11583(new_n11978, new_n13931, new_n13932);
xor_4  g11584(new_n11978, new_n7975, new_n13933);
nand_5 g11585(new_n7975, new_n7907, new_n13934);
nand_5 g11586(new_n8048, new_n7976, new_n13935);
and_5  g11587(new_n13935, new_n13934, new_n13936);
or_5   g11588(new_n13936, new_n13933, new_n13937);
and_5  g11589(new_n13937, new_n13932, n2582);
xor_4  g11590(new_n4295, new_n4285, n2602);
nor_5  g11591(n22201, n2420, new_n13940);
and_5  g11592(new_n13940, new_n8236, new_n13941);
and_5  g11593(new_n13941, new_n8234, new_n13942);
and_5  g11594(new_n13942, new_n8230, new_n13943);
xor_4  g11595(new_n13943, new_n8226, new_n13944);
xor_4  g11596(new_n13944, new_n3971_1, new_n13945);
xor_4  g11597(new_n13942, new_n8230, new_n13946);
or_5   g11598(new_n13946, new_n3974, new_n13947);
xor_4  g11599(new_n13941, new_n8234, new_n13948);
nor_5  g11600(new_n13948, new_n3976, new_n13949);
not_10 g11601(new_n13949, new_n13950);
xor_4  g11602(new_n13948, new_n3976, new_n13951_1);
xor_4  g11603(new_n13940, new_n8236, new_n13952);
nand_5 g11604(new_n13952, new_n3981, new_n13953);
xor_4  g11605(new_n13952, new_n3981, new_n13954);
xor_4  g11606(n22201, n2420, new_n13955);
or_5   g11607(new_n13955, new_n3985, new_n13956);
and_5  g11608(new_n2554, n22201, new_n13957);
not_10 g11609(new_n13957, new_n13958);
xor_4  g11610(new_n13955, new_n3985, new_n13959);
nand_5 g11611(new_n13959, new_n13958, new_n13960);
and_5  g11612(new_n13960, new_n13956, new_n13961);
nand_5 g11613(new_n13961, new_n13954, new_n13962);
and_5  g11614(new_n13962, new_n13953, new_n13963);
and_5  g11615(new_n13963, new_n13951_1, new_n13964);
not_10 g11616(new_n13964, new_n13965);
and_5  g11617(new_n13965, new_n13950, new_n13966);
xnor_4 g11618(new_n13946, new_n3974, new_n13967);
or_5   g11619(new_n13967, new_n13966, new_n13968);
and_5  g11620(new_n13968, new_n13947, new_n13969);
xnor_4 g11621(new_n13969, new_n13945, new_n13970);
not_10 g11622(new_n13970, new_n13971);
xor_4  g11623(new_n8224, n7678, new_n13972);
or_5   g11624(new_n8228, n3785, new_n13973);
xor_4  g11625(new_n8228, n3785, new_n13974);
not_10 g11626(new_n13974, new_n13975);
or_5   g11627(new_n8232, n20250, new_n13976);
xor_4  g11628(new_n8232, n20250, new_n13977);
or_5   g11629(new_n8238, new_n4377, new_n13978);
nand_5 g11630(new_n8238, new_n4377, new_n13979);
and_5  g11631(new_n8243, new_n4382, new_n13980);
or_5   g11632(new_n2549, new_n4386, new_n13981);
xor_4  g11633(new_n8243, new_n4382, new_n13982);
and_5  g11634(new_n13982, new_n13981, new_n13983);
nor_5  g11635(new_n13983, new_n13980, new_n13984);
nand_5 g11636(new_n13984, new_n13979, new_n13985);
and_5  g11637(new_n13985, new_n13978, new_n13986);
nand_5 g11638(new_n13986, new_n13977, new_n13987);
and_5  g11639(new_n13987, new_n13976, new_n13988);
or_5   g11640(new_n13988, new_n13975, new_n13989);
and_5  g11641(new_n13989, new_n13973, new_n13990);
xor_4  g11642(new_n13990, new_n13972, new_n13991);
xor_4  g11643(new_n13991, new_n13971, new_n13992);
xor_4  g11644(new_n13988, new_n13975, new_n13993);
xor_4  g11645(new_n13967, new_n13966, new_n13994);
nand_5 g11646(new_n13994, new_n13993, new_n13995);
not_10 g11647(new_n13993, new_n13996);
xnor_4 g11648(new_n13994, new_n13996, new_n13997);
xor_4  g11649(new_n13963, new_n13951_1, new_n13998);
xor_4  g11650(new_n13986, new_n13977, new_n13999);
nand_5 g11651(new_n13999, new_n13998, new_n14000);
not_10 g11652(new_n13998, new_n14001);
xnor_4 g11653(new_n13999, new_n14001, new_n14002);
xor_4  g11654(new_n13961, new_n13954, new_n14003);
xor_4  g11655(new_n8238, new_n4377, new_n14004_1);
xor_4  g11656(new_n14004_1, new_n13984, new_n14005);
and_5  g11657(new_n14005, new_n14003, new_n14006);
xor_4  g11658(new_n13959, new_n13958, new_n14007);
xor_4  g11659(new_n13982, new_n13981, new_n14008);
nand_5 g11660(new_n14008, new_n14007, new_n14009);
xor_4  g11661(new_n2549, new_n4386, new_n14010);
xor_4  g11662(new_n2554, n22201, new_n14011);
and_5  g11663(new_n14011, new_n14010, new_n14012);
xor_4  g11664(new_n14008, new_n14007, new_n14013);
not_10 g11665(new_n14013, new_n14014);
or_5   g11666(new_n14014, new_n14012, new_n14015);
and_5  g11667(new_n14015, new_n14009, new_n14016);
xor_4  g11668(new_n14005, new_n14003, new_n14017);
and_5  g11669(new_n14017, new_n14016, new_n14018);
nor_5  g11670(new_n14018, new_n14006, new_n14019);
nand_5 g11671(new_n14019, new_n14002, new_n14020);
nand_5 g11672(new_n14020, new_n14000, new_n14021);
nand_5 g11673(new_n14021, new_n13997, new_n14022);
nand_5 g11674(new_n14022, new_n13995, new_n14023);
xnor_4 g11675(new_n14023, new_n13992, n2619);
nor_5  g11676(new_n5969, n12900, new_n14025);
xor_4  g11677(new_n5969, n12900, new_n14026);
not_10 g11678(new_n14026, new_n14027);
or_5   g11679(new_n5974, n20411, new_n14028);
xor_4  g11680(new_n5974, n20411, new_n14029);
not_10 g11681(new_n14029, new_n14030);
or_5   g11682(new_n5980_1, n17069, new_n14031);
xor_4  g11683(new_n5980_1, n17069, new_n14032);
not_10 g11684(new_n14032, new_n14033);
or_5   g11685(new_n5986, n15918, new_n14034);
nor_5  g11686(new_n5992, n17784, new_n14035);
not_10 g11687(new_n14035, new_n14036_1);
xor_4  g11688(new_n5992, n17784, new_n14037);
nand_5 g11689(new_n5998, n14323, new_n14038);
or_5   g11690(new_n13344, new_n13335, new_n14039);
and_5  g11691(new_n14039, new_n14038, new_n14040);
and_5  g11692(new_n14040, new_n14037, new_n14041);
not_10 g11693(new_n14041, new_n14042);
and_5  g11694(new_n14042, new_n14036_1, new_n14043);
xnor_4 g11695(new_n5986, n15918, new_n14044);
or_5   g11696(new_n14044, new_n14043, new_n14045);
and_5  g11697(new_n14045, new_n14034, new_n14046);
or_5   g11698(new_n14046, new_n14033, new_n14047);
and_5  g11699(new_n14047, new_n14031, new_n14048);
or_5   g11700(new_n14048, new_n14030, new_n14049);
and_5  g11701(new_n14049, new_n14028, new_n14050);
nor_5  g11702(new_n14050, new_n14027, new_n14051);
nor_5  g11703(new_n14051, new_n14025, new_n14052);
xor_4  g11704(new_n5922, n10650, new_n14053);
xnor_4 g11705(new_n14053, new_n14052, new_n14054);
not_10 g11706(new_n14054, new_n14055);
or_5   g11707(new_n14055, n6456, new_n14056);
xnor_4 g11708(new_n14055, n6456, new_n14057);
xor_4  g11709(new_n14050, new_n14027, new_n14058);
not_10 g11710(new_n14058, new_n14059_1);
or_5   g11711(new_n14059_1, n4085, new_n14060);
xnor_4 g11712(new_n14059_1, n4085, new_n14061);
xor_4  g11713(new_n14048, new_n14030, new_n14062);
not_10 g11714(new_n14062, new_n14063);
or_5   g11715(new_n14063, n26725, new_n14064);
xnor_4 g11716(new_n14063, n26725, new_n14065);
not_10 g11717(n11980, new_n14066);
xor_4  g11718(new_n14046, new_n14033, new_n14067);
nand_5 g11719(new_n14067, new_n14066, new_n14068);
xor_4  g11720(new_n14067, n11980, new_n14069);
not_10 g11721(n3253, new_n14070);
xor_4  g11722(new_n14044, new_n14043, new_n14071_1);
nand_5 g11723(new_n14071_1, new_n14070, new_n14072);
xor_4  g11724(new_n14071_1, new_n14070, new_n14073);
xor_4  g11725(new_n14040, new_n14037, new_n14074);
not_10 g11726(new_n14074, new_n14075);
and_5  g11727(new_n14075, n7759, new_n14076);
xnor_4 g11728(new_n14075, n7759, new_n14077);
nand_5 g11729(new_n13345, n12562, new_n14078);
nand_5 g11730(new_n13360, new_n13347, new_n14079);
and_5  g11731(new_n14079, new_n14078, new_n14080);
nor_5  g11732(new_n14080, new_n14077, new_n14081_1);
nor_5  g11733(new_n14081_1, new_n14076, new_n14082);
nand_5 g11734(new_n14082, new_n14073, new_n14083);
and_5  g11735(new_n14083, new_n14072, new_n14084);
or_5   g11736(new_n14084, new_n14069, new_n14085);
and_5  g11737(new_n14085, new_n14068, new_n14086);
or_5   g11738(new_n14086, new_n14065, new_n14087);
and_5  g11739(new_n14087, new_n14064, new_n14088);
or_5   g11740(new_n14088, new_n14061, new_n14089);
and_5  g11741(new_n14089, new_n14060, new_n14090_1);
or_5   g11742(new_n14090_1, new_n14057, new_n14091);
and_5  g11743(new_n14091, new_n14056, new_n14092);
not_10 g11744(new_n14052, new_n14093);
nor_5  g11745(new_n5922, n10650, new_n14094);
nor_5  g11746(new_n14094, new_n14093, new_n14095_1);
and_5  g11747(new_n5921, new_n5910, new_n14096);
and_5  g11748(new_n5922, n10650, new_n14097);
nor_5  g11749(new_n14097, new_n14096, new_n14098);
not_10 g11750(new_n14098, new_n14099);
nor_5  g11751(new_n14099, new_n14095_1, new_n14100);
and_5  g11752(new_n14100, new_n14092, new_n14101);
or_5   g11753(new_n14101, new_n13063, new_n14102);
xor_4  g11754(new_n14101, new_n13063, new_n14103);
not_10 g11755(new_n14103, new_n14104);
xor_4  g11756(new_n14100, new_n14092, new_n14105);
or_5   g11757(new_n14105, new_n13067, new_n14106);
xnor_4 g11758(new_n14105, new_n13066, new_n14107_1);
xor_4  g11759(new_n14090_1, new_n14057, new_n14108);
nand_5 g11760(new_n14108, new_n13072, new_n14109);
xor_4  g11761(new_n14108, new_n13072, new_n14110);
xor_4  g11762(new_n14088, new_n14061, new_n14111);
nand_5 g11763(new_n14111, new_n13077, new_n14112);
xor_4  g11764(new_n14111, new_n13077, new_n14113);
not_10 g11765(new_n13082_1, new_n14114);
xor_4  g11766(new_n14086, new_n14065, new_n14115);
nand_5 g11767(new_n14115, new_n14114, new_n14116);
xnor_4 g11768(new_n14115, new_n13082_1, new_n14117);
not_10 g11769(new_n14117, new_n14118);
xor_4  g11770(new_n14084, new_n14069, new_n14119);
nand_5 g11771(new_n14119, new_n13088, new_n14120);
xor_4  g11772(new_n14119, new_n13088, new_n14121_1);
not_10 g11773(new_n14073, new_n14122);
xnor_4 g11774(new_n14082, new_n14122, new_n14123);
not_10 g11775(new_n14123, new_n14124);
or_5   g11776(new_n14124, new_n13093, new_n14125);
xnor_4 g11777(new_n14123, new_n13093, new_n14126_1);
not_10 g11778(new_n14126_1, new_n14127);
xor_4  g11779(new_n14080, new_n14077, new_n14128);
or_5   g11780(new_n14128, new_n13099, new_n14129);
xor_4  g11781(new_n14128, new_n13099, new_n14130_1);
not_10 g11782(new_n14130_1, new_n14131);
or_5   g11783(new_n13361, new_n13105, new_n14132);
or_5   g11784(new_n13376, new_n13363, new_n14133);
and_5  g11785(new_n14133, new_n14132, new_n14134);
or_5   g11786(new_n14134, new_n14131, new_n14135);
and_5  g11787(new_n14135, new_n14129, new_n14136_1);
or_5   g11788(new_n14136_1, new_n14127, new_n14137);
nand_5 g11789(new_n14137, new_n14125, new_n14138);
nand_5 g11790(new_n14138, new_n14121_1, new_n14139);
and_5  g11791(new_n14139, new_n14120, new_n14140);
or_5   g11792(new_n14140, new_n14118, new_n14141);
nand_5 g11793(new_n14141, new_n14116, new_n14142);
nand_5 g11794(new_n14142, new_n14113, new_n14143);
nand_5 g11795(new_n14143, new_n14112, new_n14144);
nand_5 g11796(new_n14144, new_n14110, new_n14145);
nand_5 g11797(new_n14145, new_n14109, new_n14146);
nand_5 g11798(new_n14146, new_n14107_1, new_n14147_1);
and_5  g11799(new_n14147_1, new_n14106, new_n14148_1);
or_5   g11800(new_n14148_1, new_n14104, new_n14149);
and_5  g11801(new_n14149, new_n14102, n2661);
xnor_4 g11802(new_n11375_1, new_n11373, n2693);
xnor_4 g11803(new_n13854, new_n7338, new_n14152);
not_10 g11804(new_n14152, new_n14153);
or_5   g11805(new_n13872, new_n7344, new_n14154);
xnor_4 g11806(new_n13872, new_n7343, new_n14155);
not_10 g11807(new_n14155, new_n14156);
or_5   g11808(new_n13881, new_n7348, new_n14157);
nor_5  g11809(new_n13877, new_n7350, new_n14158);
xor_4  g11810(new_n13881, new_n7348, new_n14159);
nand_5 g11811(new_n14159, new_n14158, new_n14160);
and_5  g11812(new_n14160, new_n14157, new_n14161);
or_5   g11813(new_n14161, new_n14156, new_n14162);
and_5  g11814(new_n14162, new_n14154, new_n14163);
xor_4  g11815(new_n14163, new_n14153, new_n14164);
not_10 g11816(new_n14164, new_n14165);
xor_4  g11817(n8309, n4665, new_n14166);
or_5   g11818(new_n10286, n19005, new_n14167);
or_5   g11819(n19144, new_n2858_1, new_n14168);
and_5  g11820(n12593, new_n2860_1, new_n14169);
and_5  g11821(new_n10288, n4326, new_n14170);
not_10 g11822(new_n14170, new_n14171);
and_5  g11823(n13714, new_n2865, new_n14172);
and_5  g11824(new_n14172, new_n14171, new_n14173);
nor_5  g11825(new_n14173, new_n14169, new_n14174_1);
not_10 g11826(new_n14174_1, new_n14175);
nand_5 g11827(new_n14175, new_n14168, new_n14176);
and_5  g11828(new_n14176, new_n14167, new_n14177);
xor_4  g11829(new_n14177, new_n14166, new_n14178);
xor_4  g11830(new_n14178, new_n14165, new_n14179);
xor_4  g11831(new_n14161, new_n14156, new_n14180);
not_10 g11832(new_n14180, new_n14181);
xnor_4 g11833(n19144, n19005, new_n14182);
xor_4  g11834(new_n14182, new_n14175, new_n14183);
and_5  g11835(new_n14183, new_n14181, new_n14184);
not_10 g11836(new_n14184, new_n14185);
xor_4  g11837(new_n14183, new_n14181, new_n14186);
xor_4  g11838(n13714, n5438, new_n14187);
xor_4  g11839(new_n13877, new_n7350, new_n14188);
and_5  g11840(new_n14188, new_n14187, new_n14189);
not_10 g11841(new_n14189, new_n14190_1);
xnor_4 g11842(n12593, n4326, new_n14191);
xor_4  g11843(new_n14191, new_n14172, new_n14192);
and_5  g11844(new_n14192, new_n14190_1, new_n14193);
xor_4  g11845(new_n14159, new_n14158, new_n14194);
not_10 g11846(new_n14194, new_n14195);
xor_4  g11847(new_n14192, new_n14190_1, new_n14196);
and_5  g11848(new_n14196, new_n14195, new_n14197);
nor_5  g11849(new_n14197, new_n14193, new_n14198);
not_10 g11850(new_n14198, new_n14199);
and_5  g11851(new_n14199, new_n14186, new_n14200);
not_10 g11852(new_n14200, new_n14201);
and_5  g11853(new_n14201, new_n14185, new_n14202);
xor_4  g11854(new_n14202, new_n14179, n2703);
xnor_4 g11855(new_n13208, new_n13195, n2706);
and_5  g11856(new_n6236, n1831, new_n14205);
xnor_4 g11857(n3320, n1831, new_n14206);
not_10 g11858(new_n14206, new_n14207);
not_10 g11859(n13137, new_n14208);
or_5   g11860(new_n14208, n1288, new_n14209);
xnor_4 g11861(n13137, n1288, new_n14210);
not_10 g11862(new_n14210, new_n14211_1);
not_10 g11863(n18452, new_n14212);
or_5   g11864(new_n14212, n1752, new_n14213);
xnor_4 g11865(n18452, n1752, new_n14214);
not_10 g11866(new_n14214, new_n14215);
not_10 g11867(n21317, new_n14216);
or_5   g11868(new_n14216, n13110, new_n14217);
xor_4  g11869(n21317, n13110, new_n14218);
or_5   g11870(n25694, new_n4000_1, new_n14219);
xor_4  g11871(n25694, n12398, new_n14220);
or_5   g11872(new_n4001, n15424, new_n14221);
xnor_4 g11873(n19789, n15424, new_n14222_1);
or_5   g11874(n20169, new_n4012, new_n14223);
or_5   g11875(new_n12445, new_n12432, new_n14224);
and_5  g11876(new_n14224, new_n14223, new_n14225);
nand_5 g11877(new_n14225, new_n14222_1, new_n14226);
and_5  g11878(new_n14226, new_n14221, new_n14227);
or_5   g11879(new_n14227, new_n14220, new_n14228);
and_5  g11880(new_n14228, new_n14219, new_n14229);
or_5   g11881(new_n14229, new_n14218, new_n14230_1);
and_5  g11882(new_n14230_1, new_n14217, new_n14231);
or_5   g11883(new_n14231, new_n14215, new_n14232);
and_5  g11884(new_n14232, new_n14213, new_n14233);
or_5   g11885(new_n14233, new_n14211_1, new_n14234);
and_5  g11886(new_n14234, new_n14209, new_n14235);
nor_5  g11887(new_n14235, new_n14207, new_n14236);
nor_5  g11888(new_n14236, new_n14205, new_n14237);
not_10 g11889(n19539, new_n14238);
and_5  g11890(new_n14238, n1483, new_n14239);
not_10 g11891(new_n14239, new_n14240);
nor_5  g11892(new_n11480, new_n11464, new_n14241);
not_10 g11893(new_n14241, new_n14242);
and_5  g11894(new_n14242, new_n14240, new_n14243);
not_10 g11895(new_n11481_1, new_n14244);
and_5  g11896(new_n6509, new_n6500, new_n14245);
and_5  g11897(new_n14245, new_n12604, new_n14246);
xor_4  g11898(new_n14246, new_n12601, new_n14247);
not_10 g11899(new_n14247, new_n14248);
and_5  g11900(new_n14248, new_n12551, new_n14249);
xor_4  g11901(new_n14248, new_n12551, new_n14250);
xor_4  g11902(new_n14245, new_n12604, new_n14251);
not_10 g11903(new_n14251, new_n14252);
or_5   g11904(new_n14252, new_n12555, new_n14253);
and_5  g11905(new_n14252, new_n12555, new_n14254);
not_10 g11906(new_n6550, new_n14255);
nor_5  g11907(new_n14255, new_n6513_1, new_n14256);
nor_5  g11908(new_n14256, new_n6512, new_n14257);
or_5   g11909(new_n14257, new_n14254, new_n14258);
and_5  g11910(new_n14258, new_n14253, new_n14259);
and_5  g11911(new_n14259, new_n14250, new_n14260);
or_5   g11912(new_n14260, new_n14249, new_n14261);
not_10 g11913(n5140, new_n14262);
not_10 g11914(n10018, new_n14263);
and_5  g11915(new_n14246, new_n12601, new_n14264);
xor_4  g11916(new_n14264, new_n14263, new_n14265);
not_10 g11917(new_n14265, new_n14266);
xor_4  g11918(new_n14266, new_n14262, new_n14267_1);
xor_4  g11919(new_n14267_1, new_n14261, new_n14268);
and_5  g11920(new_n14268, new_n14244, new_n14269);
xnor_4 g11921(new_n14268, new_n14244, new_n14270);
not_10 g11922(new_n11547, new_n14271_1);
xor_4  g11923(new_n14259, new_n14250, new_n14272);
nand_5 g11924(new_n14272, new_n14271_1, new_n14273);
xor_4  g11925(new_n14272, new_n14271_1, new_n14274);
xor_4  g11926(new_n14252, n3349, new_n14275_1);
xor_4  g11927(new_n14275_1, new_n14257, new_n14276);
nand_5 g11928(new_n14276, new_n11552, new_n14277_1);
xnor_4 g11929(new_n14276, new_n11552, new_n14278);
or_5   g11930(new_n6551, new_n6498, new_n14279);
or_5   g11931(new_n6592, new_n6552, new_n14280);
and_5  g11932(new_n14280, new_n14279, new_n14281);
or_5   g11933(new_n14281, new_n14278, new_n14282);
and_5  g11934(new_n14282, new_n14277_1, new_n14283);
nand_5 g11935(new_n14283, new_n14274, new_n14284);
and_5  g11936(new_n14284, new_n14273, new_n14285);
nor_5  g11937(new_n14285, new_n14270, new_n14286);
or_5   g11938(new_n14286, new_n14269, new_n14287);
nand_5 g11939(new_n14264, new_n14263, new_n14288);
and_5  g11940(new_n14266, new_n14262, new_n14289);
or_5   g11941(new_n14266, new_n14262, new_n14290);
and_5  g11942(new_n14290, new_n14261, new_n14291);
or_5   g11943(new_n14291, new_n14289, new_n14292);
and_5  g11944(new_n14292, new_n14288, new_n14293);
nor_5  g11945(new_n14293, new_n14287, new_n14294_1);
and_5  g11946(new_n14294_1, new_n14243, new_n14295);
and_5  g11947(new_n14293, new_n14287, new_n14296);
not_10 g11948(new_n14296, new_n14297);
nor_5  g11949(new_n14297, new_n14243, new_n14298);
nor_5  g11950(new_n14298, new_n14295, new_n14299);
not_10 g11951(new_n14299, new_n14300);
xnor_4 g11952(new_n14300, new_n14237, new_n14301);
xor_4  g11953(new_n14293, new_n14287, new_n14302);
xnor_4 g11954(new_n14302, new_n14243, new_n14303);
and_5  g11955(new_n14303, new_n14237, new_n14304);
nor_5  g11956(new_n14303, new_n14237, new_n14305);
not_10 g11957(new_n14305, new_n14306);
xor_4  g11958(new_n14235, new_n14207, new_n14307);
not_10 g11959(new_n14307, new_n14308);
xor_4  g11960(new_n14285, new_n14270, new_n14309);
and_5  g11961(new_n14309, new_n14308, new_n14310_1);
xor_4  g11962(new_n14309, new_n14308, new_n14311);
not_10 g11963(new_n14311, new_n14312);
xor_4  g11964(new_n14233, new_n14211_1, new_n14313);
not_10 g11965(new_n14313, new_n14314);
xor_4  g11966(new_n14283, new_n14274, new_n14315);
and_5  g11967(new_n14315, new_n14314, new_n14316);
xor_4  g11968(new_n14315, new_n14314, new_n14317);
not_10 g11969(new_n14317, new_n14318);
xor_4  g11970(new_n14231, new_n14215, new_n14319);
xor_4  g11971(new_n14281, new_n14278, new_n14320);
nor_5  g11972(new_n14320, new_n14319, new_n14321);
xor_4  g11973(new_n14320, new_n14319, new_n14322);
not_10 g11974(new_n14322, new_n14323_1);
xor_4  g11975(new_n14229, new_n14218, new_n14324);
nor_5  g11976(new_n14324, new_n6593, new_n14325);
xor_4  g11977(new_n14227, new_n14220, new_n14326_1);
nor_5  g11978(new_n14326_1, new_n6595, new_n14327);
xor_4  g11979(new_n14326_1, new_n6595, new_n14328);
not_10 g11980(new_n14328, new_n14329);
xor_4  g11981(new_n14225, new_n14222_1, new_n14330);
nor_5  g11982(new_n14330, new_n6600, new_n14331);
xor_4  g11983(new_n14330, new_n6600, new_n14332);
and_5  g11984(new_n12446_1, new_n6605, new_n14333);
not_10 g11985(new_n12464, new_n14334);
and_5  g11986(new_n14334, new_n12447, new_n14335);
nor_5  g11987(new_n14335, new_n14333, new_n14336);
not_10 g11988(new_n14336, new_n14337);
and_5  g11989(new_n14337, new_n14332, new_n14338);
nor_5  g11990(new_n14338, new_n14331, new_n14339);
nor_5  g11991(new_n14339, new_n14329, new_n14340);
nor_5  g11992(new_n14340, new_n14327, new_n14341);
xor_4  g11993(new_n14324, new_n6593, new_n14342_1);
not_10 g11994(new_n14342_1, new_n14343);
nor_5  g11995(new_n14343, new_n14341, new_n14344);
nor_5  g11996(new_n14344, new_n14325, new_n14345_1);
nor_5  g11997(new_n14345_1, new_n14323_1, new_n14346);
nor_5  g11998(new_n14346, new_n14321, new_n14347);
nor_5  g11999(new_n14347, new_n14318, new_n14348);
nor_5  g12000(new_n14348, new_n14316, new_n14349);
nor_5  g12001(new_n14349, new_n14312, new_n14350);
nor_5  g12002(new_n14350, new_n14310_1, new_n14351);
and_5  g12003(new_n14351, new_n14306, new_n14352);
nor_5  g12004(new_n14352, new_n14304, new_n14353_1);
xor_4  g12005(new_n14353_1, new_n14301, n2711);
xor_4  g12006(n10611, n2680, new_n14355);
or_5   g12007(n2783, new_n9298, new_n14356);
or_5   g12008(new_n9328, n1667, new_n14357);
and_5  g12009(new_n9330, n7339, new_n14358);
nor_5  g12010(new_n9330, n7339, new_n14359);
not_10 g12011(new_n14359, new_n14360);
and_5  g12012(n26808, new_n9333, new_n14361);
and_5  g12013(new_n14361, new_n14360, new_n14362);
nor_5  g12014(new_n14362, new_n14358, new_n14363);
not_10 g12015(new_n14363, new_n14364_1);
nand_5 g12016(new_n14364_1, new_n14357, new_n14365);
and_5  g12017(new_n14365, new_n14356, new_n14366);
xor_4  g12018(new_n14366, new_n14355, new_n14367);
xnor_4 g12019(new_n14367, new_n9237, new_n14368);
xnor_4 g12020(n2783, n1667, new_n14369);
xor_4  g12021(new_n14369, new_n14364_1, new_n14370);
nand_5 g12022(new_n14370, new_n9241, new_n14371);
xnor_4 g12023(new_n14370, new_n9245, new_n14372);
xnor_4 g12024(n26808, n18, new_n14373);
nor_5  g12025(new_n14373, new_n9249, new_n14374);
xnor_4 g12026(n15490, n7339, new_n14375_1);
xnor_4 g12027(new_n14375_1, new_n14361, new_n14376);
or_5   g12028(new_n14376, new_n14374, new_n14377);
xor_4  g12029(new_n14376, new_n14374, new_n14378);
nand_5 g12030(new_n14378, new_n9255, new_n14379);
nand_5 g12031(new_n14379, new_n14377, new_n14380);
nand_5 g12032(new_n14380, new_n14372, new_n14381);
nand_5 g12033(new_n14381, new_n14371, new_n14382);
xnor_4 g12034(new_n14382, new_n14368, n2761);
xnor_4 g12035(n25120, n8526, new_n14384);
or_5   g12036(n8363, n2816, new_n14385);
xnor_4 g12037(n8363, n2816, new_n14386);
or_5   g12038(n20359, n14680, new_n14387);
xnor_4 g12039(n20359, n14680, new_n14388);
or_5   g12040(n17250, n4409, new_n14389);
or_5   g12041(new_n9554_1, new_n9532, new_n14390);
and_5  g12042(new_n14390, new_n14389, new_n14391);
or_5   g12043(new_n14391, new_n14388, new_n14392);
and_5  g12044(new_n14392, new_n14387, new_n14393);
or_5   g12045(new_n14393, new_n14386, new_n14394);
and_5  g12046(new_n14394, new_n14385, new_n14395);
xor_4  g12047(new_n14395, new_n14384, new_n14396);
and_5  g12048(new_n14396, new_n7250, new_n14397);
xor_4  g12049(new_n14396, new_n7250, new_n14398);
xor_4  g12050(new_n14393, new_n14386, new_n14399);
or_5   g12051(new_n14399, new_n11171, new_n14400);
xor_4  g12052(new_n14391, new_n14388, new_n14401);
nand_5 g12053(new_n14401, new_n11175, new_n14402);
xor_4  g12054(new_n14401, new_n11175, new_n14403);
or_5   g12055(new_n9555, new_n11179, new_n14404);
xor_4  g12056(new_n9555, new_n11179, new_n14405);
not_10 g12057(new_n14405, new_n14406);
or_5   g12058(new_n9558_1, new_n11183, new_n14407);
xor_4  g12059(new_n9558_1, new_n11183, new_n14408);
not_10 g12060(new_n14408, new_n14409);
or_5   g12061(new_n9562, new_n11187, new_n14410);
xor_4  g12062(new_n9562, new_n11187, new_n14411);
not_10 g12063(new_n14411, new_n14412_1);
or_5   g12064(new_n9566, new_n11190, new_n14413);
xor_4  g12065(new_n9566, new_n11190, new_n14414_1);
not_10 g12066(new_n14414_1, new_n14415);
or_5   g12067(new_n9570, new_n7268_1, new_n14416);
and_5  g12068(new_n9572, new_n7272, new_n14417);
and_5  g12069(new_n9574, n8581, new_n14418);
not_10 g12070(new_n14418, new_n14419);
xor_4  g12071(new_n9572, new_n7272, new_n14420);
and_5  g12072(new_n14420, new_n14419, new_n14421);
nor_5  g12073(new_n14421, new_n14417, new_n14422);
xor_4  g12074(new_n9570, new_n7268_1, new_n14423);
nand_5 g12075(new_n14423, new_n14422, new_n14424);
and_5  g12076(new_n14424, new_n14416, new_n14425);
or_5   g12077(new_n14425, new_n14415, new_n14426);
and_5  g12078(new_n14426, new_n14413, new_n14427);
or_5   g12079(new_n14427, new_n14412_1, new_n14428);
and_5  g12080(new_n14428, new_n14410, new_n14429);
or_5   g12081(new_n14429, new_n14409, new_n14430);
and_5  g12082(new_n14430, new_n14407, new_n14431);
or_5   g12083(new_n14431, new_n14406, new_n14432);
and_5  g12084(new_n14432, new_n14404, new_n14433);
nand_5 g12085(new_n14433, new_n14403, new_n14434);
and_5  g12086(new_n14434, new_n14402, new_n14435);
xor_4  g12087(new_n14399, new_n11171, new_n14436);
nand_5 g12088(new_n14436, new_n14435, new_n14437);
and_5  g12089(new_n14437, new_n14400, new_n14438);
and_5  g12090(new_n14438, new_n14398, new_n14439);
nor_5  g12091(new_n14439, new_n14397, new_n14440_1);
nor_5  g12092(n25120, n8526, new_n14441);
nor_5  g12093(new_n14395, new_n14384, new_n14442);
nor_5  g12094(new_n14442, new_n14441, new_n14443);
and_5  g12095(new_n14443, new_n14440_1, new_n14444);
not_10 g12096(n11898, new_n14445);
not_10 g12097(n19941, new_n14446);
not_10 g12098(n1099, new_n14447);
and_5  g12099(new_n3734, new_n3725_1, new_n14448);
and_5  g12100(new_n14448, new_n14447, new_n14449);
and_5  g12101(new_n14449, new_n14446, new_n14450);
xor_4  g12102(new_n14450, new_n14445, new_n14451);
nor_5  g12103(new_n14451, new_n4856, new_n14452);
not_10 g12104(new_n14452, new_n14453);
xor_4  g12105(new_n14451, new_n4857, new_n14454);
xor_4  g12106(new_n14449, new_n14446, new_n14455);
or_5   g12107(new_n14455, new_n4861, new_n14456);
xnor_4 g12108(new_n14455, new_n4862, new_n14457_1);
not_10 g12109(new_n14457_1, new_n14458);
xor_4  g12110(new_n14448, new_n14447, new_n14459);
or_5   g12111(new_n14459, new_n4865, new_n14460);
xor_4  g12112(new_n14459, new_n4866, new_n14461);
or_5   g12113(new_n4869, new_n3735, new_n14462);
xnor_4 g12114(new_n4870, new_n3735, new_n14463);
not_10 g12115(new_n14463, new_n14464_1);
or_5   g12116(new_n4873, new_n3737, new_n14465);
xor_4  g12117(new_n4873, new_n3737, new_n14466);
not_10 g12118(new_n14466, new_n14467);
or_5   g12119(new_n4876, new_n3741, new_n14468);
xor_4  g12120(new_n4876, new_n3741, new_n14469);
not_10 g12121(new_n14469, new_n14470);
or_5   g12122(new_n4879, new_n3745, new_n14471_1);
xnor_4 g12123(new_n4880, new_n3745, new_n14472);
or_5   g12124(new_n4883, new_n3747, new_n14473);
xnor_4 g12125(new_n4884, new_n3747, new_n14474);
not_10 g12126(n25435, new_n14475_1);
and_5  g12127(new_n4890, new_n14475_1, new_n14476);
not_10 g12128(new_n14476, new_n14477);
or_5   g12129(new_n14477, n13319, new_n14478);
nand_5 g12130(new_n14477, new_n3751, new_n14479);
and_5  g12131(new_n14479, new_n14478, new_n14480);
nand_5 g12132(new_n14480, new_n4888, new_n14481);
nand_5 g12133(new_n14481, new_n14478, new_n14482);
nand_5 g12134(new_n14482, new_n14474, new_n14483);
nand_5 g12135(new_n14483, new_n14473, new_n14484);
nand_5 g12136(new_n14484, new_n14472, new_n14485);
and_5  g12137(new_n14485, new_n14471_1, new_n14486);
or_5   g12138(new_n14486, new_n14470, new_n14487);
and_5  g12139(new_n14487, new_n14468, new_n14488);
or_5   g12140(new_n14488, new_n14467, new_n14489);
and_5  g12141(new_n14489, new_n14465, new_n14490);
or_5   g12142(new_n14490, new_n14464_1, new_n14491);
and_5  g12143(new_n14491, new_n14462, new_n14492);
or_5   g12144(new_n14492, new_n14461, new_n14493);
and_5  g12145(new_n14493, new_n14460, new_n14494);
or_5   g12146(new_n14494, new_n14458, new_n14495);
and_5  g12147(new_n14495, new_n14456, new_n14496);
nor_5  g12148(new_n14496, new_n14454, new_n14497);
not_10 g12149(new_n14497, new_n14498);
and_5  g12150(new_n14498, new_n14453, new_n14499);
and_5  g12151(new_n14450, new_n14445, new_n14500);
not_10 g12152(new_n14500, new_n14501);
nor_5  g12153(new_n14501, new_n4916, new_n14502);
and_5  g12154(new_n14502, new_n14499, new_n14503);
and_5  g12155(new_n14501, new_n4916, new_n14504);
not_10 g12156(new_n14504, new_n14505);
nor_5  g12157(new_n14505, new_n14499, new_n14506);
nor_5  g12158(new_n14506, new_n14503, new_n14507);
nand_5 g12159(new_n14507, new_n14444, new_n14508);
or_5   g12160(new_n14507, new_n14444, new_n14509);
xor_4  g12161(new_n14443, new_n14440_1, new_n14510_1);
xor_4  g12162(new_n14500, new_n4916, new_n14511);
xor_4  g12163(new_n14511, new_n14499, new_n14512);
nor_5  g12164(new_n14512, new_n14510_1, new_n14513);
not_10 g12165(new_n14510_1, new_n14514);
xnor_4 g12166(new_n14512, new_n14514, new_n14515);
xor_4  g12167(new_n14438, new_n14398, new_n14516);
xor_4  g12168(new_n14496, new_n14454, new_n14517);
and_5  g12169(new_n14517, new_n14516, new_n14518);
xor_4  g12170(new_n14517, new_n14516, new_n14519);
not_10 g12171(new_n14519, new_n14520);
xor_4  g12172(new_n14494, new_n14458, new_n14521);
not_10 g12173(new_n14521, new_n14522);
xor_4  g12174(new_n14436, new_n14435, new_n14523);
nor_5  g12175(new_n14523, new_n14522, new_n14524);
not_10 g12176(new_n14524, new_n14525);
xor_4  g12177(new_n14523, new_n14522, new_n14526);
xor_4  g12178(new_n14433, new_n14403, new_n14527);
xor_4  g12179(new_n14492, new_n14461, new_n14528);
and_5  g12180(new_n14528, new_n14527, new_n14529);
xor_4  g12181(new_n14528, new_n14527, new_n14530);
not_10 g12182(new_n14530, new_n14531);
xnor_4 g12183(new_n14490, new_n14463, new_n14532);
not_10 g12184(new_n14532, new_n14533);
xor_4  g12185(new_n14431, new_n14406, new_n14534);
nor_5  g12186(new_n14534, new_n14533, new_n14535);
not_10 g12187(new_n14535, new_n14536);
xor_4  g12188(new_n14534, new_n14533, new_n14537);
xor_4  g12189(new_n14488, new_n14467, new_n14538);
not_10 g12190(new_n14538, new_n14539);
xor_4  g12191(new_n14429, new_n14409, new_n14540);
nor_5  g12192(new_n14540, new_n14539, new_n14541_1);
xnor_4 g12193(new_n14540, new_n14538, new_n14542);
not_10 g12194(new_n14542, new_n14543);
xor_4  g12195(new_n14486, new_n14470, new_n14544);
not_10 g12196(new_n14544, new_n14545);
xor_4  g12197(new_n14427, new_n14412_1, new_n14546_1);
nor_5  g12198(new_n14546_1, new_n14545, new_n14547_1);
xnor_4 g12199(new_n14546_1, new_n14544, new_n14548);
not_10 g12200(new_n14548, new_n14549);
xor_4  g12201(new_n14484, new_n14472, new_n14550);
not_10 g12202(new_n14550, new_n14551);
xor_4  g12203(new_n14425, new_n14415, new_n14552);
nor_5  g12204(new_n14552, new_n14551, new_n14553);
not_10 g12205(new_n14553, new_n14554);
xor_4  g12206(new_n14552, new_n14551, new_n14555);
xnor_4 g12207(new_n14482, new_n14474, new_n14556);
xor_4  g12208(new_n14423, new_n14422, new_n14557);
and_5  g12209(new_n14557, new_n14556, new_n14558);
xor_4  g12210(new_n14557, new_n14556, new_n14559);
xor_4  g12211(new_n14420, new_n14419, new_n14560);
xnor_4 g12212(new_n14480, new_n4887, new_n14561);
nand_5 g12213(new_n14561, new_n14560, new_n14562);
xor_4  g12214(new_n9574, n8581, new_n14563);
not_10 g12215(new_n14563, new_n14564);
xor_4  g12216(new_n4890, new_n14475_1, new_n14565);
nor_5  g12217(new_n14565, new_n14564, new_n14566);
not_10 g12218(new_n14566, new_n14567);
xor_4  g12219(new_n14561, new_n14560, new_n14568);
nand_5 g12220(new_n14568, new_n14567, new_n14569);
and_5  g12221(new_n14569, new_n14562, new_n14570_1);
and_5  g12222(new_n14570_1, new_n14559, new_n14571);
nor_5  g12223(new_n14571, new_n14558, new_n14572);
and_5  g12224(new_n14572, new_n14555, new_n14573);
not_10 g12225(new_n14573, new_n14574);
and_5  g12226(new_n14574, new_n14554, new_n14575_1);
nor_5  g12227(new_n14575_1, new_n14549, new_n14576_1);
nor_5  g12228(new_n14576_1, new_n14547_1, new_n14577);
nor_5  g12229(new_n14577, new_n14543, new_n14578);
nor_5  g12230(new_n14578, new_n14541_1, new_n14579);
not_10 g12231(new_n14579, new_n14580);
and_5  g12232(new_n14580, new_n14537, new_n14581);
not_10 g12233(new_n14581, new_n14582);
and_5  g12234(new_n14582, new_n14536, new_n14583);
nor_5  g12235(new_n14583, new_n14531, new_n14584);
nor_5  g12236(new_n14584, new_n14529, new_n14585);
not_10 g12237(new_n14585, new_n14586);
and_5  g12238(new_n14586, new_n14526, new_n14587);
not_10 g12239(new_n14587, new_n14588);
and_5  g12240(new_n14588, new_n14525, new_n14589);
nor_5  g12241(new_n14589, new_n14520, new_n14590);
nor_5  g12242(new_n14590, new_n14518, new_n14591);
not_10 g12243(new_n14591, new_n14592);
and_5  g12244(new_n14592, new_n14515, new_n14593_1);
nor_5  g12245(new_n14593_1, new_n14513, new_n14594);
and_5  g12246(new_n14594, new_n14509, new_n14595);
nor_5  g12247(new_n14595, new_n14503, new_n14596);
and_5  g12248(new_n14596, new_n14508, n2774);
and_5  g12249(new_n9634, new_n7798, new_n14598);
and_5  g12250(new_n14598, new_n7795, new_n14599);
and_5  g12251(new_n14599, new_n7792, new_n14600);
and_5  g12252(new_n14600, new_n7789, new_n14601);
and_5  g12253(new_n14601, new_n7785, new_n14602);
xor_4  g12254(new_n14602, new_n7782, new_n14603_1);
xor_4  g12255(new_n14603_1, new_n4923, new_n14604);
xor_4  g12256(new_n14601, new_n7785, new_n14605);
nor_5  g12257(new_n14605, n2659, new_n14606);
xor_4  g12258(new_n14605, new_n4927, new_n14607);
xor_4  g12259(new_n14600, new_n7789, new_n14608);
or_5   g12260(new_n14608, n24327, new_n14609);
xor_4  g12261(new_n14608, new_n4931, new_n14610);
xor_4  g12262(new_n14599, new_n7792, new_n14611);
or_5   g12263(new_n14611, n22198, new_n14612);
xor_4  g12264(new_n14598, new_n7795, new_n14613);
nand_5 g12265(new_n14613, n20826, new_n14614);
xor_4  g12266(new_n14613, new_n4939_1, new_n14615);
nand_5 g12267(new_n9635_1, n7305, new_n14616);
or_5   g12268(new_n9648_1, new_n9637, new_n14617);
and_5  g12269(new_n14617, new_n14616, new_n14618);
or_5   g12270(new_n14618, new_n14615, new_n14619);
and_5  g12271(new_n14619, new_n14614, new_n14620);
xor_4  g12272(new_n14611, n22198, new_n14621);
nand_5 g12273(new_n14621, new_n14620, new_n14622);
and_5  g12274(new_n14622, new_n14612, new_n14623);
or_5   g12275(new_n14623, new_n14610, new_n14624);
and_5  g12276(new_n14624, new_n14609, new_n14625);
nor_5  g12277(new_n14625, new_n14607, new_n14626);
nor_5  g12278(new_n14626, new_n14606, new_n14627);
xor_4  g12279(new_n14627, new_n14604, new_n14628);
xor_4  g12280(new_n14628, new_n3475, new_n14629);
xor_4  g12281(new_n14625, new_n14607, new_n14630);
or_5   g12282(new_n14630, new_n3480_1, new_n14631);
xor_4  g12283(new_n14623, new_n14610, new_n14632);
and_5  g12284(new_n14632, new_n3485, new_n14633_1);
xnor_4 g12285(new_n14632, new_n3485, new_n14634);
xor_4  g12286(new_n14621, new_n14620, new_n14635);
nand_5 g12287(new_n14635, new_n3490, new_n14636_1);
xnor_4 g12288(new_n14635, new_n3490, new_n14637);
xor_4  g12289(new_n14618, new_n14615, new_n14638);
or_5   g12290(new_n14638, new_n3495, new_n14639);
xnor_4 g12291(new_n14638, new_n3494, new_n14640);
or_5   g12292(new_n9650, new_n3500, new_n14641);
xnor_4 g12293(new_n9649, new_n3500, new_n14642);
not_10 g12294(new_n14642, new_n14643);
nand_5 g12295(new_n9668, new_n3504, new_n14644);
xnor_4 g12296(new_n9668, new_n3503, new_n14645);
not_10 g12297(new_n14645, new_n14646);
nand_5 g12298(new_n9672, new_n3508, new_n14647);
and_5  g12299(new_n9675, new_n3510, new_n14648);
xnor_4 g12300(new_n9673, new_n3508, new_n14649);
nand_5 g12301(new_n14649, new_n14648, new_n14650);
and_5  g12302(new_n14650, new_n14647, new_n14651);
or_5   g12303(new_n14651, new_n14646, new_n14652);
and_5  g12304(new_n14652, new_n14644, new_n14653);
or_5   g12305(new_n14653, new_n14643, new_n14654);
and_5  g12306(new_n14654, new_n14641, new_n14655);
nand_5 g12307(new_n14655, new_n14640, new_n14656);
and_5  g12308(new_n14656, new_n14639, new_n14657);
or_5   g12309(new_n14657, new_n14637, new_n14658);
and_5  g12310(new_n14658, new_n14636_1, new_n14659);
nor_5  g12311(new_n14659, new_n14634, new_n14660);
nor_5  g12312(new_n14660, new_n14633_1, new_n14661);
xor_4  g12313(new_n14630, new_n3480_1, new_n14662);
nand_5 g12314(new_n14662, new_n14661, new_n14663);
and_5  g12315(new_n14663, new_n14631, new_n14664);
xor_4  g12316(new_n14664, new_n14629, new_n14665);
not_10 g12317(new_n14665, new_n14666);
xor_4  g12318(new_n3603, new_n3533, new_n14667);
and_5  g12319(new_n3607, n13719, new_n14668);
nor_5  g12320(new_n3607, n13719, new_n14669);
nor_5  g12321(new_n3611, n442, new_n14670);
xor_4  g12322(new_n3611, n442, new_n14671);
not_10 g12323(new_n14671, new_n14672);
or_5   g12324(new_n3615, n9172, new_n14673);
xor_4  g12325(new_n3615, n9172, new_n14674);
not_10 g12326(new_n14674, new_n14675);
or_5   g12327(new_n3618_1, n4913, new_n14676);
xor_4  g12328(new_n3618_1, new_n3549, new_n14677);
or_5   g12329(new_n3623, n604, new_n14678);
and_5  g12330(new_n3627, new_n3558, new_n14679);
not_10 g12331(new_n14679, new_n14680_1);
xor_4  g12332(new_n3627, new_n3558, new_n14681);
not_10 g12333(new_n14681, new_n14682);
or_5   g12334(new_n3632, n16521, new_n14683);
nand_5 g12335(n21993, n7139, new_n14684_1);
xor_4  g12336(new_n3632, n16521, new_n14685);
nand_5 g12337(new_n14685, new_n14684_1, new_n14686);
and_5  g12338(new_n14686, new_n14683, new_n14687);
nor_5  g12339(new_n14687, new_n14682, new_n14688);
not_10 g12340(new_n14688, new_n14689);
and_5  g12341(new_n14689, new_n14680_1, new_n14690);
xor_4  g12342(new_n3623, new_n3553, new_n14691);
or_5   g12343(new_n14691, new_n14690, new_n14692_1);
and_5  g12344(new_n14692_1, new_n14678, new_n14693);
or_5   g12345(new_n14693, new_n14677, new_n14694);
and_5  g12346(new_n14694, new_n14676, new_n14695);
or_5   g12347(new_n14695, new_n14675, new_n14696);
and_5  g12348(new_n14696, new_n14673, new_n14697);
nor_5  g12349(new_n14697, new_n14672, new_n14698);
nor_5  g12350(new_n14698, new_n14670, new_n14699);
not_10 g12351(new_n14699, new_n14700);
nor_5  g12352(new_n14700, new_n14669, new_n14701_1);
nor_5  g12353(new_n14701_1, new_n14668, new_n14702_1);
xor_4  g12354(new_n14702_1, new_n14667, new_n14703);
xor_4  g12355(new_n14703, new_n14666, new_n14704_1);
xor_4  g12356(new_n14662, new_n14661, new_n14705);
xor_4  g12357(new_n3607, new_n3537, new_n14706);
xor_4  g12358(new_n14706, new_n14700, new_n14707);
and_5  g12359(new_n14707, new_n14705, new_n14708);
not_10 g12360(new_n14705, new_n14709);
xnor_4 g12361(new_n14707, new_n14709, new_n14710);
xor_4  g12362(new_n14697, new_n14672, new_n14711);
xor_4  g12363(new_n14659, new_n14634, new_n14712);
nand_5 g12364(new_n14712, new_n14711, new_n14713);
xor_4  g12365(new_n14712, new_n14711, new_n14714);
not_10 g12366(new_n14714, new_n14715);
xor_4  g12367(new_n14695, new_n14675, new_n14716);
xor_4  g12368(new_n14657, new_n14637, new_n14717);
nand_5 g12369(new_n14717, new_n14716, new_n14718);
xor_4  g12370(new_n14717, new_n14716, new_n14719);
xor_4  g12371(new_n14693, new_n14677, new_n14720);
xor_4  g12372(new_n14655, new_n14640, new_n14721);
nor_5  g12373(new_n14721, new_n14720, new_n14722);
xor_4  g12374(new_n14691, new_n14690, new_n14723);
xor_4  g12375(new_n14653, new_n14643, new_n14724);
not_10 g12376(new_n14724, new_n14725);
nor_5  g12377(new_n14725, new_n14723, new_n14726);
xor_4  g12378(new_n14724, new_n14723, new_n14727);
xor_4  g12379(new_n14687, new_n14681, new_n14728);
xor_4  g12380(new_n14651, new_n14646, new_n14729);
nand_5 g12381(new_n14729, new_n14728, new_n14730);
xor_4  g12382(new_n14729, new_n14728, new_n14731);
xor_4  g12383(new_n14649, new_n14648, new_n14732);
or_5   g12384(new_n14732, new_n14685, new_n14733);
not_10 g12385(new_n14732, new_n14734_1);
xor_4  g12386(new_n14685, new_n14684_1, new_n14735);
nor_5  g12387(new_n14735, new_n14734_1, new_n14736);
xor_4  g12388(n21993, n7139, new_n14737);
xor_4  g12389(new_n9675, new_n3510, new_n14738);
and_5  g12390(new_n14738, new_n14737, new_n14739);
or_5   g12391(new_n14739, new_n14736, new_n14740);
and_5  g12392(new_n14740, new_n14733, new_n14741);
nand_5 g12393(new_n14741, new_n14731, new_n14742);
and_5  g12394(new_n14742, new_n14730, new_n14743);
nor_5  g12395(new_n14743, new_n14727, new_n14744);
or_5   g12396(new_n14744, new_n14726, new_n14745);
xor_4  g12397(new_n14721, new_n14720, new_n14746_1);
and_5  g12398(new_n14746_1, new_n14745, new_n14747);
nor_5  g12399(new_n14747, new_n14722, new_n14748);
nand_5 g12400(new_n14748, new_n14719, new_n14749);
and_5  g12401(new_n14749, new_n14718, new_n14750);
or_5   g12402(new_n14750, new_n14715, new_n14751);
and_5  g12403(new_n14751, new_n14713, new_n14752);
and_5  g12404(new_n14752, new_n14710, new_n14753);
nor_5  g12405(new_n14753, new_n14708, new_n14754);
xnor_4 g12406(new_n14754, new_n14704_1, n2779);
nor_5  g12407(new_n10542, n25751, new_n14756);
not_10 g12408(n25751, new_n14757);
xor_4  g12409(new_n10542, new_n14757, new_n14758);
or_5   g12410(new_n10545, n26053, new_n14759);
not_10 g12411(n26053, new_n14760);
xor_4  g12412(new_n10545, new_n14760, new_n14761);
or_5   g12413(new_n10548, n7917, new_n14762);
not_10 g12414(n7917, new_n14763_1);
xor_4  g12415(new_n10548, new_n14763_1, new_n14764);
or_5   g12416(new_n10551, n17302, new_n14765);
not_10 g12417(n17302, new_n14766);
xor_4  g12418(new_n10551, new_n14766, new_n14767);
or_5   g12419(new_n10553, n2013, new_n14768);
not_10 g12420(n2013, new_n14769);
xor_4  g12421(new_n10553, new_n14769, new_n14770);
or_5   g12422(new_n10556, n23755, new_n14771);
nor_5  g12423(new_n10559, n19163, new_n14772_1);
not_10 g12424(n19163, new_n14773);
xor_4  g12425(new_n10559, new_n14773, new_n14774);
or_5   g12426(new_n5868, n22358, new_n14775);
nand_5 g12427(n25926, n9646, new_n14776);
xor_4  g12428(new_n5868, n22358, new_n14777);
nand_5 g12429(new_n14777, new_n14776, new_n14778);
and_5  g12430(new_n14778, new_n14775, new_n14779);
nor_5  g12431(new_n14779, new_n14774, new_n14780);
or_5   g12432(new_n14780, new_n14772_1, new_n14781);
xor_4  g12433(new_n10556, n23755, new_n14782);
nand_5 g12434(new_n14782, new_n14781, new_n14783);
and_5  g12435(new_n14783, new_n14771, new_n14784);
or_5   g12436(new_n14784, new_n14770, new_n14785);
and_5  g12437(new_n14785, new_n14768, new_n14786);
or_5   g12438(new_n14786, new_n14767, new_n14787);
and_5  g12439(new_n14787, new_n14765, new_n14788);
or_5   g12440(new_n14788, new_n14764, new_n14789);
and_5  g12441(new_n14789, new_n14762, new_n14790_1);
or_5   g12442(new_n14790_1, new_n14761, new_n14791);
and_5  g12443(new_n14791, new_n14759, new_n14792);
nor_5  g12444(new_n14792, new_n14758, new_n14793);
or_5   g12445(new_n14793, new_n14756, new_n14794);
not_10 g12446(n25586, new_n14795);
xor_4  g12447(new_n10540_1, new_n14795, new_n14796);
xor_4  g12448(new_n14796, new_n14794, new_n14797);
xor_4  g12449(new_n14797, n4514, new_n14798);
xor_4  g12450(new_n14792, new_n14758, new_n14799);
or_5   g12451(new_n14799, n3984, new_n14800);
xor_4  g12452(new_n14799, new_n11756, new_n14801_1);
xor_4  g12453(new_n14790_1, new_n14761, new_n14802);
or_5   g12454(new_n14802, n19652, new_n14803);
xor_4  g12455(new_n14802, new_n11759, new_n14804);
xor_4  g12456(new_n14788, new_n14764, new_n14805);
or_5   g12457(new_n14805, n3366, new_n14806);
xor_4  g12458(new_n14786, new_n14767, new_n14807);
nor_5  g12459(new_n14807, n26565, new_n14808);
xor_4  g12460(new_n14807, new_n11765, new_n14809);
xor_4  g12461(new_n14784, new_n14770, new_n14810);
or_5   g12462(new_n14810, n3959, new_n14811);
xor_4  g12463(new_n14810, new_n11768, new_n14812);
xor_4  g12464(new_n14782, new_n14781, new_n14813);
or_5   g12465(new_n14813, n11566, new_n14814);
xor_4  g12466(new_n14813, new_n11771_1, new_n14815);
xor_4  g12467(new_n14779, new_n14774, new_n14816);
or_5   g12468(new_n14816, n26744, new_n14817);
xor_4  g12469(new_n14777, new_n14776, new_n14818);
nor_5  g12470(new_n14818, n26625, new_n14819_1);
or_5   g12471(new_n6631_1, new_n6630_1, new_n14820);
xor_4  g12472(new_n14818, n26625, new_n14821);
and_5  g12473(new_n14821, new_n14820, new_n14822);
or_5   g12474(new_n14822, new_n14819_1, new_n14823);
xor_4  g12475(new_n14816, n26744, new_n14824);
nand_5 g12476(new_n14824, new_n14823, new_n14825);
and_5  g12477(new_n14825, new_n14817, new_n14826_1);
or_5   g12478(new_n14826_1, new_n14815, new_n14827_1);
and_5  g12479(new_n14827_1, new_n14814, new_n14828);
or_5   g12480(new_n14828, new_n14812, new_n14829);
and_5  g12481(new_n14829, new_n14811, new_n14830);
nor_5  g12482(new_n14830, new_n14809, new_n14831);
or_5   g12483(new_n14831, new_n14808, new_n14832);
xor_4  g12484(new_n14805, n3366, new_n14833);
nand_5 g12485(new_n14833, new_n14832, new_n14834);
and_5  g12486(new_n14834, new_n14806, new_n14835);
or_5   g12487(new_n14835, new_n14804, new_n14836);
and_5  g12488(new_n14836, new_n14803, new_n14837);
or_5   g12489(new_n14837, new_n14801_1, new_n14838);
and_5  g12490(new_n14838, new_n14800, new_n14839_1);
xor_4  g12491(new_n14839_1, new_n14798, new_n14840);
nand_5 g12492(new_n14840, new_n10658, new_n14841);
xor_4  g12493(new_n14840, new_n10655, new_n14842);
not_10 g12494(new_n10661, new_n14843);
xor_4  g12495(new_n14837, new_n14801_1, new_n14844);
or_5   g12496(new_n14844, new_n14843, new_n14845);
xor_4  g12497(new_n14844, new_n10661, new_n14846);
xor_4  g12498(new_n14835, new_n14804, new_n14847);
or_5   g12499(new_n14847, new_n10666, new_n14848);
xor_4  g12500(new_n14847, new_n10665, new_n14849_1);
not_10 g12501(new_n10670, new_n14850);
xor_4  g12502(new_n14833, new_n14832, new_n14851);
or_5   g12503(new_n14851, new_n14850, new_n14852);
xor_4  g12504(new_n14851, new_n10670, new_n14853);
xor_4  g12505(new_n14830, new_n14809, new_n14854);
or_5   g12506(new_n14854, new_n10675, new_n14855);
xor_4  g12507(new_n14854, new_n10674, new_n14856);
not_10 g12508(new_n10679, new_n14857);
xor_4  g12509(new_n14828, new_n14812, new_n14858);
or_5   g12510(new_n14858, new_n14857, new_n14859);
xor_4  g12511(new_n14858, new_n10679, new_n14860);
xor_4  g12512(new_n14826_1, new_n14815, new_n14861);
or_5   g12513(new_n14861, new_n10685, new_n14862);
xor_4  g12514(new_n14861, new_n10684, new_n14863);
xor_4  g12515(new_n14824, new_n14823, new_n14864);
or_5   g12516(new_n14864, new_n10691, new_n14865);
xnor_4 g12517(new_n14864, new_n10691, new_n14866);
xor_4  g12518(new_n14821, new_n14820, new_n14867);
or_5   g12519(new_n14867, new_n5864, new_n14868);
nor_5  g12520(new_n6632, new_n6629, new_n14869);
and_5  g12521(new_n14867, new_n5866, new_n14870);
or_5   g12522(new_n14870, new_n14869, new_n14871);
and_5  g12523(new_n14871, new_n14868, new_n14872);
or_5   g12524(new_n14872, new_n14866, new_n14873);
and_5  g12525(new_n14873, new_n14865, new_n14874);
or_5   g12526(new_n14874, new_n14863, new_n14875);
and_5  g12527(new_n14875, new_n14862, new_n14876);
or_5   g12528(new_n14876, new_n14860, new_n14877);
and_5  g12529(new_n14877, new_n14859, new_n14878);
or_5   g12530(new_n14878, new_n14856, new_n14879);
and_5  g12531(new_n14879, new_n14855, new_n14880);
or_5   g12532(new_n14880, new_n14853, new_n14881);
and_5  g12533(new_n14881, new_n14852, new_n14882);
or_5   g12534(new_n14882, new_n14849_1, new_n14883);
and_5  g12535(new_n14883, new_n14848, new_n14884);
or_5   g12536(new_n14884, new_n14846, new_n14885);
and_5  g12537(new_n14885, new_n14845, new_n14886);
or_5   g12538(new_n14886, new_n14842, new_n14887);
and_5  g12539(new_n14887, new_n14841, new_n14888);
xor_4  g12540(new_n14888, new_n10650_1, new_n14889);
and_5  g12541(new_n14797, n4514, new_n14890);
and_5  g12542(new_n14839_1, new_n14798, new_n14891_1);
or_5   g12543(new_n14891_1, new_n14890, new_n14892);
and_5  g12544(new_n10540_1, new_n14795, new_n14893);
or_5   g12545(new_n14893, new_n14794, new_n14894);
nor_5  g12546(new_n10540_1, new_n14795, new_n14895);
nor_5  g12547(new_n14895, new_n10537, new_n14896);
and_5  g12548(new_n14896, new_n14894, new_n14897);
xor_4  g12549(new_n14897, new_n14892, new_n14898);
xor_4  g12550(new_n14898, new_n14889, n2826);
nand_5 g12551(new_n6278, n5140, new_n14900);
xor_4  g12552(new_n6278, new_n14262, new_n14901);
nand_5 g12553(new_n6285, n6204, new_n14902);
xor_4  g12554(new_n6285, new_n12551, new_n14903);
nand_5 g12555(new_n6292, n3349, new_n14904);
xor_4  g12556(new_n6292, new_n12555, new_n14905);
nand_5 g12557(new_n6296, n1742, new_n14906);
xor_4  g12558(new_n6296, new_n6499, new_n14907);
nand_5 g12559(new_n6300, n4858, new_n14908);
nor_5  g12560(new_n6305, n8244, new_n14909);
xor_4  g12561(new_n6305, n8244, new_n14910);
or_5   g12562(new_n6306, new_n6525, new_n14911);
xor_4  g12563(new_n6306, new_n6525, new_n14912);
or_5   g12564(new_n6309, n15167, new_n14913);
or_5   g12565(new_n6312, new_n12573, new_n14914);
and_5  g12566(new_n6314, n8656, new_n14915);
xor_4  g12567(new_n6312, new_n12573, new_n14916);
nand_5 g12568(new_n14916, new_n14915, new_n14917);
and_5  g12569(new_n14917, new_n14914, new_n14918);
xor_4  g12570(new_n6309, n15167, new_n14919);
nand_5 g12571(new_n14919, new_n14918, new_n14920);
and_5  g12572(new_n14920, new_n14913, new_n14921);
nand_5 g12573(new_n14921, new_n14912, new_n14922);
and_5  g12574(new_n14922, new_n14911, new_n14923);
and_5  g12575(new_n14923, new_n14910, new_n14924);
nor_5  g12576(new_n14924, new_n14909, new_n14925);
xor_4  g12577(new_n6300, n4858, new_n14926);
nand_5 g12578(new_n14926, new_n14925, new_n14927);
and_5  g12579(new_n14927, new_n14908, new_n14928);
or_5   g12580(new_n14928, new_n14907, new_n14929);
and_5  g12581(new_n14929, new_n14906, new_n14930);
or_5   g12582(new_n14930, new_n14905, new_n14931_1);
and_5  g12583(new_n14931_1, new_n14904, new_n14932);
or_5   g12584(new_n14932, new_n14903, new_n14933);
and_5  g12585(new_n14933, new_n14902, new_n14934);
or_5   g12586(new_n14934, new_n14901, new_n14935);
and_5  g12587(new_n14935, new_n14900, new_n14936);
or_5   g12588(new_n14936, new_n6235, new_n14937);
nor_5  g12589(new_n2592, new_n2557, new_n14938);
nor_5  g12590(new_n2648, new_n2594, new_n14939);
or_5   g12591(new_n14939, new_n14938, new_n14940);
nor_5  g12592(n20040, n9396, new_n14941);
not_10 g12593(new_n14941, new_n14942);
nor_5  g12594(new_n2591, new_n2558, new_n14943);
not_10 g12595(new_n14943, new_n14944_1);
and_5  g12596(new_n14944_1, new_n14942, new_n14945);
and_5  g12597(new_n14945, new_n14940, new_n14946);
not_10 g12598(new_n14946, new_n14947);
xor_4  g12599(new_n14947, new_n14937, new_n14948);
xor_4  g12600(new_n14936, new_n6235, new_n14949);
not_10 g12601(new_n14949, new_n14950);
xor_4  g12602(new_n14945, new_n14940, new_n14951);
and_5  g12603(new_n14951, new_n14950, new_n14952);
xor_4  g12604(new_n14951, new_n14950, new_n14953);
xnor_4 g12605(new_n14934, new_n14901, new_n14954_1);
and_5  g12606(new_n14954_1, new_n2649, new_n14955);
xor_4  g12607(new_n14954_1, new_n2649, new_n14956);
not_10 g12608(new_n14956, new_n14957);
xnor_4 g12609(new_n14932, new_n14903, new_n14958);
and_5  g12610(new_n14958, new_n2776, new_n14959);
xor_4  g12611(new_n14958, new_n2776, new_n14960);
not_10 g12612(new_n14960, new_n14961);
xor_4  g12613(new_n14930, new_n14905, new_n14962);
nor_5  g12614(new_n14962, new_n2781, new_n14963);
xnor_4 g12615(new_n14962, new_n2780, new_n14964);
not_10 g12616(new_n14964, new_n14965);
xor_4  g12617(new_n14928, new_n14907, new_n14966);
nor_5  g12618(new_n14966, new_n2787, new_n14967);
not_10 g12619(new_n14967, new_n14968);
xor_4  g12620(new_n14966, new_n2787, new_n14969);
xor_4  g12621(new_n14926, new_n14925, new_n14970);
nor_5  g12622(new_n14970, new_n2791, new_n14971);
xor_4  g12623(new_n14970, new_n2791, new_n14972);
not_10 g12624(new_n14972, new_n14973);
xor_4  g12625(new_n14923, new_n14910, new_n14974);
and_5  g12626(new_n14974, new_n2798, new_n14975);
not_10 g12627(new_n14975, new_n14976);
xor_4  g12628(new_n14974, new_n2798, new_n14977_1);
xor_4  g12629(new_n14921, new_n14912, new_n14978);
nor_5  g12630(new_n14978, new_n2803, new_n14979);
xnor_4 g12631(new_n14978, new_n2802, new_n14980);
not_10 g12632(new_n14980, new_n14981);
xor_4  g12633(new_n14919, new_n14918, new_n14982);
and_5  g12634(new_n14982, new_n2807, new_n14983);
xor_4  g12635(new_n14982, new_n2807, new_n14984);
not_10 g12636(new_n14984, new_n14985);
xor_4  g12637(new_n14916, new_n14915, new_n14986);
nor_5  g12638(new_n14986, new_n2811, new_n14987);
not_10 g12639(new_n14987, new_n14988);
xor_4  g12640(new_n6314, n8656, new_n14989_1);
nor_5  g12641(new_n14989_1, new_n2813, new_n14990);
xor_4  g12642(new_n14986, new_n2811, new_n14991);
and_5  g12643(new_n14991, new_n14990, new_n14992);
not_10 g12644(new_n14992, new_n14993);
and_5  g12645(new_n14993, new_n14988, new_n14994);
nor_5  g12646(new_n14994, new_n14985, new_n14995);
nor_5  g12647(new_n14995, new_n14983, new_n14996);
nor_5  g12648(new_n14996, new_n14981, new_n14997);
nor_5  g12649(new_n14997, new_n14979, new_n14998);
not_10 g12650(new_n14998, new_n14999);
and_5  g12651(new_n14999, new_n14977_1, new_n15000);
not_10 g12652(new_n15000, new_n15001);
and_5  g12653(new_n15001, new_n14976, new_n15002_1);
nor_5  g12654(new_n15002_1, new_n14973, new_n15003);
nor_5  g12655(new_n15003, new_n14971, new_n15004_1);
not_10 g12656(new_n15004_1, new_n15005);
and_5  g12657(new_n15005, new_n14969, new_n15006);
not_10 g12658(new_n15006, new_n15007);
and_5  g12659(new_n15007, new_n14968, new_n15008);
nor_5  g12660(new_n15008, new_n14965, new_n15009);
nor_5  g12661(new_n15009, new_n14963, new_n15010);
nor_5  g12662(new_n15010, new_n14961, new_n15011_1);
nor_5  g12663(new_n15011_1, new_n14959, new_n15012);
nor_5  g12664(new_n15012, new_n14957, new_n15013);
nor_5  g12665(new_n15013, new_n14955, new_n15014);
not_10 g12666(new_n15014, new_n15015);
and_5  g12667(new_n15015, new_n14953, new_n15016);
nor_5  g12668(new_n15016, new_n14952, new_n15017);
xnor_4 g12669(new_n15017, new_n14948, n2853);
xor_4  g12670(n7099, n2035, new_n15019_1);
or_5   g12671(new_n12060, n5213, new_n15020);
xor_4  g12672(n12811, n5213, new_n15021);
or_5   g12673(n4665, new_n12064, new_n15022);
xnor_4 g12674(n4665, n1118, new_n15023);
or_5   g12675(n25974, new_n2858_1, new_n15024);
nand_5 g12676(n25974, new_n2858_1, new_n15025);
not_10 g12677(n1630, new_n15026);
and_5  g12678(n4326, new_n15026, new_n15027);
and_5  g12679(new_n2860_1, n1630, new_n15028);
not_10 g12680(new_n15028, new_n15029);
and_5  g12681(n5438, new_n12069, new_n15030);
and_5  g12682(new_n15030, new_n15029, new_n15031_1);
nor_5  g12683(new_n15031_1, new_n15027, new_n15032);
not_10 g12684(new_n15032, new_n15033_1);
nand_5 g12685(new_n15033_1, new_n15025, new_n15034);
and_5  g12686(new_n15034, new_n15024, new_n15035);
nand_5 g12687(new_n15035, new_n15023, new_n15036);
and_5  g12688(new_n15036, new_n15022, new_n15037);
or_5   g12689(new_n15037, new_n15021, new_n15038);
and_5  g12690(new_n15038, new_n15020, new_n15039);
xor_4  g12691(new_n15039, new_n15019_1, new_n15040);
and_5  g12692(new_n4225, new_n4220, new_n15041);
xor_4  g12693(new_n15041, new_n6088, new_n15042);
xor_4  g12694(new_n15042, n5337, new_n15043);
and_5  g12695(new_n4226, n626, new_n15044);
nor_5  g12696(new_n4245, new_n4228, new_n15045);
nor_5  g12697(new_n15045, new_n15044, new_n15046);
xor_4  g12698(new_n15046, new_n15043, new_n15047);
xnor_4 g12699(new_n15047, new_n11285, new_n15048);
not_10 g12700(new_n15048, new_n15049);
or_5   g12701(new_n4247, new_n4219, new_n15050);
or_5   g12702(new_n4273, new_n4248, new_n15051);
and_5  g12703(new_n15051, new_n15050, new_n15052_1);
xor_4  g12704(new_n15052_1, new_n15049, new_n15053_1);
not_10 g12705(new_n15053_1, new_n15054);
xnor_4 g12706(new_n15054, new_n15040, new_n15055);
xor_4  g12707(new_n15037, new_n15021, new_n15056);
or_5   g12708(new_n15056, new_n4274, new_n15057);
xor_4  g12709(new_n15035, new_n15023, new_n15058);
or_5   g12710(new_n15058, new_n4277, new_n15059);
xor_4  g12711(new_n15058, new_n4277, new_n15060);
not_10 g12712(new_n15060, new_n15061);
xnor_4 g12713(n25974, n19005, new_n15062);
xor_4  g12714(new_n15062, new_n15033_1, new_n15063);
nand_5 g12715(new_n15063, new_n4282, new_n15064);
xnor_4 g12716(new_n15063, new_n4282, new_n15065);
not_10 g12717(new_n4292, new_n15066);
xnor_4 g12718(n5438, n1451, new_n15067);
or_5   g12719(new_n15067, new_n15066, new_n15068);
xnor_4 g12720(n4326, n1630, new_n15069);
xor_4  g12721(new_n15069, new_n15030, new_n15070);
nor_5  g12722(new_n15070, new_n15068, new_n15071);
not_10 g12723(new_n15071, new_n15072);
xor_4  g12724(new_n15070, new_n15068, new_n15073);
and_5  g12725(new_n15073, new_n4286, new_n15074);
not_10 g12726(new_n15074, new_n15075);
and_5  g12727(new_n15075, new_n15072, new_n15076);
not_10 g12728(new_n15076, new_n15077_1);
or_5   g12729(new_n15077_1, new_n15065, new_n15078);
and_5  g12730(new_n15078, new_n15064, new_n15079);
or_5   g12731(new_n15079, new_n15061, new_n15080);
and_5  g12732(new_n15080, new_n15059, new_n15081);
xor_4  g12733(new_n15056, new_n4274, new_n15082_1);
not_10 g12734(new_n15082_1, new_n15083);
or_5   g12735(new_n15083, new_n15081, new_n15084);
and_5  g12736(new_n15084, new_n15057, new_n15085);
xor_4  g12737(new_n15085, new_n15055, n2860);
xnor_4 g12738(new_n14140, new_n14118, n2887);
and_5  g12739(new_n15041, new_n6088, new_n15088);
and_5  g12740(new_n15088, new_n6083, new_n15089);
and_5  g12741(new_n15089, new_n6078, new_n15090);
and_5  g12742(new_n15090, new_n6073, new_n15091);
xor_4  g12743(new_n15091, new_n6035, new_n15092);
nor_5  g12744(new_n15092, n21784, new_n15093);
xor_4  g12745(new_n15090, new_n6073, new_n15094_1);
and_5  g12746(new_n15094_1, n5521, new_n15095);
nor_5  g12747(new_n15094_1, n5521, new_n15096);
xor_4  g12748(new_n15089, new_n6078, new_n15097);
nor_5  g12749(new_n15097, n11926, new_n15098);
xor_4  g12750(new_n15097, n11926, new_n15099);
xor_4  g12751(new_n15088, new_n6083, new_n15100);
nand_5 g12752(new_n15100, n4325, new_n15101);
nor_5  g12753(new_n15100, n4325, new_n15102);
and_5  g12754(new_n15042, n5337, new_n15103);
nor_5  g12755(new_n15042, n5337, new_n15104);
nor_5  g12756(new_n15046, new_n15104, new_n15105);
nor_5  g12757(new_n15105, new_n15103, new_n15106);
or_5   g12758(new_n15106, new_n15102, new_n15107);
and_5  g12759(new_n15107, new_n15101, new_n15108);
and_5  g12760(new_n15108, new_n15099, new_n15109);
nor_5  g12761(new_n15109, new_n15098, new_n15110);
not_10 g12762(new_n15110, new_n15111);
nor_5  g12763(new_n15111, new_n15096, new_n15112);
nor_5  g12764(new_n15112, new_n15095, new_n15113);
or_5   g12765(new_n15113, new_n15093, new_n15114);
nand_5 g12766(new_n15091, new_n6035, new_n15115);
nand_5 g12767(new_n15092, n21784, new_n15116);
and_5  g12768(new_n15116, new_n15115, new_n15117);
and_5  g12769(new_n15117, new_n15114, new_n15118_1);
xor_4  g12770(new_n15118_1, new_n11259, new_n15119);
xor_4  g12771(new_n15092, new_n12092, new_n15120);
xor_4  g12772(new_n15120, new_n15113, new_n15121);
nand_5 g12773(new_n15121, new_n11264, new_n15122);
xor_4  g12774(new_n15121, new_n11264, new_n15123);
xor_4  g12775(new_n15094_1, new_n12093, new_n15124);
xor_4  g12776(new_n15124, new_n15111, new_n15125);
or_5   g12777(new_n15125, new_n11269, new_n15126);
xor_4  g12778(new_n15125, new_n11269, new_n15127);
not_10 g12779(new_n15127, new_n15128_1);
xor_4  g12780(new_n15108, new_n15099, new_n15129);
nand_5 g12781(new_n15129, new_n11275_1, new_n15130);
xor_4  g12782(new_n15100, n4325, new_n15131);
xnor_4 g12783(new_n15131, new_n15106, new_n15132);
and_5  g12784(new_n15132, new_n11279, new_n15133);
xor_4  g12785(new_n15132, new_n11279, new_n15134);
not_10 g12786(new_n15134, new_n15135);
not_10 g12787(new_n15047, new_n15136);
nand_5 g12788(new_n15136, new_n11285, new_n15137);
or_5   g12789(new_n15052_1, new_n15049, new_n15138);
and_5  g12790(new_n15138, new_n15137, new_n15139_1);
nor_5  g12791(new_n15139_1, new_n15135, new_n15140);
nor_5  g12792(new_n15140, new_n15133, new_n15141);
xnor_4 g12793(new_n15129, new_n11274, new_n15142);
nand_5 g12794(new_n15142, new_n15141, new_n15143);
and_5  g12795(new_n15143, new_n15130, new_n15144);
or_5   g12796(new_n15144, new_n15128_1, new_n15145_1);
and_5  g12797(new_n15145_1, new_n15126, new_n15146_1);
nand_5 g12798(new_n15146_1, new_n15123, new_n15147);
and_5  g12799(new_n15147, new_n15122, new_n15148);
xor_4  g12800(new_n15148, new_n15119, new_n15149);
not_10 g12801(n8827, new_n15150);
not_10 g12802(n18035, new_n15151);
and_5  g12803(new_n4170, new_n4165_1, new_n15152);
and_5  g12804(new_n15152, new_n10766, new_n15153);
and_5  g12805(new_n15153, new_n10762, new_n15154);
and_5  g12806(new_n15154, new_n10743, new_n15155);
and_5  g12807(new_n15155, new_n15151, new_n15156);
and_5  g12808(new_n15156, new_n15150, new_n15157);
xor_4  g12809(new_n15156, new_n15150, new_n15158);
nor_5  g12810(new_n15158, n11898, new_n15159);
xor_4  g12811(new_n15155, new_n15151, new_n15160);
nor_5  g12812(new_n15160, n19941, new_n15161);
xor_4  g12813(new_n15160, new_n14446, new_n15162);
xor_4  g12814(new_n15154, new_n10743, new_n15163);
or_5   g12815(new_n15163, n1099, new_n15164);
xor_4  g12816(new_n15163, new_n14447, new_n15165_1);
xor_4  g12817(new_n15153, new_n10762, new_n15166);
or_5   g12818(new_n15166, n2113, new_n15167_1);
xor_4  g12819(new_n15152, new_n10766, new_n15168);
nor_5  g12820(new_n15168, n21134, new_n15169);
xor_4  g12821(new_n15168, new_n3726, new_n15170);
or_5   g12822(new_n4171, n6369, new_n15171);
nand_5 g12823(new_n4189, new_n4172_1, new_n15172);
and_5  g12824(new_n15172, new_n15171, new_n15173);
nor_5  g12825(new_n15173, new_n15170, new_n15174);
or_5   g12826(new_n15174, new_n15169, new_n15175);
xor_4  g12827(new_n15166, n2113, new_n15176_1);
nand_5 g12828(new_n15176_1, new_n15175, new_n15177);
and_5  g12829(new_n15177, new_n15167_1, new_n15178);
or_5   g12830(new_n15178, new_n15165_1, new_n15179);
and_5  g12831(new_n15179, new_n15164, new_n15180_1);
nor_5  g12832(new_n15180_1, new_n15162, new_n15181);
nor_5  g12833(new_n15181, new_n15161, new_n15182_1);
and_5  g12834(new_n15158, n11898, new_n15183);
nor_5  g12835(new_n15183, new_n15182_1, new_n15184);
nor_5  g12836(new_n15184, new_n15159, new_n15185);
nor_5  g12837(new_n15185, new_n15157, new_n15186);
xnor_4 g12838(new_n15186, new_n15149, new_n15187);
xor_4  g12839(new_n15146_1, new_n15123, new_n15188);
not_10 g12840(new_n15188, new_n15189);
xor_4  g12841(new_n15158, new_n14445, new_n15190);
xor_4  g12842(new_n15190, new_n15182_1, new_n15191);
and_5  g12843(new_n15191, new_n15189, new_n15192);
xor_4  g12844(new_n15191, new_n15189, new_n15193);
xor_4  g12845(new_n15180_1, new_n15162, new_n15194);
xnor_4 g12846(new_n15144, new_n15127, new_n15195);
and_5  g12847(new_n15195, new_n15194, new_n15196);
xor_4  g12848(new_n15195, new_n15194, new_n15197);
not_10 g12849(new_n15197, new_n15198);
xor_4  g12850(new_n15178, new_n15165_1, new_n15199);
xor_4  g12851(new_n15142, new_n15141, new_n15200);
and_5  g12852(new_n15200, new_n15199, new_n15201);
xor_4  g12853(new_n15200, new_n15199, new_n15202);
not_10 g12854(new_n15202, new_n15203);
xor_4  g12855(new_n15139_1, new_n15135, new_n15204);
not_10 g12856(new_n15204, new_n15205_1);
xor_4  g12857(new_n15176_1, new_n15175, new_n15206);
and_5  g12858(new_n15206, new_n15205_1, new_n15207);
not_10 g12859(new_n15207, new_n15208);
xor_4  g12860(new_n15206, new_n15205_1, new_n15209);
not_10 g12861(new_n15209, new_n15210);
xor_4  g12862(new_n15173, new_n15170, new_n15211);
and_5  g12863(new_n15211, new_n15054, new_n15212);
not_10 g12864(new_n15212, new_n15213);
xor_4  g12865(new_n15211, new_n15054, new_n15214);
nor_5  g12866(new_n4274, new_n4191, new_n15215);
not_10 g12867(new_n15215, new_n15216);
and_5  g12868(new_n4299, new_n4275, new_n15217);
not_10 g12869(new_n15217, new_n15218);
and_5  g12870(new_n15218, new_n15216, new_n15219);
not_10 g12871(new_n15219, new_n15220);
and_5  g12872(new_n15220, new_n15214, new_n15221);
not_10 g12873(new_n15221, new_n15222);
and_5  g12874(new_n15222, new_n15213, new_n15223);
nor_5  g12875(new_n15223, new_n15210, new_n15224);
not_10 g12876(new_n15224, new_n15225);
and_5  g12877(new_n15225, new_n15208, new_n15226);
nor_5  g12878(new_n15226, new_n15203, new_n15227);
nor_5  g12879(new_n15227, new_n15201, new_n15228);
nor_5  g12880(new_n15228, new_n15198, new_n15229);
nor_5  g12881(new_n15229, new_n15196, new_n15230_1);
not_10 g12882(new_n15230_1, new_n15231);
and_5  g12883(new_n15231, new_n15193, new_n15232);
nor_5  g12884(new_n15232, new_n15192, new_n15233);
xor_4  g12885(new_n15233, new_n15187, n2929);
xor_4  g12886(n22793, n767, new_n15235);
or_5   g12887(n8439, new_n11221, new_n15236);
xor_4  g12888(n8439, n7330, new_n15237);
or_5   g12889(n25523, new_n11222, new_n15238);
xor_4  g12890(n25523, n22492, new_n15239);
or_5   g12891(new_n11223_1, n5579, new_n15240);
xor_4  g12892(n12821, n5579, new_n15241_1);
or_5   g12893(n23430, new_n4192, new_n15242);
xnor_4 g12894(n23430, n3468, new_n15243);
or_5   g12895(n18558, new_n2656, new_n15244);
or_5   g12896(new_n13853, new_n13842, new_n15245);
and_5  g12897(new_n15245, new_n15244, new_n15246);
nand_5 g12898(new_n15246, new_n15243, new_n15247);
and_5  g12899(new_n15247, new_n15242, new_n15248);
or_5   g12900(new_n15248, new_n15241_1, new_n15249);
and_5  g12901(new_n15249, new_n15240, new_n15250);
or_5   g12902(new_n15250, new_n15239, new_n15251);
and_5  g12903(new_n15251, new_n15238, new_n15252);
or_5   g12904(new_n15252, new_n15237, new_n15253);
and_5  g12905(new_n15253, new_n15236, new_n15254);
xor_4  g12906(new_n15254, new_n15235, new_n15255_1);
xor_4  g12907(new_n15255_1, new_n7316, new_n15256);
not_10 g12908(new_n15256, new_n15257);
xor_4  g12909(new_n15252, new_n15237, new_n15258_1);
nand_5 g12910(new_n15258_1, new_n7321, new_n15259);
xor_4  g12911(new_n15258_1, new_n7321, new_n15260);
xor_4  g12912(new_n15250, new_n15239, new_n15261);
or_5   g12913(new_n15261, new_n7326, new_n15262);
xor_4  g12914(new_n15261, new_n7326, new_n15263);
not_10 g12915(new_n15263, new_n15264);
xor_4  g12916(new_n15248, new_n15241_1, new_n15265);
or_5   g12917(new_n15265, new_n7330_1, new_n15266);
xor_4  g12918(new_n15265, new_n7330_1, new_n15267);
xor_4  g12919(new_n15246, new_n15243, new_n15268);
nand_5 g12920(new_n15268, new_n7334, new_n15269);
xor_4  g12921(new_n15268, new_n7334, new_n15270);
not_10 g12922(new_n15270, new_n15271_1);
or_5   g12923(new_n13854, new_n12366, new_n15272);
or_5   g12924(new_n14163, new_n14153, new_n15273);
and_5  g12925(new_n15273, new_n15272, new_n15274);
or_5   g12926(new_n15274, new_n15271_1, new_n15275_1);
and_5  g12927(new_n15275_1, new_n15269, new_n15276);
nand_5 g12928(new_n15276, new_n15267, new_n15277);
and_5  g12929(new_n15277, new_n15266, new_n15278);
or_5   g12930(new_n15278, new_n15264, new_n15279);
and_5  g12931(new_n15279, new_n15262, new_n15280);
nand_5 g12932(new_n15280, new_n15260, new_n15281);
and_5  g12933(new_n15281, new_n15259, new_n15282);
xor_4  g12934(new_n15282, new_n15257, new_n15283);
xor_4  g12935(n22379, n15077, new_n15284);
or_5   g12936(n3710, new_n2837, new_n15285);
xnor_4 g12937(n3710, n1662, new_n15286);
not_10 g12938(new_n15286, new_n15287);
or_5   g12939(n26318, new_n2841, new_n15288);
xnor_4 g12940(n26318, n12875, new_n15289_1);
not_10 g12941(new_n15289_1, new_n15290);
or_5   g12942(n26054, new_n2845, new_n15291);
xnor_4 g12943(n26054, n2035, new_n15292);
not_10 g12944(new_n15292, new_n15293);
or_5   g12945(n19081, new_n2849, new_n15294);
or_5   g12946(new_n8921, n5213, new_n15295);
and_5  g12947(n8309, new_n2853_1, new_n15296);
nor_5  g12948(new_n14177, new_n14166, new_n15297);
nor_5  g12949(new_n15297, new_n15296, new_n15298);
nand_5 g12950(new_n15298, new_n15295, new_n15299);
and_5  g12951(new_n15299, new_n15294, new_n15300_1);
or_5   g12952(new_n15300_1, new_n15293, new_n15301);
and_5  g12953(new_n15301, new_n15291, new_n15302);
or_5   g12954(new_n15302, new_n15290, new_n15303);
and_5  g12955(new_n15303, new_n15288, new_n15304);
or_5   g12956(new_n15304, new_n15287, new_n15305);
and_5  g12957(new_n15305, new_n15285, new_n15306);
xor_4  g12958(new_n15306, new_n15284, new_n15307_1);
xor_4  g12959(new_n15307_1, new_n15283, new_n15308);
not_10 g12960(new_n15308, new_n15309);
xor_4  g12961(new_n15304, new_n15287, new_n15310);
xor_4  g12962(new_n15280, new_n15260, new_n15311);
nor_5  g12963(new_n15311, new_n15310, new_n15312);
xor_4  g12964(new_n15311, new_n15310, new_n15313);
not_10 g12965(new_n15313, new_n15314);
xor_4  g12966(new_n15302, new_n15290, new_n15315);
xor_4  g12967(new_n15278, new_n15264, new_n15316);
not_10 g12968(new_n15316, new_n15317);
nor_5  g12969(new_n15317, new_n15315, new_n15318);
not_10 g12970(new_n15318, new_n15319);
xor_4  g12971(new_n15317, new_n15315, new_n15320);
xor_4  g12972(new_n15300_1, new_n15293, new_n15321);
xor_4  g12973(new_n15276, new_n15267, new_n15322);
not_10 g12974(new_n15322, new_n15323);
nor_5  g12975(new_n15323, new_n15321, new_n15324);
not_10 g12976(new_n15324, new_n15325);
xor_4  g12977(new_n15274, new_n15271_1, new_n15326);
xnor_4 g12978(n19081, n5213, new_n15327_1);
xor_4  g12979(new_n15327_1, new_n15298, new_n15328);
nor_5  g12980(new_n15328, new_n15326, new_n15329);
not_10 g12981(new_n15329, new_n15330);
not_10 g12982(new_n15326, new_n15331);
xnor_4 g12983(new_n15328, new_n15331, new_n15332_1);
and_5  g12984(new_n14178, new_n14165, new_n15333);
not_10 g12985(new_n15333, new_n15334);
not_10 g12986(new_n14202, new_n15335);
and_5  g12987(new_n15335, new_n14179, new_n15336);
not_10 g12988(new_n15336, new_n15337);
and_5  g12989(new_n15337, new_n15334, new_n15338);
not_10 g12990(new_n15338, new_n15339);
and_5  g12991(new_n15339, new_n15332_1, new_n15340);
not_10 g12992(new_n15340, new_n15341);
and_5  g12993(new_n15341, new_n15330, new_n15342);
not_10 g12994(new_n15342, new_n15343);
xor_4  g12995(new_n15323, new_n15321, new_n15344);
and_5  g12996(new_n15344, new_n15343, new_n15345_1);
not_10 g12997(new_n15345_1, new_n15346);
and_5  g12998(new_n15346, new_n15325, new_n15347);
not_10 g12999(new_n15347, new_n15348);
and_5  g13000(new_n15348, new_n15320, new_n15349);
not_10 g13001(new_n15349, new_n15350);
and_5  g13002(new_n15350, new_n15319, new_n15351);
nor_5  g13003(new_n15351, new_n15314, new_n15352);
nor_5  g13004(new_n15352, new_n15312, new_n15353_1);
xnor_4 g13005(new_n15353_1, new_n15309, n2948);
xor_4  g13006(new_n14743, new_n14727, n2961);
xnor_4 g13007(new_n11586, new_n11560, n2971);
xnor_4 g13008(new_n2538, new_n2519, n3010);
xor_4  g13009(new_n6767, new_n6759, n3017);
xor_4  g13010(new_n11965_1, new_n9199, new_n15359);
xor_4  g13011(new_n15359, new_n11969, n3020);
xor_4  g13012(new_n6177, new_n6152, n3067);
xor_4  g13013(n23541, n19234, new_n15362);
xor_4  g13014(n27134, n4588, new_n15363);
xor_4  g13015(new_n15363, new_n15362, new_n15364);
not_10 g13016(new_n15364, new_n15365);
xor_4  g13017(new_n15365, new_n10144, n3076);
nor_5  g13018(n15490, n18, new_n15367);
and_5  g13019(new_n15367, new_n9328, new_n15368);
xor_4  g13020(new_n15368, new_n9324, new_n15369);
xor_4  g13021(new_n15369, new_n6634_1, new_n15370);
xor_4  g13022(new_n15367, new_n9328, new_n15371);
nand_5 g13023(new_n15371, n19680, new_n15372);
xor_4  g13024(new_n15371, n19680, new_n15373);
xor_4  g13025(n15490, n18, new_n15374);
or_5   g13026(new_n15374, n2809, new_n15375);
nand_5 g13027(n15508, n18, new_n15376);
xor_4  g13028(new_n15374, n2809, new_n15377);
nand_5 g13029(new_n15377, new_n15376, new_n15378_1);
and_5  g13030(new_n15378_1, new_n15375, new_n15379);
nand_5 g13031(new_n15379, new_n15373, new_n15380);
and_5  g13032(new_n15380, new_n15372, new_n15381);
xor_4  g13033(new_n15381, new_n15370, new_n15382_1);
xor_4  g13034(new_n15382_1, new_n10887, new_n15383);
xor_4  g13035(new_n15379, new_n15373, new_n15384);
nand_5 g13036(new_n15384, new_n10890, new_n15385);
xor_4  g13037(new_n15384, new_n10890, new_n15386);
or_5   g13038(new_n15377, new_n5848, new_n15387);
xor_4  g13039(new_n15377, new_n15376, new_n15388);
nor_5  g13040(new_n15388, new_n5849, new_n15389);
xor_4  g13041(n15508, n18, new_n15390);
and_5  g13042(new_n15390, new_n5831, new_n15391);
or_5   g13043(new_n15391, new_n15389, new_n15392);
and_5  g13044(new_n15392, new_n15387, new_n15393);
nand_5 g13045(new_n15393, new_n15386, new_n15394);
and_5  g13046(new_n15394, new_n15385, new_n15395);
xor_4  g13047(new_n15395, new_n15383, n3089);
xor_4  g13048(new_n5224, new_n5222, n3125);
xnor_4 g13049(n21839, n19282, new_n15398);
or_5   g13050(n27089, n12657, new_n15399);
or_5   g13051(new_n2950, new_n2915, new_n15400);
and_5  g13052(new_n15400, new_n15399, new_n15401);
xor_4  g13053(new_n15401, new_n15398, new_n15402);
nor_5  g13054(new_n15402, new_n11229, new_n15403);
not_10 g13055(new_n15403, new_n15404);
xnor_4 g13056(new_n15402, new_n11229, new_n15405);
or_5   g13057(new_n11232, new_n2951, new_n15406);
nor_5  g13058(new_n11235, new_n2954, new_n15407_1);
xnor_4 g13059(new_n11235, new_n2955, new_n15408);
nand_5 g13060(new_n11239, new_n2959, new_n15409);
xor_4  g13061(new_n11239, new_n2960, new_n15410);
nand_5 g13062(new_n11242, new_n2965, new_n15411);
or_5   g13063(new_n13633, new_n13615, new_n15412);
and_5  g13064(new_n15412, new_n15411, new_n15413);
or_5   g13065(new_n15413, new_n15410, new_n15414);
and_5  g13066(new_n15414, new_n15409, new_n15415);
and_5  g13067(new_n15415, new_n15408, new_n15416);
or_5   g13068(new_n15416, new_n15407_1, new_n15417);
not_10 g13069(new_n2951, new_n15418);
xnor_4 g13070(new_n11232, new_n15418, new_n15419);
nand_5 g13071(new_n15419, new_n15417, new_n15420);
and_5  g13072(new_n15420, new_n15406, new_n15421);
nor_5  g13073(new_n15421, new_n15405, new_n15422);
not_10 g13074(new_n15422, new_n15423);
and_5  g13075(new_n15423, new_n15404, new_n15424_1);
nor_5  g13076(n21839, n19282, new_n15425);
nor_5  g13077(new_n15401, new_n15398, new_n15426);
nor_5  g13078(new_n15426, new_n15425, new_n15427);
nor_5  g13079(new_n15427, new_n11231, new_n15428_1);
and_5  g13080(new_n15428_1, new_n15424_1, new_n15429);
and_5  g13081(new_n15427, new_n11231, new_n15430);
not_10 g13082(new_n15430, new_n15431);
nor_5  g13083(new_n15431, new_n15424_1, new_n15432);
nor_5  g13084(new_n15432, new_n15429, new_n15433);
xor_4  g13085(new_n15433, new_n12188, new_n15434);
xnor_4 g13086(new_n15427, new_n11231, new_n15435_1);
xor_4  g13087(new_n15435_1, new_n15424_1, new_n15436);
nor_5  g13088(new_n15436, new_n11658, new_n15437);
xor_4  g13089(new_n15436, new_n11658, new_n15438_1);
xor_4  g13090(new_n15421, new_n15405, new_n15439);
and_5  g13091(new_n15439, new_n12251, new_n15440);
xnor_4 g13092(new_n15439, new_n11672, new_n15441);
not_10 g13093(new_n15441, new_n15442);
xor_4  g13094(new_n15419, new_n15417, new_n15443);
and_5  g13095(new_n15443, new_n11680, new_n15444);
not_10 g13096(new_n15444, new_n15445);
xor_4  g13097(new_n15443, new_n11680, new_n15446);
xor_4  g13098(new_n15415, new_n15408, new_n15447);
and_5  g13099(new_n15447, new_n11682_1, new_n15448);
xor_4  g13100(new_n15447, new_n11682_1, new_n15449);
not_10 g13101(new_n15449, new_n15450);
xor_4  g13102(new_n15413, new_n15410, new_n15451);
nor_5  g13103(new_n15451, new_n11688, new_n15452);
not_10 g13104(new_n15452, new_n15453);
xor_4  g13105(new_n15451, new_n11688, new_n15454);
nor_5  g13106(new_n13634, new_n11693, new_n15455);
nor_5  g13107(new_n13662, new_n13636, new_n15456);
nor_5  g13108(new_n15456, new_n15455, new_n15457);
not_10 g13109(new_n15457, new_n15458);
and_5  g13110(new_n15458, new_n15454, new_n15459);
not_10 g13111(new_n15459, new_n15460);
and_5  g13112(new_n15460, new_n15453, new_n15461);
nor_5  g13113(new_n15461, new_n15450, new_n15462);
nor_5  g13114(new_n15462, new_n15448, new_n15463);
not_10 g13115(new_n15463, new_n15464);
and_5  g13116(new_n15464, new_n15446, new_n15465_1);
not_10 g13117(new_n15465_1, new_n15466);
and_5  g13118(new_n15466, new_n15445, new_n15467_1);
nor_5  g13119(new_n15467_1, new_n15442, new_n15468);
nor_5  g13120(new_n15468, new_n15440, new_n15469);
not_10 g13121(new_n15469, new_n15470_1);
and_5  g13122(new_n15470_1, new_n15438_1, new_n15471);
nor_5  g13123(new_n15471, new_n15437, new_n15472);
xor_4  g13124(new_n15472, new_n15434, n3126);
xnor_4 g13125(new_n12305, new_n12263, n3208);
xor_4  g13126(new_n14568, new_n14566, n3219);
xnor_4 g13127(new_n14994, new_n14985, n3235);
xnor_4 g13128(new_n11448, new_n11435, n3244);
not_10 g13129(n15146, new_n15478);
or_5   g13130(new_n15478, n5532, new_n15479);
not_10 g13131(new_n10105, new_n15480);
not_10 g13132(n11579, new_n15481_1);
or_5   g13133(new_n15481_1, n3962, new_n15482);
not_10 g13134(new_n10102, new_n15483);
not_10 g13135(n21, new_n15484);
or_5   g13136(n23513, new_n15484, new_n15485);
not_10 g13137(new_n10085, new_n15486);
not_10 g13138(new_n10134, new_n15487);
nand_5 g13139(new_n13867, new_n15487, new_n15488);
not_10 g13140(n1682, new_n15489);
or_5   g13141(n6427, new_n15489, new_n15490_1);
and_5  g13142(new_n15490_1, new_n15488, new_n15491);
or_5   g13143(new_n15491, new_n15486, new_n15492);
and_5  g13144(new_n15492, new_n15485, new_n15493);
or_5   g13145(new_n15493, new_n15483, new_n15494);
and_5  g13146(new_n15494, new_n15482, new_n15495);
or_5   g13147(new_n15495, new_n15480, new_n15496_1);
and_5  g13148(new_n15496_1, new_n15479, new_n15497);
xnor_4 g13149(new_n15497, new_n10108, new_n15498);
xor_4  g13150(new_n15498, new_n15258_1, new_n15499);
not_10 g13151(new_n15499, new_n15500);
xnor_4 g13152(new_n15495, new_n10105, new_n15501_1);
or_5   g13153(new_n15501_1, new_n15261, new_n15502);
xor_4  g13154(new_n15501_1, new_n15261, new_n15503);
not_10 g13155(new_n15503, new_n15504);
xnor_4 g13156(new_n15493, new_n10102, new_n15505);
or_5   g13157(new_n15505, new_n15265, new_n15506_1);
xor_4  g13158(new_n15505, new_n15265, new_n15507);
not_10 g13159(new_n15507, new_n15508_1);
xor_4  g13160(new_n15491, new_n15486, new_n15509);
or_5   g13161(new_n15509, new_n15268, new_n15510);
xor_4  g13162(new_n15509, new_n15268, new_n15511);
or_5   g13163(new_n13869, new_n13854, new_n15512);
nand_5 g13164(new_n13889, new_n13870, new_n15513);
and_5  g13165(new_n15513, new_n15512, new_n15514);
nand_5 g13166(new_n15514, new_n15511, new_n15515);
and_5  g13167(new_n15515, new_n15510, new_n15516);
or_5   g13168(new_n15516, new_n15508_1, new_n15517);
and_5  g13169(new_n15517, new_n15506_1, new_n15518);
or_5   g13170(new_n15518, new_n15504, new_n15519);
and_5  g13171(new_n15519, new_n15502, new_n15520);
xor_4  g13172(new_n15520, new_n15500, new_n15521);
nor_5  g13173(n23541, n16247, new_n15522);
and_5  g13174(new_n15522, new_n2622, new_n15523);
and_5  g13175(new_n15523, new_n2617, new_n15524);
and_5  g13176(new_n15524, new_n2613, new_n15525);
and_5  g13177(new_n15525, new_n2608, new_n15526);
and_5  g13178(new_n15526, new_n2605, new_n15527);
xor_4  g13179(new_n15527, new_n2600, new_n15528);
xor_4  g13180(new_n15528, n18345, new_n15529);
not_10 g13181(new_n15529, new_n15530);
xor_4  g13182(new_n15526, new_n2605, new_n15531);
or_5   g13183(new_n15531, n13190, new_n15532);
xor_4  g13184(new_n15531, n13190, new_n15533);
not_10 g13185(new_n15533, new_n15534);
xor_4  g13186(new_n15525, new_n2608, new_n15535);
or_5   g13187(new_n15535, n3460, new_n15536);
xor_4  g13188(new_n15535, n3460, new_n15537);
not_10 g13189(new_n15537, new_n15538);
xor_4  g13190(new_n15524, new_n2613, new_n15539_1);
or_5   g13191(new_n15539_1, n5226, new_n15540);
xor_4  g13192(new_n15539_1, n5226, new_n15541);
not_10 g13193(new_n15541, new_n15542);
xor_4  g13194(new_n15523, new_n2617, new_n15543);
or_5   g13195(new_n15543, n17664, new_n15544);
xor_4  g13196(new_n15522, new_n2622, new_n15545);
nor_5  g13197(new_n15545, n23369, new_n15546_1);
not_10 g13198(new_n15546_1, new_n15547);
xor_4  g13199(new_n15545, new_n8866, new_n15548);
xor_4  g13200(n23541, n16247, new_n15549);
or_5   g13201(new_n15549, n1136, new_n15550);
nand_5 g13202(n23541, n19234, new_n15551);
xor_4  g13203(new_n15549, n1136, new_n15552);
nand_5 g13204(new_n15552, new_n15551, new_n15553);
and_5  g13205(new_n15553, new_n15550, new_n15554);
nor_5  g13206(new_n15554, new_n15548, new_n15555_1);
not_10 g13207(new_n15555_1, new_n15556);
and_5  g13208(new_n15556, new_n15547, new_n15557);
xor_4  g13209(new_n15543, new_n9746, new_n15558_1);
or_5   g13210(new_n15558_1, new_n15557, new_n15559_1);
and_5  g13211(new_n15559_1, new_n15544, new_n15560);
or_5   g13212(new_n15560, new_n15542, new_n15561);
and_5  g13213(new_n15561, new_n15540, new_n15562);
or_5   g13214(new_n15562, new_n15538, new_n15563);
and_5  g13215(new_n15563, new_n15536, new_n15564);
or_5   g13216(new_n15564, new_n15534, new_n15565);
and_5  g13217(new_n15565, new_n15532, new_n15566);
xor_4  g13218(new_n15566, new_n15530, new_n15567);
xor_4  g13219(new_n15567, new_n15521, new_n15568);
not_10 g13220(new_n15568, new_n15569);
xor_4  g13221(new_n15564, new_n15534, new_n15570_1);
xor_4  g13222(new_n15518, new_n15504, new_n15571);
and_5  g13223(new_n15571, new_n15570_1, new_n15572);
xor_4  g13224(new_n15562, new_n15538, new_n15573_1);
xor_4  g13225(new_n15516, new_n15508_1, new_n15574);
and_5  g13226(new_n15574, new_n15573_1, new_n15575);
xor_4  g13227(new_n15574, new_n15573_1, new_n15576);
not_10 g13228(new_n15576, new_n15577);
xor_4  g13229(new_n15560, new_n15542, new_n15578);
not_10 g13230(new_n15578, new_n15579);
xor_4  g13231(new_n15514, new_n15511, new_n15580);
not_10 g13232(new_n15580, new_n15581);
nor_5  g13233(new_n15581, new_n15579, new_n15582);
xor_4  g13234(new_n15543, n17664, new_n15583);
xnor_4 g13235(new_n15583, new_n15557, new_n15584);
not_10 g13236(new_n15584, new_n15585);
nor_5  g13237(new_n15585, new_n13890, new_n15586);
not_10 g13238(new_n15586, new_n15587);
xor_4  g13239(new_n15585, new_n13890, new_n15588_1);
xnor_4 g13240(new_n15554, new_n15548, new_n15589);
and_5  g13241(new_n15589, new_n13910, new_n15590_1);
xor_4  g13242(new_n15554, new_n15548, new_n15591);
xnor_4 g13243(new_n15591, new_n13910, new_n15592);
xor_4  g13244(new_n15552, new_n15551, new_n15593);
nand_5 g13245(new_n15593, new_n13923_1, new_n15594);
nand_5 g13246(new_n15362, new_n13916, new_n15595);
xor_4  g13247(new_n15593, new_n13923_1, new_n15596);
nand_5 g13248(new_n15596, new_n15595, new_n15597);
and_5  g13249(new_n15597, new_n15594, new_n15598_1);
and_5  g13250(new_n15598_1, new_n15592, new_n15599);
nor_5  g13251(new_n15599, new_n15590_1, new_n15600);
and_5  g13252(new_n15600, new_n15588_1, new_n15601);
not_10 g13253(new_n15601, new_n15602_1);
and_5  g13254(new_n15602_1, new_n15587, new_n15603);
not_10 g13255(new_n15603, new_n15604);
xor_4  g13256(new_n15581, new_n15579, new_n15605);
and_5  g13257(new_n15605, new_n15604, new_n15606);
nor_5  g13258(new_n15606, new_n15582, new_n15607);
nor_5  g13259(new_n15607, new_n15577, new_n15608);
nor_5  g13260(new_n15608, new_n15575, new_n15609);
xor_4  g13261(new_n15571, new_n15570_1, new_n15610);
not_10 g13262(new_n15610, new_n15611);
nor_5  g13263(new_n15611, new_n15609, new_n15612);
nor_5  g13264(new_n15612, new_n15572, new_n15613);
xnor_4 g13265(new_n15613, new_n15569, n3263);
xnor_4 g13266(new_n12525, new_n12509, n3289);
xor_4  g13267(n21832, n5211, new_n15616);
nand_5 g13268(n26913, n12956, new_n15617);
or_5   g13269(n26913, n12956, new_n15618);
nor_5  g13270(n18295, n16223, new_n15619);
nor_5  g13271(new_n5057, new_n5052, new_n15620);
nor_5  g13272(new_n15620, new_n15619, new_n15621);
nand_5 g13273(new_n15621, new_n15618, new_n15622);
and_5  g13274(new_n15622, new_n15617, new_n15623);
xor_4  g13275(new_n15623, new_n15616, new_n15624);
xor_4  g13276(new_n15624, n18537, new_n15625);
not_10 g13277(new_n15625, new_n15626);
xor_4  g13278(n26913, n12956, new_n15627);
xor_4  g13279(new_n15627, new_n15621, new_n15628);
not_10 g13280(new_n15628, new_n15629);
or_5   g13281(new_n15629, n7057, new_n15630);
xor_4  g13282(new_n15629, n7057, new_n15631);
not_10 g13283(new_n15631, new_n15632);
or_5   g13284(new_n5058, n8381, new_n15633);
or_5   g13285(new_n5069, new_n5060_1, new_n15634);
and_5  g13286(new_n15634, new_n15633, new_n15635);
or_5   g13287(new_n15635, new_n15632, new_n15636_1);
and_5  g13288(new_n15636_1, new_n15630, new_n15637);
xor_4  g13289(new_n15637, new_n15626, new_n15638);
not_10 g13290(new_n15638, new_n15639);
xor_4  g13291(new_n14638, n21649, new_n15640);
nand_5 g13292(new_n9650, new_n5183, new_n15641);
xor_4  g13293(new_n9650, n18274, new_n15642);
or_5   g13294(new_n9668, n3828, new_n15643);
and_5  g13295(new_n9673, new_n5189, new_n15644);
nand_5 g13296(new_n9675, n21654, new_n15645);
xor_4  g13297(new_n9673, new_n5189, new_n15646);
and_5  g13298(new_n15646, new_n15645, new_n15647);
or_5   g13299(new_n15647, new_n15644, new_n15648);
xor_4  g13300(new_n9668, n3828, new_n15649);
nand_5 g13301(new_n15649, new_n15648, new_n15650);
and_5  g13302(new_n15650, new_n15643, new_n15651);
or_5   g13303(new_n15651, new_n15642, new_n15652_1);
and_5  g13304(new_n15652_1, new_n15641, new_n15653);
xor_4  g13305(new_n15653, new_n15640, new_n15654);
xor_4  g13306(new_n15654, new_n15639, new_n15655);
not_10 g13307(new_n15655, new_n15656);
xnor_4 g13308(new_n15635, new_n15631, new_n15657);
xor_4  g13309(new_n15651, new_n15642, new_n15658);
nand_5 g13310(new_n15658, new_n15657, new_n15659);
not_10 g13311(new_n15657, new_n15660);
xnor_4 g13312(new_n15658, new_n15660, new_n15661);
not_10 g13313(new_n15661, new_n15662_1);
xor_4  g13314(new_n15649, new_n15648, new_n15663);
nand_5 g13315(new_n15663, new_n5070, new_n15664);
xor_4  g13316(new_n15646, new_n15645, new_n15665);
nand_5 g13317(new_n15665, new_n5098_1, new_n15666);
xor_4  g13318(new_n9675, n21654, new_n15667);
and_5  g13319(new_n15667, new_n5100, new_n15668);
xor_4  g13320(new_n15665, new_n5098_1, new_n15669);
not_10 g13321(new_n15669, new_n15670);
or_5   g13322(new_n15670, new_n15668, new_n15671);
and_5  g13323(new_n15671, new_n15666, new_n15672);
xnor_4 g13324(new_n15663, new_n5071, new_n15673);
not_10 g13325(new_n15673, new_n15674);
or_5   g13326(new_n15674, new_n15672, new_n15675);
and_5  g13327(new_n15675, new_n15664, new_n15676);
or_5   g13328(new_n15676, new_n15662_1, new_n15677);
and_5  g13329(new_n15677, new_n15659, new_n15678);
xnor_4 g13330(new_n15678, new_n15656, n3301);
xor_4  g13331(new_n10929, n3030, new_n15680);
not_10 g13332(n19515, new_n15681);
or_5   g13333(new_n10923, new_n15681, new_n15682);
xor_4  g13334(new_n10923, n19515, new_n15683);
or_5   g13335(new_n10917, new_n13893, new_n15684);
xor_4  g13336(new_n10917, new_n13893, new_n15685);
or_5   g13337(new_n10910, n12209, new_n15686);
nand_5 g13338(new_n13670, new_n13669, new_n15687);
and_5  g13339(new_n15687, new_n15686, new_n15688);
nand_5 g13340(new_n15688, new_n15685, new_n15689);
and_5  g13341(new_n15689, new_n15684, new_n15690);
or_5   g13342(new_n15690, new_n15683, new_n15691);
and_5  g13343(new_n15691, new_n15682, new_n15692);
xor_4  g13344(new_n15692, new_n15680, new_n15693);
xor_4  g13345(new_n15693, new_n10211, new_n15694);
xor_4  g13346(new_n15690, new_n15683, new_n15695);
nand_5 g13347(new_n15695, new_n10217, new_n15696);
xor_4  g13348(new_n15695, new_n10217, new_n15697);
not_10 g13349(new_n15697, new_n15698);
xor_4  g13350(new_n15688, new_n15685, new_n15699);
nand_5 g13351(new_n15699, new_n10222, new_n15700);
xor_4  g13352(new_n15699, new_n10222, new_n15701);
not_10 g13353(new_n15701, new_n15702);
not_10 g13354(new_n13671, new_n15703);
nand_5 g13355(new_n15703, new_n10228, new_n15704);
or_5   g13356(new_n13673, new_n13667, new_n15705);
and_5  g13357(new_n15705, new_n15704, new_n15706);
or_5   g13358(new_n15706, new_n15702, new_n15707);
and_5  g13359(new_n15707, new_n15700, new_n15708);
or_5   g13360(new_n15708, new_n15698, new_n15709);
and_5  g13361(new_n15709, new_n15696, new_n15710);
xor_4  g13362(new_n15710, new_n15694, n3316);
xnor_4 g13363(new_n13657, new_n13644, n3332);
and_5  g13364(new_n8092, new_n7250, new_n15713);
xor_4  g13365(new_n8092, n17458, new_n15714);
or_5   g13366(new_n8098, n1222, new_n15715);
xor_4  g13367(new_n8098, new_n11171, new_n15716_1);
or_5   g13368(new_n8104, n25240, new_n15717);
or_5   g13369(new_n10740, new_n10721, new_n15718);
and_5  g13370(new_n15718, new_n15717, new_n15719);
or_5   g13371(new_n15719, new_n15716_1, new_n15720);
and_5  g13372(new_n15720, new_n15715, new_n15721);
nor_5  g13373(new_n15721, new_n15714, new_n15722);
nor_5  g13374(new_n15722, new_n15713, new_n15723);
nand_5 g13375(new_n15723, new_n8162, new_n15724);
nor_5  g13376(new_n13159, new_n15150, new_n15725);
nor_5  g13377(new_n13169, new_n13160, new_n15726);
or_5   g13378(new_n15726, new_n15725, new_n15727);
nor_5  g13379(n23166, n11898, new_n15728);
not_10 g13380(new_n15728, new_n15729);
and_5  g13381(new_n13158, new_n13151, new_n15730);
not_10 g13382(new_n15730, new_n15731);
and_5  g13383(new_n15731, new_n15729, new_n15732);
and_5  g13384(new_n15732, new_n15727, new_n15733);
not_10 g13385(new_n15733, new_n15734);
xor_4  g13386(new_n15734, new_n15724, new_n15735);
xor_4  g13387(new_n15723, new_n8162, new_n15736);
not_10 g13388(new_n15736, new_n15737);
xor_4  g13389(new_n15732, new_n15727, new_n15738);
and_5  g13390(new_n15738, new_n15737, new_n15739);
xor_4  g13391(new_n15738, new_n15737, new_n15740);
xor_4  g13392(new_n15721, new_n15714, new_n15741);
nor_5  g13393(new_n15741, new_n13170, new_n15742);
xor_4  g13394(new_n15741, new_n13170, new_n15743_1);
xor_4  g13395(new_n15719, new_n15716_1, new_n15744);
nand_5 g13396(new_n15744, new_n13174, new_n15745);
or_5   g13397(new_n10783, new_n10742, new_n15746);
nand_5 g13398(new_n10808, new_n10784, new_n15747);
and_5  g13399(new_n15747, new_n15746, new_n15748);
xor_4  g13400(new_n15744, new_n13174, new_n15749_1);
not_10 g13401(new_n15749_1, new_n15750);
or_5   g13402(new_n15750, new_n15748, new_n15751);
and_5  g13403(new_n15751, new_n15745, new_n15752);
and_5  g13404(new_n15752, new_n15743_1, new_n15753);
nor_5  g13405(new_n15753, new_n15742, new_n15754);
and_5  g13406(new_n15754, new_n15740, new_n15755);
nor_5  g13407(new_n15755, new_n15739, new_n15756);
xnor_4 g13408(new_n15756, new_n15735, n3340);
xor_4  g13409(n13851, n5077, new_n15758);
or_5   g13410(n24937, new_n10762, new_n15759);
xor_4  g13411(n24937, n15546, new_n15760);
or_5   g13412(new_n10766, n5098, new_n15761_1);
xor_4  g13413(n26452, n5098, new_n15762_1);
or_5   g13414(new_n4165_1, n3030, new_n15763);
xnor_4 g13415(n19905, n3030, new_n15764);
or_5   g13416(new_n15681, n17035, new_n15765);
or_5   g13417(new_n13905, new_n13892, new_n15766_1);
and_5  g13418(new_n15766_1, new_n15765, new_n15767);
nand_5 g13419(new_n15767, new_n15764, new_n15768);
and_5  g13420(new_n15768, new_n15763, new_n15769);
or_5   g13421(new_n15769, new_n15762_1, new_n15770);
and_5  g13422(new_n15770, new_n15761_1, new_n15771);
or_5   g13423(new_n15771, new_n15760, new_n15772);
and_5  g13424(new_n15772, new_n15759, new_n15773);
xor_4  g13425(new_n15773, new_n15758, new_n15774);
xnor_4 g13426(new_n15774, new_n15521, new_n15775);
xnor_4 g13427(new_n15771, new_n15760, new_n15776);
nand_5 g13428(new_n15776, new_n15571, new_n15777);
xor_4  g13429(new_n15771, new_n15760, new_n15778);
xnor_4 g13430(new_n15778, new_n15571, new_n15779);
not_10 g13431(new_n15779, new_n15780_1);
xnor_4 g13432(new_n15769, new_n15762_1, new_n15781);
nand_5 g13433(new_n15781, new_n15574, new_n15782);
xor_4  g13434(new_n15769, new_n15762_1, new_n15783);
xor_4  g13435(new_n15783, new_n15574, new_n15784);
xor_4  g13436(new_n15767, new_n15764, new_n15785);
and_5  g13437(new_n15785, new_n15581, new_n15786);
xor_4  g13438(new_n15785, new_n15581, new_n15787);
or_5   g13439(new_n13907, new_n13890, new_n15788);
or_5   g13440(new_n13929, new_n13909, new_n15789);
and_5  g13441(new_n15789, new_n15788, new_n15790);
and_5  g13442(new_n15790, new_n15787, new_n15791);
nor_5  g13443(new_n15791, new_n15786, new_n15792);
not_10 g13444(new_n15792, new_n15793_1);
or_5   g13445(new_n15793_1, new_n15784, new_n15794);
and_5  g13446(new_n15794, new_n15782, new_n15795);
or_5   g13447(new_n15795, new_n15780_1, new_n15796);
and_5  g13448(new_n15796, new_n15777, new_n15797);
xor_4  g13449(new_n15797, new_n15775, n3343);
and_5  g13450(new_n15527, new_n2600, new_n15799);
and_5  g13451(new_n15799, new_n2595, new_n15800);
and_5  g13452(new_n15800, new_n2557, new_n15801);
xor_4  g13453(new_n15800, new_n2557, new_n15802);
nor_5  g13454(new_n15802, n20040, new_n15803);
xor_4  g13455(new_n15799, new_n2595, new_n15804);
nor_5  g13456(new_n15804, n19531, new_n15805);
xor_4  g13457(new_n15804, n19531, new_n15806);
not_10 g13458(new_n15806, new_n15807);
or_5   g13459(new_n15528, n18345, new_n15808);
or_5   g13460(new_n15566, new_n15530, new_n15809);
and_5  g13461(new_n15809, new_n15808, new_n15810);
nor_5  g13462(new_n15810, new_n15807, new_n15811);
nor_5  g13463(new_n15811, new_n15805, new_n15812_1);
and_5  g13464(new_n15802, n20040, new_n15813);
nor_5  g13465(new_n15813, new_n15812_1, new_n15814);
nor_5  g13466(new_n15814, new_n15803, new_n15815_1);
nor_5  g13467(new_n15815_1, new_n15801, new_n15816_1);
xor_4  g13468(new_n15802, n20040, new_n15817);
xnor_4 g13469(new_n15817, new_n15812_1, new_n15818);
or_5   g13470(new_n15818, new_n14266, new_n15819);
and_5  g13471(new_n15818, new_n14266, new_n15820);
xor_4  g13472(new_n15810, new_n15807, new_n15821);
not_10 g13473(new_n15821, new_n15822);
and_5  g13474(new_n15822, new_n14247, new_n15823);
xor_4  g13475(new_n15822, new_n14247, new_n15824);
not_10 g13476(new_n15824, new_n15825);
not_10 g13477(new_n15567, new_n15826);
nand_5 g13478(new_n15826, new_n14251, new_n15827);
xor_4  g13479(new_n15826, new_n14251, new_n15828);
not_10 g13480(new_n15828, new_n15829);
not_10 g13481(new_n15570_1, new_n15830);
nand_5 g13482(new_n15830, new_n6510, new_n15831_1);
xor_4  g13483(new_n15830, new_n6510, new_n15832);
not_10 g13484(new_n15573_1, new_n15833);
nand_5 g13485(new_n15833, new_n6516, new_n15834);
and_5  g13486(new_n15579, new_n6521, new_n15835);
not_10 g13487(new_n15835, new_n15836);
xor_4  g13488(new_n15579, new_n6521, new_n15837);
nand_5 g13489(new_n15584, new_n6527, new_n15838);
xnor_4 g13490(new_n15584, new_n6526, new_n15839);
or_5   g13491(new_n15591, new_n6531, new_n15840);
xnor_4 g13492(new_n15591, new_n6530, new_n15841);
not_10 g13493(new_n6535, new_n15842);
nand_5 g13494(new_n15593, new_n15842, new_n15843);
and_5  g13495(new_n15362, n4939, new_n15844);
not_10 g13496(new_n15844, new_n15845);
xnor_4 g13497(new_n15593, new_n6535, new_n15846_1);
nand_5 g13498(new_n15846_1, new_n15845, new_n15847);
and_5  g13499(new_n15847, new_n15843, new_n15848);
nand_5 g13500(new_n15848, new_n15841, new_n15849);
and_5  g13501(new_n15849, new_n15840, new_n15850);
nand_5 g13502(new_n15850, new_n15839, new_n15851);
and_5  g13503(new_n15851, new_n15838, new_n15852);
and_5  g13504(new_n15852, new_n15837, new_n15853);
not_10 g13505(new_n15853, new_n15854);
and_5  g13506(new_n15854, new_n15836, new_n15855);
xor_4  g13507(new_n15833, new_n6517, new_n15856);
or_5   g13508(new_n15856, new_n15855, new_n15857);
nand_5 g13509(new_n15857, new_n15834, new_n15858);
nand_5 g13510(new_n15858, new_n15832, new_n15859_1);
and_5  g13511(new_n15859_1, new_n15831_1, new_n15860);
or_5   g13512(new_n15860, new_n15829, new_n15861);
and_5  g13513(new_n15861, new_n15827, new_n15862);
nor_5  g13514(new_n15862, new_n15825, new_n15863);
nor_5  g13515(new_n15863, new_n15823, new_n15864);
or_5   g13516(new_n15864, new_n15820, new_n15865);
and_5  g13517(new_n15865, new_n14288, new_n15866);
and_5  g13518(new_n15866, new_n15819, new_n15867);
xnor_4 g13519(new_n15867, new_n15816_1, new_n15868);
not_10 g13520(new_n15868, new_n15869_1);
not_10 g13521(new_n12598, new_n15870);
or_5   g13522(new_n12696, n10250, new_n15871);
xor_4  g13523(new_n12696, n10250, new_n15872);
not_10 g13524(new_n15872, new_n15873);
or_5   g13525(new_n12702_1, n7674, new_n15874);
xor_4  g13526(new_n12702_1, n7674, new_n15875);
not_10 g13527(new_n15875, new_n15876);
or_5   g13528(new_n12708, n6397, new_n15877);
xor_4  g13529(new_n12708, n6397, new_n15878);
not_10 g13530(new_n15878, new_n15879);
or_5   g13531(new_n12714, n19196, new_n15880);
xor_4  g13532(new_n12714, n19196, new_n15881);
not_10 g13533(new_n15881, new_n15882);
or_5   g13534(new_n12720, n23586, new_n15883);
xor_4  g13535(new_n12720, n23586, new_n15884_1);
not_10 g13536(new_n15884_1, new_n15885_1);
or_5   g13537(new_n12726, n21226, new_n15886);
xor_4  g13538(new_n12726, n21226, new_n15887);
not_10 g13539(new_n15887, new_n15888);
or_5   g13540(new_n12732, n4426, new_n15889_1);
xor_4  g13541(new_n12732, n4426, new_n15890);
not_10 g13542(new_n15890, new_n15891);
or_5   g13543(new_n12741, n20036, new_n15892);
xor_4  g13544(new_n12741, n20036, new_n15893);
nand_5 g13545(new_n12749, n11192, new_n15894);
or_5   g13546(new_n12745, n9380, new_n15895);
xor_4  g13547(new_n12749, n11192, new_n15896);
nand_5 g13548(new_n15896, new_n15895, new_n15897);
and_5  g13549(new_n15897, new_n15894, new_n15898);
nand_5 g13550(new_n15898, new_n15893, new_n15899);
and_5  g13551(new_n15899, new_n15892, new_n15900);
or_5   g13552(new_n15900, new_n15891, new_n15901);
and_5  g13553(new_n15901, new_n15889_1, new_n15902);
or_5   g13554(new_n15902, new_n15888, new_n15903);
and_5  g13555(new_n15903, new_n15886, new_n15904);
or_5   g13556(new_n15904, new_n15885_1, new_n15905);
and_5  g13557(new_n15905, new_n15883, new_n15906);
or_5   g13558(new_n15906, new_n15882, new_n15907);
and_5  g13559(new_n15907, new_n15880, new_n15908);
or_5   g13560(new_n15908, new_n15879, new_n15909);
and_5  g13561(new_n15909, new_n15877, new_n15910);
or_5   g13562(new_n15910, new_n15876, new_n15911);
and_5  g13563(new_n15911, new_n15874, new_n15912);
or_5   g13564(new_n15912, new_n15873, new_n15913);
and_5  g13565(new_n15913, new_n15871, new_n15914);
xor_4  g13566(new_n15914, new_n15870, new_n15915);
nor_5  g13567(new_n15915, new_n15869_1, new_n15916);
xor_4  g13568(new_n15912, new_n15873, new_n15917_1);
not_10 g13569(new_n15917_1, new_n15918_1);
xor_4  g13570(new_n15818, new_n14266, new_n15919);
xnor_4 g13571(new_n15919, new_n15864, new_n15920);
nor_5  g13572(new_n15920, new_n15918_1, new_n15921);
xor_4  g13573(new_n15920, new_n15918_1, new_n15922_1);
xor_4  g13574(new_n15910, new_n15876, new_n15923);
not_10 g13575(new_n15923, new_n15924);
xor_4  g13576(new_n15862, new_n15825, new_n15925);
nor_5  g13577(new_n15925, new_n15924, new_n15926);
not_10 g13578(new_n15925, new_n15927);
xnor_4 g13579(new_n15927, new_n15924, new_n15928);
xor_4  g13580(new_n15908, new_n15879, new_n15929);
not_10 g13581(new_n15929, new_n15930);
xnor_4 g13582(new_n15860, new_n15828, new_n15931);
nor_5  g13583(new_n15931, new_n15930, new_n15932);
not_10 g13584(new_n15931, new_n15933);
xnor_4 g13585(new_n15933, new_n15930, new_n15934);
xor_4  g13586(new_n15906, new_n15882, new_n15935);
not_10 g13587(new_n15935, new_n15936_1);
xor_4  g13588(new_n15858, new_n15832, new_n15937);
nor_5  g13589(new_n15937, new_n15936_1, new_n15938);
not_10 g13590(new_n15937, new_n15939);
xnor_4 g13591(new_n15939, new_n15936_1, new_n15940);
xor_4  g13592(new_n15904, new_n15885_1, new_n15941);
not_10 g13593(new_n15941, new_n15942);
xor_4  g13594(new_n15856, new_n15855, new_n15943);
nor_5  g13595(new_n15943, new_n15942, new_n15944);
xor_4  g13596(new_n15943, new_n15942, new_n15945);
xor_4  g13597(new_n15902, new_n15888, new_n15946);
not_10 g13598(new_n15946, new_n15947_1);
xor_4  g13599(new_n15852, new_n15837, new_n15948);
nor_5  g13600(new_n15948, new_n15947_1, new_n15949);
not_10 g13601(new_n15948, new_n15950);
xnor_4 g13602(new_n15950, new_n15947_1, new_n15951);
xor_4  g13603(new_n15900, new_n15891, new_n15952);
xor_4  g13604(new_n15850, new_n15839, new_n15953);
and_5  g13605(new_n15953, new_n15952, new_n15954);
xor_4  g13606(new_n15953, new_n15952, new_n15955);
xor_4  g13607(new_n15898, new_n15893, new_n15956_1);
not_10 g13608(new_n15956_1, new_n15957);
xor_4  g13609(new_n15848, new_n15841, new_n15958_1);
nor_5  g13610(new_n15958_1, new_n15957, new_n15959);
xor_4  g13611(new_n15846_1, new_n15845, new_n15960);
not_10 g13612(new_n15960, new_n15961);
xor_4  g13613(new_n15896, new_n15895, new_n15962);
and_5  g13614(new_n15962, new_n15961, new_n15963);
xor_4  g13615(new_n15362, new_n12618, new_n15964);
xor_4  g13616(new_n12745, n9380, new_n15965);
nor_5  g13617(new_n15965, new_n15964, new_n15966);
xor_4  g13618(new_n15962, new_n15961, new_n15967_1);
and_5  g13619(new_n15967_1, new_n15966, new_n15968);
nor_5  g13620(new_n15968, new_n15963, new_n15969);
not_10 g13621(new_n15958_1, new_n15970);
xnor_4 g13622(new_n15970, new_n15957, new_n15971);
and_5  g13623(new_n15971, new_n15969, new_n15972);
nor_5  g13624(new_n15972, new_n15959, new_n15973);
not_10 g13625(new_n15973, new_n15974);
and_5  g13626(new_n15974, new_n15955, new_n15975);
nor_5  g13627(new_n15975, new_n15954, new_n15976);
not_10 g13628(new_n15976, new_n15977);
and_5  g13629(new_n15977, new_n15951, new_n15978);
nor_5  g13630(new_n15978, new_n15949, new_n15979_1);
not_10 g13631(new_n15979_1, new_n15980);
and_5  g13632(new_n15980, new_n15945, new_n15981);
nor_5  g13633(new_n15981, new_n15944, new_n15982);
not_10 g13634(new_n15982, new_n15983);
and_5  g13635(new_n15983, new_n15940, new_n15984);
nor_5  g13636(new_n15984, new_n15938, new_n15985);
not_10 g13637(new_n15985, new_n15986_1);
and_5  g13638(new_n15986_1, new_n15934, new_n15987);
nor_5  g13639(new_n15987, new_n15932, new_n15988);
not_10 g13640(new_n15988, new_n15989);
and_5  g13641(new_n15989, new_n15928, new_n15990);
nor_5  g13642(new_n15990, new_n15926, new_n15991);
not_10 g13643(new_n15991, new_n15992);
and_5  g13644(new_n15992, new_n15922_1, new_n15993);
nor_5  g13645(new_n15993, new_n15921, new_n15994);
xor_4  g13646(new_n15915, new_n15869_1, new_n15995);
not_10 g13647(new_n15995, new_n15996);
nor_5  g13648(new_n15996, new_n15994, new_n15997);
nor_5  g13649(new_n15997, new_n15916, new_n15998);
not_10 g13650(new_n15816_1, new_n15999);
and_5  g13651(new_n15867, new_n15999, new_n16000);
and_5  g13652(new_n15914, new_n15870, new_n16001);
xnor_4 g13653(new_n16001, new_n16000, new_n16002);
xor_4  g13654(new_n16002, new_n15998, n3390);
not_10 g13655(new_n6616, new_n16004);
xor_4  g13656(new_n6617, new_n16004, n3426);
xor_4  g13657(new_n4749, new_n4747_1, n3451);
xnor_4 g13658(new_n12423, new_n12403, n3459);
not_10 g13659(new_n14011, new_n16008);
xor_4  g13660(n6773, n583, new_n16009);
xor_4  g13661(new_n16009, new_n12439, new_n16010);
nor_5  g13662(new_n16010, new_n16008, new_n16011);
nor_5  g13663(new_n16009, new_n12439, new_n16012);
or_5   g13664(new_n16012, n6729, new_n16013_1);
nand_5 g13665(n21687, n6729, new_n16014);
or_5   g13666(new_n16009, new_n16014, new_n16015);
and_5  g13667(new_n16015, new_n16013_1, new_n16016);
nand_5 g13668(n6773, n583, new_n16017);
xor_4  g13669(n22173, n17090, new_n16018);
xor_4  g13670(new_n16018, new_n16017, new_n16019);
xor_4  g13671(new_n16019, new_n16016, new_n16020);
xor_4  g13672(new_n16020, new_n14007, new_n16021);
xor_4  g13673(new_n16021, new_n16011, n3502);
xnor_4 g13674(new_n11066, new_n11025_1, n3516);
not_10 g13675(n18145, new_n16024);
not_10 g13676(n10712, new_n16025);
not_10 g13677(n25126, new_n16026);
not_10 g13678(n19608, new_n16027);
not_10 g13679(n1689, new_n16028);
nor_5  g13680(n24129, n22274, new_n16029_1);
and_5  g13681(new_n16029_1, new_n16028, new_n16030);
and_5  g13682(new_n16030, new_n16027, new_n16031);
and_5  g13683(new_n16031, new_n16026, new_n16032);
and_5  g13684(new_n16032, new_n16025, new_n16033);
xor_4  g13685(new_n16033, new_n16024, new_n16034);
xor_4  g13686(new_n16034, n15761, new_n16035);
xor_4  g13687(new_n16032, new_n16025, new_n16036);
or_5   g13688(new_n16036, new_n10479, new_n16037);
xor_4  g13689(new_n16036, n11201, new_n16038);
xor_4  g13690(new_n16031, new_n16026, new_n16039);
or_5   g13691(new_n16039, new_n10482, new_n16040);
xor_4  g13692(new_n16039, n18690, new_n16041);
xor_4  g13693(new_n16030, new_n16027, new_n16042);
or_5   g13694(new_n16042, new_n10485, new_n16043);
xor_4  g13695(new_n16042, n12153, new_n16044);
not_10 g13696(n13044, new_n16045);
xor_4  g13697(new_n16029_1, new_n16028, new_n16046);
or_5   g13698(new_n16046, new_n16045, new_n16047);
xor_4  g13699(new_n16046, n13044, new_n16048);
not_10 g13700(n18745, new_n16049);
xor_4  g13701(n24129, n22274, new_n16050);
or_5   g13702(new_n16050, new_n16049, new_n16051);
nor_5  g13703(n24129, new_n5858, new_n16052);
xor_4  g13704(new_n16050, new_n16049, new_n16053);
nand_5 g13705(new_n16053, new_n16052, new_n16054);
and_5  g13706(new_n16054, new_n16051, new_n16055);
or_5   g13707(new_n16055, new_n16048, new_n16056);
and_5  g13708(new_n16056, new_n16047, new_n16057);
or_5   g13709(new_n16057, new_n16044, new_n16058);
and_5  g13710(new_n16058, new_n16043, new_n16059);
or_5   g13711(new_n16059, new_n16041, new_n16060_1);
and_5  g13712(new_n16060_1, new_n16040, new_n16061);
or_5   g13713(new_n16061, new_n16038, new_n16062_1);
and_5  g13714(new_n16062_1, new_n16037, new_n16063);
xor_4  g13715(new_n16063, new_n16035, new_n16064);
xnor_4 g13716(new_n16064, new_n6884, new_n16065);
xor_4  g13717(new_n16061, new_n16038, new_n16066);
nand_5 g13718(new_n16066, new_n6889, new_n16067);
xnor_4 g13719(new_n16066, new_n6889, new_n16068_1);
xor_4  g13720(new_n16059, new_n16041, new_n16069);
nand_5 g13721(new_n16069, new_n6894, new_n16070);
xnor_4 g13722(new_n16069, new_n6894, new_n16071);
xor_4  g13723(new_n16057, new_n16044, new_n16072);
nand_5 g13724(new_n16072, new_n6900, new_n16073);
xnor_4 g13725(new_n16072, new_n6899, new_n16074);
xor_4  g13726(new_n16055, new_n16048, new_n16075);
or_5   g13727(new_n16075, new_n4120, new_n16076);
xnor_4 g13728(new_n16075, new_n4120, new_n16077);
xor_4  g13729(new_n16053, new_n16052, new_n16078);
or_5   g13730(new_n16078, new_n4131, new_n16079);
xnor_4 g13731(n24129, n16167, new_n16080_1);
nor_5  g13732(new_n16080_1, new_n4136, new_n16081);
xor_4  g13733(new_n16078, new_n4131, new_n16082);
nand_5 g13734(new_n16082, new_n16081, new_n16083);
and_5  g13735(new_n16083, new_n16079, new_n16084);
or_5   g13736(new_n16084, new_n16077, new_n16085);
and_5  g13737(new_n16085, new_n16076, new_n16086);
nand_5 g13738(new_n16086, new_n16074, new_n16087);
and_5  g13739(new_n16087, new_n16073, new_n16088);
or_5   g13740(new_n16088, new_n16071, new_n16089);
and_5  g13741(new_n16089, new_n16070, new_n16090);
or_5   g13742(new_n16090, new_n16068_1, new_n16091);
and_5  g13743(new_n16091, new_n16067, new_n16092);
xor_4  g13744(new_n16092, new_n16065, new_n16093);
xor_4  g13745(new_n16093, new_n10603, new_n16094);
xor_4  g13746(new_n16090, new_n16068_1, new_n16095);
nand_5 g13747(new_n16095, new_n10608, new_n16096);
xor_4  g13748(new_n16095, new_n10608, new_n16097);
not_10 g13749(new_n16097, new_n16098_1);
xor_4  g13750(new_n16088, new_n16071, new_n16099);
nand_5 g13751(new_n16099, new_n10614_1, new_n16100);
xor_4  g13752(new_n16099, new_n10614_1, new_n16101);
not_10 g13753(new_n16101, new_n16102);
xor_4  g13754(new_n16086, new_n16074, new_n16103);
nand_5 g13755(new_n16103, new_n10621, new_n16104);
xor_4  g13756(new_n16084, new_n16077, new_n16105);
or_5   g13757(new_n16105, new_n10624, new_n16106);
xor_4  g13758(new_n16105, new_n10624, new_n16107);
not_10 g13759(new_n16107, new_n16108);
xor_4  g13760(new_n16082, new_n16081, new_n16109);
or_5   g13761(new_n16109, new_n5870, new_n16110_1);
xnor_4 g13762(new_n16080_1, new_n4135, new_n16111);
and_5  g13763(new_n16111, new_n5856, new_n16112);
xor_4  g13764(new_n16109, new_n5870, new_n16113);
not_10 g13765(new_n16113, new_n16114);
or_5   g13766(new_n16114, new_n16112, new_n16115);
and_5  g13767(new_n16115, new_n16110_1, new_n16116);
or_5   g13768(new_n16116, new_n16108, new_n16117);
and_5  g13769(new_n16117, new_n16106, new_n16118);
xnor_4 g13770(new_n16103, new_n10619, new_n16119);
not_10 g13771(new_n16119, new_n16120);
or_5   g13772(new_n16120, new_n16118, new_n16121);
and_5  g13773(new_n16121, new_n16104, new_n16122);
or_5   g13774(new_n16122, new_n16102, new_n16123);
and_5  g13775(new_n16123, new_n16100, new_n16124);
or_5   g13776(new_n16124, new_n16098_1, new_n16125);
and_5  g13777(new_n16125, new_n16096, new_n16126);
xor_4  g13778(new_n16126, new_n16094, n3528);
xor_4  g13779(new_n9286, new_n9204, n3555);
and_5  g13780(new_n2709, new_n2666, new_n16129);
nor_5  g13781(new_n2773, new_n2711_1, new_n16130);
nor_5  g13782(new_n16130, new_n16129, new_n16131);
not_10 g13783(new_n16131, new_n16132);
nand_5 g13784(new_n2665, new_n2650, new_n16133);
nor_5  g13785(new_n10338, new_n16133, new_n16134);
and_5  g13786(new_n16134, new_n16132, new_n16135);
and_5  g13787(new_n10338, new_n16133, new_n16136);
and_5  g13788(new_n16136, new_n16131, new_n16137);
nor_5  g13789(new_n16137, new_n16135, new_n16138);
nor_5  g13790(new_n16138, new_n14946, new_n16139);
xor_4  g13791(new_n16138, new_n14947, new_n16140);
xnor_4 g13792(new_n10338, new_n16133, new_n16141);
xor_4  g13793(new_n16141, new_n16132, new_n16142_1);
nor_5  g13794(new_n16142_1, new_n14951, new_n16143);
xor_4  g13795(new_n16142_1, new_n14951, new_n16144);
not_10 g13796(new_n16144, new_n16145);
nor_5  g13797(new_n2774_1, new_n2649, new_n16146);
not_10 g13798(new_n16146, new_n16147);
and_5  g13799(new_n2833, new_n2775, new_n16148);
not_10 g13800(new_n16148, new_n16149);
and_5  g13801(new_n16149, new_n16147, new_n16150);
nor_5  g13802(new_n16150, new_n16145, new_n16151);
nor_5  g13803(new_n16151, new_n16143, new_n16152);
nor_5  g13804(new_n16152, new_n16140, new_n16153);
nor_5  g13805(new_n16153, new_n16139, new_n16154);
nor_5  g13806(new_n16154, new_n16135, n3561);
xnor_4 g13807(n16439, n14680, new_n16156);
not_10 g13808(new_n16156, new_n16157);
nand_5 g13809(n17250, new_n4364, new_n16158_1);
or_5   g13810(new_n10831, new_n10811, new_n16159);
and_5  g13811(new_n16159, new_n16158_1, new_n16160);
xor_4  g13812(new_n16160, new_n16157, new_n16161);
not_10 g13813(new_n16161, new_n16162);
not_10 g13814(n1654, new_n16163);
xor_4  g13815(new_n9860, new_n16163, new_n16164);
or_5   g13816(new_n9863, n13783, new_n16165);
or_5   g13817(new_n10846, new_n10835, new_n16166);
and_5  g13818(new_n16166, new_n16165, new_n16167_1);
xor_4  g13819(new_n16167_1, new_n16164, new_n16168);
xnor_4 g13820(new_n16168, new_n16162, new_n16169);
or_5   g13821(new_n10847, new_n10833, new_n16170);
or_5   g13822(new_n10878, new_n10848, new_n16171);
and_5  g13823(new_n16171, new_n16170, new_n16172);
xor_4  g13824(new_n16172, new_n16169, new_n16173);
xnor_4 g13825(new_n16173, new_n5667, new_n16174);
nand_5 g13826(new_n10879, new_n5672, new_n16175);
nand_5 g13827(new_n10904, new_n10880, new_n16176);
and_5  g13828(new_n16176, new_n16175, new_n16177);
xor_4  g13829(new_n16177, new_n16174, n3563);
xor_4  g13830(new_n6170, new_n6169, n3617);
xor_4  g13831(n22253, n8305, new_n16180);
not_10 g13832(n1255, new_n16181);
or_5   g13833(n12861, new_n16181, new_n16182);
xor_4  g13834(n12861, n1255, new_n16183);
not_10 g13835(n9512, new_n16184);
or_5   g13836(n13333, new_n16184, new_n16185_1);
xor_4  g13837(n13333, n9512, new_n16186);
not_10 g13838(n16608, new_n16187);
or_5   g13839(new_n16187, n2210, new_n16188);
and_5  g13840(n21735, new_n12953, new_n16189);
nor_5  g13841(new_n4637, new_n4612, new_n16190);
or_5   g13842(new_n16190, new_n16189, new_n16191);
xnor_4 g13843(n16608, n2210, new_n16192);
nand_5 g13844(new_n16192, new_n16191, new_n16193);
and_5  g13845(new_n16193, new_n16188, new_n16194);
or_5   g13846(new_n16194, new_n16186, new_n16195);
and_5  g13847(new_n16195, new_n16185_1, new_n16196_1);
or_5   g13848(new_n16196_1, new_n16183, new_n16197);
and_5  g13849(new_n16197, new_n16182, new_n16198);
xor_4  g13850(new_n16198, new_n16180, new_n16199);
xor_4  g13851(new_n16199, new_n11545, new_n16200);
xor_4  g13852(new_n16196_1, new_n16183, new_n16201);
or_5   g13853(new_n16201, new_n11548_1, new_n16202);
xor_4  g13854(new_n16201, new_n11548_1, new_n16203);
not_10 g13855(new_n16203, new_n16204);
xor_4  g13856(new_n16194, new_n16186, new_n16205);
or_5   g13857(new_n16205, new_n11554, new_n16206_1);
xor_4  g13858(new_n16192, new_n16191, new_n16207);
and_5  g13859(new_n16207, new_n11557, new_n16208);
xnor_4 g13860(new_n16207, new_n11557, new_n16209);
nand_5 g13861(new_n4731_1, new_n4638, new_n16210);
nand_5 g13862(new_n4767, new_n4732, new_n16211);
and_5  g13863(new_n16211, new_n16210, new_n16212);
nor_5  g13864(new_n16212, new_n16209, new_n16213);
nor_5  g13865(new_n16213, new_n16208, new_n16214);
xor_4  g13866(new_n16205, new_n11554, new_n16215_1);
nand_5 g13867(new_n16215_1, new_n16214, new_n16216);
and_5  g13868(new_n16216, new_n16206_1, new_n16217_1);
or_5   g13869(new_n16217_1, new_n16204, new_n16218_1);
and_5  g13870(new_n16218_1, new_n16202, new_n16219_1);
xor_4  g13871(new_n16219_1, new_n16200, n3642);
xnor_4 g13872(n16544, n4319, new_n16221);
or_5   g13873(n23463, n6814, new_n16222);
xnor_4 g13874(n23463, n6814, new_n16223_1);
or_5   g13875(n19701, n13074, new_n16224);
xnor_4 g13876(n19701, n13074, new_n16225);
or_5   g13877(n23529, n10739, new_n16226);
xnor_4 g13878(n23529, n10739, new_n16227);
or_5   g13879(n24620, n21753, new_n16228);
xnor_4 g13880(n24620, n21753, new_n16229);
or_5   g13881(n21832, n5211, new_n16230_1);
nand_5 g13882(new_n15623, new_n15616, new_n16231);
and_5  g13883(new_n16231, new_n16230_1, new_n16232);
or_5   g13884(new_n16232, new_n16229, new_n16233);
and_5  g13885(new_n16233, new_n16228, new_n16234);
or_5   g13886(new_n16234, new_n16227, new_n16235);
and_5  g13887(new_n16235, new_n16226, new_n16236);
or_5   g13888(new_n16236, new_n16225, new_n16237);
and_5  g13889(new_n16237, new_n16224, new_n16238);
or_5   g13890(new_n16238, new_n16223_1, new_n16239);
and_5  g13891(new_n16239, new_n16222, new_n16240);
xor_4  g13892(new_n16240, new_n16221, new_n16241);
xor_4  g13893(new_n16241, n3324, new_n16242);
not_10 g13894(new_n16242, new_n16243_1);
xor_4  g13895(new_n16238, new_n16223_1, new_n16244);
or_5   g13896(new_n16244, n17911, new_n16245);
xor_4  g13897(new_n16244, n17911, new_n16246);
not_10 g13898(new_n16246, new_n16247_1);
xor_4  g13899(new_n16236, new_n16225, new_n16248);
or_5   g13900(new_n16248, n21997, new_n16249);
xor_4  g13901(new_n16248, n21997, new_n16250);
not_10 g13902(new_n16250, new_n16251);
xor_4  g13903(new_n16234, new_n16227, new_n16252);
or_5   g13904(new_n16252, n25119, new_n16253);
xor_4  g13905(new_n16252, n25119, new_n16254);
xor_4  g13906(new_n16232, new_n16229, new_n16255);
nand_5 g13907(new_n16255, n1163, new_n16256);
or_5   g13908(new_n15624, n18537, new_n16257);
or_5   g13909(new_n15637, new_n15626, new_n16258);
and_5  g13910(new_n16258, new_n16257, new_n16259);
xor_4  g13911(new_n16255, n1163, new_n16260);
nand_5 g13912(new_n16260, new_n16259, new_n16261);
and_5  g13913(new_n16261, new_n16256, new_n16262);
nand_5 g13914(new_n16262, new_n16254, new_n16263);
and_5  g13915(new_n16263, new_n16253, new_n16264);
or_5   g13916(new_n16264, new_n16251, new_n16265);
and_5  g13917(new_n16265, new_n16249, new_n16266);
or_5   g13918(new_n16266, new_n16247_1, new_n16267);
and_5  g13919(new_n16267, new_n16245, new_n16268);
xor_4  g13920(new_n16268, new_n16243_1, new_n16269);
not_10 g13921(new_n16269, new_n16270);
xor_4  g13922(n23250, n16507, new_n16271);
not_10 g13923(n11455, new_n16272);
or_5   g13924(n22470, new_n16272, new_n16273);
xor_4  g13925(n22470, n11455, new_n16274);
not_10 g13926(n3945, new_n16275_1);
or_5   g13927(n19116, new_n16275_1, new_n16276);
xor_4  g13928(n19116, n3945, new_n16277);
not_10 g13929(n5255, new_n16278);
or_5   g13930(n6861, new_n16278, new_n16279_1);
xor_4  g13931(n6861, n5255, new_n16280);
or_5   g13932(new_n5179, n19357, new_n16281);
xor_4  g13933(n21649, n19357, new_n16282);
or_5   g13934(new_n5183, n2328, new_n16283);
nand_5 g13935(n15053, new_n5187, new_n16284);
or_5   g13936(new_n5090, new_n5086, new_n16285);
and_5  g13937(new_n16285, new_n16284, new_n16286);
xnor_4 g13938(n18274, n2328, new_n16287);
nand_5 g13939(new_n16287, new_n16286, new_n16288);
and_5  g13940(new_n16288, new_n16283, new_n16289);
or_5   g13941(new_n16289, new_n16282, new_n16290);
and_5  g13942(new_n16290, new_n16281, new_n16291);
or_5   g13943(new_n16291, new_n16280, new_n16292);
and_5  g13944(new_n16292, new_n16279_1, new_n16293);
or_5   g13945(new_n16293, new_n16277, new_n16294);
and_5  g13946(new_n16294, new_n16276, new_n16295);
or_5   g13947(new_n16295, new_n16274, new_n16296);
and_5  g13948(new_n16296, new_n16273, new_n16297);
xor_4  g13949(new_n16297, new_n16271, new_n16298);
or_5   g13950(new_n16298, n4967, new_n16299);
not_10 g13951(n4967, new_n16300);
xor_4  g13952(new_n16298, new_n16300, new_n16301);
xor_4  g13953(new_n16295, new_n16274, new_n16302);
or_5   g13954(new_n16302, n15602, new_n16303);
xor_4  g13955(new_n16293, new_n16277, new_n16304);
nand_5 g13956(new_n16304, n8694, new_n16305);
xor_4  g13957(new_n16291, new_n16280, new_n16306);
or_5   g13958(new_n16306, n12380, new_n16307);
not_10 g13959(n12380, new_n16308);
xor_4  g13960(new_n16306, new_n16308, new_n16309);
xor_4  g13961(new_n16289, new_n16282, new_n16310);
or_5   g13962(new_n16310, n8943, new_n16311);
not_10 g13963(n8943, new_n16312);
xor_4  g13964(new_n16310, new_n16312, new_n16313);
not_10 g13965(new_n16313, new_n16314);
xor_4  g13966(new_n16287, new_n16286, new_n16315);
nand_5 g13967(new_n16315, n8255, new_n16316);
nor_5  g13968(new_n5091, new_n5085, new_n16317);
and_5  g13969(new_n5092, new_n5084, new_n16318);
or_5   g13970(new_n16318, new_n16317, new_n16319);
not_10 g13971(new_n16315, new_n16320);
xnor_4 g13972(new_n16320, n8255, new_n16321);
nand_5 g13973(new_n16321, new_n16319, new_n16322_1);
and_5  g13974(new_n16322_1, new_n16316, new_n16323);
nand_5 g13975(new_n16323, new_n16314, new_n16324);
and_5  g13976(new_n16324, new_n16311, new_n16325);
or_5   g13977(new_n16325, new_n16309, new_n16326);
and_5  g13978(new_n16326, new_n16307, new_n16327_1);
not_10 g13979(n8694, new_n16328);
xor_4  g13980(new_n16304, new_n16328, new_n16329);
not_10 g13981(new_n16329, new_n16330);
nand_5 g13982(new_n16330, new_n16327_1, new_n16331);
and_5  g13983(new_n16331, new_n16305, new_n16332);
xor_4  g13984(new_n16302, n15602, new_n16333);
nand_5 g13985(new_n16333, new_n16332, new_n16334);
and_5  g13986(new_n16334, new_n16303, new_n16335);
or_5   g13987(new_n16335, new_n16301, new_n16336);
and_5  g13988(new_n16336, new_n16299, new_n16337);
not_10 g13989(n13419, new_n16338);
xor_4  g13990(n6659, n5101, new_n16339);
not_10 g13991(n23250, new_n16340);
or_5   g13992(new_n16340, n16507, new_n16341);
or_5   g13993(new_n16297, new_n16271, new_n16342);
and_5  g13994(new_n16342, new_n16341, new_n16343);
xor_4  g13995(new_n16343, new_n16339, new_n16344);
xor_4  g13996(new_n16344, new_n16338, new_n16345);
xor_4  g13997(new_n16345, new_n16337, new_n16346);
xnor_4 g13998(new_n16346, new_n16270, new_n16347);
xor_4  g13999(new_n16266, new_n16247_1, new_n16348);
xor_4  g14000(new_n16335, new_n16301, new_n16349);
nand_5 g14001(new_n16349, new_n16348, new_n16350_1);
not_10 g14002(new_n16348, new_n16351);
xnor_4 g14003(new_n16349, new_n16351, new_n16352);
not_10 g14004(new_n16352, new_n16353);
xor_4  g14005(new_n16264, new_n16251, new_n16354);
xor_4  g14006(new_n16333, new_n16332, new_n16355);
nand_5 g14007(new_n16355, new_n16354, new_n16356);
not_10 g14008(new_n16354, new_n16357);
xnor_4 g14009(new_n16355, new_n16357, new_n16358);
not_10 g14010(new_n16358, new_n16359);
xor_4  g14011(new_n16262, new_n16254, new_n16360);
not_10 g14012(new_n16360, new_n16361);
xor_4  g14013(new_n16330, new_n16327_1, new_n16362);
or_5   g14014(new_n16362, new_n16361, new_n16363);
xor_4  g14015(new_n16362, new_n16361, new_n16364);
not_10 g14016(new_n16364, new_n16365);
xor_4  g14017(new_n16325, new_n16309, new_n16366);
not_10 g14018(new_n16366, new_n16367_1);
xor_4  g14019(new_n16260, new_n16259, new_n16368);
or_5   g14020(new_n16368, new_n16367_1, new_n16369);
xor_4  g14021(new_n16368, new_n16367_1, new_n16370);
xor_4  g14022(new_n16323, new_n16314, new_n16371);
nand_5 g14023(new_n16371, new_n15638, new_n16372);
xnor_4 g14024(new_n16371, new_n15639, new_n16373);
not_10 g14025(new_n16373, new_n16374);
xor_4  g14026(new_n16321, new_n16319, new_n16375);
or_5   g14027(new_n16375, new_n15660, new_n16376_1);
xor_4  g14028(new_n16375, new_n15660, new_n16377);
not_10 g14029(new_n16377, new_n16378);
or_5   g14030(new_n5093, new_n5071, new_n16379_1);
or_5   g14031(new_n5105, new_n5095, new_n16380);
and_5  g14032(new_n16380, new_n16379_1, new_n16381);
or_5   g14033(new_n16381, new_n16378, new_n16382);
and_5  g14034(new_n16382, new_n16376_1, new_n16383);
or_5   g14035(new_n16383, new_n16374, new_n16384);
nand_5 g14036(new_n16384, new_n16372, new_n16385);
nand_5 g14037(new_n16385, new_n16370, new_n16386);
and_5  g14038(new_n16386, new_n16369, new_n16387);
or_5   g14039(new_n16387, new_n16365, new_n16388);
and_5  g14040(new_n16388, new_n16363, new_n16389);
or_5   g14041(new_n16389, new_n16359, new_n16390);
and_5  g14042(new_n16390, new_n16356, new_n16391);
or_5   g14043(new_n16391, new_n16353, new_n16392);
and_5  g14044(new_n16392, new_n16350_1, new_n16393);
xor_4  g14045(new_n16393, new_n16347, n3649);
nor_5  g14046(n26625, n14230, new_n16395);
and_5  g14047(new_n16395, new_n11774, new_n16396_1);
and_5  g14048(new_n16396_1, new_n11771_1, new_n16397);
and_5  g14049(new_n16397, new_n11768, new_n16398_1);
and_5  g14050(new_n16398_1, new_n11765, new_n16399);
xor_4  g14051(new_n16399, new_n11762, new_n16400);
xor_4  g14052(new_n16400, n26191, new_n16401);
xor_4  g14053(new_n16398_1, new_n11765, new_n16402);
nand_5 g14054(new_n16402, new_n11663, new_n16403);
xor_4  g14055(new_n16402, n26512, new_n16404);
xor_4  g14056(new_n16397, new_n11768, new_n16405);
nand_5 g14057(new_n16405, new_n9738, new_n16406_1);
xor_4  g14058(new_n16405, n19575, new_n16407_1);
xor_4  g14059(new_n16396_1, new_n11771_1, new_n16408);
nand_5 g14060(new_n16408, new_n9739, new_n16409);
xor_4  g14061(new_n16408, n15378, new_n16410);
xor_4  g14062(new_n16395, new_n11774, new_n16411);
nand_5 g14063(new_n16411, new_n9740, new_n16412);
not_10 g14064(n22591, new_n16413);
xor_4  g14065(n26625, n14230, new_n16414);
or_5   g14066(new_n16414, new_n16413, new_n16415);
and_5  g14067(n26167, new_n6630_1, new_n16416);
xor_4  g14068(new_n16414, new_n16413, new_n16417);
nand_5 g14069(new_n16417, new_n16416, new_n16418);
and_5  g14070(new_n16418, new_n16415, new_n16419_1);
xor_4  g14071(new_n16411, new_n9740, new_n16420);
nand_5 g14072(new_n16420, new_n16419_1, new_n16421);
and_5  g14073(new_n16421, new_n16412, new_n16422);
or_5   g14074(new_n16422, new_n16410, new_n16423);
and_5  g14075(new_n16423, new_n16409, new_n16424_1);
or_5   g14076(new_n16424_1, new_n16407_1, new_n16425);
and_5  g14077(new_n16425, new_n16406_1, new_n16426);
or_5   g14078(new_n16426, new_n16404, new_n16427);
and_5  g14079(new_n16427, new_n16403, new_n16428_1);
xor_4  g14080(new_n16428_1, new_n16401, new_n16429);
xor_4  g14081(new_n16429, n7917, new_n16430);
xor_4  g14082(new_n16426, new_n16404, new_n16431);
nand_5 g14083(new_n16431, new_n14766, new_n16432);
xor_4  g14084(new_n16431, new_n14766, new_n16433_1);
xor_4  g14085(new_n16424_1, new_n16407_1, new_n16434);
or_5   g14086(new_n16434, new_n14769, new_n16435);
xor_4  g14087(new_n16434, n2013, new_n16436);
not_10 g14088(n23755, new_n16437);
xor_4  g14089(new_n16422, new_n16410, new_n16438);
or_5   g14090(new_n16438, new_n16437, new_n16439_1);
xor_4  g14091(new_n16438, n23755, new_n16440_1);
xor_4  g14092(new_n16420, new_n16419_1, new_n16441);
or_5   g14093(new_n16441, new_n14773, new_n16442);
xor_4  g14094(new_n16441, n19163, new_n16443);
xor_4  g14095(new_n16417, new_n16416, new_n16444);
nand_5 g14096(new_n16444, n22358, new_n16445_1);
or_5   g14097(new_n16444, n22358, new_n16446);
xnor_4 g14098(n26167, n14230, new_n16447);
and_5  g14099(new_n16447, n9646, new_n16448);
nand_5 g14100(new_n16448, new_n16446, new_n16449);
and_5  g14101(new_n16449, new_n16445_1, new_n16450);
or_5   g14102(new_n16450, new_n16443, new_n16451);
and_5  g14103(new_n16451, new_n16442, new_n16452);
or_5   g14104(new_n16452, new_n16440_1, new_n16453);
and_5  g14105(new_n16453, new_n16439_1, new_n16454);
or_5   g14106(new_n16454, new_n16436, new_n16455);
and_5  g14107(new_n16455, new_n16435, new_n16456);
nand_5 g14108(new_n16456, new_n16433_1, new_n16457);
and_5  g14109(new_n16457, new_n16432, new_n16458);
xor_4  g14110(new_n16458, new_n16430, new_n16459);
xor_4  g14111(new_n16459, new_n6934, new_n16460_1);
xor_4  g14112(new_n16456, new_n16433_1, new_n16461);
or_5   g14113(new_n16461, new_n6940, new_n16462);
xor_4  g14114(new_n16461, new_n6940, new_n16463);
not_10 g14115(new_n16463, new_n16464);
xor_4  g14116(new_n16454, new_n16436, new_n16465);
nand_5 g14117(new_n16465, new_n6944, new_n16466);
xor_4  g14118(new_n16465, new_n6944, new_n16467);
not_10 g14119(new_n16467, new_n16468);
xor_4  g14120(new_n16452, new_n16440_1, new_n16469);
nand_5 g14121(new_n16469, new_n6949, new_n16470);
xor_4  g14122(new_n16469, new_n6949, new_n16471);
not_10 g14123(new_n16471, new_n16472);
xor_4  g14124(new_n16450, new_n16443, new_n16473);
nand_5 g14125(new_n16473, new_n6959, new_n16474);
xnor_4 g14126(new_n16473, new_n6956, new_n16475);
xor_4  g14127(new_n16444, n22358, new_n16476_1);
xor_4  g14128(new_n16476_1, new_n16448, new_n16477);
nor_5  g14129(new_n16477, new_n6963, new_n16478);
xor_4  g14130(new_n16447, n9646, new_n16479);
nor_5  g14131(new_n16479, new_n6967_1, new_n16480);
xor_4  g14132(new_n16477, new_n6963, new_n16481_1);
and_5  g14133(new_n16481_1, new_n16480, new_n16482_1);
nor_5  g14134(new_n16482_1, new_n16478, new_n16483);
nand_5 g14135(new_n16483, new_n16475, new_n16484);
and_5  g14136(new_n16484, new_n16474, new_n16485);
or_5   g14137(new_n16485, new_n16472, new_n16486);
and_5  g14138(new_n16486, new_n16470, new_n16487);
or_5   g14139(new_n16487, new_n16468, new_n16488);
and_5  g14140(new_n16488, new_n16466, new_n16489);
or_5   g14141(new_n16489, new_n16464, new_n16490);
and_5  g14142(new_n16490, new_n16462, new_n16491);
xor_4  g14143(new_n16491, new_n16460_1, n3665);
xor_4  g14144(new_n5859, new_n5857, n3679);
nor_5  g14145(n16521, n7139, new_n16494);
and_5  g14146(new_n16494, new_n3558, new_n16495);
and_5  g14147(new_n16495, new_n3553, new_n16496);
and_5  g14148(new_n16496, new_n3549, new_n16497);
and_5  g14149(new_n16497, new_n3545, new_n16498);
and_5  g14150(new_n16498, new_n3541_1, new_n16499);
and_5  g14151(new_n16499, new_n3537, new_n16500);
xor_4  g14152(new_n16500, new_n3533, new_n16501);
xnor_4 g14153(new_n16501, new_n5972, new_n16502_1);
xor_4  g14154(new_n16499, new_n3537, new_n16503);
nand_5 g14155(new_n16503, new_n5975, new_n16504);
xnor_4 g14156(new_n16503, new_n5977, new_n16505);
xor_4  g14157(new_n16498, new_n3541_1, new_n16506_1);
or_5   g14158(new_n16506_1, new_n5981, new_n16507_1);
xor_4  g14159(new_n16506_1, new_n5983, new_n16508);
xor_4  g14160(new_n16497, new_n3545, new_n16509);
or_5   g14161(new_n16509, new_n5987, new_n16510);
xor_4  g14162(new_n16509, new_n5989, new_n16511);
xor_4  g14163(new_n16496, new_n3549, new_n16512);
or_5   g14164(new_n16512, new_n5993, new_n16513);
xor_4  g14165(new_n16512, new_n5995, new_n16514);
xor_4  g14166(new_n16495, new_n3553, new_n16515);
or_5   g14167(new_n16515, new_n5999, new_n16516_1);
xor_4  g14168(new_n16515, new_n6001, new_n16517_1);
xor_4  g14169(new_n16494, new_n3558, new_n16518);
or_5   g14170(new_n16518, new_n6004, new_n16519);
xor_4  g14171(new_n16518, new_n6006, new_n16520);
nand_5 g14172(new_n16494, new_n6009, new_n16521_1);
nor_5  g14173(new_n6009, n7139, new_n16522);
xor_4  g14174(new_n16522, n16521, new_n16523);
nand_5 g14175(new_n16523, new_n6013, new_n16524_1);
and_5  g14176(new_n16524_1, new_n16521_1, new_n16525);
or_5   g14177(new_n16525, new_n16520, new_n16526);
and_5  g14178(new_n16526, new_n16519, new_n16527_1);
or_5   g14179(new_n16527_1, new_n16517_1, new_n16528);
and_5  g14180(new_n16528, new_n16516_1, new_n16529);
or_5   g14181(new_n16529, new_n16514, new_n16530);
and_5  g14182(new_n16530, new_n16513, new_n16531);
or_5   g14183(new_n16531, new_n16511, new_n16532);
and_5  g14184(new_n16532, new_n16510, new_n16533);
or_5   g14185(new_n16533, new_n16508, new_n16534);
and_5  g14186(new_n16534, new_n16507_1, new_n16535);
nand_5 g14187(new_n16535, new_n16505, new_n16536);
nand_5 g14188(new_n16536, new_n16504, new_n16537);
xor_4  g14189(new_n16537, new_n16502_1, new_n16538);
not_10 g14190(new_n16538, new_n16539);
xor_4  g14191(new_n6074, new_n4923, new_n16540);
or_5   g14192(new_n6079, new_n4927, new_n16541);
xor_4  g14193(new_n6079, new_n4927, new_n16542);
not_10 g14194(new_n16542, new_n16543);
or_5   g14195(new_n6084_1, new_n4931, new_n16544_1);
or_5   g14196(new_n8650, new_n8624, new_n16545);
and_5  g14197(new_n16545, new_n16544_1, new_n16546);
or_5   g14198(new_n16546, new_n16543, new_n16547);
and_5  g14199(new_n16547, new_n16541, new_n16548);
xor_4  g14200(new_n16548, new_n16540, new_n16549);
xor_4  g14201(new_n16549, new_n16539, new_n16550);
xor_4  g14202(new_n16546, new_n16543, new_n16551);
xor_4  g14203(new_n16535, new_n16505, new_n16552);
nor_5  g14204(new_n16552, new_n16551, new_n16553);
xor_4  g14205(new_n16552, new_n16551, new_n16554_1);
not_10 g14206(new_n16554_1, new_n16555);
not_10 g14207(new_n8651, new_n16556);
xor_4  g14208(new_n16533, new_n16508, new_n16557);
and_5  g14209(new_n16557, new_n16556, new_n16558);
xnor_4 g14210(new_n16557, new_n8651, new_n16559);
not_10 g14211(new_n16559, new_n16560);
xor_4  g14212(new_n16531, new_n16511, new_n16561);
and_5  g14213(new_n16561, new_n8684, new_n16562);
xnor_4 g14214(new_n16561, new_n8683, new_n16563);
not_10 g14215(new_n16563, new_n16564);
not_10 g14216(new_n8690, new_n16565);
xor_4  g14217(new_n16529, new_n16514, new_n16566);
and_5  g14218(new_n16566, new_n16565, new_n16567);
xnor_4 g14219(new_n16566, new_n8690, new_n16568);
not_10 g14220(new_n16568, new_n16569);
xnor_4 g14221(new_n16527_1, new_n16517_1, new_n16570);
nor_5  g14222(new_n16570, new_n8695, new_n16571);
not_10 g14223(new_n16571, new_n16572);
xor_4  g14224(new_n16570, new_n8695, new_n16573);
xor_4  g14225(new_n16525, new_n16520, new_n16574);
nor_5  g14226(new_n16574, new_n8704, new_n16575);
xnor_4 g14227(new_n16574, new_n8701, new_n16576);
xor_4  g14228(new_n16523, new_n6013, new_n16577);
nand_5 g14229(new_n16577, new_n8706, new_n16578);
xor_4  g14230(new_n6009, n7139, new_n16579);
and_5  g14231(new_n16579, new_n8711, new_n16580);
xor_4  g14232(new_n16577, new_n8706, new_n16581);
not_10 g14233(new_n16581, new_n16582);
or_5   g14234(new_n16582, new_n16580, new_n16583_1);
and_5  g14235(new_n16583_1, new_n16578, new_n16584_1);
and_5  g14236(new_n16584_1, new_n16576, new_n16585);
nor_5  g14237(new_n16585, new_n16575, new_n16586);
and_5  g14238(new_n16586, new_n16573, new_n16587);
not_10 g14239(new_n16587, new_n16588);
and_5  g14240(new_n16588, new_n16572, new_n16589_1);
nor_5  g14241(new_n16589_1, new_n16569, new_n16590);
nor_5  g14242(new_n16590, new_n16567, new_n16591);
nor_5  g14243(new_n16591, new_n16564, new_n16592);
nor_5  g14244(new_n16592, new_n16562, new_n16593);
nor_5  g14245(new_n16593, new_n16560, new_n16594);
nor_5  g14246(new_n16594, new_n16558, new_n16595);
nor_5  g14247(new_n16595, new_n16555, new_n16596_1);
nor_5  g14248(new_n16596_1, new_n16553, new_n16597);
xor_4  g14249(new_n16597, new_n16550, n3725);
nor_5  g14250(n11220, n3425, new_n16599);
not_10 g14251(new_n16599, new_n16600);
nor_5  g14252(new_n13308, new_n13305, new_n16601);
not_10 g14253(new_n16601, new_n16602);
and_5  g14254(new_n16602, new_n16600, new_n16603);
or_5   g14255(n7335, n2160, new_n16604);
or_5   g14256(new_n13302, new_n13299, new_n16605);
and_5  g14257(new_n16605, new_n16604, new_n16606);
xnor_4 g14258(new_n16606, new_n16603, new_n16607);
nor_5  g14259(new_n13310, new_n13303, new_n16608_1);
nor_5  g14260(new_n13315, new_n13312, new_n16609);
nor_5  g14261(new_n16609, new_n16608_1, new_n16610);
xor_4  g14262(new_n16610, new_n16607, new_n16611);
not_10 g14263(new_n16611, new_n16612);
xor_4  g14264(new_n16612, new_n15118_1, new_n16613);
nor_5  g14265(new_n15121, new_n13316, new_n16614);
xnor_4 g14266(new_n15121, new_n13317, new_n16615);
and_5  g14267(new_n15125, new_n5426, new_n16616);
xnor_4 g14268(new_n15125, new_n5426, new_n16617_1);
or_5   g14269(new_n15129, new_n5430_1, new_n16618);
not_10 g14270(new_n15132, new_n16619);
nand_5 g14271(new_n16619, new_n5434, new_n16620);
xnor_4 g14272(new_n15132, new_n5434, new_n16621);
not_10 g14273(new_n16621, new_n16622);
nand_5 g14274(new_n15047, new_n5439_1, new_n16623);
xor_4  g14275(new_n15047, new_n5439_1, new_n16624);
not_10 g14276(new_n16624, new_n16625);
or_5   g14277(new_n5445, new_n4246, new_n16626);
nor_5  g14278(new_n5449, new_n4252, new_n16627);
xor_4  g14279(new_n5449, new_n4251, new_n16628);
or_5   g14280(new_n5454, new_n4256_1, new_n16629);
xor_4  g14281(new_n5454, new_n4255, new_n16630_1);
or_5   g14282(new_n5457, new_n4259, new_n16631);
or_5   g14283(new_n5458, new_n4239, new_n16632);
not_10 g14284(new_n4261, new_n16633);
nor_5  g14285(new_n5463, new_n16633, new_n16634);
nand_5 g14286(new_n16634, new_n16632, new_n16635);
and_5  g14287(new_n16635, new_n16631, new_n16636);
or_5   g14288(new_n16636, new_n16630_1, new_n16637);
and_5  g14289(new_n16637, new_n16629, new_n16638);
nor_5  g14290(new_n16638, new_n16628, new_n16639);
or_5   g14291(new_n16639, new_n16627, new_n16640_1);
xor_4  g14292(new_n5445, new_n4246, new_n16641);
not_10 g14293(new_n16641, new_n16642);
or_5   g14294(new_n16642, new_n16640_1, new_n16643);
and_5  g14295(new_n16643, new_n16626, new_n16644);
or_5   g14296(new_n16644, new_n16625, new_n16645);
and_5  g14297(new_n16645, new_n16623, new_n16646);
or_5   g14298(new_n16646, new_n16622, new_n16647);
and_5  g14299(new_n16647, new_n16620, new_n16648);
xor_4  g14300(new_n15129, new_n5430_1, new_n16649);
nand_5 g14301(new_n16649, new_n16648, new_n16650);
and_5  g14302(new_n16650, new_n16618, new_n16651);
nor_5  g14303(new_n16651, new_n16617_1, new_n16652);
nor_5  g14304(new_n16652, new_n16616, new_n16653);
and_5  g14305(new_n16653, new_n16615, new_n16654);
nor_5  g14306(new_n16654, new_n16614, new_n16655);
not_10 g14307(new_n16655, new_n16656_1);
xnor_4 g14308(new_n16656_1, new_n16613, n3733);
xnor_4 g14309(new_n10975, n24937, new_n16658);
nand_5 g14310(new_n10979, n5098, new_n16659);
xnor_4 g14311(new_n10979, n5098, new_n16660);
not_10 g14312(n3030, new_n16661);
or_5   g14313(new_n10929, new_n16661, new_n16662);
or_5   g14314(new_n15692, new_n15680, new_n16663);
and_5  g14315(new_n16663, new_n16662, new_n16664);
or_5   g14316(new_n16664, new_n16660, new_n16665);
and_5  g14317(new_n16665, new_n16659, new_n16666);
xor_4  g14318(new_n16666, new_n16658, new_n16667);
xnor_4 g14319(new_n16667, new_n10199, new_n16668);
xor_4  g14320(new_n16664, new_n16660, new_n16669);
or_5   g14321(new_n16669, new_n10205, new_n16670);
xnor_4 g14322(new_n16669, new_n10205, new_n16671);
or_5   g14323(new_n15693, new_n10211, new_n16672);
nand_5 g14324(new_n15710, new_n15694, new_n16673);
and_5  g14325(new_n16673, new_n16672, new_n16674_1);
or_5   g14326(new_n16674_1, new_n16671, new_n16675);
and_5  g14327(new_n16675, new_n16670, new_n16676);
xor_4  g14328(new_n16676, new_n16668, n3755);
xor_4  g14329(new_n9270, new_n9229, n3758);
not_10 g14330(n2570, new_n16679);
not_10 g14331(n19033, new_n16680);
not_10 g14332(n655, new_n16681);
and_5  g14333(new_n16033, new_n16024, new_n16682_1);
and_5  g14334(new_n16682_1, new_n16681, new_n16683);
and_5  g14335(new_n16683, new_n16680, new_n16684_1);
xor_4  g14336(new_n16684_1, new_n16679, new_n16685);
xor_4  g14337(new_n16685, n14692, new_n16686);
xor_4  g14338(new_n16683, new_n16680, new_n16687);
or_5   g14339(new_n16687, new_n10470, new_n16688_1);
xor_4  g14340(new_n16687, n4100, new_n16689);
xor_4  g14341(new_n16682_1, new_n16681, new_n16690);
or_5   g14342(new_n16690, new_n10473, new_n16691);
xor_4  g14343(new_n16690, n21957, new_n16692);
or_5   g14344(new_n16034, new_n10476, new_n16693);
or_5   g14345(new_n16063, new_n16035, new_n16694);
and_5  g14346(new_n16694, new_n16693, new_n16695);
or_5   g14347(new_n16695, new_n16692, new_n16696);
and_5  g14348(new_n16696, new_n16691, new_n16697);
or_5   g14349(new_n16697, new_n16689, new_n16698);
and_5  g14350(new_n16698, new_n16688_1, new_n16699);
xor_4  g14351(new_n16699, new_n16686, new_n16700);
and_5  g14352(new_n16700, new_n12195, new_n16701);
xor_4  g14353(new_n16700, new_n12194, new_n16702);
xor_4  g14354(new_n16697, new_n16689, new_n16703);
nand_5 g14355(new_n16703, new_n6876, new_n16704);
xnor_4 g14356(new_n16703, new_n6876, new_n16705);
xor_4  g14357(new_n16695, new_n16692, new_n16706);
nand_5 g14358(new_n16706, new_n6879, new_n16707);
xnor_4 g14359(new_n16706, new_n6879, new_n16708);
nand_5 g14360(new_n16064, new_n6884, new_n16709);
or_5   g14361(new_n16092, new_n16065, new_n16710);
and_5  g14362(new_n16710, new_n16709, new_n16711);
or_5   g14363(new_n16711, new_n16708, new_n16712);
and_5  g14364(new_n16712, new_n16707, new_n16713);
or_5   g14365(new_n16713, new_n16705, new_n16714);
and_5  g14366(new_n16714, new_n16704, new_n16715);
nor_5  g14367(new_n16715, new_n16702, new_n16716);
nor_5  g14368(new_n16716, new_n16701, new_n16717);
and_5  g14369(new_n16684_1, new_n16679, new_n16718);
not_10 g14370(n14692, new_n16719);
nor_5  g14371(new_n16685, new_n16719, new_n16720);
nor_5  g14372(new_n16699, new_n16686, new_n16721);
nor_5  g14373(new_n16721, new_n16720, new_n16722_1);
xnor_4 g14374(new_n16722_1, new_n16718, new_n16723);
xor_4  g14375(new_n16723, new_n12241, new_n16724);
xor_4  g14376(new_n16724, new_n16717, new_n16725);
nor_5  g14377(new_n16725, new_n10584, new_n16726);
xor_4  g14378(new_n16725, new_n10584, new_n16727);
xor_4  g14379(new_n16715, new_n16702, new_n16728);
and_5  g14380(new_n16728, new_n10588_1, new_n16729);
xor_4  g14381(new_n16728, new_n10588_1, new_n16730);
xor_4  g14382(new_n16713, new_n16705, new_n16731);
and_5  g14383(new_n16731, new_n10592, new_n16732);
xor_4  g14384(new_n16731, new_n10592, new_n16733_1);
not_10 g14385(new_n16733_1, new_n16734);
xor_4  g14386(new_n16711, new_n16708, new_n16735);
nand_5 g14387(new_n16735, new_n10597, new_n16736);
xor_4  g14388(new_n16735, new_n10597, new_n16737);
or_5   g14389(new_n16093, new_n10603, new_n16738);
nand_5 g14390(new_n16126, new_n16094, new_n16739);
and_5  g14391(new_n16739, new_n16738, new_n16740);
nand_5 g14392(new_n16740, new_n16737, new_n16741);
and_5  g14393(new_n16741, new_n16736, new_n16742);
nor_5  g14394(new_n16742, new_n16734, new_n16743_1);
nor_5  g14395(new_n16743_1, new_n16732, new_n16744);
not_10 g14396(new_n16744, new_n16745);
and_5  g14397(new_n16745, new_n16730, new_n16746);
nor_5  g14398(new_n16746, new_n16729, new_n16747);
not_10 g14399(new_n16747, new_n16748);
and_5  g14400(new_n16748, new_n16727, new_n16749);
nor_5  g14401(new_n16749, new_n16726, new_n16750);
not_10 g14402(new_n16750, new_n16751);
or_5   g14403(new_n16723, new_n12241, new_n16752);
nand_5 g14404(new_n16722_1, new_n16718, new_n16753);
nand_5 g14405(new_n16723, new_n12241, new_n16754);
nand_5 g14406(new_n16754, new_n16717, new_n16755);
and_5  g14407(new_n16755, new_n16753, new_n16756);
and_5  g14408(new_n16756, new_n16752, new_n16757);
xnor_4 g14409(new_n16757, new_n16751, n3760);
xnor_4 g14410(new_n3930, new_n3906, n3781);
xor_4  g14411(new_n13821, new_n13795, n3794);
and_5  g14412(new_n11073, new_n5024_1, new_n16761);
not_10 g14413(new_n16761, new_n16762);
nand_5 g14414(new_n16762, new_n5029, new_n16763);
and_5  g14415(new_n16761, new_n4796, new_n16764);
not_10 g14416(new_n16764, new_n16765);
nand_5 g14417(new_n16765, new_n16763, new_n16766);
nand_5 g14418(new_n11072, new_n6009, new_n16767);
and_5  g14419(new_n6009, new_n5948, new_n16768);
nor_5  g14420(new_n6013, new_n6009, new_n16769);
nor_5  g14421(new_n16769, new_n16768, new_n16770);
xor_4  g14422(new_n16770, new_n13354, new_n16771);
xor_4  g14423(new_n16771, new_n16767, new_n16772);
xor_4  g14424(new_n16772, new_n16766, n3842);
xnor_4 g14425(new_n12518, new_n9070, n3850);
xnor_4 g14426(new_n15073, new_n4288, n3869);
xnor_4 g14427(n21749, n919, new_n16776);
or_5   g14428(n25316, n7769, new_n16777);
and_5  g14429(n21138, n20385, new_n16778);
xnor_4 g14430(n25316, n7769, new_n16779);
or_5   g14431(new_n16779, new_n16778, new_n16780);
and_5  g14432(new_n16780, new_n16777, new_n16781);
xor_4  g14433(new_n16781, new_n16776, new_n16782);
xor_4  g14434(new_n16782, n19584, new_n16783);
not_10 g14435(n15332, new_n16784);
xor_4  g14436(n21138, n20385, new_n16785);
nor_5  g14437(new_n16785, new_n16784, new_n16786);
or_5   g14438(new_n16786, n5060, new_n16787);
xnor_4 g14439(new_n16779, new_n16778, new_n16788);
xor_4  g14440(new_n16786, n5060, new_n16789);
nand_5 g14441(new_n16789, new_n16788, new_n16790);
and_5  g14442(new_n16790, new_n16787, new_n16791);
xor_4  g14443(new_n16791, new_n16783, new_n16792);
xor_4  g14444(new_n16792, new_n15970, new_n16793);
xor_4  g14445(new_n16789, new_n16788, new_n16794);
or_5   g14446(new_n16794, new_n15961, new_n16795);
xor_4  g14447(new_n16785, new_n16784, new_n16796);
or_5   g14448(new_n16796, new_n15964, new_n16797);
xor_4  g14449(new_n16794, new_n15961, new_n16798_1);
nand_5 g14450(new_n16798_1, new_n16797, new_n16799);
nand_5 g14451(new_n16799, new_n16795, new_n16800);
xnor_4 g14452(new_n16800, new_n16793, n3871);
xor_4  g14453(new_n16584_1, new_n16576, n3891);
not_10 g14454(new_n6384, new_n16803);
xor_4  g14455(n10250, n2570, new_n16804);
or_5   g14456(n19033, new_n12199, new_n16805);
xor_4  g14457(n19033, n7674, new_n16806);
or_5   g14458(new_n12202, n655, new_n16807);
xor_4  g14459(n6397, n655, new_n16808);
or_5   g14460(new_n12205, n18145, new_n16809);
xor_4  g14461(n19196, n18145, new_n16810);
not_10 g14462(n23586, new_n16811);
or_5   g14463(new_n16811, n10712, new_n16812_1);
xor_4  g14464(n23586, n10712, new_n16813);
not_10 g14465(n21226, new_n16814);
or_5   g14466(n25126, new_n16814, new_n16815);
xor_4  g14467(n25126, n21226, new_n16816);
or_5   g14468(n19608, new_n12210, new_n16817);
or_5   g14469(n20036, new_n16028, new_n16818_1);
or_5   g14470(new_n4128, new_n4121, new_n16819);
and_5  g14471(new_n16819, new_n16818_1, new_n16820);
xnor_4 g14472(n19608, n4426, new_n16821);
nand_5 g14473(new_n16821, new_n16820, new_n16822);
and_5  g14474(new_n16822, new_n16817, new_n16823);
or_5   g14475(new_n16823, new_n16816, new_n16824_1);
and_5  g14476(new_n16824_1, new_n16815, new_n16825);
or_5   g14477(new_n16825, new_n16813, new_n16826);
and_5  g14478(new_n16826, new_n16812_1, new_n16827);
or_5   g14479(new_n16827, new_n16810, new_n16828);
and_5  g14480(new_n16828, new_n16809, new_n16829);
or_5   g14481(new_n16829, new_n16808, new_n16830);
and_5  g14482(new_n16830, new_n16807, new_n16831);
or_5   g14483(new_n16831, new_n16806, new_n16832);
and_5  g14484(new_n16832, new_n16805, new_n16833);
xor_4  g14485(new_n16833, new_n16804, new_n16834_1);
xnor_4 g14486(new_n16834_1, new_n12194, new_n16835);
xor_4  g14487(new_n16831, new_n16806, new_n16836);
or_5   g14488(new_n16836, new_n6877, new_n16837_1);
xor_4  g14489(new_n16836, new_n6876, new_n16838);
xor_4  g14490(new_n16829, new_n16808, new_n16839);
or_5   g14491(new_n16839, new_n6880, new_n16840);
xor_4  g14492(new_n16839, new_n6879, new_n16841_1);
xor_4  g14493(new_n16827, new_n16810, new_n16842);
or_5   g14494(new_n16842, new_n6885, new_n16843);
xor_4  g14495(new_n16842, new_n6884, new_n16844);
xor_4  g14496(new_n16825, new_n16813, new_n16845);
or_5   g14497(new_n16845, new_n6890, new_n16846);
xor_4  g14498(new_n16845, new_n6889, new_n16847);
xor_4  g14499(new_n16823, new_n16816, new_n16848);
or_5   g14500(new_n16848, new_n6895, new_n16849);
xor_4  g14501(new_n16848, new_n6894, new_n16850);
xor_4  g14502(new_n16821, new_n16820, new_n16851);
or_5   g14503(new_n16851, new_n6899, new_n16852);
xnor_4 g14504(new_n16851, new_n6899, new_n16853);
nand_5 g14505(new_n4129, new_n4120, new_n16854);
nand_5 g14506(new_n4141, new_n4130, new_n16855);
and_5  g14507(new_n16855, new_n16854, new_n16856);
or_5   g14508(new_n16856, new_n16853, new_n16857);
and_5  g14509(new_n16857, new_n16852, new_n16858);
or_5   g14510(new_n16858, new_n16850, new_n16859);
and_5  g14511(new_n16859, new_n16849, new_n16860);
or_5   g14512(new_n16860, new_n16847, new_n16861);
and_5  g14513(new_n16861, new_n16846, new_n16862);
or_5   g14514(new_n16862, new_n16844, new_n16863);
and_5  g14515(new_n16863, new_n16843, new_n16864);
or_5   g14516(new_n16864, new_n16841_1, new_n16865);
and_5  g14517(new_n16865, new_n16840, new_n16866);
or_5   g14518(new_n16866, new_n16838, new_n16867);
and_5  g14519(new_n16867, new_n16837_1, new_n16868);
xor_4  g14520(new_n16868, new_n16835, new_n16869);
xor_4  g14521(new_n16869, new_n16803, new_n16870);
not_10 g14522(new_n16870, new_n16871);
not_10 g14523(new_n6391, new_n16872);
xor_4  g14524(new_n16866, new_n16838, new_n16873);
and_5  g14525(new_n16873, new_n16872, new_n16874);
xnor_4 g14526(new_n16873, new_n6391, new_n16875);
not_10 g14527(new_n16875, new_n16876);
not_10 g14528(new_n6396, new_n16877);
xor_4  g14529(new_n16864, new_n16841_1, new_n16878);
and_5  g14530(new_n16878, new_n16877, new_n16879);
xnor_4 g14531(new_n16878, new_n6396, new_n16880);
not_10 g14532(new_n16880, new_n16881);
not_10 g14533(new_n6399, new_n16882);
xor_4  g14534(new_n16862, new_n16844, new_n16883);
and_5  g14535(new_n16883, new_n16882, new_n16884);
xor_4  g14536(new_n16883, new_n16882, new_n16885_1);
not_10 g14537(new_n16885_1, new_n16886);
xor_4  g14538(new_n16860, new_n16847, new_n16887);
and_5  g14539(new_n16887, new_n6406, new_n16888);
xnor_4 g14540(new_n16887, new_n6405, new_n16889);
not_10 g14541(new_n16889, new_n16890);
not_10 g14542(new_n6412, new_n16891);
xor_4  g14543(new_n16858, new_n16850, new_n16892);
and_5  g14544(new_n16892, new_n16891, new_n16893);
xnor_4 g14545(new_n16892, new_n6412, new_n16894);
not_10 g14546(new_n16894, new_n16895);
xor_4  g14547(new_n16856, new_n16853, new_n16896);
and_5  g14548(new_n16896, new_n6417, new_n16897);
xor_4  g14549(new_n16896, new_n6417, new_n16898);
not_10 g14550(new_n16898, new_n16899);
nor_5  g14551(new_n4150_1, new_n4143, new_n16900);
not_10 g14552(new_n16900, new_n16901);
not_10 g14553(new_n4163, new_n16902);
and_5  g14554(new_n16902, new_n4151_1, new_n16903);
not_10 g14555(new_n16903, new_n16904);
and_5  g14556(new_n16904, new_n16901, new_n16905_1);
nor_5  g14557(new_n16905_1, new_n16899, new_n16906);
nor_5  g14558(new_n16906, new_n16897, new_n16907);
nor_5  g14559(new_n16907, new_n16895, new_n16908);
nor_5  g14560(new_n16908, new_n16893, new_n16909);
nor_5  g14561(new_n16909, new_n16890, new_n16910);
nor_5  g14562(new_n16910, new_n16888, new_n16911_1);
nor_5  g14563(new_n16911_1, new_n16886, new_n16912);
nor_5  g14564(new_n16912, new_n16884, new_n16913);
nor_5  g14565(new_n16913, new_n16881, new_n16914);
nor_5  g14566(new_n16914, new_n16879, new_n16915);
nor_5  g14567(new_n16915, new_n16876, new_n16916);
nor_5  g14568(new_n16916, new_n16874, new_n16917);
xnor_4 g14569(new_n16917, new_n16871, n3932);
xnor_4 g14570(new_n3924, new_n3922, n3934);
xnor_4 g14571(new_n4100_1, new_n4098, n3971);
nor_5  g14572(n8581, n5026, new_n16921);
and_5  g14573(new_n16921, new_n7268_1, new_n16922);
and_5  g14574(new_n16922, new_n11190, new_n16923);
and_5  g14575(new_n16923, new_n11187, new_n16924);
and_5  g14576(new_n16924, new_n11183, new_n16925);
and_5  g14577(new_n16925, new_n11179, new_n16926);
and_5  g14578(new_n16926, new_n11175, new_n16927);
xor_4  g14579(new_n16927, new_n11171, new_n16928);
xor_4  g14580(new_n16928, new_n8954, new_n16929);
xor_4  g14581(new_n16926, new_n11175, new_n16930);
or_5   g14582(new_n16930, n3710, new_n16931);
xor_4  g14583(new_n16930, n3710, new_n16932);
xor_4  g14584(new_n16925, new_n11179, new_n16933);
nand_5 g14585(new_n16933, n26318, new_n16934);
or_5   g14586(new_n16933, n26318, new_n16935);
xor_4  g14587(new_n16924, new_n11183, new_n16936);
nor_5  g14588(new_n16936, n26054, new_n16937);
xor_4  g14589(new_n16936, new_n8917, new_n16938);
xor_4  g14590(new_n16923, new_n11187, new_n16939);
or_5   g14591(new_n16939, n19081, new_n16940);
xor_4  g14592(new_n16939, new_n8921, new_n16941);
xor_4  g14593(new_n16922, new_n11190, new_n16942);
or_5   g14594(new_n16942, n8309, new_n16943);
xor_4  g14595(new_n16921, new_n7268_1, new_n16944);
nor_5  g14596(new_n16944, n19144, new_n16945);
xor_4  g14597(new_n16944, new_n10286, new_n16946);
xor_4  g14598(n8581, n5026, new_n16947);
or_5   g14599(new_n16947, n12593, new_n16948);
nand_5 g14600(n13714, n8581, new_n16949);
xor_4  g14601(new_n16947, n12593, new_n16950);
nand_5 g14602(new_n16950, new_n16949, new_n16951_1);
and_5  g14603(new_n16951_1, new_n16948, new_n16952);
nor_5  g14604(new_n16952, new_n16946, new_n16953);
or_5   g14605(new_n16953, new_n16945, new_n16954_1);
xor_4  g14606(new_n16942, n8309, new_n16955);
nand_5 g14607(new_n16955, new_n16954_1, new_n16956);
and_5  g14608(new_n16956, new_n16943, new_n16957);
or_5   g14609(new_n16957, new_n16941, new_n16958);
and_5  g14610(new_n16958, new_n16940, new_n16959);
nor_5  g14611(new_n16959, new_n16938, new_n16960);
nor_5  g14612(new_n16960, new_n16937, new_n16961);
nand_5 g14613(new_n16961, new_n16935, new_n16962);
and_5  g14614(new_n16962, new_n16934, new_n16963);
nand_5 g14615(new_n16963, new_n16932, new_n16964);
and_5  g14616(new_n16964, new_n16931, new_n16965);
xor_4  g14617(new_n16965, new_n16929, new_n16966);
xor_4  g14618(new_n16966, new_n5592, new_n16967);
xor_4  g14619(new_n16963, new_n16932, new_n16968_1);
or_5   g14620(new_n16968_1, new_n5593_1, new_n16969);
xor_4  g14621(new_n16968_1, n23913, new_n16970);
xor_4  g14622(new_n16933, n26318, new_n16971_1);
xor_4  g14623(new_n16971_1, new_n16961, new_n16972);
not_10 g14624(new_n16972, new_n16973);
or_5   g14625(new_n16973, new_n5594, new_n16974);
xor_4  g14626(new_n16973, n22554, new_n16975);
xor_4  g14627(new_n16959, new_n16938, new_n16976);
or_5   g14628(new_n16976, new_n5595, new_n16977);
xor_4  g14629(new_n16976, n20429, new_n16978);
xor_4  g14630(new_n16957, new_n16941, new_n16979);
or_5   g14631(new_n16979, new_n5596, new_n16980);
xor_4  g14632(new_n16979, n3909, new_n16981);
xor_4  g14633(new_n16955, new_n16954_1, new_n16982);
or_5   g14634(new_n16982, new_n5597, new_n16983);
xor_4  g14635(new_n16982, n23974, new_n16984);
xor_4  g14636(new_n16952, new_n16946, new_n16985);
or_5   g14637(new_n16985, new_n5598, new_n16986);
xor_4  g14638(new_n16985, n2146, new_n16987);
xor_4  g14639(new_n16950, new_n16949, new_n16988_1);
or_5   g14640(new_n16988_1, new_n8181, new_n16989_1);
xor_4  g14641(n13714, n8581, new_n16990);
and_5  g14642(new_n16990, n583, new_n16991);
xor_4  g14643(new_n16988_1, new_n8181, new_n16992);
nand_5 g14644(new_n16992, new_n16991, new_n16993);
and_5  g14645(new_n16993, new_n16989_1, new_n16994_1);
or_5   g14646(new_n16994_1, new_n16987, new_n16995);
and_5  g14647(new_n16995, new_n16986, new_n16996);
or_5   g14648(new_n16996, new_n16984, new_n16997);
and_5  g14649(new_n16997, new_n16983, new_n16998);
or_5   g14650(new_n16998, new_n16981, new_n16999);
and_5  g14651(new_n16999, new_n16980, new_n17000);
or_5   g14652(new_n17000, new_n16978, new_n17001);
and_5  g14653(new_n17001, new_n16977, new_n17002);
or_5   g14654(new_n17002, new_n16975, new_n17003);
and_5  g14655(new_n17003, new_n16974, new_n17004);
or_5   g14656(new_n17004, new_n16970, new_n17005);
and_5  g14657(new_n17005, new_n16969, new_n17006_1);
xor_4  g14658(new_n17006_1, new_n16967, new_n17007);
xnor_4 g14659(new_n17007, new_n8282, new_n17008);
not_10 g14660(new_n17008, new_n17009);
xor_4  g14661(new_n17004, new_n16970, new_n17010);
or_5   g14662(new_n17010, new_n8287, new_n17011);
xor_4  g14663(new_n17010, new_n8287, new_n17012);
not_10 g14664(new_n17012, new_n17013);
xor_4  g14665(new_n17002, new_n16975, new_n17014);
or_5   g14666(new_n17014, new_n8292, new_n17015);
xor_4  g14667(new_n17014, new_n8292, new_n17016);
not_10 g14668(new_n17016, new_n17017);
xor_4  g14669(new_n17000, new_n16978, new_n17018);
or_5   g14670(new_n17018, new_n8297, new_n17019);
xor_4  g14671(new_n17018, new_n8297, new_n17020);
not_10 g14672(new_n17020, new_n17021);
xor_4  g14673(new_n16998, new_n16981, new_n17022);
or_5   g14674(new_n17022, new_n8303, new_n17023);
xor_4  g14675(new_n17022, new_n8303, new_n17024);
not_10 g14676(new_n17024, new_n17025);
xor_4  g14677(new_n16996, new_n16984, new_n17026);
or_5   g14678(new_n17026, new_n8308, new_n17027);
xor_4  g14679(new_n17026, new_n8308, new_n17028);
not_10 g14680(new_n17028, new_n17029);
xor_4  g14681(new_n16994_1, new_n16987, new_n17030);
or_5   g14682(new_n17030, new_n8310, new_n17031);
xor_4  g14683(new_n16992, new_n16991, new_n17032);
or_5   g14684(new_n17032, new_n8318, new_n17033);
xor_4  g14685(new_n16990, n583, new_n17034);
and_5  g14686(new_n17034, new_n2547_1, new_n17035_1);
xnor_4 g14687(new_n17032, new_n8317, new_n17036);
not_10 g14688(new_n17036, new_n17037_1);
or_5   g14689(new_n17037_1, new_n17035_1, new_n17038);
and_5  g14690(new_n17038, new_n17033, new_n17039);
xor_4  g14691(new_n17030, new_n8310, new_n17040);
not_10 g14692(new_n17040, new_n17041);
or_5   g14693(new_n17041, new_n17039, new_n17042);
and_5  g14694(new_n17042, new_n17031, new_n17043);
or_5   g14695(new_n17043, new_n17029, new_n17044);
and_5  g14696(new_n17044, new_n17027, new_n17045);
or_5   g14697(new_n17045, new_n17025, new_n17046);
and_5  g14698(new_n17046, new_n17023, new_n17047);
or_5   g14699(new_n17047, new_n17021, new_n17048);
and_5  g14700(new_n17048, new_n17019, new_n17049);
or_5   g14701(new_n17049, new_n17017, new_n17050);
and_5  g14702(new_n17050, new_n17015, new_n17051);
or_5   g14703(new_n17051, new_n17013, new_n17052);
and_5  g14704(new_n17052, new_n17011, new_n17053);
xnor_4 g14705(new_n17053, new_n17009, n3983);
xor_4  g14706(n13714, n583, new_n17055);
xor_4  g14707(new_n17055, n6611, new_n17056);
not_10 g14708(new_n17056, new_n17057);
and_5  g14709(new_n17057, new_n6702, new_n17058);
nand_5 g14710(new_n17055, n6611, new_n17059);
nand_5 g14711(n13714, n583, new_n17060);
xor_4  g14712(n22173, n12593, new_n17061);
xor_4  g14713(new_n17061, new_n17060, new_n17062);
xor_4  g14714(new_n17062, new_n9175, new_n17063);
xor_4  g14715(new_n17063, new_n17059, new_n17064);
xor_4  g14716(new_n17064, new_n17058, new_n17065);
xor_4  g14717(new_n17065, new_n6698, n4000);
xor_4  g14718(n26823, n20179, new_n17067);
or_5   g14719(n19228, new_n3188, new_n17068_1);
xor_4  g14720(n19228, n4812, new_n17069_1);
or_5   g14721(new_n3189, n15539, new_n17070_1);
xor_4  g14722(n24278, n15539, new_n17071);
or_5   g14723(new_n3190, n8052, new_n17072);
or_5   g14724(n24618, new_n7532, new_n17073);
and_5  g14725(n10158, new_n3241, new_n17074);
and_5  g14726(new_n11459, new_n11458, new_n17075_1);
nor_5  g14727(new_n17075_1, new_n17074, new_n17076);
nand_5 g14728(new_n17076, new_n17073, new_n17077_1);
and_5  g14729(new_n17077_1, new_n17072, new_n17078);
or_5   g14730(new_n17078, new_n17071, new_n17079);
and_5  g14731(new_n17079, new_n17070_1, new_n17080);
or_5   g14732(new_n17080, new_n17069_1, new_n17081);
and_5  g14733(new_n17081, new_n17068_1, new_n17082);
xor_4  g14734(new_n17082, new_n17067, new_n17083);
xor_4  g14735(new_n17083, new_n7444, new_n17084_1);
xor_4  g14736(new_n17080, new_n17069_1, new_n17085);
nor_5  g14737(new_n17085, new_n7450, new_n17086);
not_10 g14738(new_n17086, new_n17087);
xor_4  g14739(new_n17085, new_n7450, new_n17088);
xor_4  g14740(new_n17078, new_n17071, new_n17089);
nor_5  g14741(new_n17089, new_n7455, new_n17090_1);
not_10 g14742(new_n17090_1, new_n17091);
xnor_4 g14743(n24618, n8052, new_n17092);
xor_4  g14744(new_n17092, new_n17076, new_n17093);
nor_5  g14745(new_n17093, new_n7463, new_n17094);
xor_4  g14746(new_n17093, new_n7463, new_n17095_1);
nor_5  g14747(new_n11460, new_n11457, new_n17096);
and_5  g14748(new_n11461, new_n7472, new_n17097);
nor_5  g14749(new_n17097, new_n17096, new_n17098);
and_5  g14750(new_n17098, new_n17095_1, new_n17099);
nor_5  g14751(new_n17099, new_n17094, new_n17100);
not_10 g14752(new_n17100, new_n17101);
xor_4  g14753(new_n17089, new_n7455, new_n17102);
and_5  g14754(new_n17102, new_n17101, new_n17103);
not_10 g14755(new_n17103, new_n17104_1);
and_5  g14756(new_n17104_1, new_n17091, new_n17105);
not_10 g14757(new_n17105, new_n17106_1);
and_5  g14758(new_n17106_1, new_n17088, new_n17107);
not_10 g14759(new_n17107, new_n17108);
and_5  g14760(new_n17108, new_n17087, new_n17109);
xor_4  g14761(new_n17109, new_n17084_1, n4010);
xor_4  g14762(n11220, n2160, new_n17111);
not_10 g14763(n10763, new_n17112);
or_5   g14764(n22379, new_n17112, new_n17113);
xor_4  g14765(n22379, n10763, new_n17114);
not_10 g14766(n7437, new_n17115);
or_5   g14767(new_n17115, n1662, new_n17116);
xor_4  g14768(n7437, n1662, new_n17117);
or_5   g14769(new_n12052, n12875, new_n17118);
and_5  g14770(n7099, new_n2845, new_n17119_1);
nor_5  g14771(new_n15039, new_n15019_1, new_n17120);
or_5   g14772(new_n17120, new_n17119_1, new_n17121);
xnor_4 g14773(n20700, n12875, new_n17122);
nand_5 g14774(new_n17122, new_n17121, new_n17123);
and_5  g14775(new_n17123, new_n17118, new_n17124);
or_5   g14776(new_n17124, new_n17117, new_n17125);
and_5  g14777(new_n17125, new_n17116, new_n17126);
or_5   g14778(new_n17126, new_n17114, new_n17127);
and_5  g14779(new_n17127, new_n17113, new_n17128);
xor_4  g14780(new_n17128, new_n17111, new_n17129);
xnor_4 g14781(new_n17129, new_n15189, new_n17130_1);
not_10 g14782(new_n15195, new_n17131);
xor_4  g14783(new_n17126, new_n17114, new_n17132);
or_5   g14784(new_n17132, new_n17131, new_n17133);
xor_4  g14785(new_n17132, new_n17131, new_n17134);
not_10 g14786(new_n15200, new_n17135);
xor_4  g14787(new_n17124, new_n17117, new_n17136);
or_5   g14788(new_n17136, new_n17135, new_n17137);
xor_4  g14789(new_n17122, new_n17121, new_n17138_1);
and_5  g14790(new_n17138_1, new_n15204, new_n17139);
xor_4  g14791(new_n17138_1, new_n15205_1, new_n17140);
nand_5 g14792(new_n15053_1, new_n15040, new_n17141);
nand_5 g14793(new_n15085, new_n15055, new_n17142);
and_5  g14794(new_n17142, new_n17141, new_n17143);
nor_5  g14795(new_n17143, new_n17140, new_n17144);
nor_5  g14796(new_n17144, new_n17139, new_n17145);
xor_4  g14797(new_n17136, new_n17135, new_n17146);
nand_5 g14798(new_n17146, new_n17145, new_n17147);
nand_5 g14799(new_n17147, new_n17137, new_n17148);
nand_5 g14800(new_n17148, new_n17134, new_n17149);
and_5  g14801(new_n17149, new_n17133, new_n17150);
xor_4  g14802(new_n17150, new_n17130_1, n4014);
xor_4  g14803(new_n14455, new_n12917_1, new_n17152);
or_5   g14804(new_n14459, n26224, new_n17153);
xor_4  g14805(new_n14459, new_n12918, new_n17154);
or_5   g14806(new_n3735, n19327, new_n17155);
or_5   g14807(new_n3766, new_n3736, new_n17156);
and_5  g14808(new_n17156, new_n17155, new_n17157);
or_5   g14809(new_n17157, new_n17154, new_n17158);
and_5  g14810(new_n17158, new_n17153, new_n17159);
xor_4  g14811(new_n17159, new_n17152, new_n17160);
xor_4  g14812(new_n17160, n647, new_n17161);
xor_4  g14813(new_n17157, new_n17154, new_n17162);
or_5   g14814(new_n17162, new_n5912, new_n17163_1);
xor_4  g14815(new_n17162, n20409, new_n17164);
or_5   g14816(new_n3767, new_n5913, new_n17165);
or_5   g14817(new_n3802, new_n3768, new_n17166);
and_5  g14818(new_n17166, new_n17165, new_n17167);
or_5   g14819(new_n17167, new_n17164, new_n17168_1);
and_5  g14820(new_n17168_1, new_n17163_1, new_n17169);
xor_4  g14821(new_n17169, new_n17161, new_n17170);
xnor_4 g14822(new_n17170, new_n12120, new_n17171);
xor_4  g14823(new_n17167, new_n17164, new_n17172);
or_5   g14824(new_n17172, new_n12128, new_n17173);
xnor_4 g14825(new_n17172, new_n12127, new_n17174);
not_10 g14826(new_n17174, new_n17175);
or_5   g14827(new_n12135, new_n3803, new_n17176);
not_10 g14828(new_n3896, new_n17177);
or_5   g14829(new_n3934_1, new_n17177, new_n17178);
and_5  g14830(new_n17178, new_n17176, new_n17179);
or_5   g14831(new_n17179, new_n17175, new_n17180);
and_5  g14832(new_n17180, new_n17173, new_n17181);
xor_4  g14833(new_n17181, new_n17171, n4071);
xnor_4 g14834(new_n13206, new_n13198_1, n4088);
nand_5 g14835(new_n13319_1, new_n13318, new_n17184);
nor_5  g14836(new_n13320, n5025, new_n17185);
and_5  g14837(new_n13320, n5025, new_n17186);
nor_5  g14838(new_n13325, new_n17186, new_n17187);
or_5   g14839(new_n17187, new_n17185, new_n17188);
and_5  g14840(new_n17188, new_n17184, new_n17189);
not_10 g14841(new_n16603, new_n17190);
nor_5  g14842(new_n16606, new_n17190, new_n17191);
and_5  g14843(new_n16606, new_n17190, new_n17192);
not_10 g14844(new_n16610, new_n17193);
nor_5  g14845(new_n17193, new_n17192, new_n17194);
nor_5  g14846(new_n17194, new_n17191, new_n17195);
and_5  g14847(new_n17195, new_n17189, new_n17196);
nor_5  g14848(new_n17189, new_n16612, new_n17197);
and_5  g14849(new_n17189, new_n16612, new_n17198);
nor_5  g14850(new_n13326, new_n13317, new_n17199);
nor_5  g14851(new_n13330, new_n13327, new_n17200);
nor_5  g14852(new_n17200, new_n17199, new_n17201);
not_10 g14853(new_n17201, new_n17202_1);
nor_5  g14854(new_n17202_1, new_n17198, new_n17203);
nor_5  g14855(new_n17203, new_n17197, new_n17204);
or_5   g14856(new_n17204, new_n17196, new_n17205);
nor_5  g14857(new_n17195, new_n17189, new_n17206);
or_5   g14858(new_n17206, new_n17203, new_n17207);
and_5  g14859(new_n17207, new_n17205, n4089);
and_5  g14860(new_n12357, new_n7519, new_n17209);
xor_4  g14861(new_n17209, new_n7515, new_n17210);
xor_4  g14862(new_n17210, n3228, new_n17211);
nor_5  g14863(new_n12358, n5302, new_n17212);
xor_4  g14864(new_n12358, n5302, new_n17213);
nand_5 g14865(new_n12360, n25738, new_n17214);
or_5   g14866(new_n12360, n25738, new_n17215);
nor_5  g14867(new_n8733, n21471, new_n17216);
and_5  g14868(new_n8751, new_n8734, new_n17217);
nor_5  g14869(new_n17217, new_n17216, new_n17218);
nand_5 g14870(new_n17218, new_n17215, new_n17219_1);
and_5  g14871(new_n17219_1, new_n17214, new_n17220);
and_5  g14872(new_n17220, new_n17213, new_n17221);
nor_5  g14873(new_n17221, new_n17212, new_n17222);
xnor_4 g14874(new_n17222, new_n17211, new_n17223);
not_10 g14875(new_n17223, new_n17224);
xor_4  g14876(new_n17224, n13775, new_n17225);
not_10 g14877(new_n17225, new_n17226);
xor_4  g14878(new_n17220, new_n17213, new_n17227);
nand_5 g14879(new_n17227, new_n8806_1, new_n17228);
xor_4  g14880(new_n17227, new_n8806_1, new_n17229);
xor_4  g14881(new_n12360, n25738, new_n17230);
xor_4  g14882(new_n17230, new_n17218, new_n17231);
nand_5 g14883(new_n17231, n19042, new_n17232_1);
and_5  g14884(new_n8753, n19472, new_n17233);
and_5  g14885(new_n8774, new_n8754, new_n17234);
or_5   g14886(new_n17234, new_n17233, new_n17235);
xor_4  g14887(new_n17231, n19042, new_n17236_1);
nand_5 g14888(new_n17236_1, new_n17235, new_n17237);
and_5  g14889(new_n17237, new_n17232_1, new_n17238);
nand_5 g14890(new_n17238, new_n17229, new_n17239);
and_5  g14891(new_n17239, new_n17228, new_n17240);
xor_4  g14892(new_n17240, new_n17226, new_n17241);
not_10 g14893(new_n17241, new_n17242);
xor_4  g14894(new_n7626, n11736, new_n17243_1);
nand_5 g14895(new_n2451, n23200, new_n17244);
xor_4  g14896(new_n2451, new_n5492, new_n17245);
nand_5 g14897(new_n2455, n17959, new_n17246);
xor_4  g14898(new_n2455, new_n5496, new_n17247);
nand_5 g14899(new_n2461, n7566, new_n17248);
or_5   g14900(new_n6727, new_n6714, new_n17249);
and_5  g14901(new_n17249, new_n17248, new_n17250_1);
or_5   g14902(new_n17250_1, new_n17247, new_n17251_1);
and_5  g14903(new_n17251_1, new_n17246, new_n17252);
or_5   g14904(new_n17252, new_n17245, new_n17253);
and_5  g14905(new_n17253, new_n17244, new_n17254);
xor_4  g14906(new_n17254, new_n17243_1, new_n17255);
xor_4  g14907(new_n17255, new_n17242, new_n17256);
xor_4  g14908(new_n17238, new_n17229, new_n17257);
not_10 g14909(new_n17257, new_n17258);
xor_4  g14910(new_n17252, new_n17245, new_n17259);
or_5   g14911(new_n17259, new_n17258, new_n17260);
xor_4  g14912(new_n17259, new_n17258, new_n17261);
not_10 g14913(new_n17261, new_n17262);
xnor_4 g14914(new_n17250_1, new_n17247, new_n17263_1);
not_10 g14915(new_n17263_1, new_n17264);
xor_4  g14916(new_n17236_1, new_n17235, new_n17265);
or_5   g14917(new_n17265, new_n17264, new_n17266);
or_5   g14918(new_n8775, new_n6728, new_n17267);
not_10 g14919(new_n8776, new_n17268);
or_5   g14920(new_n8795, new_n17268, new_n17269);
and_5  g14921(new_n17269, new_n17267, new_n17270);
xor_4  g14922(new_n17265, new_n17264, new_n17271);
not_10 g14923(new_n17271, new_n17272);
or_5   g14924(new_n17272, new_n17270, new_n17273);
and_5  g14925(new_n17273, new_n17266, new_n17274);
or_5   g14926(new_n17274, new_n17262, new_n17275);
and_5  g14927(new_n17275, new_n17260, new_n17276);
xor_4  g14928(new_n17276, new_n17256, n4103);
nor_5  g14929(new_n15118_1, new_n13062, new_n17278);
not_10 g14930(new_n17278, new_n17279);
xor_4  g14931(new_n15118_1, new_n13062, new_n17280);
or_5   g14932(new_n15121, new_n12989, new_n17281);
nor_5  g14933(new_n15125, new_n12995, new_n17282);
not_10 g14934(new_n17282, new_n17283);
xnor_4 g14935(new_n15125, new_n12995, new_n17284);
nand_5 g14936(new_n15129, new_n13001, new_n17285_1);
xnor_4 g14937(new_n15129, new_n13001, new_n17286);
or_5   g14938(new_n15132, new_n13007, new_n17287);
xor_4  g14939(new_n16619, new_n13007, new_n17288);
nand_5 g14940(new_n15047, new_n13013, new_n17289);
and_5  g14941(new_n13018, new_n4247, new_n17290);
xnor_4 g14942(new_n13018, new_n4246, new_n17291);
or_5   g14943(new_n13023, new_n4252, new_n17292);
xnor_4 g14944(new_n13023, new_n4251, new_n17293);
nand_5 g14945(new_n13026_1, new_n4256_1, new_n17294);
xor_4  g14946(new_n13027, new_n4256_1, new_n17295);
nand_5 g14947(new_n13032, new_n4259, new_n17296);
and_5  g14948(new_n13034, new_n4261, new_n17297);
not_10 g14949(new_n17297, new_n17298);
xor_4  g14950(new_n13032, new_n4259, new_n17299);
nand_5 g14951(new_n17299, new_n17298, new_n17300);
and_5  g14952(new_n17300, new_n17296, new_n17301);
or_5   g14953(new_n17301, new_n17295, new_n17302_1);
and_5  g14954(new_n17302_1, new_n17294, new_n17303);
nand_5 g14955(new_n17303, new_n17293, new_n17304);
and_5  g14956(new_n17304, new_n17292, new_n17305);
and_5  g14957(new_n17305, new_n17291, new_n17306);
or_5   g14958(new_n17306, new_n17290, new_n17307);
xor_4  g14959(new_n15047, new_n13013, new_n17308);
nand_5 g14960(new_n17308, new_n17307, new_n17309);
and_5  g14961(new_n17309, new_n17289, new_n17310);
or_5   g14962(new_n17310, new_n17288, new_n17311);
and_5  g14963(new_n17311, new_n17287, new_n17312);
or_5   g14964(new_n17312, new_n17286, new_n17313);
and_5  g14965(new_n17313, new_n17285_1, new_n17314);
nor_5  g14966(new_n17314, new_n17284, new_n17315);
not_10 g14967(new_n17315, new_n17316);
and_5  g14968(new_n17316, new_n17283, new_n17317);
xnor_4 g14969(new_n15121, new_n12989, new_n17318);
or_5   g14970(new_n17318, new_n17317, new_n17319);
and_5  g14971(new_n17319, new_n17281, new_n17320_1);
and_5  g14972(new_n17320_1, new_n17280, new_n17321);
not_10 g14973(new_n17321, new_n17322);
and_5  g14974(new_n17322, new_n17279, new_n17323);
and_5  g14975(new_n5922, n6456, new_n17324);
not_10 g14976(new_n17324, new_n17325);
nor_5  g14977(new_n5922, n6456, new_n17326);
nor_5  g14978(new_n5969, n4085, new_n17327);
xor_4  g14979(new_n5969, n4085, new_n17328);
not_10 g14980(new_n17328, new_n17329);
or_5   g14981(new_n5974, n26725, new_n17330);
xor_4  g14982(new_n5974, n26725, new_n17331);
not_10 g14983(new_n17331, new_n17332);
or_5   g14984(new_n5980_1, n11980, new_n17333);
xor_4  g14985(new_n5980_1, n11980, new_n17334);
not_10 g14986(new_n17334, new_n17335);
or_5   g14987(new_n5986, n3253, new_n17336);
xor_4  g14988(new_n5986, n3253, new_n17337_1);
not_10 g14989(new_n17337_1, new_n17338);
or_5   g14990(new_n5992, n7759, new_n17339);
xor_4  g14991(new_n5992, n7759, new_n17340);
not_10 g14992(new_n17340, new_n17341);
or_5   g14993(new_n5998, n12562, new_n17342);
nor_5  g14994(new_n6003, n7949, new_n17343);
xor_4  g14995(new_n6003, new_n13350, new_n17344_1);
or_5   g14996(new_n6014, n24374, new_n17345);
nand_5 g14997(n20658, n14575, new_n17346);
xor_4  g14998(new_n6014, n24374, new_n17347);
nand_5 g14999(new_n17347, new_n17346, new_n17348);
and_5  g15000(new_n17348, new_n17345, new_n17349);
nor_5  g15001(new_n17349, new_n17344_1, new_n17350);
or_5   g15002(new_n17350, new_n17343, new_n17351_1);
xor_4  g15003(new_n5998, n12562, new_n17352);
nand_5 g15004(new_n17352, new_n17351_1, new_n17353);
and_5  g15005(new_n17353, new_n17342, new_n17354);
or_5   g15006(new_n17354, new_n17341, new_n17355);
and_5  g15007(new_n17355, new_n17339, new_n17356);
or_5   g15008(new_n17356, new_n17338, new_n17357);
and_5  g15009(new_n17357, new_n17336, new_n17358);
or_5   g15010(new_n17358, new_n17335, new_n17359_1);
and_5  g15011(new_n17359_1, new_n17333, new_n17360);
or_5   g15012(new_n17360, new_n17332, new_n17361);
and_5  g15013(new_n17361, new_n17330, new_n17362);
nor_5  g15014(new_n17362, new_n17329, new_n17363);
nor_5  g15015(new_n17363, new_n17327, new_n17364);
not_10 g15016(new_n17364, new_n17365);
nor_5  g15017(new_n17365, new_n17326, new_n17366);
nor_5  g15018(new_n17366, new_n14096, new_n17367);
and_5  g15019(new_n17367, new_n17325, new_n17368);
not_10 g15020(new_n17368, new_n17369);
nor_5  g15021(new_n17369, new_n17323, new_n17370);
xor_4  g15022(new_n17320_1, new_n17280, new_n17371);
nor_5  g15023(new_n17371, new_n17368, new_n17372);
xor_4  g15024(new_n17371, new_n17368, new_n17373);
not_10 g15025(new_n17373, new_n17374);
xor_4  g15026(new_n15121, new_n12989, new_n17375);
xnor_4 g15027(new_n17375, new_n17317, new_n17376);
xor_4  g15028(new_n5922, n6456, new_n17377);
xor_4  g15029(new_n17377, new_n17365, new_n17378);
and_5  g15030(new_n17378, new_n17376, new_n17379);
xor_4  g15031(new_n17378, new_n17376, new_n17380);
xor_4  g15032(new_n17362, new_n17329, new_n17381);
xor_4  g15033(new_n17314, new_n17284, new_n17382);
and_5  g15034(new_n17382, new_n17381, new_n17383);
xor_4  g15035(new_n17382, new_n17381, new_n17384);
xor_4  g15036(new_n17360, new_n17332, new_n17385);
xor_4  g15037(new_n17312, new_n17286, new_n17386);
and_5  g15038(new_n17386, new_n17385, new_n17387_1);
xor_4  g15039(new_n17386, new_n17385, new_n17388);
xor_4  g15040(new_n17358, new_n17335, new_n17389);
xor_4  g15041(new_n17310, new_n17288, new_n17390);
and_5  g15042(new_n17390, new_n17389, new_n17391_1);
xor_4  g15043(new_n17390, new_n17389, new_n17392_1);
xor_4  g15044(new_n17356, new_n17338, new_n17393);
xor_4  g15045(new_n17308, new_n17307, new_n17394);
and_5  g15046(new_n17394, new_n17393, new_n17395);
xor_4  g15047(new_n17394, new_n17393, new_n17396);
xor_4  g15048(new_n17354, new_n17341, new_n17397);
xor_4  g15049(new_n17305, new_n17291, new_n17398);
and_5  g15050(new_n17398, new_n17397, new_n17399);
xor_4  g15051(new_n17398, new_n17397, new_n17400);
xor_4  g15052(new_n17303, new_n17293, new_n17401);
not_10 g15053(new_n17401, new_n17402);
xor_4  g15054(new_n17352, new_n17351_1, new_n17403);
and_5  g15055(new_n17403, new_n17402, new_n17404);
xor_4  g15056(new_n17403, new_n17402, new_n17405);
xor_4  g15057(new_n17349, new_n17344_1, new_n17406);
xor_4  g15058(new_n17301, new_n17295, new_n17407);
nor_5  g15059(new_n17407, new_n17406, new_n17408);
xor_4  g15060(new_n17407, new_n17406, new_n17409);
xor_4  g15061(new_n17299, new_n17298, new_n17410);
not_10 g15062(new_n17410, new_n17411);
or_5   g15063(new_n17411, new_n17347, new_n17412);
xor_4  g15064(new_n17347, new_n17346, new_n17413);
nor_5  g15065(new_n17413, new_n17410, new_n17414);
xor_4  g15066(n20658, n14575, new_n17415);
xor_4  g15067(new_n13034, new_n4261, new_n17416);
and_5  g15068(new_n17416, new_n17415, new_n17417);
or_5   g15069(new_n17417, new_n17414, new_n17418);
and_5  g15070(new_n17418, new_n17412, new_n17419);
and_5  g15071(new_n17419, new_n17409, new_n17420);
nor_5  g15072(new_n17420, new_n17408, new_n17421_1);
and_5  g15073(new_n17421_1, new_n17405, new_n17422);
nor_5  g15074(new_n17422, new_n17404, new_n17423);
not_10 g15075(new_n17423, new_n17424);
and_5  g15076(new_n17424, new_n17400, new_n17425);
nor_5  g15077(new_n17425, new_n17399, new_n17426);
not_10 g15078(new_n17426, new_n17427);
and_5  g15079(new_n17427, new_n17396, new_n17428);
nor_5  g15080(new_n17428, new_n17395, new_n17429);
not_10 g15081(new_n17429, new_n17430);
and_5  g15082(new_n17430, new_n17392_1, new_n17431);
nor_5  g15083(new_n17431, new_n17391_1, new_n17432_1);
not_10 g15084(new_n17432_1, new_n17433);
and_5  g15085(new_n17433, new_n17388, new_n17434);
nor_5  g15086(new_n17434, new_n17387_1, new_n17435);
not_10 g15087(new_n17435, new_n17436_1);
and_5  g15088(new_n17436_1, new_n17384, new_n17437);
nor_5  g15089(new_n17437, new_n17383, new_n17438);
not_10 g15090(new_n17438, new_n17439);
and_5  g15091(new_n17439, new_n17380, new_n17440_1);
nor_5  g15092(new_n17440_1, new_n17379, new_n17441);
nor_5  g15093(new_n17441, new_n17374, new_n17442);
nor_5  g15094(new_n17442, new_n17372, new_n17443);
or_5   g15095(new_n17443, new_n17370, new_n17444);
and_5  g15096(new_n17369, new_n17323, new_n17445);
or_5   g15097(new_n17445, new_n17442, new_n17446);
and_5  g15098(new_n17446, new_n17444, n4123);
xor_4  g15099(new_n13582, new_n8007, new_n17448);
nand_5 g15100(new_n13586, new_n8014, new_n17449);
xnor_4 g15101(new_n13587, new_n8014, new_n17450_1);
or_5   g15102(new_n13591, new_n8031_1, new_n17451);
xor_4  g15103(new_n13591, new_n8031_1, new_n17452);
and_5  g15104(new_n13602_1, new_n8022, new_n17453);
and_5  g15105(new_n9951, new_n8024, new_n17454);
xnor_4 g15106(new_n13602_1, new_n8021, new_n17455);
and_5  g15107(new_n17455, new_n17454, new_n17456);
nor_5  g15108(new_n17456, new_n17453, new_n17457);
nand_5 g15109(new_n17457, new_n17452, new_n17458_1);
nand_5 g15110(new_n17458_1, new_n17451, new_n17459);
nand_5 g15111(new_n17459, new_n17450_1, new_n17460);
and_5  g15112(new_n17460, new_n17449, new_n17461_1);
xor_4  g15113(new_n17461_1, new_n17448, n4134);
xor_4  g15114(new_n9282, new_n9211, n4146);
xnor_4 g15115(new_n15695, new_n14552, new_n17464);
not_10 g15116(new_n14557, new_n17465);
nor_5  g15117(new_n15699, new_n17465, new_n17466_1);
xnor_4 g15118(new_n15699, new_n14557, new_n17467);
nand_5 g15119(new_n14560, new_n15703, new_n17468);
or_5   g15120(new_n14563, new_n13666, new_n17469);
xnor_4 g15121(new_n14560, new_n13671, new_n17470);
not_10 g15122(new_n17470, new_n17471);
or_5   g15123(new_n17471, new_n17469, new_n17472);
and_5  g15124(new_n17472, new_n17468, new_n17473);
and_5  g15125(new_n17473, new_n17467, new_n17474);
nor_5  g15126(new_n17474, new_n17466_1, new_n17475);
xnor_4 g15127(new_n17475, new_n17464, n4150);
xor_4  g15128(new_n12809, new_n12807, n4151);
xnor_4 g15129(new_n13143, new_n13074_1, n4152);
xor_4  g15130(new_n6183_1, new_n6142, n4153);
and_5  g15131(n25972, new_n12189, new_n17480);
not_10 g15132(new_n17480, new_n17481);
nor_5  g15133(new_n8845, new_n8797, new_n17482);
not_10 g15134(new_n17482, new_n17483);
and_5  g15135(new_n17483, new_n17481, new_n17484);
xor_4  g15136(new_n17484, new_n12486, new_n17485);
nand_5 g15137(new_n17484, new_n12490, new_n17486);
nor_5  g15138(new_n17484, new_n12490, new_n17487);
and_5  g15139(new_n9019, new_n8846, new_n17488);
not_10 g15140(new_n17488, new_n17489);
and_5  g15141(new_n9087, new_n9020, new_n17490);
not_10 g15142(new_n17490, new_n17491);
and_5  g15143(new_n17491, new_n17489, new_n17492);
or_5   g15144(new_n17492, new_n17487, new_n17493_1);
and_5  g15145(new_n17493_1, new_n17486, new_n17494);
xor_4  g15146(new_n17494, new_n17485, n4165);
xnor_4 g15147(new_n11752, new_n11719, n4172);
xor_4  g15148(new_n11571, new_n4754, n4173);
xnor_4 g15149(new_n6623, new_n6602, n4176);
xnor_4 g15150(new_n9256, new_n9255, n4186);
xnor_4 g15151(new_n17047, new_n17021, n4204);
not_10 g15152(new_n11657, new_n17501);
or_5   g15153(new_n11619, new_n11979, new_n17502);
xor_4  g15154(new_n11619, new_n11979, new_n17503);
not_10 g15155(new_n17503, new_n17504);
or_5   g15156(new_n6805, new_n5541, new_n17505);
or_5   g15157(new_n6846, new_n6807, new_n17506);
and_5  g15158(new_n17506, new_n17505, new_n17507);
or_5   g15159(new_n17507, new_n17504, new_n17508);
and_5  g15160(new_n17508, new_n17502, new_n17509);
nor_5  g15161(new_n17509, new_n17501, new_n17510);
and_5  g15162(new_n16399, new_n11762, new_n17511);
and_5  g15163(new_n17511, new_n11759, new_n17512);
xor_4  g15164(new_n17512, new_n11756, new_n17513);
and_5  g15165(new_n17513, new_n11660, new_n17514);
xor_4  g15166(new_n17513, new_n11660, new_n17515);
xor_4  g15167(new_n17511, new_n11759, new_n17516);
or_5   g15168(new_n17516, new_n11661, new_n17517);
nand_5 g15169(new_n16400, new_n11662, new_n17518);
or_5   g15170(new_n16428_1, new_n16401, new_n17519);
and_5  g15171(new_n17519, new_n17518, new_n17520);
xor_4  g15172(new_n17516, new_n11661, new_n17521);
nand_5 g15173(new_n17521, new_n17520, new_n17522);
and_5  g15174(new_n17522, new_n17517, new_n17523);
and_5  g15175(new_n17523, new_n17515, new_n17524_1);
nor_5  g15176(new_n17524_1, new_n17514, new_n17525);
and_5  g15177(new_n17512, new_n11756, new_n17526);
xor_4  g15178(new_n17526, new_n11843_1, new_n17527);
xor_4  g15179(new_n17527, new_n11659, new_n17528);
xor_4  g15180(new_n17528, new_n17525, new_n17529_1);
and_5  g15181(new_n17529_1, n25586, new_n17530);
xor_4  g15182(new_n17529_1, n25586, new_n17531);
not_10 g15183(new_n17531, new_n17532);
xor_4  g15184(new_n17523, new_n17515, new_n17533);
or_5   g15185(new_n17533, new_n14757, new_n17534);
xor_4  g15186(new_n17533, new_n14757, new_n17535);
xor_4  g15187(new_n17521, new_n17520, new_n17536);
or_5   g15188(new_n17536, n26053, new_n17537);
xor_4  g15189(new_n17536, new_n14760, new_n17538);
nand_5 g15190(new_n16429, new_n14763_1, new_n17539);
or_5   g15191(new_n16458, new_n16430, new_n17540);
and_5  g15192(new_n17540, new_n17539, new_n17541);
or_5   g15193(new_n17541, new_n17538, new_n17542);
and_5  g15194(new_n17542, new_n17537, new_n17543);
nand_5 g15195(new_n17543, new_n17535, new_n17544);
and_5  g15196(new_n17544, new_n17534, new_n17545);
nor_5  g15197(new_n17545, new_n17532, new_n17546);
nor_5  g15198(new_n17546, new_n17530, new_n17547);
not_10 g15199(new_n17547, new_n17548);
and_5  g15200(new_n17526, new_n11843_1, new_n17549);
nor_5  g15201(new_n17527, new_n11659, new_n17550);
nor_5  g15202(new_n17550, new_n17525, new_n17551);
and_5  g15203(new_n17551, new_n17549, new_n17552);
not_10 g15204(new_n17552, new_n17553);
nor_5  g15205(new_n17553, new_n17548, new_n17554);
nand_5 g15206(new_n17527, new_n11659, new_n17555);
xnor_4 g15207(new_n17551, new_n17549, new_n17556);
and_5  g15208(new_n17556, new_n17555, new_n17557_1);
and_5  g15209(new_n17557_1, new_n17548, new_n17558);
and_5  g15210(new_n17558, new_n17553, new_n17559);
nor_5  g15211(new_n17559, new_n17554, new_n17560);
or_5   g15212(new_n17560, new_n17510, new_n17561);
xor_4  g15213(new_n17557_1, new_n17548, new_n17562);
xnor_4 g15214(new_n17509, new_n11657, new_n17563);
not_10 g15215(new_n17563, new_n17564);
and_5  g15216(new_n17564, new_n17562, new_n17565);
xor_4  g15217(new_n17564, new_n17562, new_n17566);
xor_4  g15218(new_n17545, new_n17532, new_n17567);
xor_4  g15219(new_n17507, new_n17504, new_n17568);
not_10 g15220(new_n17568, new_n17569);
and_5  g15221(new_n17569, new_n17567, new_n17570);
xor_4  g15222(new_n17569, new_n17567, new_n17571);
not_10 g15223(new_n6847, new_n17572);
xor_4  g15224(new_n17543, new_n17535, new_n17573);
and_5  g15225(new_n17573, new_n17572, new_n17574);
xor_4  g15226(new_n17573, new_n17572, new_n17575);
xor_4  g15227(new_n17541, new_n17538, new_n17576);
nor_5  g15228(new_n17576, new_n6928, new_n17577);
or_5   g15229(new_n16459, new_n6934, new_n17578);
not_10 g15230(new_n16460_1, new_n17579);
or_5   g15231(new_n16491, new_n17579, new_n17580);
and_5  g15232(new_n17580, new_n17578, new_n17581);
xor_4  g15233(new_n17576, new_n6928, new_n17582);
not_10 g15234(new_n17582, new_n17583_1);
nor_5  g15235(new_n17583_1, new_n17581, new_n17584);
nor_5  g15236(new_n17584, new_n17577, new_n17585);
not_10 g15237(new_n17585, new_n17586);
and_5  g15238(new_n17586, new_n17575, new_n17587);
nor_5  g15239(new_n17587, new_n17574, new_n17588);
not_10 g15240(new_n17588, new_n17589);
and_5  g15241(new_n17589, new_n17571, new_n17590);
nor_5  g15242(new_n17590, new_n17570, new_n17591);
not_10 g15243(new_n17591, new_n17592_1);
and_5  g15244(new_n17592_1, new_n17566, new_n17593);
nor_5  g15245(new_n17593, new_n17565, new_n17594);
nand_5 g15246(new_n17594, new_n17561, new_n17595);
and_5  g15247(new_n17560, new_n17510, new_n17596);
nor_5  g15248(new_n17596, new_n17554, new_n17597);
and_5  g15249(new_n17597, new_n17595, n4205);
and_5  g15250(new_n13503, new_n4935, new_n17599);
and_5  g15251(new_n17599, new_n4931, new_n17600);
xor_4  g15252(new_n17600, new_n4927, new_n17601);
xor_4  g15253(new_n17601, new_n8349, new_n17602);
xor_4  g15254(new_n17599, new_n4931, new_n17603);
or_5   g15255(new_n17603, n24638, new_n17604);
xor_4  g15256(new_n17603, new_n8350, new_n17605);
or_5   g15257(new_n13504, n21674, new_n17606);
or_5   g15258(new_n13526, new_n13505, new_n17607);
and_5  g15259(new_n17607, new_n17606, new_n17608);
or_5   g15260(new_n17608, new_n17605, new_n17609);
and_5  g15261(new_n17609, new_n17604, new_n17610);
xor_4  g15262(new_n17610, new_n17602, new_n17611);
xor_4  g15263(new_n17611, new_n7844, new_n17612);
not_10 g15264(new_n7850, new_n17613);
xor_4  g15265(new_n17608, new_n17605, new_n17614);
or_5   g15266(new_n17614, new_n17613, new_n17615);
xnor_4 g15267(new_n17614, new_n7850, new_n17616);
not_10 g15268(new_n7855, new_n17617);
nand_5 g15269(new_n13527, new_n17617, new_n17618);
or_5   g15270(new_n13553, new_n13529, new_n17619);
and_5  g15271(new_n17619, new_n17618, new_n17620);
nand_5 g15272(new_n17620, new_n17616, new_n17621);
and_5  g15273(new_n17621, new_n17615, new_n17622);
xor_4  g15274(new_n17622, new_n17612, new_n17623);
xor_4  g15275(n21997, n5400, new_n17624);
not_10 g15276(n23923, new_n17625);
or_5   g15277(n25119, new_n17625, new_n17626);
xor_4  g15278(n25119, n23923, new_n17627);
nand_5 g15279(new_n8654, n329, new_n17628);
or_5   g15280(new_n13576, new_n13555, new_n17629);
and_5  g15281(new_n17629, new_n17628, new_n17630);
or_5   g15282(new_n17630, new_n17627, new_n17631);
and_5  g15283(new_n17631, new_n17626, new_n17632);
xor_4  g15284(new_n17632, new_n17624, new_n17633);
xnor_4 g15285(new_n17633, new_n17623, new_n17634);
xor_4  g15286(new_n17630, new_n17627, new_n17635);
xor_4  g15287(new_n17620, new_n17616, new_n17636);
nand_5 g15288(new_n17636, new_n17635, new_n17637);
xor_4  g15289(new_n17636, new_n17635, new_n17638_1);
not_10 g15290(new_n13577, new_n17639);
nand_5 g15291(new_n17639, new_n13554, new_n17640);
or_5   g15292(new_n13613, new_n13579, new_n17641);
and_5  g15293(new_n17641, new_n17640, new_n17642);
nand_5 g15294(new_n17642, new_n17638_1, new_n17643);
and_5  g15295(new_n17643, new_n17637, new_n17644);
xor_4  g15296(new_n17644, new_n17634, n4215);
not_10 g15297(n3582, new_n17646);
and_5  g15298(new_n14602, new_n7782, new_n17647);
xor_4  g15299(new_n17647, new_n17646, new_n17648);
xor_4  g15300(new_n17648, n3740, new_n17649);
nand_5 g15301(new_n14603_1, n2858, new_n17650);
or_5   g15302(new_n14603_1, n2858, new_n17651);
nand_5 g15303(new_n14627, new_n17651, new_n17652);
and_5  g15304(new_n17652, new_n17650, new_n17653);
xnor_4 g15305(new_n17653, new_n17649, new_n17654);
and_5  g15306(new_n9857, new_n4304, new_n17655);
xor_4  g15307(new_n17655, new_n4301, new_n17656);
xor_4  g15308(new_n17656, n22626, new_n17657);
nor_5  g15309(new_n9858, n14440, new_n17658);
xor_4  g15310(new_n9858, n14440, new_n17659);
not_10 g15311(new_n17659, new_n17660);
or_5   g15312(new_n9860, n1654, new_n17661);
or_5   g15313(new_n16167_1, new_n16164, new_n17662);
and_5  g15314(new_n17662, new_n17661, new_n17663);
nor_5  g15315(new_n17663, new_n17660, new_n17664_1);
nor_5  g15316(new_n17664_1, new_n17658, new_n17665);
xnor_4 g15317(new_n17665, new_n17657, new_n17666);
not_10 g15318(new_n17666, new_n17667);
xor_4  g15319(new_n17667, new_n17654, new_n17668);
xor_4  g15320(new_n17663, new_n17660, new_n17669);
or_5   g15321(new_n17669, new_n14628, new_n17670);
nand_5 g15322(new_n16168, new_n14630, new_n17671);
xor_4  g15323(new_n16168, new_n14630, new_n17672);
not_10 g15324(new_n17672, new_n17673);
nand_5 g15325(new_n14632, new_n10847, new_n17674);
xor_4  g15326(new_n14632, new_n10847, new_n17675);
not_10 g15327(new_n17675, new_n17676);
nand_5 g15328(new_n14635, new_n10849, new_n17677);
xnor_4 g15329(new_n14635, new_n10850, new_n17678);
nand_5 g15330(new_n14638, new_n10857, new_n17679);
xnor_4 g15331(new_n14638, new_n10857, new_n17680);
or_5   g15332(new_n9665, new_n9650, new_n17681);
not_10 g15333(new_n9666, new_n17682);
or_5   g15334(new_n9681, new_n17682, new_n17683);
and_5  g15335(new_n17683, new_n17681, new_n17684);
or_5   g15336(new_n17684, new_n17680, new_n17685);
and_5  g15337(new_n17685, new_n17679, new_n17686);
nand_5 g15338(new_n17686, new_n17678, new_n17687_1);
and_5  g15339(new_n17687_1, new_n17677, new_n17688);
or_5   g15340(new_n17688, new_n17676, new_n17689);
and_5  g15341(new_n17689, new_n17674, new_n17690);
or_5   g15342(new_n17690, new_n17673, new_n17691);
and_5  g15343(new_n17691, new_n17671, new_n17692);
not_10 g15344(new_n17669, new_n17693);
xnor_4 g15345(new_n17693, new_n14628, new_n17694);
nand_5 g15346(new_n17694, new_n17692, new_n17695);
and_5  g15347(new_n17695, new_n17670, new_n17696);
xor_4  g15348(new_n17696, new_n17668, new_n17697);
not_10 g15349(new_n17697, new_n17698);
not_10 g15350(n23166, new_n17699);
and_5  g15351(new_n15368, new_n9324, new_n17700);
and_5  g15352(new_n17700, new_n9321, new_n17701);
and_5  g15353(new_n17701, new_n9318_1, new_n17702);
and_5  g15354(new_n17702, new_n9315, new_n17703);
and_5  g15355(new_n17703, new_n9312, new_n17704);
and_5  g15356(new_n17704, new_n9309, new_n17705);
xor_4  g15357(new_n17705, new_n17699, new_n17706);
xor_4  g15358(new_n17706, new_n7908, new_n17707);
xor_4  g15359(new_n17704, new_n9309, new_n17708);
nor_5  g15360(new_n17708, n26408, new_n17709);
xor_4  g15361(new_n17708, n26408, new_n17710);
not_10 g15362(new_n17710, new_n17711);
xor_4  g15363(new_n17703, new_n9312, new_n17712);
or_5   g15364(new_n17712, n18227, new_n17713);
xor_4  g15365(new_n17712, n18227, new_n17714);
not_10 g15366(new_n17714, new_n17715);
xor_4  g15367(new_n17702, new_n9315, new_n17716);
or_5   g15368(new_n17716, n7377, new_n17717);
xor_4  g15369(new_n17716, n7377, new_n17718);
not_10 g15370(new_n17718, new_n17719);
xor_4  g15371(new_n17701, new_n9318_1, new_n17720);
or_5   g15372(new_n17720, n11630, new_n17721_1);
xor_4  g15373(new_n17700, new_n9321, new_n17722);
nor_5  g15374(new_n17722, n13453, new_n17723);
xor_4  g15375(new_n17722, n13453, new_n17724);
nand_5 g15376(new_n15369, n7421, new_n17725);
or_5   g15377(new_n15381, new_n15370, new_n17726);
and_5  g15378(new_n17726, new_n17725, new_n17727);
and_5  g15379(new_n17727, new_n17724, new_n17728);
or_5   g15380(new_n17728, new_n17723, new_n17729);
xor_4  g15381(new_n17720, n11630, new_n17730);
nand_5 g15382(new_n17730, new_n17729, new_n17731);
and_5  g15383(new_n17731, new_n17721_1, new_n17732);
or_5   g15384(new_n17732, new_n17719, new_n17733);
and_5  g15385(new_n17733, new_n17717, new_n17734);
or_5   g15386(new_n17734, new_n17715, new_n17735_1);
and_5  g15387(new_n17735_1, new_n17713, new_n17736);
nor_5  g15388(new_n17736, new_n17711, new_n17737);
nor_5  g15389(new_n17737, new_n17709, new_n17738_1);
xor_4  g15390(new_n17738_1, new_n17707, new_n17739);
xnor_4 g15391(new_n17739, new_n17698, new_n17740);
xor_4  g15392(new_n17736, new_n17711, new_n17741);
not_10 g15393(new_n17741, new_n17742);
xor_4  g15394(new_n17694, new_n17692, new_n17743);
nor_5  g15395(new_n17743, new_n17742, new_n17744);
xor_4  g15396(new_n17743, new_n17742, new_n17745);
not_10 g15397(new_n17745, new_n17746_1);
xor_4  g15398(new_n17734, new_n17715, new_n17747);
not_10 g15399(new_n17747, new_n17748);
xor_4  g15400(new_n17690, new_n17673, new_n17749_1);
not_10 g15401(new_n17749_1, new_n17750);
nor_5  g15402(new_n17750, new_n17748, new_n17751);
not_10 g15403(new_n17751, new_n17752);
xor_4  g15404(new_n17750, new_n17748, new_n17753);
xor_4  g15405(new_n17732, new_n17719, new_n17754);
not_10 g15406(new_n17754, new_n17755);
xor_4  g15407(new_n17688, new_n17676, new_n17756);
not_10 g15408(new_n17756, new_n17757);
nor_5  g15409(new_n17757, new_n17755, new_n17758);
not_10 g15410(new_n17758, new_n17759);
xor_4  g15411(new_n17757, new_n17755, new_n17760);
xor_4  g15412(new_n17686, new_n17678, new_n17761);
xor_4  g15413(new_n17730, new_n17729, new_n17762);
and_5  g15414(new_n17762, new_n17761, new_n17763);
not_10 g15415(new_n17761, new_n17764);
xnor_4 g15416(new_n17762, new_n17764, new_n17765);
xor_4  g15417(new_n17727, new_n17724, new_n17766);
not_10 g15418(new_n17766, new_n17767);
xor_4  g15419(new_n17684, new_n17680, new_n17768);
nor_5  g15420(new_n17768, new_n17767, new_n17769);
xnor_4 g15421(new_n17768, new_n17766, new_n17770);
not_10 g15422(new_n17770, new_n17771);
not_10 g15423(new_n15382_1, new_n17772);
and_5  g15424(new_n17772, new_n9683, new_n17773);
xor_4  g15425(new_n17772, new_n9683, new_n17774);
and_5  g15426(new_n15384, new_n9699_1, new_n17775);
xor_4  g15427(new_n15384, new_n9700, new_n17776);
or_5   g15428(new_n15388, new_n9712, new_n17777);
and_5  g15429(new_n15390, new_n9706, new_n17778);
xor_4  g15430(new_n15388, new_n9712, new_n17779);
nand_5 g15431(new_n17779, new_n17778, new_n17780);
and_5  g15432(new_n17780, new_n17777, new_n17781);
nor_5  g15433(new_n17781, new_n17776, new_n17782);
nor_5  g15434(new_n17782, new_n17775, new_n17783);
and_5  g15435(new_n17783, new_n17774, new_n17784_1);
nor_5  g15436(new_n17784_1, new_n17773, new_n17785);
nor_5  g15437(new_n17785, new_n17771, new_n17786);
nor_5  g15438(new_n17786, new_n17769, new_n17787);
not_10 g15439(new_n17787, new_n17788);
and_5  g15440(new_n17788, new_n17765, new_n17789);
nor_5  g15441(new_n17789, new_n17763, new_n17790);
not_10 g15442(new_n17790, new_n17791);
and_5  g15443(new_n17791, new_n17760, new_n17792);
not_10 g15444(new_n17792, new_n17793);
and_5  g15445(new_n17793, new_n17759, new_n17794);
not_10 g15446(new_n17794, new_n17795);
and_5  g15447(new_n17795, new_n17753, new_n17796);
not_10 g15448(new_n17796, new_n17797);
and_5  g15449(new_n17797, new_n17752, new_n17798);
nor_5  g15450(new_n17798, new_n17746_1, new_n17799);
nor_5  g15451(new_n17799, new_n17744, new_n17800);
xor_4  g15452(new_n17800, new_n17740, n4221);
xor_4  g15453(new_n10760, new_n7910, new_n17802);
or_5   g15454(new_n10763_1, new_n7911, new_n17803);
xor_4  g15455(new_n10763_1, n7377, new_n17804);
or_5   g15456(new_n10767, new_n7912, new_n17805);
and_5  g15457(new_n10770, n13453, new_n17806);
nor_5  g15458(new_n13246, new_n13243, new_n17807);
or_5   g15459(new_n17807, new_n17806, new_n17808);
xor_4  g15460(new_n10767, new_n7912, new_n17809);
nand_5 g15461(new_n17809, new_n17808, new_n17810);
and_5  g15462(new_n17810, new_n17805, new_n17811);
or_5   g15463(new_n17811, new_n17804, new_n17812);
and_5  g15464(new_n17812, new_n17803, new_n17813);
xor_4  g15465(new_n17813, new_n17802, new_n17814);
xor_4  g15466(new_n17814, new_n16551, new_n17815);
not_10 g15467(new_n17815, new_n17816);
xor_4  g15468(new_n17811, new_n17804, new_n17817);
nand_5 g15469(new_n17817, new_n16556, new_n17818);
xnor_4 g15470(new_n17817, new_n8651, new_n17819);
not_10 g15471(new_n17819, new_n17820_1);
xor_4  g15472(new_n17809, new_n17808, new_n17821);
nand_5 g15473(new_n17821, new_n8684, new_n17822);
xnor_4 g15474(new_n17821, new_n8683, new_n17823);
not_10 g15475(new_n17823, new_n17824);
nand_5 g15476(new_n13247, new_n16565, new_n17825);
xnor_4 g15477(new_n13247, new_n8690, new_n17826);
not_10 g15478(new_n17826, new_n17827);
not_10 g15479(new_n6663, new_n17828);
or_5   g15480(new_n8695, new_n17828, new_n17829);
xnor_4 g15481(new_n8695, new_n6663, new_n17830);
not_10 g15482(new_n17830, new_n17831);
not_10 g15483(new_n6692, new_n17832);
or_5   g15484(new_n8701, new_n17832, new_n17833);
xnor_4 g15485(new_n8704, new_n17832, new_n17834);
nand_5 g15486(new_n8706, new_n6697, new_n17835);
nor_5  g15487(new_n8711, new_n6701, new_n17836);
xnor_4 g15488(new_n8707, new_n6697, new_n17837);
nand_5 g15489(new_n17837, new_n17836, new_n17838);
nand_5 g15490(new_n17838, new_n17835, new_n17839);
nand_5 g15491(new_n17839, new_n17834, new_n17840);
and_5  g15492(new_n17840, new_n17833, new_n17841);
or_5   g15493(new_n17841, new_n17831, new_n17842);
and_5  g15494(new_n17842, new_n17829, new_n17843);
or_5   g15495(new_n17843, new_n17827, new_n17844);
and_5  g15496(new_n17844, new_n17825, new_n17845);
or_5   g15497(new_n17845, new_n17824, new_n17846);
and_5  g15498(new_n17846, new_n17822, new_n17847);
or_5   g15499(new_n17847, new_n17820_1, new_n17848);
and_5  g15500(new_n17848, new_n17818, new_n17849);
xnor_4 g15501(new_n17849, new_n17816, n4224);
xor_4  g15502(new_n10895, new_n10894, n4231);
xor_4  g15503(new_n14451, n9934, new_n17852);
nor_5  g15504(new_n14455, n18496, new_n17853);
nor_5  g15505(new_n17159, new_n17152, new_n17854);
nor_5  g15506(new_n17854, new_n17853, new_n17855_1);
xnor_4 g15507(new_n17855_1, new_n17852, new_n17856);
not_10 g15508(new_n17856, new_n17857);
xor_4  g15509(new_n17857, n2979, new_n17858);
nor_5  g15510(new_n17160, new_n5911_1, new_n17859);
nor_5  g15511(new_n17169, new_n17161, new_n17860);
nor_5  g15512(new_n17860, new_n17859, new_n17861);
not_10 g15513(new_n17861, new_n17862);
xor_4  g15514(new_n17862, new_n17858, new_n17863);
xor_4  g15515(new_n17863, new_n12117, new_n17864);
or_5   g15516(new_n17170, new_n12121_1, new_n17865);
not_10 g15517(new_n17171, new_n17866);
or_5   g15518(new_n17181, new_n17866, new_n17867);
nand_5 g15519(new_n17867, new_n17865, new_n17868);
xnor_4 g15520(new_n17868, new_n17864, n4266);
xnor_4 g15521(new_n6979, new_n6948, n4340);
xnor_4 g15522(new_n16769, new_n6006, new_n17871);
xnor_4 g15523(new_n17871, new_n13348, new_n17872);
or_5   g15524(new_n16770, new_n13354, new_n17873);
nand_5 g15525(new_n16771, new_n16767, new_n17874);
and_5  g15526(new_n17874, new_n17873, new_n17875);
xor_4  g15527(new_n17875, new_n17872, new_n17876);
xnor_4 g15528(new_n17876, new_n5019, new_n17877_1);
or_5   g15529(new_n16772, new_n16766, new_n17878);
and_5  g15530(new_n17878, new_n16765, new_n17879);
xor_4  g15531(new_n17879, new_n17877_1, n4374);
xnor_4 g15532(new_n11391_1, new_n11341, n4401);
xor_4  g15533(new_n13294, new_n13293, n4424);
not_10 g15534(n1881, new_n17883);
nor_5  g15535(new_n10964, new_n17883, new_n17884);
xor_4  g15536(new_n10964, new_n17883, new_n17885);
not_10 g15537(n5834, new_n17886);
nand_5 g15538(new_n10957, new_n17886, new_n17887);
xor_4  g15539(new_n10957, new_n17886, new_n17888);
nand_5 g15540(new_n10971, n13851, new_n17889_1);
xnor_4 g15541(new_n10971, n13851, new_n17890);
nand_5 g15542(new_n10975, n24937, new_n17891);
or_5   g15543(new_n16666, new_n16658, new_n17892);
and_5  g15544(new_n17892, new_n17891, new_n17893);
or_5   g15545(new_n17893, new_n17890, new_n17894);
and_5  g15546(new_n17894, new_n17889_1, new_n17895);
nand_5 g15547(new_n17895, new_n17888, new_n17896);
and_5  g15548(new_n17896, new_n17887, new_n17897);
and_5  g15549(new_n17897, new_n17885, new_n17898);
or_5   g15550(new_n17898, new_n17884, new_n17899);
nor_5  g15551(n8827, n4306, new_n17900);
nor_5  g15552(new_n10963, new_n10960, new_n17901);
nor_5  g15553(new_n17901, new_n17900, new_n17902);
xor_4  g15554(new_n17902, new_n17899, new_n17903);
xnor_4 g15555(new_n17903, new_n10174, new_n17904);
not_10 g15556(new_n17904, new_n17905);
xor_4  g15557(new_n17897, new_n17885, new_n17906);
and_5  g15558(new_n17906, new_n10181, new_n17907);
xor_4  g15559(new_n17906, new_n10181, new_n17908);
not_10 g15560(new_n17908, new_n17909);
xor_4  g15561(new_n17895, new_n17888, new_n17910);
nor_5  g15562(new_n17910, new_n10186, new_n17911_1);
not_10 g15563(new_n17911_1, new_n17912_1);
xor_4  g15564(new_n17893, new_n17890, new_n17913);
nor_5  g15565(new_n17913, new_n10193, new_n17914);
xnor_4 g15566(new_n17913, new_n10193, new_n17915);
or_5   g15567(new_n16667, new_n10199, new_n17916);
or_5   g15568(new_n16676, new_n16668, new_n17917);
and_5  g15569(new_n17917, new_n17916, new_n17918);
nor_5  g15570(new_n17918, new_n17915, new_n17919);
nor_5  g15571(new_n17919, new_n17914, new_n17920);
xnor_4 g15572(new_n17910, new_n10185, new_n17921);
and_5  g15573(new_n17921, new_n17920, new_n17922);
not_10 g15574(new_n17922, new_n17923);
and_5  g15575(new_n17923, new_n17912_1, new_n17924);
nor_5  g15576(new_n17924, new_n17909, new_n17925);
nor_5  g15577(new_n17925, new_n17907, new_n17926);
xnor_4 g15578(new_n17926, new_n17905, n4432);
xnor_4 g15579(new_n15083, new_n15081, n4441);
nor_5  g15580(n27120, n23065, new_n17929);
and_5  g15581(new_n17929, new_n8823, new_n17930);
and_5  g15582(new_n17930, new_n8818, new_n17931_1);
and_5  g15583(new_n17931_1, new_n8814, new_n17932);
and_5  g15584(new_n17932, new_n8810, new_n17933);
and_5  g15585(new_n17933, new_n8806_1, new_n17934);
xor_4  g15586(new_n17934, new_n8802, new_n17935);
xor_4  g15587(new_n17935, new_n17224, new_n17936);
xor_4  g15588(new_n17933, n1293, new_n17937);
nand_5 g15589(new_n17937, new_n17227, new_n17938);
xnor_4 g15590(new_n17937, new_n17227, new_n17939);
xor_4  g15591(new_n17932, new_n8810, new_n17940);
or_5   g15592(new_n17940, new_n17231, new_n17941);
xor_4  g15593(new_n17931_1, new_n8814, new_n17942);
nor_5  g15594(new_n17942, new_n8753, new_n17943);
xor_4  g15595(new_n17942, new_n8753, new_n17944);
xor_4  g15596(new_n17930, new_n8818, new_n17945);
nand_5 g15597(new_n17945, new_n8755, new_n17946);
xor_4  g15598(new_n17945, new_n8755, new_n17947);
xor_4  g15599(new_n17929, new_n8823, new_n17948_1);
or_5   g15600(new_n17948_1, new_n8757, new_n17949);
xnor_4 g15601(new_n17948_1, new_n8757, new_n17950);
xor_4  g15602(n27120, n23065, new_n17951);
or_5   g15603(new_n17951, new_n8763, new_n17952);
and_5  g15604(new_n17952, new_n8766, new_n17953);
or_5   g15605(new_n17953, new_n17950, new_n17954_1);
and_5  g15606(new_n17954_1, new_n17949, new_n17955);
nand_5 g15607(new_n17955, new_n17947, new_n17956_1);
and_5  g15608(new_n17956_1, new_n17946, new_n17957);
and_5  g15609(new_n17957, new_n17944, new_n17958);
or_5   g15610(new_n17958, new_n17943, new_n17959_1);
xor_4  g15611(new_n17940, new_n17231, new_n17960);
nand_5 g15612(new_n17960, new_n17959_1, new_n17961);
and_5  g15613(new_n17961, new_n17941, new_n17962);
or_5   g15614(new_n17962, new_n17939, new_n17963_1);
and_5  g15615(new_n17963_1, new_n17938, new_n17964);
xor_4  g15616(new_n17964, new_n17936, new_n17965);
and_5  g15617(new_n12322, new_n8913, new_n17966);
xor_4  g15618(new_n17966, new_n8961, new_n17967);
xor_4  g15619(new_n17967, new_n5377, new_n17968_1);
or_5   g15620(new_n12323, new_n5382, new_n17969);
not_10 g15621(new_n12324_1, new_n17970);
or_5   g15622(new_n12353, new_n17970, new_n17971);
and_5  g15623(new_n17971, new_n17969, new_n17972);
xor_4  g15624(new_n17972, new_n17968_1, new_n17973);
xor_4  g15625(new_n17973, new_n17965, new_n17974);
not_10 g15626(new_n17974, new_n17975);
xor_4  g15627(new_n17962, new_n17939, new_n17976_1);
and_5  g15628(new_n17976_1, new_n12354, new_n17977);
xor_4  g15629(new_n17976_1, new_n12354, new_n17978);
not_10 g15630(new_n17978, new_n17979);
xor_4  g15631(new_n17960, new_n17959_1, new_n17980);
and_5  g15632(new_n17980, new_n12390, new_n17981);
not_10 g15633(new_n17981, new_n17982);
xor_4  g15634(new_n17980, new_n12390, new_n17983);
xor_4  g15635(new_n17957, new_n17944, new_n17984);
nor_5  g15636(new_n17984, new_n12393, new_n17985);
not_10 g15637(new_n12399, new_n17986);
xor_4  g15638(new_n17955, new_n17947, new_n17987);
or_5   g15639(new_n17987, new_n17986, new_n17988);
xor_4  g15640(new_n17987, new_n12399, new_n17989);
xor_4  g15641(new_n17953, new_n17950, new_n17990);
nor_5  g15642(new_n17990, new_n12404, new_n17991);
and_5  g15643(new_n17990, new_n12404, new_n17992);
not_10 g15644(new_n17992, new_n17993);
xnor_4 g15645(new_n17951, new_n8767, new_n17994);
and_5  g15646(new_n17994, new_n12413, new_n17995);
not_10 g15647(new_n8783, new_n17996);
nor_5  g15648(new_n12416, new_n17996, new_n17997);
xor_4  g15649(new_n17994, new_n12412, new_n17998_1);
or_5   g15650(new_n17998_1, new_n17997, new_n17999);
not_10 g15651(new_n17999, new_n18000);
nor_5  g15652(new_n18000, new_n17995, new_n18001);
and_5  g15653(new_n18001, new_n17993, new_n18002);
nor_5  g15654(new_n18002, new_n17991, new_n18003);
not_10 g15655(new_n18003, new_n18004);
or_5   g15656(new_n18004, new_n17989, new_n18005);
and_5  g15657(new_n18005, new_n17988, new_n18006);
xor_4  g15658(new_n17984, new_n12393, new_n18007);
and_5  g15659(new_n18007, new_n18006, new_n18008);
nor_5  g15660(new_n18008, new_n17985, new_n18009);
and_5  g15661(new_n18009, new_n17983, new_n18010);
not_10 g15662(new_n18010, new_n18011);
and_5  g15663(new_n18011, new_n17982, new_n18012);
nor_5  g15664(new_n18012, new_n17979, new_n18013);
nor_5  g15665(new_n18013, new_n17977, new_n18014);
xnor_4 g15666(new_n18014, new_n17975, n4451);
xor_4  g15667(n25494, n6659, new_n18016);
or_5   g15668(new_n16340, n10117, new_n18017);
xor_4  g15669(n23250, n10117, new_n18018);
or_5   g15670(n13460, new_n16272, new_n18019);
xor_4  g15671(n13460, n11455, new_n18020);
or_5   g15672(n6104, new_n16275_1, new_n18021);
xor_4  g15673(n6104, n3945, new_n18022);
or_5   g15674(new_n16278, n4119, new_n18023);
or_5   g15675(new_n5202, new_n5178, new_n18024);
and_5  g15676(new_n18024, new_n18023, new_n18025_1);
or_5   g15677(new_n18025_1, new_n18022, new_n18026);
and_5  g15678(new_n18026, new_n18021, new_n18027);
or_5   g15679(new_n18027, new_n18020, new_n18028);
and_5  g15680(new_n18028, new_n18019, new_n18029);
or_5   g15681(new_n18029, new_n18018, new_n18030);
and_5  g15682(new_n18030, new_n18017, new_n18031);
xnor_4 g15683(new_n18031, new_n18016, new_n18032);
xor_4  g15684(new_n18032, new_n13457_1, new_n18033);
xor_4  g15685(new_n18029, new_n18018, new_n18034);
not_10 g15686(new_n18034, new_n18035_1);
nand_5 g15687(new_n18035_1, new_n13463, new_n18036);
xnor_4 g15688(new_n18034, new_n13463, new_n18037);
not_10 g15689(new_n18037, new_n18038);
xnor_4 g15690(new_n18027, new_n18020, new_n18039);
nand_5 g15691(new_n18039, new_n13469, new_n18040);
xor_4  g15692(new_n18039, new_n13469, new_n18041);
xor_4  g15693(new_n18025_1, new_n18022, new_n18042);
and_5  g15694(new_n18042, new_n13475, new_n18043_1);
xnor_4 g15695(new_n18042, new_n13475, new_n18044);
nand_5 g15696(new_n5203, new_n5177, new_n18045_1);
nand_5 g15697(new_n5240, new_n5204, new_n18046);
and_5  g15698(new_n18046, new_n18045_1, new_n18047);
nor_5  g15699(new_n18047, new_n18044, new_n18048);
nor_5  g15700(new_n18048, new_n18043_1, new_n18049);
nand_5 g15701(new_n18049, new_n18041, new_n18050);
and_5  g15702(new_n18050, new_n18040, new_n18051);
or_5   g15703(new_n18051, new_n18038, new_n18052);
and_5  g15704(new_n18052, new_n18036, new_n18053);
xor_4  g15705(new_n18053, new_n18033, n4476);
not_10 g15706(n1831, new_n18055);
and_5  g15707(new_n4007, new_n4000_1, new_n18056);
and_5  g15708(new_n18056, new_n14216, new_n18057);
and_5  g15709(new_n18057, new_n14212, new_n18058);
and_5  g15710(new_n18058, new_n14208, new_n18059_1);
and_5  g15711(new_n18059_1, new_n18055, new_n18060);
xnor_4 g15712(new_n18060, new_n6273, new_n18061_1);
xor_4  g15713(new_n18059_1, new_n18055, new_n18062);
nor_5  g15714(new_n18062, new_n6280, new_n18063);
not_10 g15715(new_n18063, new_n18064);
xor_4  g15716(new_n18058, new_n14208, new_n18065);
nor_5  g15717(new_n18065, new_n6283, new_n18066);
xnor_4 g15718(new_n18065, new_n6283, new_n18067);
xor_4  g15719(new_n18057, new_n14212, new_n18068);
or_5   g15720(new_n18068, new_n6290, new_n18069);
xor_4  g15721(new_n18068, new_n6290, new_n18070);
xor_4  g15722(new_n18056, new_n14216, new_n18071_1);
nand_5 g15723(new_n18071_1, new_n6297, new_n18072);
xnor_4 g15724(new_n18071_1, new_n6297, new_n18073);
nand_5 g15725(new_n4045, new_n4008, new_n18074);
or_5   g15726(new_n4074, new_n4046, new_n18075);
and_5  g15727(new_n18075, new_n18074, new_n18076);
or_5   g15728(new_n18076, new_n18073, new_n18077);
and_5  g15729(new_n18077, new_n18072, new_n18078);
nand_5 g15730(new_n18078, new_n18070, new_n18079);
and_5  g15731(new_n18079, new_n18069, new_n18080);
nor_5  g15732(new_n18080, new_n18067, new_n18081);
or_5   g15733(new_n18081, new_n18066, new_n18082);
xor_4  g15734(new_n18062, new_n6280, new_n18083);
and_5  g15735(new_n18083, new_n18082, new_n18084);
not_10 g15736(new_n18084, new_n18085);
and_5  g15737(new_n18085, new_n18064, new_n18086);
xor_4  g15738(new_n18086, new_n18061_1, new_n18087);
xor_4  g15739(new_n18087, new_n11879, new_n18088);
xor_4  g15740(new_n18083, new_n18082, new_n18089);
and_5  g15741(new_n18089, new_n11884, new_n18090);
not_10 g15742(new_n18090, new_n18091);
xor_4  g15743(new_n18089, new_n11884, new_n18092);
not_10 g15744(new_n18092, new_n18093);
xor_4  g15745(new_n18080, new_n18067, new_n18094);
and_5  g15746(new_n18094, new_n11887, new_n18095);
not_10 g15747(new_n18095, new_n18096);
xnor_4 g15748(new_n18094, new_n11888, new_n18097);
not_10 g15749(new_n18097, new_n18098);
xor_4  g15750(new_n18078, new_n18070, new_n18099);
and_5  g15751(new_n18099, new_n11894, new_n18100);
not_10 g15752(new_n18100, new_n18101);
xnor_4 g15753(new_n18099, new_n11895, new_n18102);
not_10 g15754(new_n18102, new_n18103);
xor_4  g15755(new_n18076, new_n18073, new_n18104);
nor_5  g15756(new_n18104, new_n11902, new_n18105_1);
not_10 g15757(new_n18105_1, new_n18106);
xor_4  g15758(new_n18104, new_n11902, new_n18107);
not_10 g15759(new_n18107, new_n18108);
nor_5  g15760(new_n4075, new_n3999, new_n18109);
not_10 g15761(new_n18109, new_n18110);
not_10 g15762(new_n4076, new_n18111);
nor_5  g15763(new_n4112, new_n18111, new_n18112);
not_10 g15764(new_n18112, new_n18113);
and_5  g15765(new_n18113, new_n18110, new_n18114);
nor_5  g15766(new_n18114, new_n18108, new_n18115);
not_10 g15767(new_n18115, new_n18116);
and_5  g15768(new_n18116, new_n18106, new_n18117);
nor_5  g15769(new_n18117, new_n18103, new_n18118);
not_10 g15770(new_n18118, new_n18119);
and_5  g15771(new_n18119, new_n18101, new_n18120);
nor_5  g15772(new_n18120, new_n18098, new_n18121);
not_10 g15773(new_n18121, new_n18122);
and_5  g15774(new_n18122, new_n18096, new_n18123);
nor_5  g15775(new_n18123, new_n18093, new_n18124);
not_10 g15776(new_n18124, new_n18125);
and_5  g15777(new_n18125, new_n18091, new_n18126);
xor_4  g15778(new_n18126, new_n18088, n4478);
xnor_4 g15779(new_n12761, new_n12724, n4529);
xor_4  g15780(new_n6186, new_n6137, n4552);
xor_4  g15781(new_n6180, new_n6147, n4595);
xor_4  g15782(new_n14579, new_n14537, n4624);
not_10 g15783(new_n7833, new_n18132);
and_5  g15784(new_n17600, new_n4927, new_n18133);
xor_4  g15785(new_n18133, new_n4923, new_n18134);
nor_5  g15786(new_n18134, n14899, new_n18135);
xor_4  g15787(new_n18134, new_n8348, new_n18136);
or_5   g15788(new_n17601, n18444, new_n18137);
or_5   g15789(new_n17610, new_n17602, new_n18138);
and_5  g15790(new_n18138, new_n18137, new_n18139);
nor_5  g15791(new_n18139, new_n18136, new_n18140);
or_5   g15792(new_n18140, new_n18135, new_n18141);
and_5  g15793(new_n18133, new_n4923, new_n18142);
xor_4  g15794(new_n18142, new_n4919, new_n18143_1);
xor_4  g15795(new_n18143_1, n3506, new_n18144);
xor_4  g15796(new_n18144, new_n18141, new_n18145_1);
or_5   g15797(new_n18145_1, new_n18132, new_n18146);
xor_4  g15798(new_n18145_1, new_n7833, new_n18147);
not_10 g15799(new_n7838, new_n18148);
xor_4  g15800(new_n18139, new_n18136, new_n18149);
or_5   g15801(new_n18149, new_n18148, new_n18150);
xor_4  g15802(new_n18149, new_n7838, new_n18151_1);
or_5   g15803(new_n17611, new_n7845, new_n18152_1);
or_5   g15804(new_n17622, new_n17612, new_n18153);
and_5  g15805(new_n18153, new_n18152_1, new_n18154);
or_5   g15806(new_n18154, new_n18151_1, new_n18155);
and_5  g15807(new_n18155, new_n18150, new_n18156);
or_5   g15808(new_n18156, new_n18147, new_n18157_1);
and_5  g15809(new_n18157_1, new_n18146, new_n18158);
nand_5 g15810(new_n18142, new_n4919, new_n18159);
nand_5 g15811(new_n18143_1, n3506, new_n18160);
nor_5  g15812(new_n18143_1, n3506, new_n18161);
or_5   g15813(new_n18161, new_n18141, new_n18162);
and_5  g15814(new_n18162, new_n18160, new_n18163);
and_5  g15815(new_n18163, new_n18159, new_n18164);
xor_4  g15816(new_n18164, new_n18158, new_n18165);
xor_4  g15817(new_n18165, new_n7778, new_n18166);
xnor_4 g15818(new_n18166, new_n7975, new_n18167);
xor_4  g15819(new_n18156, new_n18147, new_n18168);
nor_5  g15820(new_n18168, new_n7981, new_n18169);
xor_4  g15821(new_n18154, new_n18151_1, new_n18170);
nor_5  g15822(new_n18170, new_n7987, new_n18171_1);
xnor_4 g15823(new_n18170, new_n7986, new_n18172);
not_10 g15824(new_n18172, new_n18173);
nor_5  g15825(new_n17623, new_n7993, new_n18174);
xnor_4 g15826(new_n17623, new_n7992_1, new_n18175);
not_10 g15827(new_n18175, new_n18176);
nor_5  g15828(new_n17636, new_n7999_1, new_n18177);
not_10 g15829(new_n18177, new_n18178);
xnor_4 g15830(new_n17636, new_n7998, new_n18179);
nor_5  g15831(new_n13554, new_n8003, new_n18180);
nand_5 g15832(new_n13582, new_n8007, new_n18181);
not_10 g15833(new_n17448, new_n18182);
or_5   g15834(new_n17461_1, new_n18182, new_n18183);
and_5  g15835(new_n18183, new_n18181, new_n18184);
xor_4  g15836(new_n13554, new_n8003, new_n18185);
and_5  g15837(new_n18185, new_n18184, new_n18186);
nor_5  g15838(new_n18186, new_n18180, new_n18187);
and_5  g15839(new_n18187, new_n18179, new_n18188);
not_10 g15840(new_n18188, new_n18189);
and_5  g15841(new_n18189, new_n18178, new_n18190);
nor_5  g15842(new_n18190, new_n18176, new_n18191);
nor_5  g15843(new_n18191, new_n18174, new_n18192);
nor_5  g15844(new_n18192, new_n18173, new_n18193_1);
nor_5  g15845(new_n18193_1, new_n18171_1, new_n18194);
xnor_4 g15846(new_n18168, new_n7980, new_n18195);
not_10 g15847(new_n18195, new_n18196);
nor_5  g15848(new_n18196, new_n18194, new_n18197);
nor_5  g15849(new_n18197, new_n18169, new_n18198);
xor_4  g15850(new_n18198, new_n18167, n4646);
xnor_4 g15851(new_n14592, new_n14515, n4674);
xor_4  g15852(n7057, n3480, new_n18201);
or_5   g15853(new_n7750, n8381, new_n18202);
or_5   g15854(n16722, new_n8663, new_n18203);
and_5  g15855(new_n5061, n11486, new_n18204);
and_5  g15856(n20235, new_n7754, new_n18205);
and_5  g15857(n13781, new_n5062_1, new_n18206);
not_10 g15858(new_n18206, new_n18207);
nor_5  g15859(new_n18207, new_n18205, new_n18208);
nor_5  g15860(new_n18208, new_n18204, new_n18209);
not_10 g15861(new_n18209, new_n18210);
nand_5 g15862(new_n18210, new_n18203, new_n18211);
and_5  g15863(new_n18211, new_n18202, new_n18212);
xor_4  g15864(new_n18212, new_n18201, new_n18213);
xnor_4 g15865(new_n18213, new_n3036, new_n18214);
xnor_4 g15866(n16722, n8381, new_n18215);
xor_4  g15867(new_n18215, new_n18210, new_n18216);
nand_5 g15868(new_n18216, new_n3041, new_n18217);
xor_4  g15869(new_n18216, new_n3041, new_n18218);
not_10 g15870(new_n3055, new_n18219);
xnor_4 g15871(n13781, n12495, new_n18220);
nor_5  g15872(new_n18220, new_n3048, new_n18221);
or_5   g15873(new_n18221, new_n18219, new_n18222);
xnor_4 g15874(new_n18221, new_n18219, new_n18223);
xnor_4 g15875(n20235, n11486, new_n18224);
xnor_4 g15876(new_n18224, new_n18207, new_n18225);
not_10 g15877(new_n18225, new_n18226);
or_5   g15878(new_n18226, new_n18223, new_n18227_1);
nand_5 g15879(new_n18227_1, new_n18222, new_n18228);
nand_5 g15880(new_n18228, new_n18218, new_n18229);
and_5  g15881(new_n18229, new_n18217, new_n18230);
xor_4  g15882(new_n18230, new_n18214, n4693);
xnor_4 g15883(new_n10897, new_n10889, n4731);
nor_5  g15884(new_n6070, new_n6035, new_n18233);
nor_5  g15885(new_n6125, new_n6072, new_n18234);
nor_5  g15886(new_n18234, new_n18233, new_n18235);
not_10 g15887(new_n18235, new_n18236);
nor_5  g15888(n21784, n3582, new_n18237);
not_10 g15889(new_n18237, new_n18238_1);
nor_5  g15890(new_n6069, new_n6036, new_n18239);
not_10 g15891(new_n18239, new_n18240);
and_5  g15892(new_n18240, new_n18238_1, new_n18241_1);
and_5  g15893(new_n18241_1, new_n18236, new_n18242);
xnor_4 g15894(new_n18242, new_n15734, new_n18243);
xor_4  g15895(new_n18241_1, new_n18236, new_n18244);
not_10 g15896(new_n18244, new_n18245);
and_5  g15897(new_n18245, new_n15738, new_n18246);
xnor_4 g15898(new_n18244, new_n15738, new_n18247);
not_10 g15899(new_n18247, new_n18248);
not_10 g15900(new_n6126, new_n18249);
and_5  g15901(new_n13170, new_n18249, new_n18250);
nor_5  g15902(new_n13220, new_n13172, new_n18251);
nor_5  g15903(new_n18251, new_n18250, new_n18252);
nor_5  g15904(new_n18252, new_n18248, new_n18253);
nor_5  g15905(new_n18253, new_n18246, new_n18254_1);
xnor_4 g15906(new_n18254_1, new_n18243, n4745);
xor_4  g15907(new_n6314, n6773, new_n18256);
xor_4  g15908(new_n18256, new_n9926_1, n4747);
xnor_4 g15909(new_n5804, new_n5803, n4766);
xnor_4 g15910(new_n14019, new_n14002, n4770);
xor_4  g15911(new_n16796, new_n15964, n4777);
xor_4  g15912(n17959, n6861, new_n18261);
nand_5 g15913(n19357, new_n5500, new_n18262);
xnor_4 g15914(n19357, n7566, new_n18263);
not_10 g15915(new_n18263, new_n18264);
nand_5 g15916(new_n5504, n2328, new_n18265);
xnor_4 g15917(n7731, n2328, new_n18266);
or_5   g15918(n15053, new_n5509, new_n18267);
nand_5 g15919(n15053, new_n5509, new_n18268);
and_5  g15920(new_n5087, n20986, new_n18269);
and_5  g15921(n25471, new_n5511, new_n18270);
not_10 g15922(new_n18270, new_n18271);
nor_5  g15923(n16502, new_n5516, new_n18272);
and_5  g15924(new_n18272, new_n18271, new_n18273);
nor_5  g15925(new_n18273, new_n18269, new_n18274_1);
not_10 g15926(new_n18274_1, new_n18275);
nand_5 g15927(new_n18275, new_n18268, new_n18276);
and_5  g15928(new_n18276, new_n18267, new_n18277);
nand_5 g15929(new_n18277, new_n18266, new_n18278);
and_5  g15930(new_n18278, new_n18265, new_n18279);
or_5   g15931(new_n18279, new_n18264, new_n18280);
and_5  g15932(new_n18280, new_n18262, new_n18281);
xor_4  g15933(new_n18281, new_n18261, new_n18282);
nor_5  g15934(n20077, n6794, new_n18283);
and_5  g15935(new_n18283, new_n6823, new_n18284);
and_5  g15936(new_n18284, new_n5561, new_n18285);
and_5  g15937(new_n18285, new_n5557, new_n18286);
xor_4  g15938(new_n18286, new_n5553, new_n18287);
xor_4  g15939(new_n18287, n11580, new_n18288_1);
xor_4  g15940(new_n18285, new_n5557, new_n18289);
or_5   g15941(new_n18289, new_n5624, new_n18290_1);
xor_4  g15942(new_n18289, n15884, new_n18291);
not_10 g15943(n6356, new_n18292);
xor_4  g15944(new_n18284, new_n5561, new_n18293);
or_5   g15945(new_n18293, new_n18292, new_n18294);
xor_4  g15946(new_n18293, n6356, new_n18295_1);
xor_4  g15947(new_n18283, new_n6823, new_n18296);
or_5   g15948(new_n18296, new_n9169, new_n18297);
xor_4  g15949(new_n18296, n27104, new_n18298);
xor_4  g15950(n20077, n6794, new_n18299);
or_5   g15951(new_n18299, new_n9175, new_n18300);
and_5  g15952(new_n5570, n6611, new_n18301_1);
xor_4  g15953(new_n18299, new_n9175, new_n18302);
nand_5 g15954(new_n18302, new_n18301_1, new_n18303);
and_5  g15955(new_n18303, new_n18300, new_n18304_1);
or_5   g15956(new_n18304_1, new_n18298, new_n18305);
and_5  g15957(new_n18305, new_n18297, new_n18306);
or_5   g15958(new_n18306, new_n18295_1, new_n18307);
and_5  g15959(new_n18307, new_n18294, new_n18308);
or_5   g15960(new_n18308, new_n18291, new_n18309);
and_5  g15961(new_n18309, new_n18290_1, new_n18310_1);
xor_4  g15962(new_n18310_1, new_n18288_1, new_n18311_1);
xnor_4 g15963(new_n18311_1, new_n16255, new_n18312);
xor_4  g15964(new_n18308, new_n18291, new_n18313);
or_5   g15965(new_n18313, new_n15624, new_n18314);
xor_4  g15966(new_n18306, new_n18295_1, new_n18315);
nand_5 g15967(new_n18315, new_n15629, new_n18316);
xnor_4 g15968(new_n18315, new_n15628, new_n18317);
xor_4  g15969(new_n18304_1, new_n18298, new_n18318);
or_5   g15970(new_n18318, new_n5058, new_n18319);
xor_4  g15971(new_n18318, new_n5058, new_n18320);
not_10 g15972(new_n18320, new_n18321);
xor_4  g15973(new_n18302, new_n18301_1, new_n18322);
or_5   g15974(new_n18322, new_n5067, new_n18323_1);
xor_4  g15975(n6794, n6611, new_n18324);
and_5  g15976(new_n18324, new_n5063, new_n18325);
xor_4  g15977(new_n18322, new_n5067, new_n18326);
nand_5 g15978(new_n18326, new_n18325, new_n18327);
and_5  g15979(new_n18327, new_n18323_1, new_n18328);
or_5   g15980(new_n18328, new_n18321, new_n18329);
and_5  g15981(new_n18329, new_n18319, new_n18330);
nand_5 g15982(new_n18330, new_n18317, new_n18331);
and_5  g15983(new_n18331, new_n18316, new_n18332_1);
xor_4  g15984(new_n18313, new_n15624, new_n18333);
nand_5 g15985(new_n18333, new_n18332_1, new_n18334);
and_5  g15986(new_n18334, new_n18314, new_n18335);
xor_4  g15987(new_n18335, new_n18312, new_n18336);
xor_4  g15988(new_n18336, new_n18282, new_n18337);
xor_4  g15989(new_n18279, new_n18264, new_n18338);
xor_4  g15990(new_n18333, new_n18332_1, new_n18339);
or_5   g15991(new_n18339, new_n18338, new_n18340);
xor_4  g15992(new_n18339, new_n18338, new_n18341);
not_10 g15993(new_n18341, new_n18342);
xor_4  g15994(new_n18330, new_n18317, new_n18343_1);
not_10 g15995(new_n18343_1, new_n18344);
xor_4  g15996(new_n18277, new_n18266, new_n18345_1);
or_5   g15997(new_n18345_1, new_n18344, new_n18346);
xor_4  g15998(new_n18345_1, new_n18344, new_n18347);
xor_4  g15999(new_n18328, new_n18321, new_n18348);
xnor_4 g16000(n15053, n12341, new_n18349);
xor_4  g16001(new_n18349, new_n18275, new_n18350_1);
not_10 g16002(new_n18350_1, new_n18351);
or_5   g16003(new_n18351, new_n18348, new_n18352);
xnor_4 g16004(new_n18350_1, new_n18348, new_n18353);
not_10 g16005(new_n18353, new_n18354);
xor_4  g16006(new_n18324, new_n5063, new_n18355);
not_10 g16007(new_n18355, new_n18356);
xnor_4 g16008(n16502, n12384, new_n18357);
nor_5  g16009(new_n18357, new_n18356, new_n18358);
xnor_4 g16010(n25471, n20986, new_n18359);
xnor_4 g16011(new_n18359, new_n18272, new_n18360);
or_5   g16012(new_n18360, new_n18358, new_n18361);
xor_4  g16013(new_n18326, new_n18325, new_n18362_1);
not_10 g16014(new_n18362_1, new_n18363);
xor_4  g16015(new_n18360, new_n18358, new_n18364);
nand_5 g16016(new_n18364, new_n18363, new_n18365);
and_5  g16017(new_n18365, new_n18361, new_n18366);
or_5   g16018(new_n18366, new_n18354, new_n18367);
nand_5 g16019(new_n18367, new_n18352, new_n18368);
nand_5 g16020(new_n18368, new_n18347, new_n18369);
and_5  g16021(new_n18369, new_n18346, new_n18370);
or_5   g16022(new_n18370, new_n18342, new_n18371);
and_5  g16023(new_n18371, new_n18340, new_n18372);
xor_4  g16024(new_n18372, new_n18337, n4785);
xnor_4 g16025(new_n14349, new_n14312, n4804);
xor_4  g16026(new_n15973, new_n15955, n4810);
and_5  g16027(n23166, new_n4449, new_n18376);
not_10 g16028(new_n18376, new_n18377_1);
nor_5  g16029(new_n9352, new_n9308_1, new_n18378);
not_10 g16030(new_n18378, new_n18379);
and_5  g16031(new_n18379, new_n18377_1, new_n18380);
and_5  g16032(new_n10966, new_n8092, new_n18381);
nor_5  g16033(new_n11014, new_n10967, new_n18382);
or_5   g16034(new_n18382, new_n18381, new_n18383);
and_5  g16035(new_n10964, new_n10958, new_n18384);
not_10 g16036(new_n18384, new_n18385);
and_5  g16037(new_n17902, new_n18385, new_n18386);
and_5  g16038(new_n18384, new_n17900, new_n18387);
nor_5  g16039(new_n18387, new_n18386, new_n18388);
xor_4  g16040(new_n18388, new_n8162, new_n18389);
xor_4  g16041(new_n18389, new_n18383, new_n18390);
and_5  g16042(new_n18390, new_n18380, new_n18391);
xnor_4 g16043(new_n18390, new_n18380, new_n18392);
and_5  g16044(new_n11015, new_n9353, new_n18393);
nor_5  g16045(new_n11070, new_n11017, new_n18394);
nor_5  g16046(new_n18394, new_n18393, new_n18395);
nor_5  g16047(new_n18395, new_n18392, new_n18396);
or_5   g16048(new_n18396, new_n18391, new_n18397);
nor_5  g16049(new_n18388, new_n8162, new_n18398);
or_5   g16050(new_n18398, new_n18383, new_n18399);
and_5  g16051(new_n18388, new_n8162, new_n18400);
nor_5  g16052(new_n18400, new_n18387, new_n18401);
and_5  g16053(new_n18401, new_n18399, new_n18402);
or_5   g16054(new_n18402, new_n18397, n4814);
xnor_4 g16055(new_n16582, new_n16580, n4850);
xor_4  g16056(new_n17429, new_n17392_1, n4891);
xnor_4 g16057(new_n17592_1, new_n17566, n4925);
xnor_4 g16058(new_n16589_1, new_n16569, n4947);
xor_4  g16059(new_n9617, new_n9615, n4952);
xor_4  g16060(n25068, n6790, new_n18409_1);
or_5   g16061(n22879, new_n8120, new_n18410);
xor_4  g16062(n22879, n2331, new_n18411);
or_5   g16063(new_n8125, n2117, new_n18412);
xnor_4 g16064(n22631, n2117, new_n18413);
or_5   g16065(n16743, new_n10045, new_n18414_1);
or_5   g16066(new_n8130_1, n5882, new_n18415);
and_5  g16067(new_n8135_1, n11775, new_n18416);
and_5  g16068(n27134, new_n8136, new_n18417);
and_5  g16069(n15258, new_n10048, new_n18418_1);
not_10 g16070(new_n18418_1, new_n18419);
and_5  g16071(new_n18419, new_n18417, new_n18420);
nor_5  g16072(new_n18420, new_n18416, new_n18421);
not_10 g16073(new_n18421, new_n18422);
nand_5 g16074(new_n18422, new_n18415, new_n18423);
and_5  g16075(new_n18423, new_n18414_1, new_n18424);
nand_5 g16076(new_n18424, new_n18413, new_n18425);
and_5  g16077(new_n18425, new_n18412, new_n18426);
or_5   g16078(new_n18426, new_n18411, new_n18427);
and_5  g16079(new_n18427, new_n18410, new_n18428);
xor_4  g16080(new_n18428, new_n18409_1, new_n18429);
xor_4  g16081(new_n18429, new_n15833, new_n18430);
xor_4  g16082(new_n18426, new_n18411, new_n18431);
or_5   g16083(new_n18431, new_n15579, new_n18432);
xor_4  g16084(new_n18431, new_n15579, new_n18433);
not_10 g16085(new_n18433, new_n18434);
xor_4  g16086(new_n18424, new_n18413, new_n18435);
or_5   g16087(new_n18435, new_n15585, new_n18436);
xnor_4 g16088(new_n18435, new_n15584, new_n18437_1);
xnor_4 g16089(n16743, n5882, new_n18438);
xor_4  g16090(new_n18438, new_n18422, new_n18439_1);
or_5   g16091(new_n18439_1, new_n15591, new_n18440);
xor_4  g16092(new_n18439_1, new_n15591, new_n18441);
not_10 g16093(new_n18441, new_n18442);
xnor_4 g16094(n15258, n11775, new_n18443);
xor_4  g16095(new_n18443, new_n18417, new_n18444_1);
or_5   g16096(new_n18444_1, new_n15593, new_n18445_1);
and_5  g16097(new_n15363, new_n15362, new_n18446);
xor_4  g16098(new_n18444_1, new_n15593, new_n18447);
nand_5 g16099(new_n18447, new_n18446, new_n18448);
and_5  g16100(new_n18448, new_n18445_1, new_n18449);
or_5   g16101(new_n18449, new_n18442, new_n18450);
and_5  g16102(new_n18450, new_n18440, new_n18451);
nand_5 g16103(new_n18451, new_n18437_1, new_n18452_1);
and_5  g16104(new_n18452_1, new_n18436, new_n18453);
or_5   g16105(new_n18453, new_n18434, new_n18454);
and_5  g16106(new_n18454, new_n18432, new_n18455);
xor_4  g16107(new_n18455, new_n18430, new_n18456);
xor_4  g16108(new_n18456, new_n15505, new_n18457);
not_10 g16109(new_n18457, new_n18458);
xnor_4 g16110(new_n18453, new_n18433, new_n18459);
not_10 g16111(new_n18459, new_n18460);
nor_5  g16112(new_n18460, new_n15509, new_n18461);
xor_4  g16113(new_n18460, new_n15509, new_n18462);
xor_4  g16114(new_n18451, new_n18437_1, new_n18463);
not_10 g16115(new_n18463, new_n18464);
nor_5  g16116(new_n18464, new_n13868, new_n18465);
xor_4  g16117(new_n18464, new_n13868, new_n18466);
xor_4  g16118(new_n18449, new_n18442, new_n18467_1);
nor_5  g16119(new_n18467_1, new_n13873, new_n18468);
xor_4  g16120(new_n18467_1, new_n13873, new_n18469);
not_10 g16121(new_n18469, new_n18470);
nor_5  g16122(new_n15365, new_n10144, new_n18471);
nor_5  g16123(new_n18471, new_n13885, new_n18472);
xor_4  g16124(new_n18471, new_n13885, new_n18473);
xor_4  g16125(new_n18447, new_n18446, new_n18474);
not_10 g16126(new_n18474, new_n18475);
and_5  g16127(new_n18475, new_n18473, new_n18476);
nor_5  g16128(new_n18476, new_n18472, new_n18477);
nor_5  g16129(new_n18477, new_n18470, new_n18478);
nor_5  g16130(new_n18478, new_n18468, new_n18479);
not_10 g16131(new_n18479, new_n18480);
and_5  g16132(new_n18480, new_n18466, new_n18481);
nor_5  g16133(new_n18481, new_n18465, new_n18482_1);
not_10 g16134(new_n18482_1, new_n18483_1);
and_5  g16135(new_n18483_1, new_n18462, new_n18484);
nor_5  g16136(new_n18484, new_n18461, new_n18485);
xnor_4 g16137(new_n18485, new_n18458, n4966);
xnor_4 g16138(new_n17921, new_n17920, n4972);
not_10 g16139(new_n7609, new_n18488);
or_5   g16140(new_n7615, n23895, new_n18489);
xor_4  g16141(new_n7615, new_n10538, new_n18490);
not_10 g16142(new_n18490, new_n18491);
nand_5 g16143(new_n7621, n17351, new_n18492);
xor_4  g16144(new_n7621, new_n5484, new_n18493);
or_5   g16145(new_n7626, new_n5488, new_n18494);
or_5   g16146(new_n17254, new_n17243_1, new_n18495);
and_5  g16147(new_n18495, new_n18494, new_n18496_1);
or_5   g16148(new_n18496_1, new_n18493, new_n18497);
and_5  g16149(new_n18497, new_n18492, new_n18498);
nand_5 g16150(new_n18498, new_n18491, new_n18499);
and_5  g16151(new_n18499, new_n18489, new_n18500);
and_5  g16152(new_n18500, new_n18488, new_n18501);
not_10 g16153(new_n18501, new_n18502);
not_10 g16154(n2978, new_n18503);
and_5  g16155(new_n17209, new_n7515, new_n18504);
and_5  g16156(new_n18504, new_n7511, new_n18505);
xor_4  g16157(new_n18505, new_n18503, new_n18506);
xor_4  g16158(new_n18506, new_n13318, new_n18507);
xor_4  g16159(new_n18504, new_n7511, new_n18508);
and_5  g16160(new_n18508, n337, new_n18509_1);
nor_5  g16161(new_n18508, n337, new_n18510);
and_5  g16162(new_n17210, n3228, new_n18511);
nor_5  g16163(new_n17210, n3228, new_n18512);
not_10 g16164(new_n17222, new_n18513_1);
nor_5  g16165(new_n18513_1, new_n18512, new_n18514);
nor_5  g16166(new_n18514, new_n18511, new_n18515_1);
nor_5  g16167(new_n18515_1, new_n18510, new_n18516);
nor_5  g16168(new_n18516, new_n18509_1, new_n18517);
xor_4  g16169(new_n18517, new_n18507, new_n18518);
or_5   g16170(new_n18518, n25972, new_n18519);
not_10 g16171(n25972, new_n18520);
xor_4  g16172(new_n18518, new_n18520, new_n18521);
xor_4  g16173(new_n18508, new_n5242, new_n18522);
xor_4  g16174(new_n18522, new_n18515_1, new_n18523);
or_5   g16175(new_n18523, n21915, new_n18524);
or_5   g16176(new_n17224, n13775, new_n18525);
or_5   g16177(new_n17240, new_n17226, new_n18526);
and_5  g16178(new_n18526, new_n18525, new_n18527);
xor_4  g16179(new_n18523, n21915, new_n18528);
not_10 g16180(new_n18528, new_n18529);
or_5   g16181(new_n18529, new_n18527, new_n18530);
and_5  g16182(new_n18530, new_n18524, new_n18531);
or_5   g16183(new_n18531, new_n18521, new_n18532);
and_5  g16184(new_n18532, new_n18519, new_n18533);
and_5  g16185(new_n18505, new_n18503, new_n18534);
not_10 g16186(new_n18534, new_n18535);
and_5  g16187(new_n18506, n7593, new_n18536);
nor_5  g16188(new_n18506, n7593, new_n18537_1);
nor_5  g16189(new_n18517, new_n18537_1, new_n18538);
nor_5  g16190(new_n18538, new_n18536, new_n18539);
and_5  g16191(new_n18539, new_n18535, new_n18540);
and_5  g16192(new_n18540, new_n18533, new_n18541);
xnor_4 g16193(new_n18500, new_n7609, new_n18542);
xor_4  g16194(new_n18540, new_n18533, new_n18543);
or_5   g16195(new_n18543, new_n18542, new_n18544);
not_10 g16196(new_n18542, new_n18545);
xor_4  g16197(new_n18543, new_n18545, new_n18546);
xor_4  g16198(new_n18498, new_n18490, new_n18547);
not_10 g16199(new_n18547, new_n18548);
xor_4  g16200(new_n18531, new_n18521, new_n18549);
nor_5  g16201(new_n18549, new_n18548, new_n18550);
xor_4  g16202(new_n18549, new_n18547, new_n18551);
xor_4  g16203(new_n18496_1, new_n18493, new_n18552);
not_10 g16204(new_n18552, new_n18553);
xnor_4 g16205(new_n18528, new_n18527, new_n18554);
or_5   g16206(new_n18554, new_n18553, new_n18555);
or_5   g16207(new_n17255, new_n17242, new_n18556);
not_10 g16208(new_n17256, new_n18557);
or_5   g16209(new_n17276, new_n18557, new_n18558_1);
and_5  g16210(new_n18558_1, new_n18556, new_n18559);
xnor_4 g16211(new_n18554, new_n18552, new_n18560);
nand_5 g16212(new_n18560, new_n18559, new_n18561);
and_5  g16213(new_n18561, new_n18555, new_n18562);
nor_5  g16214(new_n18562, new_n18551, new_n18563);
or_5   g16215(new_n18563, new_n18550, new_n18564);
or_5   g16216(new_n18564, new_n18546, new_n18565);
and_5  g16217(new_n18565, new_n18544, new_n18566);
xor_4  g16218(new_n18566, new_n18541, new_n18567);
xor_4  g16219(new_n18567, new_n18502, n5011);
and_5  g16220(n11220, new_n11219, new_n18569);
xnor_4 g16221(n11220, n2944, new_n18570);
not_10 g16222(new_n18570, new_n18571);
not_10 g16223(n22379, new_n18572_1);
or_5   g16224(new_n18572_1, n767, new_n18573);
or_5   g16225(new_n2881, new_n2836, new_n18574_1);
and_5  g16226(new_n18574_1, new_n18573, new_n18575);
nor_5  g16227(new_n18575, new_n18571, new_n18576_1);
nor_5  g16228(new_n18576_1, new_n18569, new_n18577);
not_10 g16229(new_n18577, new_n18578_1);
and_5  g16230(n16544, n2160, new_n18579);
nor_5  g16231(n16544, n2160, new_n18580);
nor_5  g16232(n10763, n6814, new_n18581);
nor_5  g16233(new_n2912, new_n2883, new_n18582_1);
nor_5  g16234(new_n18582_1, new_n18581, new_n18583_1);
not_10 g16235(new_n18583_1, new_n18584_1);
nor_5  g16236(new_n18584_1, new_n18580, new_n18585);
nor_5  g16237(new_n18585, new_n18579, new_n18586);
nor_5  g16238(new_n18586, new_n15427, new_n18587);
not_10 g16239(new_n18587, new_n18588);
xor_4  g16240(new_n18586, new_n15427, new_n18589);
not_10 g16241(new_n18589, new_n18590);
xnor_4 g16242(n16544, n2160, new_n18591);
xor_4  g16243(new_n18591, new_n18584_1, new_n18592);
nand_5 g16244(new_n18592, new_n15402, new_n18593);
xnor_4 g16245(new_n18592, new_n15402, new_n18594);
or_5   g16246(new_n15418, new_n2913, new_n18595);
or_5   g16247(new_n3008, new_n2952, new_n18596);
and_5  g16248(new_n18596, new_n18595, new_n18597);
or_5   g16249(new_n18597, new_n18594, new_n18598);
and_5  g16250(new_n18598, new_n18593, new_n18599);
nor_5  g16251(new_n18599, new_n18590, new_n18600);
not_10 g16252(new_n18600, new_n18601);
and_5  g16253(new_n18601, new_n18588, new_n18602);
or_5   g16254(new_n18602, new_n18578_1, new_n18603);
xor_4  g16255(new_n18599, new_n18590, new_n18604);
not_10 g16256(new_n18604, new_n18605);
and_5  g16257(new_n18605, new_n18578_1, new_n18606);
nor_5  g16258(new_n18605, new_n18578_1, new_n18607);
xor_4  g16259(new_n18575, new_n18571, new_n18608);
xor_4  g16260(new_n18597, new_n18594, new_n18609);
nor_5  g16261(new_n18609, new_n18608, new_n18610_1);
xor_4  g16262(new_n18609, new_n18608, new_n18611);
not_10 g16263(new_n18611, new_n18612);
nor_5  g16264(new_n3009, new_n2882, new_n18613);
nor_5  g16265(new_n3073, new_n3011, new_n18614);
nor_5  g16266(new_n18614, new_n18613, new_n18615);
nor_5  g16267(new_n18615, new_n18612, new_n18616);
nor_5  g16268(new_n18616, new_n18610_1, new_n18617);
nor_5  g16269(new_n18617, new_n18607, new_n18618);
nor_5  g16270(new_n18618, new_n18606, new_n18619);
not_10 g16271(new_n18619, new_n18620);
nand_5 g16272(new_n18620, new_n18603, new_n18621);
and_5  g16273(new_n18602, new_n18578_1, new_n18622);
or_5   g16274(new_n18622, new_n18618, new_n18623);
and_5  g16275(new_n18623, new_n18621, n5020);
not_10 g16276(n3480, new_n18625);
nor_5  g16277(n13781, n11486, new_n18626);
and_5  g16278(new_n18626, new_n7750, new_n18627);
and_5  g16279(new_n18627, new_n18625, new_n18628);
xor_4  g16280(new_n18628, new_n10855, new_n18629);
xnor_4 g16281(new_n18629, new_n2972, new_n18630);
xor_4  g16282(new_n18627, new_n18625, new_n18631);
or_5   g16283(new_n18631, new_n2977, new_n18632);
xor_4  g16284(new_n18631, new_n2978_1, new_n18633);
xor_4  g16285(new_n18626, new_n7750, new_n18634);
or_5   g16286(new_n18634, new_n2982, new_n18635_1);
xor_4  g16287(new_n18634, new_n2983, new_n18636);
xor_4  g16288(n13781, n11486, new_n18637);
or_5   g16289(new_n18637, new_n2989, new_n18638);
and_5  g16290(new_n3047, new_n7757, new_n18639);
xor_4  g16291(new_n18637, new_n2989, new_n18640);
nand_5 g16292(new_n18640, new_n18639, new_n18641);
and_5  g16293(new_n18641, new_n18638, new_n18642);
or_5   g16294(new_n18642, new_n18636, new_n18643);
and_5  g16295(new_n18643, new_n18635_1, new_n18644);
or_5   g16296(new_n18644, new_n18633, new_n18645);
and_5  g16297(new_n18645, new_n18632, new_n18646);
xnor_4 g16298(new_n18646, new_n18630, new_n18647);
xor_4  g16299(new_n18647, new_n6944, new_n18648);
not_10 g16300(new_n18648, new_n18649_1);
xor_4  g16301(new_n18644, new_n18633, new_n18650);
and_5  g16302(new_n18650, new_n6949, new_n18651);
xor_4  g16303(new_n18650, new_n6949, new_n18652);
not_10 g16304(new_n18652, new_n18653_1);
xor_4  g16305(new_n18642, new_n18636, new_n18654);
and_5  g16306(new_n18654, new_n6959, new_n18655);
xor_4  g16307(new_n18640, new_n18639, new_n18656);
and_5  g16308(new_n18656, new_n6963, new_n18657);
xor_4  g16309(new_n3047, new_n7757, new_n18658);
nor_5  g16310(new_n18658, new_n6967_1, new_n18659);
xor_4  g16311(new_n18656, new_n6963, new_n18660);
not_10 g16312(new_n18660, new_n18661);
nor_5  g16313(new_n18661, new_n18659, new_n18662);
nor_5  g16314(new_n18662, new_n18657, new_n18663);
xnor_4 g16315(new_n18654, new_n6956, new_n18664);
not_10 g16316(new_n18664, new_n18665);
nor_5  g16317(new_n18665, new_n18663, new_n18666);
nor_5  g16318(new_n18666, new_n18655, new_n18667);
nor_5  g16319(new_n18667, new_n18653_1, new_n18668);
nor_5  g16320(new_n18668, new_n18651, new_n18669);
xnor_4 g16321(new_n18669, new_n18649_1, n5024);
xnor_4 g16322(new_n3714, new_n3681, n5046);
xor_4  g16323(new_n5903_1, new_n5902, n5062);
xnor_4 g16324(new_n12820, new_n12787, n5064);
xnor_4 g16325(n12495, n11479, new_n18674);
xor_4  g16326(new_n18674, new_n2384, new_n18675);
xnor_4 g16327(n9251, n7428, new_n18676);
or_5   g16328(new_n18676, new_n18675, new_n18677);
and_5  g16329(n9251, new_n8437, new_n18678);
xnor_4 g16330(n20138, n10372, new_n18679_1);
xor_4  g16331(new_n18679_1, new_n18678, new_n18680);
xor_4  g16332(new_n18680, new_n18677, new_n18681);
nand_5 g16333(new_n18674, new_n2384, new_n18682);
nand_5 g16334(n12495, n11479, new_n18683);
xor_4  g16335(n20235, n8259, new_n18684);
xor_4  g16336(new_n18684, new_n18683, new_n18685);
xor_4  g16337(new_n18685, new_n2388_1, new_n18686);
xor_4  g16338(new_n18686, new_n18682, new_n18687);
xor_4  g16339(new_n18687, new_n18681, n5082);
xor_4  g16340(new_n14011, new_n14010, n5120);
xor_4  g16341(new_n15223, new_n15209, n5158);
xnor_4 g16342(new_n16586, new_n16573, n5168);
not_10 g16343(new_n17654, new_n18692);
xor_4  g16344(new_n18692, n6659, new_n18693_1);
nand_5 g16345(new_n14628, new_n16340, new_n18694);
xor_4  g16346(new_n14628, n23250, new_n18695);
nand_5 g16347(new_n14630, new_n16272, new_n18696);
xor_4  g16348(new_n14630, n11455, new_n18697);
nand_5 g16349(new_n14632, new_n16275_1, new_n18698);
xor_4  g16350(new_n14632, new_n16275_1, new_n18699);
nor_5  g16351(new_n14635, new_n16278, new_n18700);
xor_4  g16352(new_n14635, n5255, new_n18701);
nand_5 g16353(new_n14638, n21649, new_n18702);
nand_5 g16354(new_n15653, new_n15640, new_n18703);
and_5  g16355(new_n18703, new_n18702, new_n18704);
nor_5  g16356(new_n18704, new_n18701, new_n18705);
nor_5  g16357(new_n18705, new_n18700, new_n18706);
nand_5 g16358(new_n18706, new_n18699, new_n18707);
and_5  g16359(new_n18707, new_n18698, new_n18708_1);
or_5   g16360(new_n18708_1, new_n18697, new_n18709);
and_5  g16361(new_n18709, new_n18696, new_n18710);
or_5   g16362(new_n18710, new_n18695, new_n18711);
and_5  g16363(new_n18711, new_n18694, new_n18712);
xor_4  g16364(new_n18712, new_n18693_1, new_n18713);
xnor_4 g16365(new_n18713, new_n16270, new_n18714);
not_10 g16366(new_n18714, new_n18715);
xor_4  g16367(new_n18710, new_n18695, new_n18716);
nand_5 g16368(new_n18716, new_n16348, new_n18717);
xnor_4 g16369(new_n18716, new_n16351, new_n18718);
not_10 g16370(new_n18718, new_n18719);
xor_4  g16371(new_n18708_1, new_n18697, new_n18720);
nand_5 g16372(new_n18720, new_n16354, new_n18721_1);
xnor_4 g16373(new_n18720, new_n16357, new_n18722);
not_10 g16374(new_n18722, new_n18723);
xor_4  g16375(new_n18706, new_n18699, new_n18724);
nand_5 g16376(new_n18724, new_n16360, new_n18725_1);
xnor_4 g16377(new_n18724, new_n16361, new_n18726);
not_10 g16378(new_n18726, new_n18727);
xor_4  g16379(new_n18704, new_n18701, new_n18728);
or_5   g16380(new_n18728, new_n16368, new_n18729);
xor_4  g16381(new_n18728, new_n16368, new_n18730);
not_10 g16382(new_n18730, new_n18731);
or_5   g16383(new_n15654, new_n15639, new_n18732);
or_5   g16384(new_n15678, new_n15656, new_n18733);
and_5  g16385(new_n18733, new_n18732, new_n18734);
or_5   g16386(new_n18734, new_n18731, new_n18735);
and_5  g16387(new_n18735, new_n18729, new_n18736);
or_5   g16388(new_n18736, new_n18727, new_n18737_1);
and_5  g16389(new_n18737_1, new_n18725_1, new_n18738);
or_5   g16390(new_n18738, new_n18723, new_n18739);
and_5  g16391(new_n18739, new_n18721_1, new_n18740);
or_5   g16392(new_n18740, new_n18719, new_n18741);
and_5  g16393(new_n18741, new_n18717, new_n18742);
xnor_4 g16394(new_n18742, new_n18715, n5184);
not_10 g16395(new_n4409_1, new_n18744);
nand_5 g16396(new_n4525, new_n18744, new_n18745_1);
nor_5  g16397(new_n4610, new_n18745_1, new_n18746);
nor_5  g16398(new_n4525, new_n18744, new_n18747);
and_5  g16399(new_n4610, new_n18747, new_n18748);
or_5   g16400(new_n18748, new_n18746, n5228);
and_5  g16401(new_n3408, n1314, new_n18750);
nor_5  g16402(new_n11500, new_n11483, new_n18751_1);
nor_5  g16403(new_n18751_1, new_n18750, new_n18752);
xor_4  g16404(new_n18752, new_n7241, new_n18753);
not_10 g16405(new_n18753, new_n18754);
and_5  g16406(new_n11502, new_n7148, new_n18755);
xnor_4 g16407(new_n11501, new_n7148, new_n18756);
not_10 g16408(new_n18756, new_n18757);
and_5  g16409(new_n11524, new_n7154, new_n18758);
nor_5  g16410(new_n12822, new_n12783_1, new_n18759);
nor_5  g16411(new_n18759, new_n18758, new_n18760);
nor_5  g16412(new_n18760, new_n18757, new_n18761);
nor_5  g16413(new_n18761, new_n18755, new_n18762);
xnor_4 g16414(new_n18762, new_n18754, n5256);
xor_4  g16415(new_n6706_1, new_n6695, n5265);
xor_4  g16416(new_n17432_1, new_n17388, n5273);
xor_4  g16417(n20946, n2289, new_n18766);
or_5   g16418(new_n3186, n1112, new_n18767);
xor_4  g16419(n7751, n1112, new_n18768);
or_5   g16420(new_n3187, n20179, new_n18769);
or_5   g16421(new_n17082, new_n17067, new_n18770);
and_5  g16422(new_n18770, new_n18769, new_n18771);
or_5   g16423(new_n18771, new_n18768, new_n18772);
and_5  g16424(new_n18772, new_n18767, new_n18773);
xor_4  g16425(new_n18773, new_n18766, new_n18774);
xor_4  g16426(new_n18774, new_n7432_1, new_n18775);
xor_4  g16427(new_n18771, new_n18768, new_n18776);
nor_5  g16428(new_n18776, new_n7438, new_n18777);
not_10 g16429(new_n18777, new_n18778);
xor_4  g16430(new_n18776, new_n7438, new_n18779);
nor_5  g16431(new_n17083, new_n7444, new_n18780_1);
not_10 g16432(new_n18780_1, new_n18781);
not_10 g16433(new_n17109, new_n18782_1);
and_5  g16434(new_n18782_1, new_n17084_1, new_n18783);
not_10 g16435(new_n18783, new_n18784);
and_5  g16436(new_n18784, new_n18781, new_n18785);
not_10 g16437(new_n18785, new_n18786);
and_5  g16438(new_n18786, new_n18779, new_n18787);
not_10 g16439(new_n18787, new_n18788);
and_5  g16440(new_n18788, new_n18778, new_n18789);
xor_4  g16441(new_n18789, new_n18775, n5274);
not_10 g16442(n6513, new_n18791);
not_10 g16443(n3918, new_n18792);
nor_5  g16444(n25316, n20385, new_n18793);
and_5  g16445(new_n18793, new_n12570, new_n18794);
and_5  g16446(new_n18794, new_n18792, new_n18795);
xor_4  g16447(new_n18795, new_n18791, new_n18796);
xnor_4 g16448(new_n18796, new_n8978, new_n18797);
xor_4  g16449(new_n18794, new_n18792, new_n18798);
or_5   g16450(new_n18798, new_n8983, new_n18799);
xor_4  g16451(new_n18793, n919, new_n18800);
and_5  g16452(new_n18800, new_n8990, new_n18801);
not_10 g16453(new_n18801, new_n18802_1);
xor_4  g16454(new_n18800, new_n8990, new_n18803);
xor_4  g16455(n25316, n20385, new_n18804);
nand_5 g16456(new_n18804, new_n11366, new_n18805);
and_5  g16457(new_n8999, n20385, new_n18806);
xnor_4 g16458(new_n18804, new_n8996, new_n18807);
nand_5 g16459(new_n18807, new_n18806, new_n18808);
and_5  g16460(new_n18808, new_n18805, new_n18809);
and_5  g16461(new_n18809, new_n18803, new_n18810);
not_10 g16462(new_n18810, new_n18811);
and_5  g16463(new_n18811, new_n18802_1, new_n18812);
xor_4  g16464(new_n18798, new_n8984, new_n18813);
or_5   g16465(new_n18813, new_n18812, new_n18814);
and_5  g16466(new_n18814, new_n18799, new_n18815);
xnor_4 g16467(new_n18815, new_n18797, new_n18816);
not_10 g16468(new_n18816, new_n18817);
xor_4  g16469(new_n16848, n19472, new_n18818);
or_5   g16470(new_n16851, new_n8818, new_n18819);
xor_4  g16471(new_n16851, new_n8818, new_n18820);
not_10 g16472(new_n18820, new_n18821);
nand_5 g16473(new_n4129, n24786, new_n18822);
xor_4  g16474(new_n4129, n24786, new_n18823);
not_10 g16475(new_n18823, new_n18824);
nand_5 g16476(new_n4133, n27120, new_n18825);
or_5   g16477(new_n4137, n23065, new_n18826);
xor_4  g16478(new_n4133, n27120, new_n18827);
nand_5 g16479(new_n18827, new_n18826, new_n18828);
and_5  g16480(new_n18828, new_n18825, new_n18829);
or_5   g16481(new_n18829, new_n18824, new_n18830_1);
and_5  g16482(new_n18830_1, new_n18822, new_n18831_1);
or_5   g16483(new_n18831_1, new_n18821, new_n18832);
and_5  g16484(new_n18832, new_n18819, new_n18833);
xor_4  g16485(new_n18833, new_n18818, new_n18834);
xor_4  g16486(new_n18834, new_n18817, new_n18835);
not_10 g16487(new_n18835, new_n18836);
xor_4  g16488(new_n18831_1, new_n18821, new_n18837);
xnor_4 g16489(new_n18798, new_n8984, new_n18838);
xnor_4 g16490(new_n18838, new_n18812, new_n18839);
not_10 g16491(new_n18839, new_n18840);
nor_5  g16492(new_n18840, new_n18837, new_n18841);
xor_4  g16493(new_n18840, new_n18837, new_n18842);
not_10 g16494(new_n18842, new_n18843_1);
xor_4  g16495(new_n18829, new_n18824, new_n18844);
xor_4  g16496(new_n18809, new_n18803, new_n18845);
not_10 g16497(new_n18845, new_n18846);
nor_5  g16498(new_n18846, new_n18844, new_n18847);
xor_4  g16499(new_n18846, new_n18844, new_n18848);
not_10 g16500(new_n18848, new_n18849);
xor_4  g16501(new_n18807, new_n18806, new_n18850);
xor_4  g16502(new_n18827, new_n18826, new_n18851);
nor_5  g16503(new_n18851, new_n18850, new_n18852);
xor_4  g16504(new_n4137, n23065, new_n18853);
nor_5  g16505(new_n18853, new_n9089, new_n18854);
xor_4  g16506(new_n18851, new_n18850, new_n18855);
not_10 g16507(new_n18855, new_n18856);
nor_5  g16508(new_n18856, new_n18854, new_n18857);
nor_5  g16509(new_n18857, new_n18852, new_n18858_1);
nor_5  g16510(new_n18858_1, new_n18849, new_n18859_1);
nor_5  g16511(new_n18859_1, new_n18847, new_n18860);
nor_5  g16512(new_n18860, new_n18843_1, new_n18861);
nor_5  g16513(new_n18861, new_n18841, new_n18862);
xnor_4 g16514(new_n18862, new_n18836, n5300);
nor_5  g16515(new_n7236_1, new_n7232, new_n18864_1);
not_10 g16516(new_n18864_1, new_n18865_1);
and_5  g16517(new_n7240, new_n7237, new_n18866);
not_10 g16518(new_n18866, new_n18867);
and_5  g16519(new_n18867, new_n18865_1, new_n18868);
or_5   g16520(new_n18868, new_n18752, new_n18869);
xor_4  g16521(new_n18868, new_n18752, new_n18870);
nor_5  g16522(new_n18752, new_n7241, new_n18871);
nor_5  g16523(new_n18762, new_n18754, new_n18872);
nor_5  g16524(new_n18872, new_n18871, new_n18873);
nand_5 g16525(new_n18873, new_n18870, new_n18874);
and_5  g16526(new_n18874, new_n18869, n5325);
not_10 g16527(n23272, new_n18876);
xnor_4 g16528(n25120, n17458, new_n18877);
or_5   g16529(n8363, n1222, new_n18878);
xnor_4 g16530(n8363, n1222, new_n18879);
or_5   g16531(n25240, n14680, new_n18880_1);
xnor_4 g16532(n25240, n14680, new_n18881);
or_5   g16533(n17250, n10125, new_n18882);
xor_4  g16534(n17250, n10125, new_n18883);
nand_5 g16535(n23160, n8067, new_n18884);
or_5   g16536(n23160, n8067, new_n18885);
nor_5  g16537(n20923, n16524, new_n18886_1);
nor_5  g16538(new_n13251, new_n13248, new_n18887_1);
nor_5  g16539(new_n18887_1, new_n18886_1, new_n18888);
nand_5 g16540(new_n18888, new_n18885, new_n18889);
and_5  g16541(new_n18889, new_n18884, new_n18890);
nand_5 g16542(new_n18890, new_n18883, new_n18891);
and_5  g16543(new_n18891, new_n18882, new_n18892);
or_5   g16544(new_n18892, new_n18881, new_n18893);
and_5  g16545(new_n18893, new_n18880_1, new_n18894);
or_5   g16546(new_n18894, new_n18879, new_n18895);
and_5  g16547(new_n18895, new_n18878, new_n18896);
xor_4  g16548(new_n18896, new_n18877, new_n18897);
and_5  g16549(new_n18897, new_n18876, new_n18898);
xor_4  g16550(new_n18897, new_n18876, new_n18899);
not_10 g16551(new_n18899, new_n18900);
not_10 g16552(n11481, new_n18901_1);
xor_4  g16553(new_n18894, new_n18879, new_n18902);
nand_5 g16554(new_n18902, new_n18901_1, new_n18903);
xor_4  g16555(new_n18902, new_n18901_1, new_n18904);
not_10 g16556(new_n18904, new_n18905);
xor_4  g16557(new_n18892, new_n18881, new_n18906);
nand_5 g16558(new_n18906, new_n4360, new_n18907_1);
xor_4  g16559(new_n18906, new_n4360, new_n18908);
not_10 g16560(new_n18908, new_n18909);
xor_4  g16561(new_n18890, new_n18883, new_n18910);
nand_5 g16562(new_n18910, new_n4364, new_n18911);
xor_4  g16563(new_n18910, new_n4364, new_n18912);
not_10 g16564(new_n18912, new_n18913);
xor_4  g16565(n23160, n8067, new_n18914);
xor_4  g16566(new_n18914, new_n18888, new_n18915);
or_5   g16567(new_n18915, n7678, new_n18916);
xor_4  g16568(new_n18915, new_n4368, new_n18917);
nand_5 g16569(new_n13252, new_n10813, new_n18918);
or_5   g16570(new_n13257, new_n13254, new_n18919_1);
and_5  g16571(new_n18919_1, new_n18918, new_n18920);
or_5   g16572(new_n18920, new_n18917, new_n18921);
and_5  g16573(new_n18921, new_n18916, new_n18922);
or_5   g16574(new_n18922, new_n18913, new_n18923);
and_5  g16575(new_n18923, new_n18911, new_n18924);
or_5   g16576(new_n18924, new_n18909, new_n18925);
and_5  g16577(new_n18925, new_n18907_1, new_n18926_1);
or_5   g16578(new_n18926_1, new_n18905, new_n18927);
and_5  g16579(new_n18927, new_n18903, new_n18928);
nor_5  g16580(new_n18928, new_n18900, new_n18929);
nor_5  g16581(new_n18929, new_n18898, new_n18930);
or_5   g16582(n25120, n17458, new_n18931);
or_5   g16583(new_n18896, new_n18877, new_n18932);
and_5  g16584(new_n18932, new_n18931, new_n18933);
and_5  g16585(new_n18933, new_n18930, new_n18934);
not_10 g16586(new_n18934, new_n18935);
xnor_4 g16587(n12702, n12507, new_n18936);
or_5   g16588(n26797, n15077, new_n18937);
xnor_4 g16589(n26797, n15077, new_n18938);
or_5   g16590(n23913, n3710, new_n18939);
xnor_4 g16591(n23913, n3710, new_n18940_1);
or_5   g16592(n26318, n22554, new_n18941);
xnor_4 g16593(n26318, n22554, new_n18942);
or_5   g16594(n26054, n20429, new_n18943);
xnor_4 g16595(n26054, n20429, new_n18944);
or_5   g16596(n19081, n3909, new_n18945_1);
xnor_4 g16597(n19081, n3909, new_n18946);
or_5   g16598(n23974, n8309, new_n18947);
xor_4  g16599(n23974, n8309, new_n18948);
nand_5 g16600(n19144, n2146, new_n18949);
or_5   g16601(n19144, n2146, new_n18950);
nor_5  g16602(n22173, n12593, new_n18951);
and_5  g16603(new_n17061, new_n17060, new_n18952);
nor_5  g16604(new_n18952, new_n18951, new_n18953);
nand_5 g16605(new_n18953, new_n18950, new_n18954);
and_5  g16606(new_n18954, new_n18949, new_n18955);
nand_5 g16607(new_n18955, new_n18948, new_n18956);
and_5  g16608(new_n18956, new_n18947, new_n18957);
or_5   g16609(new_n18957, new_n18946, new_n18958);
and_5  g16610(new_n18958, new_n18945_1, new_n18959);
or_5   g16611(new_n18959, new_n18944, new_n18960);
and_5  g16612(new_n18960, new_n18943, new_n18961);
or_5   g16613(new_n18961, new_n18942, new_n18962_1);
and_5  g16614(new_n18962_1, new_n18941, new_n18963);
or_5   g16615(new_n18963, new_n18940_1, new_n18964);
and_5  g16616(new_n18964, new_n18939, new_n18965);
or_5   g16617(new_n18965, new_n18938, new_n18966);
and_5  g16618(new_n18966, new_n18937, new_n18967);
xor_4  g16619(new_n18967, new_n18936, new_n18968);
nand_5 g16620(new_n18968, new_n9141, new_n18969);
xor_4  g16621(new_n18968, n12650, new_n18970_1);
xor_4  g16622(new_n18965, new_n18938, new_n18971);
nand_5 g16623(new_n18971, new_n5608, new_n18972);
xor_4  g16624(new_n18971, n10201, new_n18973);
xor_4  g16625(new_n18963, new_n18940_1, new_n18974);
nand_5 g16626(new_n18974, new_n5612, new_n18975);
xor_4  g16627(new_n18974, n10593, new_n18976);
xor_4  g16628(new_n18961, new_n18942, new_n18977_1);
nand_5 g16629(new_n18977_1, new_n5616, new_n18978);
xor_4  g16630(new_n18959, new_n18944, new_n18979);
and_5  g16631(new_n18979, new_n5620, new_n18980);
xor_4  g16632(new_n18979, new_n5620, new_n18981);
not_10 g16633(new_n18981, new_n18982_1);
xor_4  g16634(new_n18957, new_n18946, new_n18983);
nand_5 g16635(new_n18983, new_n5624, new_n18984);
xor_4  g16636(new_n18983, n15884, new_n18985);
xor_4  g16637(new_n18955, new_n18948, new_n18986);
nand_5 g16638(new_n18986, new_n18292, new_n18987);
xor_4  g16639(n19144, n2146, new_n18988);
xor_4  g16640(new_n18988, new_n18953, new_n18989);
nand_5 g16641(new_n18989, n27104, new_n18990);
xor_4  g16642(new_n18989, n27104, new_n18991);
nand_5 g16643(new_n17062, new_n9175, new_n18992);
nand_5 g16644(new_n17063, new_n17059, new_n18993);
and_5  g16645(new_n18993, new_n18992, new_n18994);
nand_5 g16646(new_n18994, new_n18991, new_n18995);
and_5  g16647(new_n18995, new_n18990, new_n18996);
xor_4  g16648(new_n18986, new_n18292, new_n18997);
nand_5 g16649(new_n18997, new_n18996, new_n18998);
and_5  g16650(new_n18998, new_n18987, new_n18999_1);
or_5   g16651(new_n18999_1, new_n18985, new_n19000);
and_5  g16652(new_n19000, new_n18984, new_n19001);
nor_5  g16653(new_n19001, new_n18982_1, new_n19002);
or_5   g16654(new_n19002, new_n18980, new_n19003);
xor_4  g16655(new_n18977_1, new_n5616, new_n19004);
nand_5 g16656(new_n19004, new_n19003, new_n19005_1);
and_5  g16657(new_n19005_1, new_n18978, new_n19006);
or_5   g16658(new_n19006, new_n18976, new_n19007);
and_5  g16659(new_n19007, new_n18975, new_n19008);
or_5   g16660(new_n19008, new_n18973, new_n19009);
and_5  g16661(new_n19009, new_n18972, new_n19010);
or_5   g16662(new_n19010, new_n18970_1, new_n19011);
and_5  g16663(new_n19011, new_n18969, new_n19012);
or_5   g16664(n12702, n12507, new_n19013);
or_5   g16665(new_n18967, new_n18936, new_n19014);
and_5  g16666(new_n19014, new_n19013, new_n19015);
and_5  g16667(new_n19015, new_n19012, new_n19016);
xor_4  g16668(new_n19016, new_n18935, new_n19017);
xor_4  g16669(new_n18933, new_n18930, new_n19018);
not_10 g16670(new_n19018, new_n19019);
xor_4  g16671(new_n19015, new_n19012, new_n19020);
nor_5  g16672(new_n19020, new_n19019, new_n19021);
xor_4  g16673(new_n19020, new_n19019, new_n19022);
xor_4  g16674(new_n18928, new_n18900, new_n19023);
not_10 g16675(new_n19023, new_n19024);
xor_4  g16676(new_n19010, new_n18970_1, new_n19025);
and_5  g16677(new_n19025, new_n19024, new_n19026);
xnor_4 g16678(new_n19025, new_n19023, new_n19027);
xor_4  g16679(new_n18926_1, new_n18905, new_n19028);
not_10 g16680(new_n19028, new_n19029);
xor_4  g16681(new_n19008, new_n18973, new_n19030);
and_5  g16682(new_n19030, new_n19029, new_n19031);
xnor_4 g16683(new_n19030, new_n19028, new_n19032);
xor_4  g16684(new_n18924, new_n18909, new_n19033_1);
not_10 g16685(new_n19033_1, new_n19034);
xor_4  g16686(new_n19006, new_n18976, new_n19035);
and_5  g16687(new_n19035, new_n19034, new_n19036);
xnor_4 g16688(new_n19035, new_n19033_1, new_n19037);
not_10 g16689(new_n19037, new_n19038);
xor_4  g16690(new_n18922, new_n18913, new_n19039);
xnor_4 g16691(new_n19004, new_n19003, new_n19040);
or_5   g16692(new_n19040, new_n19039, new_n19041);
xor_4  g16693(new_n19004, new_n19003, new_n19042_1);
xnor_4 g16694(new_n19042_1, new_n19039, new_n19043);
not_10 g16695(new_n19043, new_n19044_1);
xor_4  g16696(new_n19001, new_n18982_1, new_n19045);
not_10 g16697(new_n19045, new_n19046);
xor_4  g16698(new_n18920, new_n18917, new_n19047);
or_5   g16699(new_n19047, new_n19046, new_n19048);
xnor_4 g16700(new_n19047, new_n19045, new_n19049);
xor_4  g16701(new_n18999_1, new_n18985, new_n19050);
not_10 g16702(new_n19050, new_n19051);
or_5   g16703(new_n19051, new_n13258, new_n19052);
xnor_4 g16704(new_n19050, new_n13258, new_n19053);
not_10 g16705(new_n19053, new_n19054);
xor_4  g16706(new_n18997, new_n18996, new_n19055);
not_10 g16707(new_n19055, new_n19056);
or_5   g16708(new_n19056, new_n6690, new_n19057);
xor_4  g16709(new_n18994, new_n18991, new_n19058);
or_5   g16710(new_n19058, new_n6693, new_n19059);
xor_4  g16711(new_n19058, new_n6693, new_n19060);
nor_5  g16712(new_n17064, new_n17058, new_n19061);
and_5  g16713(new_n17065, new_n6698, new_n19062);
nor_5  g16714(new_n19062, new_n19061, new_n19063);
nand_5 g16715(new_n19063, new_n19060, new_n19064);
and_5  g16716(new_n19064, new_n19059, new_n19065);
xnor_4 g16717(new_n19055, new_n6690, new_n19066);
not_10 g16718(new_n19066, new_n19067);
or_5   g16719(new_n19067, new_n19065, new_n19068);
and_5  g16720(new_n19068, new_n19057, new_n19069);
or_5   g16721(new_n19069, new_n19054, new_n19070);
nand_5 g16722(new_n19070, new_n19052, new_n19071);
nand_5 g16723(new_n19071, new_n19049, new_n19072);
and_5  g16724(new_n19072, new_n19048, new_n19073);
or_5   g16725(new_n19073, new_n19044_1, new_n19074);
and_5  g16726(new_n19074, new_n19041, new_n19075);
nor_5  g16727(new_n19075, new_n19038, new_n19076);
nor_5  g16728(new_n19076, new_n19036, new_n19077);
not_10 g16729(new_n19077, new_n19078);
and_5  g16730(new_n19078, new_n19032, new_n19079);
nor_5  g16731(new_n19079, new_n19031, new_n19080);
not_10 g16732(new_n19080, new_n19081_1);
and_5  g16733(new_n19081_1, new_n19027, new_n19082);
nor_5  g16734(new_n19082, new_n19026, new_n19083);
not_10 g16735(new_n19083, new_n19084);
and_5  g16736(new_n19084, new_n19022, new_n19085);
nor_5  g16737(new_n19085, new_n19021, new_n19086);
not_10 g16738(new_n19086, new_n19087);
xnor_4 g16739(new_n19087, new_n19017, n5351);
and_5  g16740(new_n16757, new_n16751, n5353);
nor_5  g16741(new_n12040, n2160, new_n19090);
nor_5  g16742(new_n12090, new_n12042, new_n19091);
nor_5  g16743(new_n19091, new_n19090, new_n19092);
not_10 g16744(new_n19092, new_n19093);
or_5   g16745(n9934, n2272, new_n19094);
or_5   g16746(new_n12039, new_n12006, new_n19095);
and_5  g16747(new_n19095, new_n19094, new_n19096);
nor_5  g16748(new_n19096, new_n19093, new_n19097);
and_5  g16749(new_n12097, new_n12092, new_n19098);
nor_5  g16750(new_n19098, new_n7310, new_n19099);
nor_5  g16751(new_n12098, new_n7313_1, new_n19100);
not_10 g16752(new_n19100, new_n19101);
nor_5  g16753(new_n12115, new_n12100, new_n19102);
not_10 g16754(new_n19102, new_n19103);
and_5  g16755(new_n19103, new_n19101, new_n19104);
not_10 g16756(new_n19104, new_n19105);
and_5  g16757(new_n19105, new_n19099, new_n19106);
not_10 g16758(new_n19106, new_n19107_1);
xnor_4 g16759(new_n19107_1, new_n19097, new_n19108);
xnor_4 g16760(new_n19096, new_n19093, new_n19109);
xor_4  g16761(new_n19098, new_n7310, new_n19110);
xor_4  g16762(new_n19110, new_n19104, new_n19111);
not_10 g16763(new_n19111, new_n19112);
nor_5  g16764(new_n19112, new_n19109, new_n19113);
xor_4  g16765(new_n19112, new_n19109, new_n19114);
not_10 g16766(new_n19114, new_n19115);
nor_5  g16767(new_n12117, new_n12091, new_n19116_1);
not_10 g16768(new_n19116_1, new_n19117);
not_10 g16769(new_n12118, new_n19118);
nor_5  g16770(new_n12185, new_n19118, new_n19119);
not_10 g16771(new_n19119, new_n19120);
and_5  g16772(new_n19120, new_n19117, new_n19121);
nor_5  g16773(new_n19121, new_n19115, new_n19122);
nor_5  g16774(new_n19122, new_n19113, new_n19123);
xor_4  g16775(new_n19123, new_n19108, n5399);
and_5  g16776(new_n17857, n2979, new_n19125_1);
and_5  g16777(new_n17862, new_n17858, new_n19126);
or_5   g16778(new_n19126, new_n19125_1, new_n19127);
and_5  g16779(new_n14451, n9934, new_n19128);
not_10 g16780(new_n19128, new_n19129);
nor_5  g16781(new_n14451, n9934, new_n19130);
not_10 g16782(new_n17855_1, new_n19131);
nor_5  g16783(new_n19131, new_n19130, new_n19132);
nor_5  g16784(new_n19132, new_n14500, new_n19133);
and_5  g16785(new_n19133, new_n19129, new_n19134);
and_5  g16786(new_n19134, new_n19127, new_n19135);
xnor_4 g16787(new_n19135, new_n19107_1, new_n19136);
xor_4  g16788(new_n19134, new_n19127, new_n19137);
or_5   g16789(new_n19137, new_n19112, new_n19138);
or_5   g16790(new_n17863, new_n12117, new_n19139);
nand_5 g16791(new_n17868, new_n17864, new_n19140);
and_5  g16792(new_n19140, new_n19139, new_n19141_1);
xor_4  g16793(new_n19137, new_n19112, new_n19142);
not_10 g16794(new_n19142, new_n19143);
or_5   g16795(new_n19143, new_n19141_1, new_n19144_1);
and_5  g16796(new_n19144_1, new_n19138, new_n19145);
xor_4  g16797(new_n19145, new_n19136, n5403);
xor_4  g16798(new_n15979_1, new_n15945, n5430);
or_5   g16799(new_n14897, new_n14892, new_n19148);
and_5  g16800(new_n14888, new_n10650_1, new_n19149);
or_5   g16801(new_n14888, new_n10650_1, new_n19150);
and_5  g16802(new_n14898, new_n19150, new_n19151);
or_5   g16803(new_n19151, new_n19149, new_n19152);
nor_5  g16804(new_n19152, new_n10509, new_n19153);
and_5  g16805(new_n19153, new_n19148, n5439);
xnor_4 g16806(new_n12527, new_n12505, n5472);
xnor_4 g16807(new_n8530, new_n8491, n5485);
xnor_4 g16808(new_n18564, new_n18546, n5524);
and_5  g16809(new_n16769, new_n6004, new_n19158);
and_5  g16810(new_n19158, new_n5999, new_n19159);
and_5  g16811(new_n19159, new_n5993, new_n19160);
and_5  g16812(new_n19160, new_n5987, new_n19161);
and_5  g16813(new_n19161, new_n5981, new_n19162);
and_5  g16814(new_n19162, new_n5975, new_n19163_1);
and_5  g16815(new_n19163_1, new_n5970, new_n19164_1);
xnor_4 g16816(new_n19164_1, new_n5966, new_n19165);
nor_5  g16817(new_n19165, new_n14055, new_n19166);
xor_4  g16818(new_n19165, new_n14054, new_n19167);
xnor_4 g16819(new_n19163_1, new_n5972, new_n19168);
or_5   g16820(new_n19168, new_n14059_1, new_n19169);
xnor_4 g16821(new_n19168, new_n14059_1, new_n19170);
xnor_4 g16822(new_n19162, new_n5977, new_n19171);
or_5   g16823(new_n19171, new_n14063, new_n19172);
xnor_4 g16824(new_n19171, new_n14063, new_n19173);
not_10 g16825(new_n14067, new_n19174_1);
xnor_4 g16826(new_n19161, new_n5983, new_n19175);
or_5   g16827(new_n19175, new_n19174_1, new_n19176_1);
xnor_4 g16828(new_n19175, new_n19174_1, new_n19177);
xor_4  g16829(new_n19160, new_n5989, new_n19178);
nand_5 g16830(new_n19178, new_n14071_1, new_n19179);
xnor_4 g16831(new_n19178, new_n14071_1, new_n19180);
xnor_4 g16832(new_n19159, new_n5995, new_n19181);
or_5   g16833(new_n19181, new_n14075, new_n19182);
xnor_4 g16834(new_n19181, new_n14075, new_n19183);
xnor_4 g16835(new_n19158, new_n6001, new_n19184);
or_5   g16836(new_n17871, new_n13348, new_n19185);
or_5   g16837(new_n17875, new_n17872, new_n19186);
and_5  g16838(new_n19186, new_n19185, new_n19187);
or_5   g16839(new_n19187, new_n19184, new_n19188);
xor_4  g16840(new_n19187, new_n19184, new_n19189);
nand_5 g16841(new_n19189, new_n13346, new_n19190);
and_5  g16842(new_n19190, new_n19188, new_n19191);
or_5   g16843(new_n19191, new_n19183, new_n19192);
and_5  g16844(new_n19192, new_n19182, new_n19193);
or_5   g16845(new_n19193, new_n19180, new_n19194);
and_5  g16846(new_n19194, new_n19179, new_n19195);
or_5   g16847(new_n19195, new_n19177, new_n19196_1);
and_5  g16848(new_n19196_1, new_n19176_1, new_n19197);
or_5   g16849(new_n19197, new_n19173, new_n19198);
and_5  g16850(new_n19198, new_n19172, new_n19199);
or_5   g16851(new_n19199, new_n19170, new_n19200);
and_5  g16852(new_n19200, new_n19169, new_n19201);
nor_5  g16853(new_n19201, new_n19167, new_n19202_1);
nor_5  g16854(new_n19202_1, new_n19166, new_n19203);
and_5  g16855(new_n19164_1, new_n5965, new_n19204);
not_10 g16856(new_n19204, new_n19205);
and_5  g16857(new_n19205, new_n13716, new_n19206);
and_5  g16858(new_n19204, new_n13714_1, new_n19207);
nor_5  g16859(new_n19207, new_n19206, new_n19208);
xor_4  g16860(new_n19208, new_n14100, new_n19209);
xor_4  g16861(new_n19209, new_n19203, new_n19210);
nor_5  g16862(new_n19210, new_n4815, new_n19211);
xor_4  g16863(new_n19210, new_n4815, new_n19212);
xor_4  g16864(new_n19201, new_n19167, new_n19213);
and_5  g16865(new_n19213, new_n4977, new_n19214);
xor_4  g16866(new_n19213, new_n4977, new_n19215);
not_10 g16867(new_n19215, new_n19216);
xor_4  g16868(new_n19199, new_n19170, new_n19217);
and_5  g16869(new_n19217, new_n4982, new_n19218);
xor_4  g16870(new_n19217, new_n4982, new_n19219);
not_10 g16871(new_n19219, new_n19220_1);
xor_4  g16872(new_n19197, new_n19173, new_n19221_1);
and_5  g16873(new_n19221_1, new_n4988, new_n19222);
xor_4  g16874(new_n19221_1, new_n4988, new_n19223_1);
not_10 g16875(new_n19223_1, new_n19224_1);
xor_4  g16876(new_n19195, new_n19177, new_n19225);
and_5  g16877(new_n19225, new_n4994, new_n19226);
xor_4  g16878(new_n19225, new_n4994, new_n19227);
not_10 g16879(new_n19227, new_n19228_1);
xor_4  g16880(new_n19193, new_n19180, new_n19229);
and_5  g16881(new_n19229, new_n5000, new_n19230);
xor_4  g16882(new_n19229, new_n5000, new_n19231);
not_10 g16883(new_n19231, new_n19232);
xor_4  g16884(new_n19191, new_n19183, new_n19233_1);
and_5  g16885(new_n19233_1, new_n5006, new_n19234_1);
xor_4  g16886(new_n19233_1, new_n5006, new_n19235);
not_10 g16887(new_n19235, new_n19236);
xnor_4 g16888(new_n19189, new_n13345, new_n19237);
and_5  g16889(new_n19237, new_n5012, new_n19238);
not_10 g16890(new_n19238, new_n19239);
xor_4  g16891(new_n19237, new_n5012, new_n19240);
nor_5  g16892(new_n17876, new_n5019, new_n19241);
nor_5  g16893(new_n17879, new_n17877_1, new_n19242);
nor_5  g16894(new_n19242, new_n19241, new_n19243);
and_5  g16895(new_n19243, new_n19240, new_n19244_1);
not_10 g16896(new_n19244_1, new_n19245);
and_5  g16897(new_n19245, new_n19239, new_n19246);
nor_5  g16898(new_n19246, new_n19236, new_n19247);
nor_5  g16899(new_n19247, new_n19234_1, new_n19248);
nor_5  g16900(new_n19248, new_n19232, new_n19249);
nor_5  g16901(new_n19249, new_n19230, new_n19250);
nor_5  g16902(new_n19250, new_n19228_1, new_n19251);
nor_5  g16903(new_n19251, new_n19226, new_n19252);
nor_5  g16904(new_n19252, new_n19224_1, new_n19253);
nor_5  g16905(new_n19253, new_n19222, new_n19254);
nor_5  g16906(new_n19254, new_n19220_1, new_n19255);
nor_5  g16907(new_n19255, new_n19218, new_n19256);
nor_5  g16908(new_n19256, new_n19216, new_n19257);
or_5   g16909(new_n19257, new_n19214, new_n19258);
and_5  g16910(new_n19258, new_n19212, new_n19259);
or_5   g16911(new_n19259, new_n19211, new_n19260);
nor_5  g16912(new_n19208, new_n14100, new_n19261);
and_5  g16913(new_n19208, new_n14100, new_n19262);
nor_5  g16914(new_n19262, new_n19203, new_n19263);
nor_5  g16915(new_n19263, new_n19261, new_n19264);
nor_5  g16916(new_n19264, new_n19207, new_n19265);
xnor_4 g16917(new_n19265, new_n19260, n5564);
xor_4  g16918(new_n6973, new_n6960, n5593);
xor_4  g16919(new_n17913, new_n14527, new_n19268);
not_10 g16920(new_n19268, new_n19269);
xnor_4 g16921(new_n16666, new_n16658, new_n19270_1);
nor_5  g16922(new_n19270_1, new_n14534, new_n19271);
xnor_4 g16923(new_n16667, new_n14534, new_n19272);
not_10 g16924(new_n19272, new_n19273);
xnor_4 g16925(new_n16664, new_n16660, new_n19274);
nor_5  g16926(new_n19274, new_n14540, new_n19275);
xnor_4 g16927(new_n16669, new_n14540, new_n19276);
not_10 g16928(new_n19276, new_n19277);
xnor_4 g16929(new_n15692, new_n15680, new_n19278);
nor_5  g16930(new_n19278, new_n14546_1, new_n19279);
xnor_4 g16931(new_n15693, new_n14546_1, new_n19280);
not_10 g16932(new_n19280, new_n19281);
xnor_4 g16933(new_n15690, new_n15683, new_n19282_1);
nor_5  g16934(new_n19282_1, new_n14552, new_n19283);
not_10 g16935(new_n19283, new_n19284);
and_5  g16936(new_n17475, new_n17464, new_n19285);
not_10 g16937(new_n19285, new_n19286);
and_5  g16938(new_n19286, new_n19284, new_n19287);
nor_5  g16939(new_n19287, new_n19281, new_n19288);
nor_5  g16940(new_n19288, new_n19279, new_n19289);
nor_5  g16941(new_n19289, new_n19277, new_n19290);
nor_5  g16942(new_n19290, new_n19275, new_n19291);
nor_5  g16943(new_n19291, new_n19273, new_n19292);
nor_5  g16944(new_n19292, new_n19271, new_n19293);
xnor_4 g16945(new_n19293, new_n19269, n5603);
xor_4  g16946(n17911, n14440, new_n19295);
not_10 g16947(n21997, new_n19296);
or_5   g16948(new_n19296, n1654, new_n19297);
xor_4  g16949(n21997, n1654, new_n19298);
or_5   g16950(new_n8652, n13783, new_n19299);
xor_4  g16951(n25119, n13783, new_n19300);
or_5   g16952(n26660, new_n8654, new_n19301);
xor_4  g16953(n26660, n1163, new_n19302);
or_5   g16954(new_n8656_1, n3018, new_n19303);
or_5   g16955(n18537, new_n10855, new_n19304);
and_5  g16956(new_n8660, n3480, new_n19305);
nor_5  g16957(new_n18212, new_n18201, new_n19306);
nor_5  g16958(new_n19306, new_n19305, new_n19307);
nand_5 g16959(new_n19307, new_n19304, new_n19308);
and_5  g16960(new_n19308, new_n19303, new_n19309);
or_5   g16961(new_n19309, new_n19302, new_n19310);
and_5  g16962(new_n19310, new_n19301, new_n19311);
or_5   g16963(new_n19311, new_n19300, new_n19312);
and_5  g16964(new_n19312, new_n19299, new_n19313);
or_5   g16965(new_n19313, new_n19298, new_n19314_1);
and_5  g16966(new_n19314_1, new_n19297, new_n19315_1);
xor_4  g16967(new_n19315_1, new_n19295, new_n19316);
xor_4  g16968(new_n19316, new_n3009, new_n19317);
xor_4  g16969(new_n19313, new_n19298, new_n19318);
or_5   g16970(new_n19318, new_n3013, new_n19319);
xor_4  g16971(new_n19318, new_n3013, new_n19320);
not_10 g16972(new_n19320, new_n19321);
xor_4  g16973(new_n19311, new_n19300, new_n19322);
not_10 g16974(new_n19322, new_n19323_1);
nand_5 g16975(new_n19323_1, new_n3019, new_n19324);
xnor_4 g16976(new_n19322, new_n3019, new_n19325);
not_10 g16977(new_n19325, new_n19326);
xnor_4 g16978(new_n19309, new_n19302, new_n19327_1);
nand_5 g16979(new_n19327_1, new_n3025, new_n19328);
xor_4  g16980(new_n19327_1, new_n3025, new_n19329);
xnor_4 g16981(n18537, n3018, new_n19330);
xnor_4 g16982(new_n19330, new_n19307, new_n19331);
nor_5  g16983(new_n19331, new_n3031, new_n19332);
nor_5  g16984(new_n18213, new_n3035, new_n19333_1);
and_5  g16985(new_n18230, new_n18214, new_n19334);
or_5   g16986(new_n19334, new_n19333_1, new_n19335);
xor_4  g16987(new_n19331, new_n3031, new_n19336);
and_5  g16988(new_n19336, new_n19335, new_n19337);
nor_5  g16989(new_n19337, new_n19332, new_n19338);
nand_5 g16990(new_n19338, new_n19329, new_n19339);
and_5  g16991(new_n19339, new_n19328, new_n19340);
or_5   g16992(new_n19340, new_n19326, new_n19341);
and_5  g16993(new_n19341, new_n19324, new_n19342);
or_5   g16994(new_n19342, new_n19321, new_n19343);
and_5  g16995(new_n19343, new_n19319, new_n19344);
xor_4  g16996(new_n19344, new_n19317, n5609);
xnor_4 g16997(new_n13660, new_n13640, n5634);
or_5   g16998(new_n3183, n2978, new_n19347);
xor_4  g16999(n3425, n2978, new_n19348_1);
or_5   g17000(n23697, new_n3184, new_n19349);
xor_4  g17001(n23697, n9967, new_n19350);
or_5   g17002(new_n3185, n2289, new_n19351);
or_5   g17003(new_n18773, new_n18766, new_n19352);
and_5  g17004(new_n19352, new_n19351, new_n19353);
or_5   g17005(new_n19353, new_n19350, new_n19354_1);
and_5  g17006(new_n19354_1, new_n19349, new_n19355);
or_5   g17007(new_n19355, new_n19348_1, new_n19356);
and_5  g17008(new_n19356, new_n19347, new_n19357_1);
nor_5  g17009(new_n19357_1, new_n7371, new_n19358);
and_5  g17010(new_n19357_1, new_n7371, new_n19359);
xor_4  g17011(new_n19355, new_n19348_1, new_n19360);
nor_5  g17012(new_n19360, new_n7420, new_n19361_1);
xor_4  g17013(new_n19360, new_n7420, new_n19362);
not_10 g17014(new_n19362, new_n19363);
xor_4  g17015(new_n19353, new_n19350, new_n19364);
nor_5  g17016(new_n19364, new_n7426, new_n19365);
not_10 g17017(new_n19365, new_n19366);
xor_4  g17018(new_n19364, new_n7426, new_n19367_1);
nor_5  g17019(new_n18774, new_n7432_1, new_n19368);
not_10 g17020(new_n19368, new_n19369);
not_10 g17021(new_n18789, new_n19370);
and_5  g17022(new_n19370, new_n18775, new_n19371);
not_10 g17023(new_n19371, new_n19372);
and_5  g17024(new_n19372, new_n19369, new_n19373);
not_10 g17025(new_n19373, new_n19374);
and_5  g17026(new_n19374, new_n19367_1, new_n19375);
not_10 g17027(new_n19375, new_n19376);
and_5  g17028(new_n19376, new_n19366, new_n19377);
nor_5  g17029(new_n19377, new_n19363, new_n19378);
nor_5  g17030(new_n19378, new_n19361_1, new_n19379);
nor_5  g17031(new_n19379, new_n19359, new_n19380);
nor_5  g17032(new_n19380, new_n19358, new_n19381);
nand_5 g17033(new_n7310, new_n7294, new_n19382);
nand_5 g17034(new_n7370, new_n7311, new_n19383);
and_5  g17035(new_n19383, new_n19382, new_n19384);
xnor_4 g17036(new_n19384, new_n19357_1, new_n19385_1);
xor_4  g17037(new_n19385_1, new_n19381, n5643);
xor_4  g17038(n18035, n5834, new_n19387);
or_5   g17039(n13851, new_n10743, new_n19388);
or_5   g17040(new_n15773, new_n15758, new_n19389_1);
and_5  g17041(new_n19389_1, new_n19388, new_n19390);
xor_4  g17042(new_n19390, new_n19387, new_n19391);
xor_4  g17043(new_n19391, new_n15283, new_n19392);
or_5   g17044(new_n15774, new_n15311, new_n19393);
xor_4  g17045(new_n15774, new_n15311, new_n19394);
not_10 g17046(new_n19394, new_n19395);
or_5   g17047(new_n15778, new_n15317, new_n19396);
xor_4  g17048(new_n15778, new_n15317, new_n19397);
or_5   g17049(new_n15783, new_n15323, new_n19398);
xor_4  g17050(new_n15783, new_n15323, new_n19399);
or_5   g17051(new_n15785, new_n15326, new_n19400);
nand_5 g17052(new_n14165, new_n13906, new_n19401_1);
xor_4  g17053(new_n14165, new_n13906, new_n19402);
nand_5 g17054(new_n14181, new_n13912_1, new_n19403);
xor_4  g17055(new_n14181, new_n13912_1, new_n19404);
and_5  g17056(new_n14188, new_n13915, new_n19405);
or_5   g17057(new_n19405, new_n13920, new_n19406);
xnor_4 g17058(new_n19405, new_n13919, new_n19407);
nand_5 g17059(new_n19407, new_n14195, new_n19408);
nand_5 g17060(new_n19408, new_n19406, new_n19409);
nand_5 g17061(new_n19409, new_n19404, new_n19410);
nand_5 g17062(new_n19410, new_n19403, new_n19411);
nand_5 g17063(new_n19411, new_n19402, new_n19412);
nand_5 g17064(new_n19412, new_n19401_1, new_n19413);
xnor_4 g17065(new_n15785, new_n15331, new_n19414_1);
nand_5 g17066(new_n19414_1, new_n19413, new_n19415);
nand_5 g17067(new_n19415, new_n19400, new_n19416);
nand_5 g17068(new_n19416, new_n19399, new_n19417);
nand_5 g17069(new_n19417, new_n19398, new_n19418);
nand_5 g17070(new_n19418, new_n19397, new_n19419);
and_5  g17071(new_n19419, new_n19396, new_n19420);
or_5   g17072(new_n19420, new_n19395, new_n19421);
and_5  g17073(new_n19421, new_n19393, new_n19422);
xor_4  g17074(new_n19422, new_n19392, n5680);
xnor_4 g17075(new_n14991, new_n14990, n5687);
xnor_4 g17076(new_n16116, new_n16108, n5700);
xor_4  g17077(new_n10713, new_n10659, n5732);
xnor_4 g17078(n23775, n8381, new_n19427);
or_5   g17079(n20235, n8259, new_n19428);
nand_5 g17080(new_n18684, new_n18683, new_n19429);
and_5  g17081(new_n19429, new_n19428, new_n19430);
xor_4  g17082(new_n19430, new_n19427, new_n19431);
xor_4  g17083(new_n19431, new_n2397, new_n19432);
or_5   g17084(new_n18685, new_n2388_1, new_n19433);
nand_5 g17085(new_n18686, new_n18682, new_n19434);
and_5  g17086(new_n19434, new_n19433, new_n19435);
xor_4  g17087(new_n19435, new_n19432, new_n19436);
not_10 g17088(new_n19436, new_n19437);
xor_4  g17089(n8869, n6385, new_n19438);
or_5   g17090(new_n2367, n10372, new_n19439);
nand_5 g17091(new_n18679_1, new_n18678, new_n19440);
and_5  g17092(new_n19440, new_n19439, new_n19441);
xor_4  g17093(new_n19441, new_n19438, new_n19442);
xor_4  g17094(new_n19442, new_n19437, new_n19443);
nor_5  g17095(new_n18680, new_n18677, new_n19444);
not_10 g17096(new_n19444, new_n19445);
and_5  g17097(new_n18687, new_n18681, new_n19446);
not_10 g17098(new_n19446, new_n19447);
and_5  g17099(new_n19447, new_n19445, new_n19448);
xor_4  g17100(new_n19448, new_n19443, n5742);
xnor_4 g17101(new_n13927, new_n13925, n5765);
xnor_4 g17102(new_n12763, new_n12718, n5776);
xnor_4 g17103(new_n2827, new_n2790, n5782);
xnor_4 g17104(n18901, n1163, new_n19453);
or_5   g17105(n18537, n4376, new_n19454_1);
xnor_4 g17106(n18537, n4376, new_n19455);
or_5   g17107(n14570, n7057, new_n19456);
xor_4  g17108(n14570, n7057, new_n19457);
not_10 g17109(new_n19457, new_n19458_1);
or_5   g17110(n23775, n8381, new_n19459);
or_5   g17111(new_n19430, new_n19427, new_n19460);
and_5  g17112(new_n19460, new_n19459, new_n19461);
or_5   g17113(new_n19461, new_n19458_1, new_n19462);
and_5  g17114(new_n19462, new_n19456, new_n19463);
or_5   g17115(new_n19463, new_n19455, new_n19464);
and_5  g17116(new_n19464, new_n19454_1, new_n19465);
xor_4  g17117(new_n19465, new_n19453, new_n19466);
xor_4  g17118(new_n19466, new_n2453, new_n19467_1);
xor_4  g17119(new_n19463, new_n19455, new_n19468);
nand_5 g17120(new_n19468, new_n2413, new_n19469);
xor_4  g17121(new_n19461, new_n19457, new_n19470);
nand_5 g17122(new_n19431, new_n2397, new_n19471);
nand_5 g17123(new_n19435, new_n19432, new_n19472_1);
and_5  g17124(new_n19472_1, new_n19471, new_n19473);
nor_5  g17125(new_n19473, new_n19470, new_n19474);
not_10 g17126(new_n19474, new_n19475);
xor_4  g17127(new_n19473, new_n19470, new_n19476);
and_5  g17128(new_n19476, new_n2464, new_n19477_1);
not_10 g17129(new_n19477_1, new_n19478);
and_5  g17130(new_n19478, new_n19475, new_n19479);
xnor_4 g17131(new_n19468, new_n2413, new_n19480);
or_5   g17132(new_n19480, new_n19479, new_n19481);
and_5  g17133(new_n19481, new_n19469, new_n19482);
xor_4  g17134(new_n19482, new_n19467_1, new_n19483);
not_10 g17135(new_n19483, new_n19484);
xor_4  g17136(n23068, n7099, new_n19485);
or_5   g17137(n19514, new_n12060, new_n19486);
xnor_4 g17138(n19514, n12811, new_n19487);
not_10 g17139(new_n19487, new_n19488);
or_5   g17140(n10053, new_n12064, new_n19489);
xnor_4 g17141(n10053, n1118, new_n19490);
or_5   g17142(n25974, new_n3817, new_n19491);
nand_5 g17143(n25974, new_n3817, new_n19492);
and_5  g17144(n9507, new_n15026, new_n19493);
and_5  g17145(new_n3823, n1630, new_n19494_1);
not_10 g17146(new_n19494_1, new_n19495);
and_5  g17147(n26979, new_n12069, new_n19496_1);
and_5  g17148(new_n19496_1, new_n19495, new_n19497);
nor_5  g17149(new_n19497, new_n19493, new_n19498);
not_10 g17150(new_n19498, new_n19499);
nand_5 g17151(new_n19499, new_n19492, new_n19500);
and_5  g17152(new_n19500, new_n19491, new_n19501);
nand_5 g17153(new_n19501, new_n19490, new_n19502);
and_5  g17154(new_n19502, new_n19489, new_n19503);
or_5   g17155(new_n19503, new_n19488, new_n19504);
and_5  g17156(new_n19504, new_n19486, new_n19505);
xor_4  g17157(new_n19505, new_n19485, new_n19506);
xnor_4 g17158(new_n19506, new_n19484, new_n19507);
xor_4  g17159(new_n19503, new_n19487, new_n19508);
xor_4  g17160(new_n19480, new_n19479, new_n19509);
nor_5  g17161(new_n19509, new_n19508, new_n19510);
xnor_4 g17162(new_n19476, new_n2404, new_n19511);
not_10 g17163(new_n19511, new_n19512);
xor_4  g17164(new_n19501, new_n19490, new_n19513);
or_5   g17165(new_n19513, new_n19512, new_n19514_1);
xor_4  g17166(new_n19513, new_n19512, new_n19515_1);
xnor_4 g17167(n25974, n8399, new_n19516);
xor_4  g17168(new_n19516, new_n19499, new_n19517);
nand_5 g17169(new_n19517, new_n19436, new_n19518);
xnor_4 g17170(new_n19517, new_n19437, new_n19519);
xnor_4 g17171(n26979, n1451, new_n19520);
nor_5  g17172(new_n19520, new_n18675, new_n19521);
not_10 g17173(new_n19521, new_n19522);
xnor_4 g17174(n9507, n1630, new_n19523_1);
xor_4  g17175(new_n19523_1, new_n19496_1, new_n19524);
nand_5 g17176(new_n19524, new_n19522, new_n19525);
not_10 g17177(new_n18687, new_n19526);
xor_4  g17178(new_n19524, new_n19522, new_n19527);
nand_5 g17179(new_n19527, new_n19526, new_n19528);
nand_5 g17180(new_n19528, new_n19525, new_n19529);
nand_5 g17181(new_n19529, new_n19519, new_n19530);
nand_5 g17182(new_n19530, new_n19518, new_n19531_1);
nand_5 g17183(new_n19531_1, new_n19515_1, new_n19532);
and_5  g17184(new_n19532, new_n19514_1, new_n19533);
xor_4  g17185(new_n19509, new_n19508, new_n19534);
and_5  g17186(new_n19534, new_n19533, new_n19535);
nor_5  g17187(new_n19535, new_n19510, new_n19536);
xnor_4 g17188(new_n19536, new_n19507, n5833);
xnor_4 g17189(new_n12759, new_n12730, n5840);
xor_4  g17190(new_n19336, new_n19335, n5841);
xnor_4 g17191(new_n13233, new_n13231, n5850);
xnor_4 g17192(new_n19411, new_n19402, n5903);
xor_4  g17193(new_n16845, new_n8810, new_n19542);
not_10 g17194(new_n19542, new_n19543);
or_5   g17195(new_n16848, new_n8814, new_n19544);
or_5   g17196(new_n18833, new_n18818, new_n19545);
and_5  g17197(new_n19545, new_n19544, new_n19546);
xor_4  g17198(new_n19546, new_n19543, new_n19547);
not_10 g17199(n26752, new_n19548);
and_5  g17200(new_n18795, new_n18791, new_n19549);
xor_4  g17201(new_n19549, new_n19548, new_n19550);
xor_4  g17202(new_n19550, new_n8973, new_n19551);
or_5   g17203(new_n18796, new_n8977, new_n19552);
nand_5 g17204(new_n18814, new_n18799, new_n19553);
nand_5 g17205(new_n19553, new_n18797, new_n19554);
and_5  g17206(new_n19554, new_n19552, new_n19555);
xor_4  g17207(new_n19555, new_n19551, new_n19556);
xnor_4 g17208(new_n19556, new_n19547, new_n19557);
not_10 g17209(new_n19557, new_n19558);
nor_5  g17210(new_n18834, new_n18817, new_n19559);
nor_5  g17211(new_n18862, new_n18836, new_n19560);
nor_5  g17212(new_n19560, new_n19559, new_n19561);
xnor_4 g17213(new_n19561, new_n19558, n5904);
xor_4  g17214(n27089, n6814, new_n19563);
or_5   g17215(new_n9150, n11841, new_n19564);
xor_4  g17216(n19701, n11841, new_n19565);
or_5   g17217(new_n9154, n10710, new_n19566);
xor_4  g17218(n23529, n10710, new_n19567);
or_5   g17219(new_n9158, n20929, new_n19568);
xor_4  g17220(n24620, n20929, new_n19569);
or_5   g17221(n8006, new_n9162, new_n19570_1);
xor_4  g17222(n8006, n5211, new_n19571);
or_5   g17223(n25074, new_n9166_1, new_n19572);
xnor_4 g17224(n25074, n12956, new_n19573);
or_5   g17225(n18295, new_n4322, new_n19574);
or_5   g17226(new_n9171, n16396, new_n19575_1);
and_5  g17227(n9399, new_n9173, new_n19576);
and_5  g17228(new_n4325_1, n6502, new_n19577);
not_10 g17229(new_n19577, new_n19578);
and_5  g17230(new_n9178, n2088, new_n19579);
and_5  g17231(new_n19579, new_n19578, new_n19580);
nor_5  g17232(new_n19580, new_n19576, new_n19581);
not_10 g17233(new_n19581, new_n19582);
nand_5 g17234(new_n19582, new_n19575_1, new_n19583);
and_5  g17235(new_n19583, new_n19574, new_n19584_1);
nand_5 g17236(new_n19584_1, new_n19573, new_n19585);
and_5  g17237(new_n19585, new_n19572, new_n19586);
or_5   g17238(new_n19586, new_n19571, new_n19587);
and_5  g17239(new_n19587, new_n19570_1, new_n19588);
or_5   g17240(new_n19588, new_n19569, new_n19589);
and_5  g17241(new_n19589, new_n19568, new_n19590);
or_5   g17242(new_n19590, new_n19567, new_n19591);
and_5  g17243(new_n19591, new_n19566, new_n19592);
or_5   g17244(new_n19592, new_n19565, new_n19593);
and_5  g17245(new_n19593, new_n19564, new_n19594);
xor_4  g17246(new_n19594, new_n19563, new_n19595);
xor_4  g17247(new_n19595, new_n10399, new_n19596);
xor_4  g17248(new_n19592, new_n19565, new_n19597);
nor_5  g17249(new_n19597, new_n10404_1, new_n19598);
xnor_4 g17250(new_n19597, new_n10403, new_n19599);
xnor_4 g17251(new_n19590, new_n19567, new_n19600);
and_5  g17252(new_n19600, new_n10410, new_n19601);
xor_4  g17253(new_n19600, new_n10410, new_n19602_1);
xor_4  g17254(new_n19588, new_n19569, new_n19603);
nor_5  g17255(new_n19603, new_n10415, new_n19604);
xor_4  g17256(new_n19586, new_n19571, new_n19605);
nor_5  g17257(new_n19605, new_n10418, new_n19606);
xor_4  g17258(new_n19605, new_n10418, new_n19607);
not_10 g17259(new_n19607, new_n19608_1);
xor_4  g17260(new_n19584_1, new_n19573, new_n19609);
nor_5  g17261(new_n19609, new_n10423, new_n19610);
xnor_4 g17262(n18295, n16396, new_n19611);
xor_4  g17263(new_n19611, new_n19582, new_n19612);
and_5  g17264(new_n19612, new_n10426, new_n19613);
not_10 g17265(new_n19613, new_n19614);
xor_4  g17266(new_n19612, new_n10426, new_n19615);
xnor_4 g17267(n15780, n2088, new_n19616);
or_5   g17268(new_n19616, new_n10432_1, new_n19617_1);
xnor_4 g17269(n9399, n6502, new_n19618_1);
xor_4  g17270(new_n19618_1, new_n19579, new_n19619);
nor_5  g17271(new_n19619, new_n19617_1, new_n19620);
xor_4  g17272(new_n19619, new_n19617_1, new_n19621);
and_5  g17273(new_n19621, new_n10438, new_n19622);
nor_5  g17274(new_n19622, new_n19620, new_n19623_1);
and_5  g17275(new_n19623_1, new_n19615, new_n19624);
not_10 g17276(new_n19624, new_n19625);
and_5  g17277(new_n19625, new_n19614, new_n19626);
xnor_4 g17278(new_n19609, new_n10422, new_n19627);
not_10 g17279(new_n19627, new_n19628);
nor_5  g17280(new_n19628, new_n19626, new_n19629);
nor_5  g17281(new_n19629, new_n19610, new_n19630);
nor_5  g17282(new_n19630, new_n19608_1, new_n19631);
nor_5  g17283(new_n19631, new_n19606, new_n19632);
not_10 g17284(new_n19632, new_n19633);
xor_4  g17285(new_n19603, new_n10415, new_n19634);
and_5  g17286(new_n19634, new_n19633, new_n19635);
nor_5  g17287(new_n19635, new_n19604, new_n19636);
not_10 g17288(new_n19636, new_n19637);
and_5  g17289(new_n19637, new_n19602_1, new_n19638);
nor_5  g17290(new_n19638, new_n19601, new_n19639);
not_10 g17291(new_n19639, new_n19640);
and_5  g17292(new_n19640, new_n19599, new_n19641_1);
nor_5  g17293(new_n19641_1, new_n19598, new_n19642);
not_10 g17294(new_n19642, new_n19643);
xnor_4 g17295(new_n19643, new_n19596, n5911);
xnor_4 g17296(new_n12152_1, new_n3921, n5936);
xnor_4 g17297(new_n10248, new_n10201_1, n5943);
xnor_4 g17298(new_n14577, new_n14543, n5964);
or_5   g17299(new_n5091, n11184, new_n19648_1);
or_5   g17300(new_n5076, n23146, new_n19649);
nor_5  g17301(new_n5079, n17968, new_n19650);
nand_5 g17302(new_n19650, new_n5082_1, new_n19651);
and_5  g17303(new_n19651, new_n19649, new_n19652_1);
or_5   g17304(new_n19652_1, new_n5092, new_n19653);
and_5  g17305(new_n19653, new_n19648_1, new_n19654);
nand_5 g17306(new_n19654, new_n16320, new_n19655);
or_5   g17307(new_n19654, new_n16321, new_n19656);
nand_5 g17308(new_n19656, n8255, new_n19657);
and_5  g17309(new_n19657, new_n19655, new_n19658);
or_5   g17310(new_n19658, new_n16310, new_n19659);
and_5  g17311(new_n19658, new_n16313, new_n19660);
or_5   g17312(new_n19660, new_n16312, new_n19661);
and_5  g17313(new_n19661, new_n19659, new_n19662);
or_5   g17314(new_n19662, new_n16306, new_n19663);
and_5  g17315(new_n19662, new_n16309, new_n19664_1);
or_5   g17316(new_n19664_1, new_n16308, new_n19665);
and_5  g17317(new_n19665, new_n19663, new_n19666);
or_5   g17318(new_n19666, new_n16304, new_n19667);
and_5  g17319(new_n19666, new_n16329, new_n19668);
or_5   g17320(new_n19668, new_n16328, new_n19669);
and_5  g17321(new_n19669, new_n19667, new_n19670);
or_5   g17322(new_n19670, new_n16302, new_n19671);
not_10 g17323(new_n16333, new_n19672);
nand_5 g17324(new_n19670, new_n19672, new_n19673);
nand_5 g17325(new_n19673, n15602, new_n19674);
and_5  g17326(new_n19674, new_n19671, new_n19675);
xnor_4 g17327(new_n19675, new_n16301, new_n19676);
xor_4  g17328(new_n19676, new_n3207, new_n19677);
xnor_4 g17329(new_n19670, new_n16333, new_n19678);
nand_5 g17330(new_n19678, new_n3213, new_n19679);
xnor_4 g17331(new_n19678, new_n3213, new_n19680_1);
xnor_4 g17332(new_n19666, new_n16330, new_n19681);
nand_5 g17333(new_n19681, new_n3218, new_n19682);
xnor_4 g17334(new_n19681, new_n3218, new_n19683);
xor_4  g17335(new_n19662, new_n16309, new_n19684);
nand_5 g17336(new_n19684, new_n3223, new_n19685);
xnor_4 g17337(new_n19684, new_n3223, new_n19686);
xor_4  g17338(new_n19658, new_n16313, new_n19687);
nand_5 g17339(new_n19687, new_n3228_1, new_n19688);
xor_4  g17340(new_n19687, new_n3228_1, new_n19689);
not_10 g17341(new_n19689, new_n19690);
xor_4  g17342(new_n19654, new_n16321, new_n19691);
nand_5 g17343(new_n19691, new_n3233, new_n19692);
xor_4  g17344(new_n19691, new_n3233, new_n19693);
not_10 g17345(new_n19693, new_n19694);
xor_4  g17346(new_n19652_1, new_n5092, new_n19695);
nand_5 g17347(new_n19695, new_n3238, new_n19696);
xor_4  g17348(new_n19695, new_n3238, new_n19697);
not_10 g17349(new_n19697, new_n19698);
not_10 g17350(new_n3246, new_n19699);
xor_4  g17351(new_n19650, new_n5082_1, new_n19700);
nand_5 g17352(new_n19700, new_n19699, new_n19701_1);
and_5  g17353(new_n5101_1, new_n3243, new_n19702);
xor_4  g17354(new_n19700, new_n19699, new_n19703);
not_10 g17355(new_n19703, new_n19704);
or_5   g17356(new_n19704, new_n19702, new_n19705);
and_5  g17357(new_n19705, new_n19701_1, new_n19706);
or_5   g17358(new_n19706, new_n19698, new_n19707);
and_5  g17359(new_n19707, new_n19696, new_n19708);
or_5   g17360(new_n19708, new_n19694, new_n19709);
and_5  g17361(new_n19709, new_n19692, new_n19710);
or_5   g17362(new_n19710, new_n19690, new_n19711);
and_5  g17363(new_n19711, new_n19688, new_n19712);
or_5   g17364(new_n19712, new_n19686, new_n19713);
and_5  g17365(new_n19713, new_n19685, new_n19714);
or_5   g17366(new_n19714, new_n19683, new_n19715);
and_5  g17367(new_n19715, new_n19682, new_n19716);
or_5   g17368(new_n19716, new_n19680_1, new_n19717);
and_5  g17369(new_n19717, new_n19679, new_n19718);
xnor_4 g17370(new_n19718, new_n19677, n5980);
xnor_4 g17371(new_n11452, new_n11429, n6012);
nor_5  g17372(new_n10341, n16544, new_n19721);
xor_4  g17373(new_n10341, n16544, new_n19722);
not_10 g17374(new_n19722, new_n19723);
or_5   g17375(new_n10344, n6814, new_n19724);
xor_4  g17376(new_n10344, n6814, new_n19725);
not_10 g17377(new_n19725, new_n19726);
or_5   g17378(new_n10349, n19701, new_n19727);
xor_4  g17379(new_n10349, n19701, new_n19728);
not_10 g17380(new_n19728, new_n19729);
or_5   g17381(new_n9494, n23529, new_n19730);
or_5   g17382(new_n9530, new_n9496, new_n19731);
and_5  g17383(new_n19731, new_n19730, new_n19732);
or_5   g17384(new_n19732, new_n19729, new_n19733);
and_5  g17385(new_n19733, new_n19727, new_n19734);
or_5   g17386(new_n19734, new_n19726, new_n19735);
and_5  g17387(new_n19735, new_n19724, new_n19736_1);
nor_5  g17388(new_n19736_1, new_n19723, new_n19737);
nor_5  g17389(new_n19737, new_n19721, new_n19738);
nand_5 g17390(new_n19738, new_n10335, new_n19739);
nand_5 g17391(new_n14396, new_n17646, new_n19740);
xor_4  g17392(new_n14396, n3582, new_n19741);
nand_5 g17393(new_n14399, new_n7782, new_n19742);
xor_4  g17394(new_n14399, n2145, new_n19743);
nand_5 g17395(new_n14401, new_n7785, new_n19744);
xor_4  g17396(new_n14401, new_n7785, new_n19745);
or_5   g17397(new_n9555, new_n7789, new_n19746);
or_5   g17398(new_n9588, new_n9557_1, new_n19747);
and_5  g17399(new_n19747, new_n19746, new_n19748);
nand_5 g17400(new_n19748, new_n19745, new_n19749_1);
and_5  g17401(new_n19749_1, new_n19744, new_n19750);
or_5   g17402(new_n19750, new_n19743, new_n19751);
and_5  g17403(new_n19751, new_n19742, new_n19752);
or_5   g17404(new_n19752, new_n19741, new_n19753);
and_5  g17405(new_n19753, new_n19740, new_n19754);
and_5  g17406(new_n19754, new_n14443, new_n19755);
not_10 g17407(new_n19755, new_n19756_1);
xor_4  g17408(new_n19756_1, new_n19739, new_n19757);
xor_4  g17409(new_n19738, new_n10335, new_n19758);
not_10 g17410(new_n19758, new_n19759);
xor_4  g17411(new_n19754, new_n14443, new_n19760);
and_5  g17412(new_n19760, new_n19759, new_n19761);
xor_4  g17413(new_n19760, new_n19759, new_n19762);
not_10 g17414(new_n19762, new_n19763);
xor_4  g17415(new_n19736_1, new_n19723, new_n19764);
not_10 g17416(new_n19764, new_n19765);
xor_4  g17417(new_n19752, new_n19741, new_n19766);
nor_5  g17418(new_n19766, new_n19765, new_n19767_1);
not_10 g17419(new_n19767_1, new_n19768);
xor_4  g17420(new_n19766, new_n19765, new_n19769);
xor_4  g17421(new_n19734, new_n19726, new_n19770_1);
not_10 g17422(new_n19770_1, new_n19771);
xor_4  g17423(new_n19750, new_n19743, new_n19772);
nor_5  g17424(new_n19772, new_n19771, new_n19773);
not_10 g17425(new_n19773, new_n19774);
xor_4  g17426(new_n19772, new_n19771, new_n19775);
xor_4  g17427(new_n19732, new_n19729, new_n19776);
not_10 g17428(new_n19776, new_n19777);
xor_4  g17429(new_n19748, new_n19745, new_n19778);
nor_5  g17430(new_n19778, new_n19777, new_n19779);
not_10 g17431(new_n19779, new_n19780_1);
xor_4  g17432(new_n19778, new_n19777, new_n19781);
and_5  g17433(new_n9589, new_n9531, new_n19782);
nor_5  g17434(new_n9631, new_n9591, new_n19783);
nor_5  g17435(new_n19783, new_n19782, new_n19784);
not_10 g17436(new_n19784, new_n19785);
and_5  g17437(new_n19785, new_n19781, new_n19786);
not_10 g17438(new_n19786, new_n19787);
and_5  g17439(new_n19787, new_n19780_1, new_n19788);
not_10 g17440(new_n19788, new_n19789_1);
and_5  g17441(new_n19789_1, new_n19775, new_n19790);
not_10 g17442(new_n19790, new_n19791);
and_5  g17443(new_n19791, new_n19774, new_n19792_1);
not_10 g17444(new_n19792_1, new_n19793);
and_5  g17445(new_n19793, new_n19769, new_n19794);
not_10 g17446(new_n19794, new_n19795);
and_5  g17447(new_n19795, new_n19768, new_n19796);
nor_5  g17448(new_n19796, new_n19763, new_n19797);
nor_5  g17449(new_n19797, new_n19761, new_n19798_1);
xnor_4 g17450(new_n19798_1, new_n19757, n6022);
xnor_4 g17451(new_n19416, new_n19399, n6031);
and_5  g17452(new_n16927, new_n11171, new_n19801);
xor_4  g17453(new_n19801, new_n7250, new_n19802);
xor_4  g17454(new_n19802, n12507, new_n19803_1);
nor_5  g17455(new_n16928, n15077, new_n19804);
nor_5  g17456(new_n16965, new_n16929, new_n19805);
nor_5  g17457(new_n19805, new_n19804, new_n19806);
not_10 g17458(new_n19806, new_n19807);
xor_4  g17459(new_n19807, new_n19803_1, new_n19808);
xor_4  g17460(new_n19808, new_n5653, new_n19809);
nand_5 g17461(new_n16966, new_n5592, new_n19810);
nand_5 g17462(new_n17006_1, new_n16967, new_n19811);
and_5  g17463(new_n19811, new_n19810, new_n19812);
xor_4  g17464(new_n19812, new_n19809, new_n19813);
xor_4  g17465(new_n19813, new_n8277, new_n19814);
not_10 g17466(new_n19814, new_n19815);
nand_5 g17467(new_n17007, new_n8279, new_n19816);
or_5   g17468(new_n17053, new_n17009, new_n19817);
and_5  g17469(new_n19817, new_n19816, new_n19818);
xnor_4 g17470(new_n19818, new_n19815, n6044);
and_5  g17471(new_n9353, new_n9307, new_n19820);
nor_5  g17472(new_n9407, new_n9354, new_n19821);
nor_5  g17473(new_n19821, new_n19820, new_n19822);
and_5  g17474(new_n9306, new_n9291, new_n19823);
xor_4  g17475(new_n18380, new_n19823, new_n19824);
xor_4  g17476(new_n19824, new_n19822, new_n19825);
nor_5  g17477(new_n19825, new_n4527, new_n19826);
xnor_4 g17478(new_n19825, new_n4528, new_n19827);
nor_5  g17479(new_n9408, new_n4538, new_n19828);
not_10 g17480(new_n19828, new_n19829);
not_10 g17481(new_n9460_1, new_n19830);
and_5  g17482(new_n19830, new_n9409, new_n19831);
not_10 g17483(new_n19831, new_n19832);
and_5  g17484(new_n19832, new_n19829, new_n19833);
not_10 g17485(new_n19833, new_n19834);
and_5  g17486(new_n19834, new_n19827, new_n19835);
nor_5  g17487(new_n19835, new_n19826, new_n19836);
nor_5  g17488(new_n18380, new_n19823, new_n19837);
and_5  g17489(new_n19837, new_n19822, new_n19838);
nand_5 g17490(new_n19838, new_n18744, new_n19839);
nor_5  g17491(new_n19839, new_n19836, new_n19840);
nor_5  g17492(new_n19838, new_n18744, new_n19841);
and_5  g17493(new_n19841, new_n19836, new_n19842);
or_5   g17494(new_n19842, new_n19840, n6046);
xnor_4 g17495(n17077, n7437, new_n19844);
not_10 g17496(new_n19844, new_n19845);
or_5   g17497(n26510, new_n12052, new_n19846);
xnor_4 g17498(n26510, n20700, new_n19847);
not_10 g17499(new_n19847, new_n19848);
or_5   g17500(n23068, new_n12056, new_n19849);
or_5   g17501(new_n19505, new_n19485, new_n19850);
and_5  g17502(new_n19850, new_n19849, new_n19851);
or_5   g17503(new_n19851, new_n19848, new_n19852);
and_5  g17504(new_n19852, new_n19846, new_n19853);
xor_4  g17505(new_n19853, new_n19845, new_n19854);
xor_4  g17506(n21997, n18483, new_n19855);
nand_5 g17507(n25119, n21934, new_n19856);
or_5   g17508(n25119, n21934, new_n19857);
nor_5  g17509(n18901, n1163, new_n19858);
nor_5  g17510(new_n19465, new_n19453, new_n19859);
nor_5  g17511(new_n19859, new_n19858, new_n19860);
nand_5 g17512(new_n19860, new_n19857, new_n19861);
and_5  g17513(new_n19861, new_n19856, new_n19862);
xor_4  g17514(new_n19862, new_n19855, new_n19863);
xor_4  g17515(new_n19863, new_n7568, new_n19864);
xor_4  g17516(n25119, n21934, new_n19865);
xor_4  g17517(new_n19865, new_n19860, new_n19866);
or_5   g17518(new_n19866, new_n2426, new_n19867);
nor_5  g17519(new_n19466, new_n2453, new_n19868);
and_5  g17520(new_n19482, new_n19467_1, new_n19869);
nor_5  g17521(new_n19869, new_n19868, new_n19870);
xor_4  g17522(new_n19866, new_n2426, new_n19871);
nand_5 g17523(new_n19871, new_n19870, new_n19872);
and_5  g17524(new_n19872, new_n19867, new_n19873_1);
xor_4  g17525(new_n19873_1, new_n19864, new_n19874);
xor_4  g17526(new_n19874, new_n19854, new_n19875);
xor_4  g17527(new_n19851, new_n19847, new_n19876);
xor_4  g17528(new_n19871, new_n19870, new_n19877);
nor_5  g17529(new_n19877, new_n19876, new_n19878);
or_5   g17530(new_n19506, new_n19483, new_n19879);
nand_5 g17531(new_n19536, new_n19507, new_n19880);
and_5  g17532(new_n19880, new_n19879, new_n19881);
not_10 g17533(new_n19877, new_n19882);
xnor_4 g17534(new_n19882, new_n19876, new_n19883);
and_5  g17535(new_n19883, new_n19881, new_n19884);
nor_5  g17536(new_n19884, new_n19878, new_n19885);
xnor_4 g17537(new_n19885, new_n19875, n6084);
xor_4  g17538(new_n19621, new_n10438, n6160);
xnor_4 g17539(new_n19628, new_n19626, n6171);
not_10 g17540(n10275, new_n19889);
or_5   g17541(n22359, new_n19889, new_n19890);
not_10 g17542(new_n10108, new_n19891);
or_5   g17543(new_n15497, new_n19891, new_n19892);
and_5  g17544(new_n19892, new_n19890, new_n19893);
xnor_4 g17545(new_n19893, new_n10111_1, new_n19894);
xor_4  g17546(n26264, n21905, new_n19895);
or_5   g17547(n22918, new_n8102, new_n19896);
xor_4  g17548(n22918, n7841, new_n19897);
or_5   g17549(n25923, new_n8108, new_n19898);
xor_4  g17550(n25923, n16812, new_n19899);
or_5   g17551(new_n8114, n6790, new_n19900);
or_5   g17552(new_n18428, new_n18409_1, new_n19901);
and_5  g17553(new_n19901, new_n19900, new_n19902);
or_5   g17554(new_n19902, new_n19899, new_n19903);
and_5  g17555(new_n19903, new_n19898, new_n19904);
or_5   g17556(new_n19904, new_n19897, new_n19905_1);
and_5  g17557(new_n19905_1, new_n19896, new_n19906);
xor_4  g17558(new_n19906, new_n19895, new_n19907);
xor_4  g17559(new_n19907, new_n15822, new_n19908);
xor_4  g17560(new_n19904, new_n19897, new_n19909_1);
or_5   g17561(new_n19909_1, new_n15826, new_n19910);
xor_4  g17562(new_n19909_1, new_n15826, new_n19911_1);
xor_4  g17563(new_n19902, new_n19899, new_n19912);
nand_5 g17564(new_n19912, new_n15830, new_n19913);
xnor_4 g17565(new_n19912, new_n15830, new_n19914);
nand_5 g17566(new_n18429, new_n15833, new_n19915);
nand_5 g17567(new_n18455, new_n18430, new_n19916_1);
and_5  g17568(new_n19916_1, new_n19915, new_n19917);
or_5   g17569(new_n19917, new_n19914, new_n19918);
and_5  g17570(new_n19918, new_n19913, new_n19919);
nand_5 g17571(new_n19919, new_n19911_1, new_n19920);
and_5  g17572(new_n19920, new_n19910, new_n19921);
xor_4  g17573(new_n19921, new_n19908, new_n19922_1);
xor_4  g17574(new_n19922_1, new_n19894, new_n19923_1);
not_10 g17575(new_n19923_1, new_n19924);
xor_4  g17576(new_n19919, new_n19911_1, new_n19925);
not_10 g17577(new_n19925, new_n19926);
nor_5  g17578(new_n19926, new_n15498, new_n19927);
xor_4  g17579(new_n19926, new_n15498, new_n19928);
xor_4  g17580(new_n19917, new_n19914, new_n19929);
nor_5  g17581(new_n19929, new_n15501_1, new_n19930_1);
xor_4  g17582(new_n19929, new_n15501_1, new_n19931);
not_10 g17583(new_n19931, new_n19932);
nor_5  g17584(new_n18456, new_n15505, new_n19933);
nor_5  g17585(new_n18485, new_n18458, new_n19934);
nor_5  g17586(new_n19934, new_n19933, new_n19935);
nor_5  g17587(new_n19935, new_n19932, new_n19936);
nor_5  g17588(new_n19936, new_n19930_1, new_n19937);
not_10 g17589(new_n19937, new_n19938);
and_5  g17590(new_n19938, new_n19928, new_n19939);
nor_5  g17591(new_n19939, new_n19927, new_n19940);
xnor_4 g17592(new_n19940, new_n19924, n6183);
xor_4  g17593(n14702, n14345, new_n19942);
or_5   g17594(new_n9318_1, n2999, new_n19943);
xor_4  g17595(n11356, n2999, new_n19944);
or_5   g17596(new_n9321, n2547, new_n19945);
xnor_4 g17597(n3164, n2547, new_n19946);
or_5   g17598(n10611, new_n9297, new_n19947);
or_5   g17599(new_n14366, new_n14355, new_n19948);
and_5  g17600(new_n19948, new_n19947, new_n19949);
nand_5 g17601(new_n19949, new_n19946, new_n19950);
and_5  g17602(new_n19950, new_n19945, new_n19951);
or_5   g17603(new_n19951, new_n19944, new_n19952);
and_5  g17604(new_n19952, new_n19943, new_n19953);
xor_4  g17605(new_n19953, new_n19942, new_n19954);
xor_4  g17606(new_n19954, new_n9220_1, new_n19955);
xor_4  g17607(new_n19951, new_n19944, new_n19956);
or_5   g17608(new_n19956, new_n9226, new_n19957);
xor_4  g17609(new_n19956, new_n9226, new_n19958);
xor_4  g17610(new_n19949, new_n19946, new_n19959);
or_5   g17611(new_n19959, new_n9232, new_n19960);
xor_4  g17612(new_n19959, new_n9232, new_n19961);
nand_5 g17613(new_n14367, new_n9236, new_n19962);
nand_5 g17614(new_n14382, new_n14368, new_n19963);
nand_5 g17615(new_n19963, new_n19962, new_n19964);
nand_5 g17616(new_n19964, new_n19961, new_n19965);
nand_5 g17617(new_n19965, new_n19960, new_n19966);
nand_5 g17618(new_n19966, new_n19958, new_n19967);
and_5  g17619(new_n19967, new_n19957, new_n19968_1);
xor_4  g17620(new_n19968_1, new_n19955, n6189);
xor_4  g17621(n20036, n15167, new_n19970);
or_5   g17622(new_n12573, n11192, new_n19971);
or_5   g17623(n21095, new_n4122, new_n19972);
and_5  g17624(new_n4125, n8656, new_n19973);
nand_5 g17625(new_n19973, new_n19972, new_n19974);
and_5  g17626(new_n19974, new_n19971, new_n19975);
xnor_4 g17627(new_n19975, new_n19970, new_n19976);
xor_4  g17628(new_n19976, new_n18467_1, new_n19977);
not_10 g17629(new_n19977, new_n19978);
xnor_4 g17630(n9380, n8656, new_n19979);
nor_5  g17631(new_n19979, new_n15365, new_n19980);
xnor_4 g17632(n21095, n11192, new_n19981);
xnor_4 g17633(new_n19981, new_n19973, new_n19982);
nor_5  g17634(new_n19982, new_n19980, new_n19983);
xor_4  g17635(new_n19982, new_n19980, new_n19984);
and_5  g17636(new_n19984, new_n18475, new_n19985);
nor_5  g17637(new_n19985, new_n19983, new_n19986);
xnor_4 g17638(new_n19986, new_n19978, n6223);
xnor_4 g17639(new_n14380, new_n14372, n6233);
xor_4  g17640(new_n19121, new_n19114, n6245);
xnor_4 g17641(new_n10441, new_n10431, n6248);
xor_4  g17642(n21839, n16544, new_n19991);
or_5   g17643(n27089, new_n9146_1, new_n19992);
or_5   g17644(new_n19594, new_n19563, new_n19993);
and_5  g17645(new_n19993, new_n19992, new_n19994);
xor_4  g17646(new_n19994, new_n19991, new_n19995);
xor_4  g17647(new_n19995, new_n10393, new_n19996);
not_10 g17648(new_n19996, new_n19997);
nor_5  g17649(new_n19595, new_n10399, new_n19998);
and_5  g17650(new_n19643, new_n19596, new_n19999);
nor_5  g17651(new_n19999, new_n19998, new_n20000);
xnor_4 g17652(new_n20000, new_n19997, n6256);
xnor_4 g17653(new_n15226, new_n15203, n6271);
nor_5  g17654(new_n11167, n13549, new_n20003);
not_10 g17655(new_n10114, new_n20004_1);
not_10 g17656(n23493, new_n20005);
or_5   g17657(new_n20005, n8405, new_n20006);
not_10 g17658(new_n10111_1, new_n20007);
or_5   g17659(new_n19893, new_n20007, new_n20008);
and_5  g17660(new_n20008, new_n20006, new_n20009);
nor_5  g17661(new_n20009, new_n20004_1, new_n20010);
nor_5  g17662(new_n20010, new_n20003, new_n20011);
or_5   g17663(n13951, new_n11219, new_n20012);
xor_4  g17664(n13951, n2944, new_n20013_1);
or_5   g17665(n22793, new_n11220_1, new_n20014);
or_5   g17666(new_n15254, new_n15235, new_n20015);
and_5  g17667(new_n20015, new_n20014, new_n20016);
or_5   g17668(new_n20016, new_n20013_1, new_n20017_1);
and_5  g17669(new_n20017_1, new_n20012, new_n20018);
and_5  g17670(new_n20018, new_n20011, new_n20019);
xor_4  g17671(new_n20016, new_n20013_1, new_n20020);
xnor_4 g17672(new_n20009, new_n10114, new_n20021);
nor_5  g17673(new_n20021, new_n20020, new_n20022);
xor_4  g17674(new_n20021, new_n20020, new_n20023);
nand_5 g17675(new_n19894, new_n15255_1, new_n20024);
xor_4  g17676(new_n19894, new_n15255_1, new_n20025);
or_5   g17677(new_n15498, new_n15258_1, new_n20026);
or_5   g17678(new_n15520, new_n15500, new_n20027);
and_5  g17679(new_n20027, new_n20026, new_n20028);
nand_5 g17680(new_n20028, new_n20025, new_n20029);
and_5  g17681(new_n20029, new_n20024, new_n20030);
and_5  g17682(new_n20030, new_n20023, new_n20031);
or_5   g17683(new_n20031, new_n20022, new_n20032);
xor_4  g17684(new_n20018, new_n20011, new_n20033_1);
and_5  g17685(new_n20033_1, new_n20032, new_n20034);
nor_5  g17686(new_n20034, new_n20019, new_n20035);
and_5  g17687(n8827, new_n17883, new_n20036_1);
not_10 g17688(new_n20036_1, new_n20037);
xnor_4 g17689(n8827, n1881, new_n20038);
not_10 g17690(new_n20038, new_n20039);
or_5   g17691(new_n15151, n5834, new_n20040_1);
or_5   g17692(new_n19390, new_n19387, new_n20041);
and_5  g17693(new_n20041, new_n20040_1, new_n20042);
nor_5  g17694(new_n20042, new_n20039, new_n20043);
not_10 g17695(new_n20043, new_n20044);
and_5  g17696(new_n20044, new_n20037, new_n20045);
not_10 g17697(new_n20045, new_n20046);
xor_4  g17698(new_n20046, new_n20035, new_n20047);
xor_4  g17699(new_n20033_1, new_n20032, new_n20048);
and_5  g17700(new_n20048, new_n20046, new_n20049);
xnor_4 g17701(new_n20048, new_n20045, new_n20050);
xor_4  g17702(new_n20042, new_n20039, new_n20051);
not_10 g17703(new_n20051, new_n20052);
xor_4  g17704(new_n20030, new_n20023, new_n20053);
nor_5  g17705(new_n20053, new_n20052, new_n20054);
xor_4  g17706(new_n20028, new_n20025, new_n20055);
or_5   g17707(new_n20055, new_n19391, new_n20056);
xor_4  g17708(new_n20055, new_n19391, new_n20057);
not_10 g17709(new_n15521, new_n20058);
and_5  g17710(new_n15774, new_n20058, new_n20059);
and_5  g17711(new_n15797, new_n15775, new_n20060);
nor_5  g17712(new_n20060, new_n20059, new_n20061_1);
nand_5 g17713(new_n20061_1, new_n20057, new_n20062);
and_5  g17714(new_n20062, new_n20056, new_n20063);
xor_4  g17715(new_n20053, new_n20052, new_n20064);
and_5  g17716(new_n20064, new_n20063, new_n20065);
nor_5  g17717(new_n20065, new_n20054, new_n20066);
and_5  g17718(new_n20066, new_n20050, new_n20067);
nor_5  g17719(new_n20067, new_n20049, new_n20068);
xor_4  g17720(new_n20068, new_n20047, n6276);
xor_4  g17721(new_n19066, new_n19065, n6308);
xnor_4 g17722(new_n17148, new_n17134, n6311);
xnor_4 g17723(new_n16909, new_n16890, n6323);
and_5  g17724(new_n5965, new_n5922, new_n20073);
not_10 g17725(new_n20073, new_n20074);
nor_5  g17726(new_n6032, new_n5968, new_n20075);
not_10 g17727(new_n20075, new_n20076);
and_5  g17728(new_n20076, new_n20074, new_n20077_1);
and_5  g17729(new_n13717, new_n14096, new_n20078);
not_10 g17730(new_n20078, new_n20079);
nor_5  g17731(new_n20079, new_n20077_1, new_n20080);
nor_5  g17732(new_n13717, new_n14096, new_n20081);
and_5  g17733(new_n20081, new_n20077_1, new_n20082);
nor_5  g17734(new_n20082, new_n20080, new_n20083);
nor_5  g17735(new_n20083, new_n18242, new_n20084);
not_10 g17736(new_n18242, new_n20085);
xor_4  g17737(new_n20083, new_n20085, new_n20086_1);
xor_4  g17738(new_n13717, new_n14096, new_n20087);
xor_4  g17739(new_n20087, new_n20077_1, new_n20088);
nor_5  g17740(new_n20088, new_n18244, new_n20089);
xor_4  g17741(new_n20088, new_n18244, new_n20090);
and_5  g17742(new_n18249, new_n6034, new_n20091);
not_10 g17743(new_n6191, new_n20092);
and_5  g17744(new_n20092, new_n6127, new_n20093);
nor_5  g17745(new_n20093, new_n20091, new_n20094);
not_10 g17746(new_n20094, new_n20095);
and_5  g17747(new_n20095, new_n20090, new_n20096_1);
nor_5  g17748(new_n20096_1, new_n20089, new_n20097);
nor_5  g17749(new_n20097, new_n20086_1, new_n20098);
nor_5  g17750(new_n20098, new_n20084, new_n20099);
nor_5  g17751(new_n20099, new_n20080, n6330);
xnor_4 g17752(new_n8726, new_n8688, n6339);
xnor_4 g17753(new_n14347, new_n14318, n6354);
not_10 g17754(new_n17323, new_n20103_1);
nor_5  g17755(new_n3199, n7335, new_n20104);
nor_5  g17756(new_n3206, n5696, new_n20105);
xnor_4 g17757(new_n3206, n5696, new_n20106);
or_5   g17758(new_n3211, n13367, new_n20107);
xor_4  g17759(new_n3212, n13367, new_n20108);
or_5   g17760(new_n3216, n932, new_n20109);
xor_4  g17761(new_n3217, n932, new_n20110);
or_5   g17762(new_n3221, n6691, new_n20111);
xor_4  g17763(new_n3222, n6691, new_n20112);
or_5   g17764(new_n3226, n3260, new_n20113);
xor_4  g17765(new_n3227, n3260, new_n20114);
or_5   g17766(new_n3231, n20489, new_n20115);
nor_5  g17767(new_n3236, n2355, new_n20116);
xor_4  g17768(new_n3237, n2355, new_n20117);
or_5   g17769(new_n3247, n11121, new_n20118);
nand_5 g17770(n16217, n12315, new_n20119);
xor_4  g17771(new_n3247, n11121, new_n20120);
nand_5 g17772(new_n20120, new_n20119, new_n20121);
and_5  g17773(new_n20121, new_n20118, new_n20122);
nor_5  g17774(new_n20122, new_n20117, new_n20123);
or_5   g17775(new_n20123, new_n20116, new_n20124);
xnor_4 g17776(new_n3232, n20489, new_n20125);
nand_5 g17777(new_n20125, new_n20124, new_n20126_1);
and_5  g17778(new_n20126_1, new_n20115, new_n20127);
or_5   g17779(new_n20127, new_n20114, new_n20128);
and_5  g17780(new_n20128, new_n20113, new_n20129);
or_5   g17781(new_n20129, new_n20112, new_n20130);
and_5  g17782(new_n20130, new_n20111, new_n20131);
or_5   g17783(new_n20131, new_n20110, new_n20132);
and_5  g17784(new_n20132, new_n20109, new_n20133);
or_5   g17785(new_n20133, new_n20108, new_n20134);
and_5  g17786(new_n20134, new_n20107, new_n20135);
nor_5  g17787(new_n20135, new_n20106, new_n20136);
or_5   g17788(new_n20136, new_n20105, new_n20137);
or_5   g17789(new_n20137, new_n20104, new_n20138_1);
nand_5 g17790(new_n3199, n7335, new_n20139);
and_5  g17791(new_n20139, new_n3204, new_n20140);
and_5  g17792(new_n20140, new_n20138_1, new_n20141);
and_5  g17793(new_n20141, new_n20103_1, new_n20142);
nor_5  g17794(new_n20141, new_n17371, new_n20143);
xor_4  g17795(new_n20141, new_n17371, new_n20144);
not_10 g17796(new_n20144, new_n20145);
xnor_4 g17797(new_n3200, n7335, new_n20146);
xor_4  g17798(new_n20146, new_n20137, new_n20147);
and_5  g17799(new_n20147, new_n17376, new_n20148);
xor_4  g17800(new_n20147, new_n17376, new_n20149_1);
xor_4  g17801(new_n20135, new_n20106, new_n20150);
and_5  g17802(new_n20150, new_n17382, new_n20151_1);
xor_4  g17803(new_n20150, new_n17382, new_n20152);
xor_4  g17804(new_n20133, new_n20108, new_n20153);
and_5  g17805(new_n20153, new_n17386, new_n20154);
xor_4  g17806(new_n20153, new_n17386, new_n20155);
xor_4  g17807(new_n20131, new_n20110, new_n20156);
and_5  g17808(new_n20156, new_n17390, new_n20157);
xor_4  g17809(new_n20156, new_n17390, new_n20158);
xor_4  g17810(new_n20129, new_n20112, new_n20159);
and_5  g17811(new_n20159, new_n17394, new_n20160);
xor_4  g17812(new_n20159, new_n17394, new_n20161);
xor_4  g17813(new_n20127, new_n20114, new_n20162);
and_5  g17814(new_n20162, new_n17398, new_n20163);
xor_4  g17815(new_n20162, new_n17398, new_n20164);
xor_4  g17816(new_n20125, new_n20124, new_n20165);
and_5  g17817(new_n20165, new_n17402, new_n20166);
xor_4  g17818(new_n20165, new_n17402, new_n20167);
xor_4  g17819(new_n20122, new_n20117, new_n20168);
nor_5  g17820(new_n20168, new_n17407, new_n20169_1);
xor_4  g17821(new_n20168, new_n17407, new_n20170);
or_5   g17822(new_n20120, new_n17411, new_n20171);
xor_4  g17823(new_n20120, new_n20119, new_n20172);
nor_5  g17824(new_n20172, new_n17410, new_n20173);
xor_4  g17825(n16217, n12315, new_n20174);
and_5  g17826(new_n20174, new_n17416, new_n20175);
or_5   g17827(new_n20175, new_n20173, new_n20176);
and_5  g17828(new_n20176, new_n20171, new_n20177);
and_5  g17829(new_n20177, new_n20170, new_n20178);
nor_5  g17830(new_n20178, new_n20169_1, new_n20179_1);
and_5  g17831(new_n20179_1, new_n20167, new_n20180);
nor_5  g17832(new_n20180, new_n20166, new_n20181);
not_10 g17833(new_n20181, new_n20182);
and_5  g17834(new_n20182, new_n20164, new_n20183);
nor_5  g17835(new_n20183, new_n20163, new_n20184);
not_10 g17836(new_n20184, new_n20185);
and_5  g17837(new_n20185, new_n20161, new_n20186);
nor_5  g17838(new_n20186, new_n20160, new_n20187_1);
not_10 g17839(new_n20187_1, new_n20188);
and_5  g17840(new_n20188, new_n20158, new_n20189);
nor_5  g17841(new_n20189, new_n20157, new_n20190);
not_10 g17842(new_n20190, new_n20191);
and_5  g17843(new_n20191, new_n20155, new_n20192);
nor_5  g17844(new_n20192, new_n20154, new_n20193);
not_10 g17845(new_n20193, new_n20194);
and_5  g17846(new_n20194, new_n20152, new_n20195);
nor_5  g17847(new_n20195, new_n20151_1, new_n20196);
not_10 g17848(new_n20196, new_n20197);
and_5  g17849(new_n20197, new_n20149_1, new_n20198);
nor_5  g17850(new_n20198, new_n20148, new_n20199);
nor_5  g17851(new_n20199, new_n20145, new_n20200);
nor_5  g17852(new_n20200, new_n20143, new_n20201);
or_5   g17853(new_n20201, new_n20142, new_n20202);
nor_5  g17854(new_n20141, new_n20103_1, new_n20203);
or_5   g17855(new_n20203, new_n20200, new_n20204);
and_5  g17856(new_n20204, new_n20202, n6375);
xnor_4 g17857(new_n19248, new_n19232, n6383);
xor_4  g17858(new_n14750, new_n14714, n6407);
xnor_4 g17859(new_n8715, new_n8714, n6431);
xnor_4 g17860(new_n16740, new_n16737, n6437);
xnor_4 g17861(new_n4160, new_n4159, n6457);
xnor_4 g17862(new_n12533, new_n12496, n6465);
nand_5 g17863(new_n17648, n3740, new_n20212);
nand_5 g17864(new_n17647, new_n17646, new_n20213_1);
nor_5  g17865(new_n17648, n3740, new_n20214);
or_5   g17866(new_n17653, new_n20214, new_n20215);
and_5  g17867(new_n20215, new_n20213_1, new_n20216);
and_5  g17868(new_n20216, new_n20212, new_n20217);
xor_4  g17869(new_n20217, new_n8478, new_n20218);
or_5   g17870(new_n18692, new_n3471, new_n20219);
xnor_4 g17871(new_n17654, new_n3471, new_n20220);
nand_5 g17872(new_n14628, new_n3475, new_n20221);
nand_5 g17873(new_n14664, new_n14629, new_n20222);
and_5  g17874(new_n20222, new_n20221, new_n20223);
nand_5 g17875(new_n20223, new_n20220, new_n20224);
and_5  g17876(new_n20224, new_n20219, new_n20225);
xor_4  g17877(new_n20225, new_n20218, new_n20226);
nor_5  g17878(new_n3600, n2743, new_n20227);
and_5  g17879(new_n3603, n7026, new_n20228);
nor_5  g17880(new_n3603, n7026, new_n20229);
nor_5  g17881(new_n14702_1, new_n20229, new_n20230);
nor_5  g17882(new_n20230, new_n20228, new_n20231);
nor_5  g17883(new_n20231, new_n20227, new_n20232);
and_5  g17884(new_n3599, new_n3584, new_n20233);
and_5  g17885(new_n3600, n2743, new_n20234);
nor_5  g17886(new_n20234, new_n20233, new_n20235_1);
not_10 g17887(new_n20235_1, new_n20236);
nor_5  g17888(new_n20236, new_n20232, new_n20237);
not_10 g17889(new_n20237, new_n20238);
xor_4  g17890(new_n20238, new_n20226, new_n20239);
xor_4  g17891(new_n20223, new_n20220, new_n20240);
not_10 g17892(n2743, new_n20241);
xor_4  g17893(new_n3600, new_n20241, new_n20242);
xor_4  g17894(new_n20242, new_n20231, new_n20243);
nor_5  g17895(new_n20243, new_n20240, new_n20244);
not_10 g17896(new_n20240, new_n20245);
xnor_4 g17897(new_n20243, new_n20245, new_n20246);
nor_5  g17898(new_n14703, new_n14666, new_n20247);
and_5  g17899(new_n14754, new_n14704_1, new_n20248);
nor_5  g17900(new_n20248, new_n20247, new_n20249);
not_10 g17901(new_n20249, new_n20250_1);
and_5  g17902(new_n20250_1, new_n20246, new_n20251);
nor_5  g17903(new_n20251, new_n20244, new_n20252);
xor_4  g17904(new_n20252, new_n20239, n6470);
xor_4  g17905(new_n11749_1, new_n11724_1, n6476);
xnor_4 g17906(new_n18736, new_n18727, n6506);
not_10 g17907(new_n9574, new_n20256);
and_5  g17908(new_n20256, new_n9572, new_n20257);
and_5  g17909(new_n20257, new_n9570, new_n20258);
and_5  g17910(new_n20258, new_n9566, new_n20259_1);
and_5  g17911(new_n20259_1, new_n9562, new_n20260);
and_5  g17912(new_n20260, new_n9558_1, new_n20261);
and_5  g17913(new_n20261, new_n9555, new_n20262);
and_5  g17914(new_n20262, new_n14401, new_n20263);
xor_4  g17915(new_n20263, new_n14399, new_n20264);
xor_4  g17916(new_n20264, new_n10343, new_n20265);
xor_4  g17917(new_n20262, new_n14401, new_n20266);
or_5   g17918(new_n20266, new_n10349, new_n20267);
xor_4  g17919(new_n20266, new_n10348, new_n20268);
xor_4  g17920(new_n20261, new_n9555, new_n20269);
or_5   g17921(new_n20269, new_n9494, new_n20270);
xor_4  g17922(new_n20269, new_n9493_1, new_n20271);
xor_4  g17923(new_n20260, new_n9558_1, new_n20272);
or_5   g17924(new_n20272, new_n9498, new_n20273);
xor_4  g17925(new_n20272, new_n9497, new_n20274);
xor_4  g17926(new_n20259_1, new_n9562, new_n20275);
or_5   g17927(new_n20275, new_n9503, new_n20276);
xor_4  g17928(new_n20275, new_n9502, new_n20277);
xor_4  g17929(new_n20258, new_n9566, new_n20278);
or_5   g17930(new_n20278, new_n9508_1, new_n20279_1);
xor_4  g17931(new_n20257, new_n9570, new_n20280);
nor_5  g17932(new_n20280, new_n9512_1, new_n20281);
xor_4  g17933(new_n20280, new_n9511, new_n20282);
and_5  g17934(new_n9574, new_n9517, new_n20283);
or_5   g17935(new_n20283, new_n9515, new_n20284);
and_5  g17936(new_n9574, new_n9544, new_n20285);
or_5   g17937(new_n20285, new_n20257, new_n20286);
nand_5 g17938(new_n20283, new_n9482, new_n20287_1);
and_5  g17939(new_n20287_1, new_n20284, new_n20288);
nand_5 g17940(new_n20288, new_n20286, new_n20289);
and_5  g17941(new_n20289, new_n20284, new_n20290);
nor_5  g17942(new_n20290, new_n20282, new_n20291);
or_5   g17943(new_n20291, new_n20281, new_n20292);
xnor_4 g17944(new_n20278, new_n9507_1, new_n20293);
nand_5 g17945(new_n20293, new_n20292, new_n20294);
and_5  g17946(new_n20294, new_n20279_1, new_n20295);
or_5   g17947(new_n20295, new_n20277, new_n20296);
and_5  g17948(new_n20296, new_n20276, new_n20297);
or_5   g17949(new_n20297, new_n20274, new_n20298);
and_5  g17950(new_n20298, new_n20273, new_n20299);
or_5   g17951(new_n20299, new_n20271, new_n20300);
and_5  g17952(new_n20300, new_n20270, new_n20301_1);
or_5   g17953(new_n20301_1, new_n20268, new_n20302);
and_5  g17954(new_n20302, new_n20267, new_n20303);
xor_4  g17955(new_n20303, new_n20265, new_n20304);
xor_4  g17956(new_n20304, new_n16966, new_n20305);
xor_4  g17957(new_n20301_1, new_n20268, new_n20306);
nand_5 g17958(new_n20306, new_n16968_1, new_n20307);
xor_4  g17959(new_n20306, new_n16968_1, new_n20308);
not_10 g17960(new_n20308, new_n20309);
xor_4  g17961(new_n20299, new_n20271, new_n20310);
nand_5 g17962(new_n20310, new_n16973, new_n20311);
xnor_4 g17963(new_n20310, new_n16972, new_n20312);
not_10 g17964(new_n20312, new_n20313);
xor_4  g17965(new_n20297, new_n20274, new_n20314);
nand_5 g17966(new_n20314, new_n16976, new_n20315);
xor_4  g17967(new_n20314, new_n16976, new_n20316);
xor_4  g17968(new_n20295, new_n20277, new_n20317);
or_5   g17969(new_n20317, new_n16979, new_n20318);
xor_4  g17970(new_n20293, new_n20292, new_n20319);
nor_5  g17971(new_n20319, new_n16982, new_n20320);
xnor_4 g17972(new_n20319, new_n16982, new_n20321);
xor_4  g17973(new_n20290, new_n20282, new_n20322);
or_5   g17974(new_n20322, new_n16985, new_n20323);
xnor_4 g17975(new_n20322, new_n16985, new_n20324);
xor_4  g17976(new_n20288, new_n20286, new_n20325);
or_5   g17977(new_n20325, new_n16988_1, new_n20326);
xor_4  g17978(new_n9574, new_n9517, new_n20327);
and_5  g17979(new_n20327, new_n16990, new_n20328);
xor_4  g17980(new_n20325, new_n16988_1, new_n20329);
nand_5 g17981(new_n20329, new_n20328, new_n20330_1);
and_5  g17982(new_n20330_1, new_n20326, new_n20331);
or_5   g17983(new_n20331, new_n20324, new_n20332);
and_5  g17984(new_n20332, new_n20323, new_n20333_1);
nor_5  g17985(new_n20333_1, new_n20321, new_n20334);
or_5   g17986(new_n20334, new_n20320, new_n20335);
xor_4  g17987(new_n20317, new_n16979, new_n20336);
nand_5 g17988(new_n20336, new_n20335, new_n20337);
and_5  g17989(new_n20337, new_n20318, new_n20338);
nand_5 g17990(new_n20338, new_n20316, new_n20339);
and_5  g17991(new_n20339, new_n20315, new_n20340);
or_5   g17992(new_n20340, new_n20313, new_n20341);
and_5  g17993(new_n20341, new_n20311, new_n20342);
or_5   g17994(new_n20342, new_n20309, new_n20343);
and_5  g17995(new_n20343, new_n20307, new_n20344);
xor_4  g17996(new_n20344, new_n20305, n6514);
not_10 g17997(new_n11614, new_n20346);
nor_5  g17998(new_n11711, new_n20346, new_n20347);
nor_5  g17999(new_n11754, new_n11713, new_n20348);
nor_5  g18000(new_n20348, new_n20347, new_n20349_1);
xor_4  g18001(new_n11669, new_n12188, new_n20350);
nand_5 g18002(new_n20350, new_n11710_1, new_n20351);
and_5  g18003(new_n11670, new_n11658, new_n20352);
nor_5  g18004(new_n11710_1, new_n20352, new_n20353);
not_10 g18005(new_n20353, new_n20354);
or_5   g18006(new_n20354, new_n20350, new_n20355_1);
nand_5 g18007(new_n20355_1, new_n20351, new_n20356);
xnor_4 g18008(new_n20356, new_n20349_1, n6542);
xnor_4 g18009(new_n15676, new_n15662_1, n6558);
xor_4  g18010(new_n18225, new_n18223, n6560);
xor_4  g18011(new_n6306, n10405, new_n20360);
nand_5 g18012(new_n6309, n11302, new_n20361);
xor_4  g18013(new_n6309, n11302, new_n20362);
nand_5 g18014(new_n6312, new_n5513, new_n20363);
nand_5 g18015(new_n6314, n6773, new_n20364);
xor_4  g18016(new_n6312, new_n5513, new_n20365);
nand_5 g18017(new_n20365, new_n20364, new_n20366_1);
and_5  g18018(new_n20366_1, new_n20363, new_n20367);
nand_5 g18019(new_n20367, new_n20362, new_n20368);
and_5  g18020(new_n20368, new_n20361, new_n20369);
xor_4  g18021(new_n20369, new_n20360, new_n20370);
xnor_4 g18022(new_n20370, new_n9914, new_n20371);
not_10 g18023(new_n20371, new_n20372);
xor_4  g18024(new_n20367, new_n20362, new_n20373);
nor_5  g18025(new_n20373, new_n9921, new_n20374);
xnor_4 g18026(new_n20373, new_n9919_1, new_n20375);
not_10 g18027(new_n20375, new_n20376);
xor_4  g18028(new_n20365, new_n20364, new_n20377);
and_5  g18029(new_n20377, new_n9930, new_n20378);
not_10 g18030(new_n20378, new_n20379);
nor_5  g18031(new_n18256, new_n9927, new_n20380);
xnor_4 g18032(new_n20377, new_n9924, new_n20381);
and_5  g18033(new_n20381, new_n20380, new_n20382);
not_10 g18034(new_n20382, new_n20383);
and_5  g18035(new_n20383, new_n20379, new_n20384);
nor_5  g18036(new_n20384, new_n20376, new_n20385_1);
nor_5  g18037(new_n20385_1, new_n20374, new_n20386);
xnor_4 g18038(new_n20386, new_n20372, n6567);
and_5  g18039(new_n13943, new_n8226, new_n20388_1);
and_5  g18040(new_n20388_1, new_n8222, new_n20389);
and_5  g18041(new_n20389, new_n8218, new_n20390);
and_5  g18042(new_n20390, new_n8214, new_n20391);
xor_4  g18043(new_n20391, new_n8210, new_n20392);
xor_4  g18044(new_n20392, new_n4468, new_n20393);
xor_4  g18045(new_n20390, new_n8214, new_n20394);
or_5   g18046(new_n20394, new_n4474, new_n20395);
xor_4  g18047(new_n20394, new_n4474, new_n20396);
not_10 g18048(new_n20396, new_n20397);
xor_4  g18049(new_n20389, new_n8218, new_n20398);
or_5   g18050(new_n20398, new_n4480, new_n20399);
xnor_4 g18051(new_n20398, new_n4479, new_n20400);
not_10 g18052(new_n20400, new_n20401);
xor_4  g18053(new_n20388_1, new_n8222, new_n20402_1);
not_10 g18054(new_n20402_1, new_n20403_1);
nand_5 g18055(new_n20403_1, new_n4486, new_n20404);
xnor_4 g18056(new_n20402_1, new_n4486, new_n20405);
not_10 g18057(new_n20405, new_n20406);
or_5   g18058(new_n13944, new_n3971_1, new_n20407);
nand_5 g18059(new_n13968, new_n13947, new_n20408);
nand_5 g18060(new_n20408, new_n13945, new_n20409_1);
and_5  g18061(new_n20409_1, new_n20407, new_n20410);
or_5   g18062(new_n20410, new_n20406, new_n20411_1);
and_5  g18063(new_n20411_1, new_n20404, new_n20412);
or_5   g18064(new_n20412, new_n20401, new_n20413);
and_5  g18065(new_n20413, new_n20399, new_n20414);
or_5   g18066(new_n20414, new_n20397, new_n20415);
and_5  g18067(new_n20415, new_n20395, new_n20416);
xor_4  g18068(new_n20416, new_n20393, new_n20417);
not_10 g18069(new_n20417, new_n20418);
xor_4  g18070(new_n8208, n23272, new_n20419);
or_5   g18071(new_n8212, n11481, new_n20420);
xor_4  g18072(new_n8212, new_n18901_1, new_n20421);
or_5   g18073(new_n8216, n16439, new_n20422);
xor_4  g18074(new_n8216, new_n4360, new_n20423);
or_5   g18075(new_n8220, n15241, new_n20424_1);
nand_5 g18076(new_n8224, n7678, new_n20425);
nand_5 g18077(new_n13990, new_n13972, new_n20426);
and_5  g18078(new_n20426, new_n20425, new_n20427);
xor_4  g18079(new_n8220, n15241, new_n20428);
nand_5 g18080(new_n20428, new_n20427, new_n20429_1);
and_5  g18081(new_n20429_1, new_n20424_1, new_n20430);
or_5   g18082(new_n20430, new_n20423, new_n20431);
and_5  g18083(new_n20431, new_n20422, new_n20432);
or_5   g18084(new_n20432, new_n20421, new_n20433);
and_5  g18085(new_n20433, new_n20420, new_n20434);
xor_4  g18086(new_n20434, new_n20419, new_n20435);
xnor_4 g18087(new_n20435, new_n20418, new_n20436_1);
xor_4  g18088(new_n20414, new_n20397, new_n20437);
xor_4  g18089(new_n20432, new_n20421, new_n20438);
nand_5 g18090(new_n20438, new_n20437, new_n20439);
not_10 g18091(new_n20437, new_n20440);
xnor_4 g18092(new_n20438, new_n20440, new_n20441_1);
xnor_4 g18093(new_n20412, new_n20400, new_n20442);
xor_4  g18094(new_n20430, new_n20423, new_n20443);
nand_5 g18095(new_n20443, new_n20442, new_n20444);
not_10 g18096(new_n20442, new_n20445_1);
xnor_4 g18097(new_n20443, new_n20445_1, new_n20446);
xnor_4 g18098(new_n20410, new_n20405, new_n20447);
xor_4  g18099(new_n20428, new_n20427, new_n20448);
nand_5 g18100(new_n20448, new_n20447, new_n20449);
not_10 g18101(new_n20447, new_n20450_1);
xnor_4 g18102(new_n20448, new_n20450_1, new_n20451);
or_5   g18103(new_n13991, new_n13971, new_n20452);
nand_5 g18104(new_n14023, new_n13992, new_n20453);
nand_5 g18105(new_n20453, new_n20452, new_n20454);
nand_5 g18106(new_n20454, new_n20451, new_n20455_1);
nand_5 g18107(new_n20455_1, new_n20449, new_n20456);
nand_5 g18108(new_n20456, new_n20446, new_n20457);
nand_5 g18109(new_n20457, new_n20444, new_n20458);
nand_5 g18110(new_n20458, new_n20441_1, new_n20459);
nand_5 g18111(new_n20459, new_n20439, new_n20460);
xnor_4 g18112(new_n20460, new_n20436_1, n6576);
xnor_4 g18113(new_n20172, new_n17411, new_n20462);
xor_4  g18114(new_n20462, new_n20175, n6587);
xor_4  g18115(new_n19080, new_n19027, n6612);
nor_5  g18116(new_n17706, new_n10964, new_n20465);
xnor_4 g18117(new_n17706, new_n10964, new_n20466);
or_5   g18118(new_n17708, new_n10957, new_n20467);
xnor_4 g18119(new_n17708, new_n10957, new_n20468);
or_5   g18120(new_n17712, new_n10950, new_n20469);
xor_4  g18121(new_n17712, new_n10971, new_n20470_1);
or_5   g18122(new_n17716, new_n10943_1, new_n20471);
xor_4  g18123(new_n17716, new_n10975, new_n20472);
or_5   g18124(new_n17720, new_n10936, new_n20473);
xor_4  g18125(new_n17720, new_n10979, new_n20474);
or_5   g18126(new_n17722, new_n10929, new_n20475);
xnor_4 g18127(new_n17722, new_n10929, new_n20476);
or_5   g18128(new_n15369, new_n10923, new_n20477);
xor_4  g18129(new_n15369, new_n10923, new_n20478_1);
nand_5 g18130(new_n15371, new_n10917, new_n20479);
and_5  g18131(new_n10906, new_n9333, new_n20480);
nand_5 g18132(new_n20480, new_n9330, new_n20481);
not_10 g18133(new_n15374, new_n20482);
or_5   g18134(new_n20480, new_n20482, new_n20483);
and_5  g18135(new_n20483, new_n20481, new_n20484);
nand_5 g18136(new_n20484, new_n10910, new_n20485);
and_5  g18137(new_n20485, new_n20481, new_n20486);
xor_4  g18138(new_n15371, new_n10917, new_n20487);
nand_5 g18139(new_n20487, new_n20486, new_n20488);
and_5  g18140(new_n20488, new_n20479, new_n20489_1);
nand_5 g18141(new_n20489_1, new_n20478_1, new_n20490_1);
and_5  g18142(new_n20490_1, new_n20477, new_n20491);
or_5   g18143(new_n20491, new_n20476, new_n20492);
and_5  g18144(new_n20492, new_n20475, new_n20493);
or_5   g18145(new_n20493, new_n20474, new_n20494);
and_5  g18146(new_n20494, new_n20473, new_n20495_1);
or_5   g18147(new_n20495_1, new_n20472, new_n20496);
and_5  g18148(new_n20496, new_n20471, new_n20497);
or_5   g18149(new_n20497, new_n20470_1, new_n20498);
and_5  g18150(new_n20498, new_n20469, new_n20499);
or_5   g18151(new_n20499, new_n20468, new_n20500);
and_5  g18152(new_n20500, new_n20467, new_n20501);
nor_5  g18153(new_n20501, new_n20466, new_n20502);
or_5   g18154(new_n20502, new_n20465, new_n20503);
and_5  g18155(new_n17705, new_n17699, new_n20504);
not_10 g18156(new_n20504, new_n20505);
or_5   g18157(new_n17902, new_n20505, new_n20506);
nor_5  g18158(new_n20506, new_n20503, new_n20507);
and_5  g18159(new_n17902, new_n20505, new_n20508);
and_5  g18160(new_n20508, new_n20503, new_n20509);
nor_5  g18161(new_n20509, new_n20507, new_n20510);
xor_4  g18162(new_n17902, new_n20505, new_n20511);
xor_4  g18163(new_n20511, new_n20503, new_n20512);
nor_5  g18164(new_n20512, new_n19760, new_n20513);
xor_4  g18165(new_n20512, new_n19760, new_n20514);
xor_4  g18166(new_n20501, new_n20466, new_n20515_1);
and_5  g18167(new_n20515_1, new_n19766, new_n20516);
xor_4  g18168(new_n20515_1, new_n19766, new_n20517);
xor_4  g18169(new_n20499, new_n20468, new_n20518);
and_5  g18170(new_n20518, new_n19772, new_n20519);
xor_4  g18171(new_n20518, new_n19772, new_n20520);
xor_4  g18172(new_n20497, new_n20470_1, new_n20521);
and_5  g18173(new_n20521, new_n19778, new_n20522);
xor_4  g18174(new_n20521, new_n19778, new_n20523);
not_10 g18175(new_n9589, new_n20524);
xor_4  g18176(new_n20495_1, new_n20472, new_n20525);
and_5  g18177(new_n20525, new_n20524, new_n20526);
xnor_4 g18178(new_n20525, new_n9589, new_n20527);
not_10 g18179(new_n9593, new_n20528);
xor_4  g18180(new_n20493, new_n20474, new_n20529);
and_5  g18181(new_n20529, new_n20528, new_n20530);
xnor_4 g18182(new_n20529, new_n9593, new_n20531);
not_10 g18183(new_n9598_1, new_n20532);
xor_4  g18184(new_n20491, new_n20476, new_n20533_1);
and_5  g18185(new_n20533_1, new_n20532, new_n20534);
xnor_4 g18186(new_n20533_1, new_n9598_1, new_n20535);
not_10 g18187(new_n9603, new_n20536);
xor_4  g18188(new_n20489_1, new_n20478_1, new_n20537);
and_5  g18189(new_n20537, new_n20536, new_n20538);
xnor_4 g18190(new_n20537, new_n9603, new_n20539);
xor_4  g18191(new_n20487, new_n20486, new_n20540);
nor_5  g18192(new_n20540, new_n9608, new_n20541);
xor_4  g18193(new_n20540, new_n9608, new_n20542);
xnor_4 g18194(new_n20484, new_n10909, new_n20543);
and_5  g18195(new_n20543, new_n9612, new_n20544);
xor_4  g18196(new_n10906, new_n9333, new_n20545);
nor_5  g18197(new_n20545, new_n9616_1, new_n20546);
not_10 g18198(new_n20546, new_n20547);
xor_4  g18199(new_n20543, new_n9612, new_n20548);
and_5  g18200(new_n20548, new_n20547, new_n20549);
or_5   g18201(new_n20549, new_n20544, new_n20550);
and_5  g18202(new_n20550, new_n20542, new_n20551);
or_5   g18203(new_n20551, new_n20541, new_n20552);
and_5  g18204(new_n20552, new_n20539, new_n20553);
or_5   g18205(new_n20553, new_n20538, new_n20554);
and_5  g18206(new_n20554, new_n20535, new_n20555);
or_5   g18207(new_n20555, new_n20534, new_n20556);
and_5  g18208(new_n20556, new_n20531, new_n20557);
or_5   g18209(new_n20557, new_n20530, new_n20558);
and_5  g18210(new_n20558, new_n20527, new_n20559);
or_5   g18211(new_n20559, new_n20526, new_n20560);
and_5  g18212(new_n20560, new_n20523, new_n20561);
or_5   g18213(new_n20561, new_n20522, new_n20562);
and_5  g18214(new_n20562, new_n20520, new_n20563);
or_5   g18215(new_n20563, new_n20519, new_n20564);
and_5  g18216(new_n20564, new_n20517, new_n20565);
or_5   g18217(new_n20565, new_n20516, new_n20566);
and_5  g18218(new_n20566, new_n20514, new_n20567);
nor_5  g18219(new_n20567, new_n20513, new_n20568);
not_10 g18220(new_n20568, new_n20569);
xor_4  g18221(new_n20569, new_n19756_1, new_n20570);
xor_4  g18222(new_n20570, new_n20510, n6628);
xnor_4 g18223(new_n2821, new_n2805, n6630);
xnor_4 g18224(n25331, n17911, new_n20573);
or_5   g18225(n21997, n18483, new_n20574);
nand_5 g18226(new_n19862, new_n19855, new_n20575);
and_5  g18227(new_n20575, new_n20574, new_n20576);
xor_4  g18228(new_n20576, new_n20573, new_n20577);
xor_4  g18229(new_n20577, new_n7577, new_n20578);
or_5   g18230(new_n19863, new_n7568, new_n20579);
nand_5 g18231(new_n19873_1, new_n19864, new_n20580);
and_5  g18232(new_n20580, new_n20579, new_n20581);
xnor_4 g18233(new_n20581, new_n20578, new_n20582_1);
not_10 g18234(new_n20582_1, new_n20583);
xor_4  g18235(n14130, n468, new_n20584);
or_5   g18236(n16482, new_n8421, new_n20585);
xor_4  g18237(n16482, n5400, new_n20586);
or_5   g18238(new_n17625, n9942, new_n20587);
and_5  g18239(new_n3413, n329, new_n20588);
xor_4  g18240(n25643, n329, new_n20589);
or_5   g18241(new_n13556, n9557, new_n20590_1);
xnor_4 g18242(n24170, n9557, new_n20591);
or_5   g18243(new_n3415, n2409, new_n20592);
xor_4  g18244(n3136, n2409, new_n20593);
or_5   g18245(n8869, new_n2361_1, new_n20594);
or_5   g18246(new_n19441, new_n19438, new_n20595);
and_5  g18247(new_n20595, new_n20594, new_n20596);
or_5   g18248(new_n20596, new_n20593, new_n20597);
and_5  g18249(new_n20597, new_n20592, new_n20598);
nand_5 g18250(new_n20598, new_n20591, new_n20599);
and_5  g18251(new_n20599, new_n20590_1, new_n20600);
nor_5  g18252(new_n20600, new_n20589, new_n20601);
or_5   g18253(new_n20601, new_n20588, new_n20602_1);
xnor_4 g18254(n23923, n9942, new_n20603);
nand_5 g18255(new_n20603, new_n20602_1, new_n20604_1);
and_5  g18256(new_n20604_1, new_n20587, new_n20605);
or_5   g18257(new_n20605, new_n20586, new_n20606);
and_5  g18258(new_n20606, new_n20585, new_n20607);
xor_4  g18259(new_n20607, new_n20584, new_n20608);
xnor_4 g18260(new_n20608, new_n20583, new_n20609_1);
xor_4  g18261(new_n20605, new_n20586, new_n20610);
or_5   g18262(new_n20610, new_n19874, new_n20611);
xor_4  g18263(new_n20610, new_n19874, new_n20612);
xor_4  g18264(new_n20603, new_n20602_1, new_n20613);
and_5  g18265(new_n20613, new_n19882, new_n20614);
xor_4  g18266(new_n20600, new_n20589, new_n20615);
or_5   g18267(new_n20615, new_n19483, new_n20616);
xnor_4 g18268(new_n20615, new_n19484, new_n20617);
xor_4  g18269(new_n20598, new_n20591, new_n20618);
not_10 g18270(new_n20618, new_n20619);
nand_5 g18271(new_n20619, new_n19509, new_n20620);
xnor_4 g18272(new_n20618, new_n19509, new_n20621);
not_10 g18273(new_n20621, new_n20622);
xor_4  g18274(new_n20596, new_n20593, new_n20623_1);
nand_5 g18275(new_n20623_1, new_n19511, new_n20624);
xnor_4 g18276(new_n20623_1, new_n19512, new_n20625);
nand_5 g18277(new_n19442, new_n19436, new_n20626);
not_10 g18278(new_n19448, new_n20627);
or_5   g18279(new_n20627, new_n19443, new_n20628);
nand_5 g18280(new_n20628, new_n20626, new_n20629_1);
nand_5 g18281(new_n20629_1, new_n20625, new_n20630);
and_5  g18282(new_n20630, new_n20624, new_n20631);
or_5   g18283(new_n20631, new_n20622, new_n20632);
nand_5 g18284(new_n20632, new_n20620, new_n20633);
nand_5 g18285(new_n20633, new_n20617, new_n20634);
and_5  g18286(new_n20634, new_n20616, new_n20635);
xor_4  g18287(new_n20613, new_n19882, new_n20636);
and_5  g18288(new_n20636, new_n20635, new_n20637);
nor_5  g18289(new_n20637, new_n20614, new_n20638);
nand_5 g18290(new_n20638, new_n20612, new_n20639);
and_5  g18291(new_n20639, new_n20611, new_n20640);
xor_4  g18292(new_n20640, new_n20609_1, n6634);
xnor_4 g18293(new_n6621, new_n6606, n6652);
xnor_4 g18294(new_n12812_1, new_n12794, n6655);
xnor_4 g18295(new_n12297, new_n12275, n6669);
xnor_4 g18296(new_n9625, new_n9606, n6671);
xor_4  g18297(new_n13819, new_n13798_1, n6673);
nor_5  g18298(new_n20356, new_n20349_1, new_n20647);
or_5   g18299(new_n11669, new_n12188, new_n20648);
nor_5  g18300(new_n20354, new_n20648, new_n20649);
or_5   g18301(new_n20649, new_n20647, n6674);
xnor_4 g18302(new_n16907, new_n16895, n6684);
xor_4  g18303(new_n12542, new_n12488, n6706);
xnor_4 g18304(n12702, n8614, new_n20653);
or_5   g18305(n26797, n15182, new_n20654);
xnor_4 g18306(n26797, n15182, new_n20655);
or_5   g18307(n27037, n23913, new_n20656);
xnor_4 g18308(n27037, n23913, new_n20657);
or_5   g18309(n22554, n8964, new_n20658_1);
xnor_4 g18310(n22554, n8964, new_n20659);
or_5   g18311(n20429, n20151, new_n20660);
xnor_4 g18312(n20429, n20151, new_n20661_1);
or_5   g18313(n7693, n3909, new_n20662);
xnor_4 g18314(n7693, n3909, new_n20663);
or_5   g18315(n23974, n10405, new_n20664);
xor_4  g18316(n23974, n10405, new_n20665);
nand_5 g18317(n11302, n2146, new_n20666);
or_5   g18318(n11302, n2146, new_n20667);
nor_5  g18319(n22173, n17090, new_n20668);
and_5  g18320(new_n16018, new_n16017, new_n20669);
nor_5  g18321(new_n20669, new_n20668, new_n20670);
nand_5 g18322(new_n20670, new_n20667, new_n20671);
and_5  g18323(new_n20671, new_n20666, new_n20672);
nand_5 g18324(new_n20672, new_n20665, new_n20673_1);
and_5  g18325(new_n20673_1, new_n20664, new_n20674);
or_5   g18326(new_n20674, new_n20663, new_n20675);
and_5  g18327(new_n20675, new_n20662, new_n20676);
or_5   g18328(new_n20676, new_n20661_1, new_n20677);
and_5  g18329(new_n20677, new_n20660, new_n20678_1);
or_5   g18330(new_n20678_1, new_n20659, new_n20679);
and_5  g18331(new_n20679, new_n20658_1, new_n20680_1);
or_5   g18332(new_n20680_1, new_n20657, new_n20681);
and_5  g18333(new_n20681, new_n20656, new_n20682);
or_5   g18334(new_n20682, new_n20655, new_n20683);
and_5  g18335(new_n20683, new_n20654, new_n20684);
xor_4  g18336(new_n20684, new_n20653, new_n20685_1);
and_5  g18337(new_n20685_1, n1831, new_n20686);
xor_4  g18338(new_n20685_1, new_n18055, new_n20687);
xor_4  g18339(new_n20682, new_n20655, new_n20688);
nand_5 g18340(new_n20688, n13137, new_n20689);
xor_4  g18341(new_n20688, new_n14208, new_n20690);
xor_4  g18342(new_n20680_1, new_n20657, new_n20691_1);
nand_5 g18343(new_n20691_1, n18452, new_n20692);
xor_4  g18344(new_n20691_1, new_n14212, new_n20693);
xor_4  g18345(new_n20678_1, new_n20659, new_n20694);
nand_5 g18346(new_n20694, n21317, new_n20695);
xor_4  g18347(new_n20694, new_n14216, new_n20696_1);
xor_4  g18348(new_n20676, new_n20661_1, new_n20697);
nand_5 g18349(new_n20697, n12398, new_n20698);
xor_4  g18350(new_n20697, new_n4000_1, new_n20699);
xor_4  g18351(new_n20674, new_n20663, new_n20700_1);
nand_5 g18352(new_n20700_1, n19789, new_n20701);
xor_4  g18353(new_n20700_1, new_n4001, new_n20702);
xor_4  g18354(new_n20672, new_n20665, new_n20703);
nand_5 g18355(new_n20703, n20169, new_n20704_1);
xor_4  g18356(new_n20703, new_n4002, new_n20705_1);
xor_4  g18357(n11302, n2146, new_n20706);
xor_4  g18358(new_n20706, new_n20670, new_n20707);
or_5   g18359(new_n20707, new_n4003, new_n20708);
xor_4  g18360(new_n20707, n8285, new_n20709_1);
nand_5 g18361(new_n16019, new_n16016, new_n20710);
and_5  g18362(new_n20710, new_n16015, new_n20711);
or_5   g18363(new_n20711, new_n20709_1, new_n20712);
and_5  g18364(new_n20712, new_n20708, new_n20713_1);
or_5   g18365(new_n20713_1, new_n20705_1, new_n20714);
and_5  g18366(new_n20714, new_n20704_1, new_n20715);
or_5   g18367(new_n20715, new_n20702, new_n20716);
and_5  g18368(new_n20716, new_n20701, new_n20717);
or_5   g18369(new_n20717, new_n20699, new_n20718);
and_5  g18370(new_n20718, new_n20698, new_n20719);
or_5   g18371(new_n20719, new_n20696_1, new_n20720);
and_5  g18372(new_n20720, new_n20695, new_n20721);
or_5   g18373(new_n20721, new_n20693, new_n20722_1);
and_5  g18374(new_n20722_1, new_n20692, new_n20723_1);
or_5   g18375(new_n20723_1, new_n20690, new_n20724);
and_5  g18376(new_n20724, new_n20689, new_n20725);
nor_5  g18377(new_n20725, new_n20687, new_n20726);
nor_5  g18378(new_n20726, new_n20686, new_n20727);
or_5   g18379(n12702, n8614, new_n20728);
or_5   g18380(new_n20684, new_n20653, new_n20729);
and_5  g18381(new_n20729, new_n20728, new_n20730);
xnor_4 g18382(new_n20730, new_n20727, new_n20731);
and_5  g18383(new_n20392, new_n4468, new_n20732);
and_5  g18384(new_n20416, new_n20393, new_n20733);
nor_5  g18385(new_n20733, new_n20732, new_n20734);
and_5  g18386(new_n20391, new_n8210, new_n20735);
xnor_4 g18387(new_n20735, new_n4448, new_n20736);
xnor_4 g18388(new_n20736, new_n20734, new_n20737);
xnor_4 g18389(new_n20737, new_n20731, new_n20738);
not_10 g18390(new_n20738, new_n20739);
xor_4  g18391(new_n20725, new_n20687, new_n20740);
and_5  g18392(new_n20740, new_n20418, new_n20741);
xor_4  g18393(new_n20740, new_n20418, new_n20742);
not_10 g18394(new_n20742, new_n20743);
xor_4  g18395(new_n20723_1, new_n20690, new_n20744);
and_5  g18396(new_n20744, new_n20437, new_n20745);
xnor_4 g18397(new_n20744, new_n20440, new_n20746);
not_10 g18398(new_n20746, new_n20747);
xor_4  g18399(new_n20721, new_n20693, new_n20748_1);
and_5  g18400(new_n20748_1, new_n20442, new_n20749);
xnor_4 g18401(new_n20748_1, new_n20445_1, new_n20750);
not_10 g18402(new_n20750, new_n20751);
xor_4  g18403(new_n20719, new_n20696_1, new_n20752);
and_5  g18404(new_n20752, new_n20447, new_n20753);
xnor_4 g18405(new_n20752, new_n20450_1, new_n20754);
not_10 g18406(new_n20754, new_n20755);
xor_4  g18407(new_n20717, new_n20699, new_n20756);
and_5  g18408(new_n20756, new_n13970, new_n20757);
xnor_4 g18409(new_n20756, new_n13971, new_n20758);
not_10 g18410(new_n20758, new_n20759);
xor_4  g18411(new_n20715, new_n20702, new_n20760);
and_5  g18412(new_n20760, new_n13994, new_n20761_1);
xor_4  g18413(new_n20760, new_n13994, new_n20762);
not_10 g18414(new_n20762, new_n20763);
xor_4  g18415(new_n20713_1, new_n20705_1, new_n20764);
and_5  g18416(new_n20764, new_n13998, new_n20765);
not_10 g18417(new_n20765, new_n20766);
xnor_4 g18418(new_n20764, new_n14001, new_n20767);
not_10 g18419(new_n14003, new_n20768);
xor_4  g18420(new_n20711, new_n20709_1, new_n20769);
nor_5  g18421(new_n20769, new_n20768, new_n20770);
nand_5 g18422(new_n16020, new_n14007, new_n20771);
not_10 g18423(new_n16011, new_n20772);
nand_5 g18424(new_n16021, new_n20772, new_n20773);
and_5  g18425(new_n20773, new_n20771, new_n20774_1);
xor_4  g18426(new_n20769, new_n20768, new_n20775);
and_5  g18427(new_n20775, new_n20774_1, new_n20776);
nor_5  g18428(new_n20776, new_n20770, new_n20777);
and_5  g18429(new_n20777, new_n20767, new_n20778);
not_10 g18430(new_n20778, new_n20779);
and_5  g18431(new_n20779, new_n20766, new_n20780);
nor_5  g18432(new_n20780, new_n20763, new_n20781);
nor_5  g18433(new_n20781, new_n20761_1, new_n20782);
nor_5  g18434(new_n20782, new_n20759, new_n20783);
nor_5  g18435(new_n20783, new_n20757, new_n20784);
nor_5  g18436(new_n20784, new_n20755, new_n20785);
nor_5  g18437(new_n20785, new_n20753, new_n20786);
nor_5  g18438(new_n20786, new_n20751, new_n20787);
nor_5  g18439(new_n20787, new_n20749, new_n20788_1);
nor_5  g18440(new_n20788_1, new_n20747, new_n20789);
nor_5  g18441(new_n20789, new_n20745, new_n20790);
nor_5  g18442(new_n20790, new_n20743, new_n20791);
nor_5  g18443(new_n20791, new_n20741, new_n20792);
xnor_4 g18444(new_n20792, new_n20739, n6707);
xor_4  g18445(new_n13370, new_n13120, n6736);
xor_4  g18446(n23895, n5101, new_n20795_1);
nand_5 g18447(new_n5484, n16507, new_n20796);
xnor_4 g18448(n17351, n16507, new_n20797);
not_10 g18449(new_n20797, new_n20798);
nand_5 g18450(n22470, new_n5488, new_n20799);
xnor_4 g18451(n22470, n11736, new_n20800);
not_10 g18452(new_n20800, new_n20801);
nand_5 g18453(new_n5492, n19116, new_n20802);
and_5  g18454(new_n5496, n6861, new_n20803_1);
not_10 g18455(new_n20803_1, new_n20804);
nor_5  g18456(new_n18281, new_n18261, new_n20805);
not_10 g18457(new_n20805, new_n20806);
and_5  g18458(new_n20806, new_n20804, new_n20807);
xor_4  g18459(n23200, n19116, new_n20808);
or_5   g18460(new_n20808, new_n20807, new_n20809);
and_5  g18461(new_n20809, new_n20802, new_n20810);
or_5   g18462(new_n20810, new_n20801, new_n20811);
and_5  g18463(new_n20811, new_n20799, new_n20812);
or_5   g18464(new_n20812, new_n20798, new_n20813);
and_5  g18465(new_n20813, new_n20796, new_n20814);
xor_4  g18466(new_n20814, new_n20795_1, new_n20815);
and_5  g18467(new_n18286, new_n5553, new_n20816);
and_5  g18468(new_n20816, new_n5549, new_n20817);
and_5  g18469(new_n20817, new_n5545, new_n20818);
and_5  g18470(new_n20818, new_n5541, new_n20819);
xor_4  g18471(new_n20819, new_n11979, new_n20820);
xor_4  g18472(new_n20820, n12650, new_n20821);
xor_4  g18473(new_n20818, new_n5541, new_n20822);
or_5   g18474(new_n20822, new_n5608, new_n20823);
xor_4  g18475(new_n20822, n10201, new_n20824);
xor_4  g18476(new_n20817, new_n5545, new_n20825);
or_5   g18477(new_n20825, new_n5612, new_n20826_1);
xor_4  g18478(new_n20825, n10593, new_n20827);
xor_4  g18479(new_n20816, new_n5549, new_n20828);
or_5   g18480(new_n20828, new_n5616, new_n20829);
xor_4  g18481(new_n20828, n18290, new_n20830);
or_5   g18482(new_n18287, new_n5620, new_n20831);
or_5   g18483(new_n18310_1, new_n18288_1, new_n20832);
and_5  g18484(new_n20832, new_n20831, new_n20833);
or_5   g18485(new_n20833, new_n20830, new_n20834);
and_5  g18486(new_n20834, new_n20829, new_n20835);
or_5   g18487(new_n20835, new_n20827, new_n20836);
and_5  g18488(new_n20836, new_n20826_1, new_n20837);
or_5   g18489(new_n20837, new_n20824, new_n20838);
and_5  g18490(new_n20838, new_n20823, new_n20839);
xor_4  g18491(new_n20839, new_n20821, new_n20840);
xnor_4 g18492(new_n20840, new_n16241, new_n20841);
xor_4  g18493(new_n20837, new_n20824, new_n20842);
or_5   g18494(new_n20842, new_n16244, new_n20843);
xor_4  g18495(new_n20835, new_n20827, new_n20844);
nand_5 g18496(new_n20844, new_n16248, new_n20845);
xor_4  g18497(new_n20844, new_n16248, new_n20846);
xor_4  g18498(new_n20833, new_n20830, new_n20847);
or_5   g18499(new_n20847, new_n16252, new_n20848);
xnor_4 g18500(new_n20847, new_n16252, new_n20849);
or_5   g18501(new_n18311_1, new_n16255, new_n20850);
or_5   g18502(new_n18335, new_n18312, new_n20851);
and_5  g18503(new_n20851, new_n20850, new_n20852);
or_5   g18504(new_n20852, new_n20849, new_n20853);
and_5  g18505(new_n20853, new_n20848, new_n20854);
nand_5 g18506(new_n20854, new_n20846, new_n20855);
and_5  g18507(new_n20855, new_n20845, new_n20856);
xor_4  g18508(new_n20842, new_n16244, new_n20857);
nand_5 g18509(new_n20857, new_n20856, new_n20858);
and_5  g18510(new_n20858, new_n20843, new_n20859);
xor_4  g18511(new_n20859, new_n20841, new_n20860);
xor_4  g18512(new_n20860, new_n20815, new_n20861);
xor_4  g18513(new_n20812, new_n20798, new_n20862);
xor_4  g18514(new_n20857, new_n20856, new_n20863);
or_5   g18515(new_n20863, new_n20862, new_n20864);
xor_4  g18516(new_n20863, new_n20862, new_n20865);
not_10 g18517(new_n20865, new_n20866);
xor_4  g18518(new_n20810, new_n20801, new_n20867);
not_10 g18519(new_n20867, new_n20868);
xor_4  g18520(new_n20854, new_n20846, new_n20869_1);
nand_5 g18521(new_n20869_1, new_n20868, new_n20870);
xor_4  g18522(new_n20869_1, new_n20868, new_n20871);
xor_4  g18523(new_n20808, new_n20807, new_n20872);
xor_4  g18524(new_n20852, new_n20849, new_n20873);
and_5  g18525(new_n20873, new_n20872, new_n20874);
xnor_4 g18526(new_n20873, new_n20872, new_n20875);
nand_5 g18527(new_n18336, new_n18282, new_n20876);
nand_5 g18528(new_n18372, new_n18337, new_n20877);
and_5  g18529(new_n20877, new_n20876, new_n20878);
nor_5  g18530(new_n20878, new_n20875, new_n20879_1);
nor_5  g18531(new_n20879_1, new_n20874, new_n20880);
nand_5 g18532(new_n20880, new_n20871, new_n20881);
and_5  g18533(new_n20881, new_n20870, new_n20882);
or_5   g18534(new_n20882, new_n20866, new_n20883);
and_5  g18535(new_n20883, new_n20864, new_n20884);
xor_4  g18536(new_n20884, new_n20861, n6791);
xnor_4 g18537(new_n3708, new_n3698, n6802);
xnor_4 g18538(new_n16591, new_n16564, n6826);
xnor_4 g18539(new_n10244_1, new_n10213, n6835);
nand_5 g18540(new_n18592, n11220, new_n20889);
not_10 g18541(n11220, new_n20890);
xor_4  g18542(new_n18592, new_n20890, new_n20891);
or_5   g18543(new_n2913, new_n18572_1, new_n20892);
xor_4  g18544(new_n2913, n22379, new_n20893);
or_5   g18545(new_n2953, new_n2837, new_n20894);
xor_4  g18546(new_n2953, n1662, new_n20895);
or_5   g18547(new_n2958, new_n2841, new_n20896);
xor_4  g18548(new_n2958, n12875, new_n20897);
or_5   g18549(new_n2964, new_n2845, new_n20898);
nand_5 g18550(new_n2970, new_n2849, new_n20899);
xor_4  g18551(new_n2970, n5213, new_n20900);
nand_5 g18552(new_n2976, new_n2853_1, new_n20901);
xor_4  g18553(new_n2976, new_n2853_1, new_n20902);
or_5   g18554(new_n2981, new_n2858_1, new_n20903);
xor_4  g18555(new_n2981, new_n2858_1, new_n20904);
and_5  g18556(new_n2991, n5438, new_n20905);
or_5   g18557(new_n20905, n4326, new_n20906);
xor_4  g18558(new_n20905, n4326, new_n20907);
nand_5 g18559(new_n20907, new_n2987, new_n20908);
and_5  g18560(new_n20908, new_n20906, new_n20909);
nand_5 g18561(new_n20909, new_n20904, new_n20910);
and_5  g18562(new_n20910, new_n20903, new_n20911);
nand_5 g18563(new_n20911, new_n20902, new_n20912);
and_5  g18564(new_n20912, new_n20901, new_n20913);
or_5   g18565(new_n20913, new_n20900, new_n20914);
and_5  g18566(new_n20914, new_n20899, new_n20915_1);
xor_4  g18567(new_n2964, new_n2845, new_n20916);
nand_5 g18568(new_n20916, new_n20915_1, new_n20917);
and_5  g18569(new_n20917, new_n20898, new_n20918);
or_5   g18570(new_n20918, new_n20897, new_n20919);
and_5  g18571(new_n20919, new_n20896, new_n20920);
or_5   g18572(new_n20920, new_n20895, new_n20921);
and_5  g18573(new_n20921, new_n20894, new_n20922);
or_5   g18574(new_n20922, new_n20893, new_n20923_1);
and_5  g18575(new_n20923_1, new_n20892, new_n20924);
or_5   g18576(new_n20924, new_n20891, new_n20925);
and_5  g18577(new_n20925, new_n20889, new_n20926);
nor_5  g18578(new_n20926, new_n18586, new_n20927);
xor_4  g18579(new_n20927, new_n18242, new_n20928);
xor_4  g18580(new_n20926, new_n18586, new_n20929_1);
nor_5  g18581(new_n20929_1, new_n18245, new_n20930);
xnor_4 g18582(new_n20929_1, new_n18244, new_n20931);
not_10 g18583(new_n20931, new_n20932);
xor_4  g18584(new_n20924, new_n20891, new_n20933);
nor_5  g18585(new_n20933, new_n18249, new_n20934);
xnor_4 g18586(new_n20933, new_n6126, new_n20935_1);
not_10 g18587(new_n20935_1, new_n20936_1);
xor_4  g18588(new_n20922, new_n20893, new_n20937);
nor_5  g18589(new_n20937, new_n13173, new_n20938);
xnor_4 g18590(new_n20937, new_n6128, new_n20939);
not_10 g18591(new_n20939, new_n20940);
xnor_4 g18592(new_n20920, new_n20895, new_n20941);
and_5  g18593(new_n20941, new_n6135, new_n20942);
xor_4  g18594(new_n20941, new_n6135, new_n20943);
not_10 g18595(new_n20943, new_n20944);
xor_4  g18596(new_n20918, new_n20897, new_n20945);
nor_5  g18597(new_n20945, new_n13181, new_n20946_1);
xnor_4 g18598(new_n20945, new_n6140, new_n20947);
not_10 g18599(new_n20947, new_n20948);
xnor_4 g18600(new_n20916, new_n20915_1, new_n20949);
and_5  g18601(new_n20949, new_n6145, new_n20950);
xor_4  g18602(new_n20949, new_n6145, new_n20951);
not_10 g18603(new_n20951, new_n20952);
xor_4  g18604(new_n20913, new_n20900, new_n20953);
and_5  g18605(new_n20953, new_n6150, new_n20954);
xor_4  g18606(new_n20953, new_n6150, new_n20955);
not_10 g18607(new_n20955, new_n20956);
xor_4  g18608(new_n20911, new_n20902, new_n20957);
and_5  g18609(new_n20957, new_n6155, new_n20958);
xor_4  g18610(new_n20957, new_n6155, new_n20959);
not_10 g18611(new_n20959, new_n20960);
xor_4  g18612(new_n20909, new_n20904, new_n20961);
nor_5  g18613(new_n20961, new_n6161, new_n20962);
xnor_4 g18614(new_n20961, new_n6160_1, new_n20963);
not_10 g18615(new_n20963, new_n20964);
xor_4  g18616(new_n20907, new_n2987, new_n20965);
and_5  g18617(new_n20965, new_n13199_1, new_n20966);
not_10 g18618(new_n20966, new_n20967);
nor_5  g18619(new_n5853, new_n6167, new_n20968);
xor_4  g18620(new_n20965, new_n13199_1, new_n20969);
and_5  g18621(new_n20969, new_n20968, new_n20970);
not_10 g18622(new_n20970, new_n20971);
and_5  g18623(new_n20971, new_n20967, new_n20972);
nor_5  g18624(new_n20972, new_n20964, new_n20973);
nor_5  g18625(new_n20973, new_n20962, new_n20974);
nor_5  g18626(new_n20974, new_n20960, new_n20975);
nor_5  g18627(new_n20975, new_n20958, new_n20976);
nor_5  g18628(new_n20976, new_n20956, new_n20977);
nor_5  g18629(new_n20977, new_n20954, new_n20978);
nor_5  g18630(new_n20978, new_n20952, new_n20979);
nor_5  g18631(new_n20979, new_n20950, new_n20980);
nor_5  g18632(new_n20980, new_n20948, new_n20981);
nor_5  g18633(new_n20981, new_n20946_1, new_n20982);
nor_5  g18634(new_n20982, new_n20944, new_n20983);
nor_5  g18635(new_n20983, new_n20942, new_n20984);
nor_5  g18636(new_n20984, new_n20940, new_n20985);
nor_5  g18637(new_n20985, new_n20938, new_n20986_1);
nor_5  g18638(new_n20986_1, new_n20936_1, new_n20987);
nor_5  g18639(new_n20987, new_n20934, new_n20988);
nor_5  g18640(new_n20988, new_n20932, new_n20989);
nor_5  g18641(new_n20989, new_n20930, new_n20990);
xnor_4 g18642(new_n20990, new_n20928, n6853);
xnor_4 g18643(new_n15206, new_n11350, new_n20992);
or_5   g18644(new_n15211, new_n11354, new_n20993);
xor_4  g18645(new_n15211, new_n11354, new_n20994);
nand_5 g18646(new_n11358, new_n4190, new_n20995);
not_10 g18647(new_n13225, new_n20996);
or_5   g18648(new_n13239, new_n20996, new_n20997);
and_5  g18649(new_n20997, new_n20995, new_n20998);
nand_5 g18650(new_n20998, new_n20994, new_n20999);
and_5  g18651(new_n20999, new_n20993, new_n21000);
xor_4  g18652(new_n21000, new_n20992, n6862);
not_10 g18653(n8305, new_n21002);
and_5  g18654(n22253, new_n21002, new_n21003);
nor_5  g18655(new_n16198, new_n16180, new_n21004);
nor_5  g18656(new_n21004, new_n21003, new_n21005);
not_10 g18657(n25296, new_n21006);
or_5   g18658(new_n21006, n23717, new_n21007);
or_5   g18659(new_n11519, new_n11504, new_n21008_1);
and_5  g18660(new_n21008_1, new_n21007, new_n21009);
nor_5  g18661(new_n21009, new_n18752, new_n21010);
nor_5  g18662(new_n11521, new_n11502, new_n21011);
not_10 g18663(new_n21011, new_n21012);
nor_5  g18664(new_n11544, new_n11522, new_n21013);
not_10 g18665(new_n21013, new_n21014);
and_5  g18666(new_n21014, new_n21012, new_n21015);
xnor_4 g18667(new_n21009, new_n18752, new_n21016);
nor_5  g18668(new_n21016, new_n21015, new_n21017_1);
nor_5  g18669(new_n21017_1, new_n21010, new_n21018);
nand_5 g18670(new_n21018, new_n21005, new_n21019);
and_5  g18671(new_n16199, new_n11545, new_n21020);
and_5  g18672(new_n16219_1, new_n16200, new_n21021);
nor_5  g18673(new_n21021, new_n21020, new_n21022);
or_5   g18674(new_n21022, new_n21018, new_n21023);
and_5  g18675(new_n21023, new_n21019, new_n21024);
xor_4  g18676(new_n21016, new_n21015, new_n21025);
or_5   g18677(new_n21025, new_n21005, new_n21026);
nand_5 g18678(new_n21025, new_n21022, new_n21027);
and_5  g18679(new_n21027, new_n21026, new_n21028);
and_5  g18680(new_n21028, new_n21024, n6863);
xnor_4 g18681(new_n6189_1, new_n6132, n6867);
xnor_4 g18682(new_n18187, new_n18179, n6965);
xor_4  g18683(new_n7492, new_n7441, n6967);
xor_4  g18684(new_n14752, new_n14710, n6975);
xor_4  g18685(new_n20329, new_n20328, n6983);
xor_4  g18686(new_n15186, new_n11336, new_n21035);
not_10 g18687(new_n21035, new_n21036);
and_5  g18688(new_n15191, new_n11338, new_n21037);
xor_4  g18689(new_n15191, new_n11338, new_n21038);
not_10 g18690(new_n21038, new_n21039);
and_5  g18691(new_n15194, new_n11342, new_n21040);
not_10 g18692(new_n21040, new_n21041);
xor_4  g18693(new_n15194, new_n11342, new_n21042);
nor_5  g18694(new_n15199, new_n11346, new_n21043);
nor_5  g18695(new_n15206, new_n11350, new_n21044);
nor_5  g18696(new_n21000, new_n20992, new_n21045);
or_5   g18697(new_n21045, new_n21044, new_n21046_1);
xor_4  g18698(new_n15199, new_n11346, new_n21047);
and_5  g18699(new_n21047, new_n21046_1, new_n21048);
nor_5  g18700(new_n21048, new_n21043, new_n21049);
and_5  g18701(new_n21049, new_n21042, new_n21050);
not_10 g18702(new_n21050, new_n21051);
and_5  g18703(new_n21051, new_n21041, new_n21052);
nor_5  g18704(new_n21052, new_n21039, new_n21053);
nor_5  g18705(new_n21053, new_n21037, new_n21054);
xnor_4 g18706(new_n21054, new_n21036, n6985);
xnor_4 g18707(new_n15010, new_n14961, n6998);
xor_4  g18708(new_n11299, new_n9064, n7032);
xor_4  g18709(new_n20190, new_n20155, n7038);
xnor_4 g18710(new_n17998_1, new_n17997, n7079);
xnor_4 g18711(new_n7474, new_n7473, n7190);
xnor_4 g18712(new_n16150, new_n16145, n7229);
xor_4  g18713(new_n8718, new_n8705, n7230);
xnor_4 g18714(new_n19414_1, new_n19413, n7233);
xnor_4 g18715(new_n13486_1, new_n13478, n7236);
xor_4  g18716(new_n16479, new_n6967_1, n7253);
and_5  g18717(new_n19801, new_n7250, new_n21066);
nor_5  g18718(new_n19802, n12507, new_n21067);
and_5  g18719(new_n19802, n12507, new_n21068);
nor_5  g18720(new_n19806, new_n21068, new_n21069);
nor_5  g18721(new_n21069, new_n21067, new_n21070);
nor_5  g18722(new_n21070, new_n21066, new_n21071);
not_10 g18723(new_n21071, new_n21072);
and_5  g18724(new_n20263, new_n14399, new_n21073);
xor_4  g18725(new_n21073, new_n14396, new_n21074);
nor_5  g18726(new_n21074, new_n10341, new_n21075);
xor_4  g18727(new_n21074, new_n10340_1, new_n21076);
or_5   g18728(new_n20264, new_n10344, new_n21077);
or_5   g18729(new_n20303, new_n20265, new_n21078_1);
and_5  g18730(new_n21078_1, new_n21077, new_n21079);
nor_5  g18731(new_n21079, new_n21076, new_n21080);
or_5   g18732(new_n21080, new_n21075, new_n21081);
and_5  g18733(new_n21073, new_n14396, new_n21082);
not_10 g18734(new_n21082, new_n21083);
and_5  g18735(new_n21083, new_n14443, new_n21084);
and_5  g18736(new_n21082, new_n14441, new_n21085);
nor_5  g18737(new_n21085, new_n21084, new_n21086);
xor_4  g18738(new_n21086, new_n10335, new_n21087);
xor_4  g18739(new_n21087, new_n21081, new_n21088);
and_5  g18740(new_n21088, new_n21072, new_n21089);
xor_4  g18741(new_n21088, new_n21072, new_n21090);
xor_4  g18742(new_n21079, new_n21076, new_n21091);
nor_5  g18743(new_n21091, new_n19808, new_n21092);
nor_5  g18744(new_n20304, new_n16966, new_n21093_1);
and_5  g18745(new_n20344, new_n20305, new_n21094_1);
or_5   g18746(new_n21094_1, new_n21093_1, new_n21095_1);
xor_4  g18747(new_n21091, new_n19808, new_n21096);
and_5  g18748(new_n21096, new_n21095_1, new_n21097);
nor_5  g18749(new_n21097, new_n21092, new_n21098);
and_5  g18750(new_n21098, new_n21090, new_n21099);
nor_5  g18751(new_n21099, new_n21089, new_n21100);
nand_5 g18752(new_n21086, new_n10335, new_n21101);
nor_5  g18753(new_n21086, new_n10335, new_n21102);
nor_5  g18754(new_n21102, new_n21081, new_n21103);
nor_5  g18755(new_n21103, new_n21085, new_n21104);
nand_5 g18756(new_n21104, new_n21101, new_n21105);
xnor_4 g18757(new_n21105, new_n21100, n7256);
or_5   g18758(new_n8894, n2416, new_n21107);
xor_4  g18759(n22764, n2416, new_n21108);
or_5   g18760(new_n8096, n21905, new_n21109);
or_5   g18761(new_n19906, new_n19895, new_n21110);
and_5  g18762(new_n21110, new_n21109, new_n21111);
or_5   g18763(new_n21111, new_n21108, new_n21112);
and_5  g18764(new_n21112, new_n21107, new_n21113);
xnor_4 g18765(new_n21111, new_n21108, new_n21114);
or_5   g18766(new_n21114, new_n15818, new_n21115);
xnor_4 g18767(new_n21114, new_n15818, new_n21116);
nand_5 g18768(new_n19907, new_n15822, new_n21117);
nand_5 g18769(new_n19921, new_n19908, new_n21118);
and_5  g18770(new_n21118, new_n21117, new_n21119);
or_5   g18771(new_n21119, new_n21116, new_n21120);
and_5  g18772(new_n21120, new_n21115, new_n21121);
xor_4  g18773(new_n21121, new_n21113, new_n21122);
xnor_4 g18774(new_n21122, new_n15816_1, new_n21123_1);
xor_4  g18775(new_n21123_1, new_n20011, new_n21124);
not_10 g18776(new_n21124, new_n21125);
xor_4  g18777(new_n21119, new_n21116, new_n21126);
nor_5  g18778(new_n21126, new_n20021, new_n21127);
xor_4  g18779(new_n21126, new_n20021, new_n21128);
not_10 g18780(new_n21128, new_n21129);
nor_5  g18781(new_n19922_1, new_n19894, new_n21130);
nor_5  g18782(new_n19940, new_n19924, new_n21131);
nor_5  g18783(new_n21131, new_n21130, new_n21132);
nor_5  g18784(new_n21132, new_n21129, new_n21133);
nor_5  g18785(new_n21133, new_n21127, new_n21134_1);
xnor_4 g18786(new_n21134_1, new_n21125, n7268);
and_5  g18787(new_n11084, new_n11075, new_n21136);
and_5  g18788(new_n21136, new_n11799, new_n21137);
and_5  g18789(new_n21137, new_n11795, new_n21138_1);
and_5  g18790(new_n21138_1, new_n11838, new_n21139);
not_10 g18791(n10514, new_n21140);
xor_4  g18792(new_n21138_1, new_n11838, new_n21141);
or_5   g18793(new_n21141, new_n21140, new_n21142);
xor_4  g18794(new_n21141, n10514, new_n21143);
not_10 g18795(n18649, new_n21144);
xor_4  g18796(new_n21137, new_n11795, new_n21145);
or_5   g18797(new_n21145, new_n21144, new_n21146);
xor_4  g18798(new_n21145, n18649, new_n21147);
not_10 g18799(n6218, new_n21148);
xor_4  g18800(new_n21136, new_n11799, new_n21149);
or_5   g18801(new_n21149, new_n21148, new_n21150);
xor_4  g18802(new_n21149, n6218, new_n21151);
not_10 g18803(n20470, new_n21152);
or_5   g18804(new_n11085, new_n21152, new_n21153);
xor_4  g18805(new_n11085, n20470, new_n21154_1);
not_10 g18806(n21222, new_n21155);
or_5   g18807(new_n11089, new_n21155, new_n21156);
xor_4  g18808(new_n11089, n21222, new_n21157_1);
not_10 g18809(n9832, new_n21158);
or_5   g18810(new_n11092, new_n21158, new_n21159);
xor_4  g18811(new_n11092, n9832, new_n21160);
not_10 g18812(n1558, new_n21161);
or_5   g18813(new_n11095, new_n21161, new_n21162);
xor_4  g18814(new_n11095, n1558, new_n21163);
not_10 g18815(n21749, new_n21164);
or_5   g18816(new_n11097, new_n21164, new_n21165);
xor_4  g18817(new_n11097, n21749, new_n21166);
not_10 g18818(n7769, new_n21167);
or_5   g18819(new_n11102, new_n21167, new_n21168_1);
and_5  g18820(n21138, new_n11100, new_n21169);
xor_4  g18821(new_n11102, new_n21167, new_n21170);
nand_5 g18822(new_n21170, new_n21169, new_n21171);
and_5  g18823(new_n21171, new_n21168_1, new_n21172);
or_5   g18824(new_n21172, new_n21166, new_n21173_1);
and_5  g18825(new_n21173_1, new_n21165, new_n21174);
or_5   g18826(new_n21174, new_n21163, new_n21175);
and_5  g18827(new_n21175, new_n21162, new_n21176_1);
or_5   g18828(new_n21176_1, new_n21160, new_n21177);
and_5  g18829(new_n21177, new_n21159, new_n21178);
or_5   g18830(new_n21178, new_n21157_1, new_n21179);
and_5  g18831(new_n21179, new_n21156, new_n21180);
or_5   g18832(new_n21180, new_n21154_1, new_n21181);
and_5  g18833(new_n21181, new_n21153, new_n21182_1);
or_5   g18834(new_n21182_1, new_n21151, new_n21183);
and_5  g18835(new_n21183, new_n21150, new_n21184);
or_5   g18836(new_n21184, new_n21147, new_n21185);
and_5  g18837(new_n21185, new_n21146, new_n21186);
or_5   g18838(new_n21186, new_n21143, new_n21187);
and_5  g18839(new_n21187, new_n21142, new_n21188);
and_5  g18840(new_n21188, new_n21139, new_n21189);
not_10 g18841(new_n21189, new_n21190);
xor_4  g18842(new_n21186, new_n21143, new_n21191);
nor_5  g18843(new_n21191, n9872, new_n21192);
not_10 g18844(new_n21192, new_n21193_1);
not_10 g18845(n9872, new_n21194);
xor_4  g18846(new_n21191, new_n21194, new_n21195);
xor_4  g18847(new_n21184, new_n21147, new_n21196);
or_5   g18848(new_n21196, n5842, new_n21197);
not_10 g18849(n5842, new_n21198);
xor_4  g18850(new_n21196, new_n21198, new_n21199);
xor_4  g18851(new_n21182_1, new_n21151, new_n21200);
or_5   g18852(new_n21200, n6379, new_n21201);
not_10 g18853(n6379, new_n21202);
xor_4  g18854(new_n21200, new_n21202, new_n21203_1);
xor_4  g18855(new_n21180, new_n21154_1, new_n21204);
or_5   g18856(new_n21204, n2102, new_n21205);
not_10 g18857(n2102, new_n21206);
xor_4  g18858(new_n21204, new_n21206, new_n21207);
xor_4  g18859(new_n21178, new_n21157_1, new_n21208);
or_5   g18860(new_n21208, n17954, new_n21209);
xor_4  g18861(new_n21176_1, new_n21160, new_n21210);
nor_5  g18862(new_n21210, n8256, new_n21211);
not_10 g18863(n8256, new_n21212);
xor_4  g18864(new_n21210, new_n21212, new_n21213);
xor_4  g18865(new_n21174, new_n21163, new_n21214);
or_5   g18866(new_n21214, n24150, new_n21215);
not_10 g18867(n24150, new_n21216);
xor_4  g18868(new_n21214, new_n21216, new_n21217);
xor_4  g18869(new_n21172, new_n21166, new_n21218);
or_5   g18870(new_n21218, n19584, new_n21219);
xor_4  g18871(new_n21218, n19584, new_n21220);
xor_4  g18872(new_n21170, new_n21169, new_n21221);
nand_5 g18873(new_n21221, n5060, new_n21222_1);
or_5   g18874(new_n21221, n5060, new_n21223);
xnor_4 g18875(n21138, n15506, new_n21224);
and_5  g18876(new_n21224, n15332, new_n21225_1);
nand_5 g18877(new_n21225_1, new_n21223, new_n21226_1);
and_5  g18878(new_n21226_1, new_n21222_1, new_n21227);
nand_5 g18879(new_n21227, new_n21220, new_n21228);
and_5  g18880(new_n21228, new_n21219, new_n21229);
or_5   g18881(new_n21229, new_n21217, new_n21230);
and_5  g18882(new_n21230, new_n21215, new_n21231);
nor_5  g18883(new_n21231, new_n21213, new_n21232);
or_5   g18884(new_n21232, new_n21211, new_n21233);
xor_4  g18885(new_n21208, n17954, new_n21234);
nand_5 g18886(new_n21234, new_n21233, new_n21235);
and_5  g18887(new_n21235, new_n21209, new_n21236);
or_5   g18888(new_n21236, new_n21207, new_n21237);
and_5  g18889(new_n21237, new_n21205, new_n21238_1);
or_5   g18890(new_n21238_1, new_n21203_1, new_n21239);
and_5  g18891(new_n21239, new_n21201, new_n21240);
or_5   g18892(new_n21240, new_n21199, new_n21241);
and_5  g18893(new_n21241, new_n21197, new_n21242);
nor_5  g18894(new_n21242, new_n21195, new_n21243);
not_10 g18895(new_n21243, new_n21244);
and_5  g18896(new_n21244, new_n21193_1, new_n21245);
nor_5  g18897(new_n21245, new_n21190, new_n21246);
nor_5  g18898(new_n21188, new_n21139, new_n21247);
and_5  g18899(new_n21247, new_n21245, new_n21248);
nor_5  g18900(new_n21248, new_n21246, new_n21249);
xor_4  g18901(new_n21249, new_n14946, new_n21250);
not_10 g18902(new_n21139, new_n21251);
xnor_4 g18903(new_n21188, new_n21251, new_n21252);
xor_4  g18904(new_n21252, new_n21245, new_n21253);
nor_5  g18905(new_n21253, new_n14951, new_n21254_1);
xor_4  g18906(new_n21253, new_n14951, new_n21255);
not_10 g18907(new_n21255, new_n21256);
xor_4  g18908(new_n21242, new_n21195, new_n21257);
nor_5  g18909(new_n21257, new_n2649, new_n21258);
xor_4  g18910(new_n21257, new_n2649, new_n21259);
not_10 g18911(new_n21259, new_n21260);
xor_4  g18912(new_n21240, new_n21199, new_n21261);
nor_5  g18913(new_n21261, new_n2776, new_n21262);
xor_4  g18914(new_n21238_1, new_n21203_1, new_n21263);
nor_5  g18915(new_n21263, new_n2780, new_n21264);
xor_4  g18916(new_n21263, new_n2780, new_n21265);
not_10 g18917(new_n21265, new_n21266);
xor_4  g18918(new_n21236, new_n21207, new_n21267);
nor_5  g18919(new_n21267, new_n2786, new_n21268);
xor_4  g18920(new_n21267, new_n2786, new_n21269);
not_10 g18921(new_n21269, new_n21270);
not_10 g18922(new_n2791, new_n21271);
xor_4  g18923(new_n21234, new_n21233, new_n21272);
nor_5  g18924(new_n21272, new_n21271, new_n21273);
xor_4  g18925(new_n21272, new_n21271, new_n21274);
not_10 g18926(new_n21274, new_n21275);
xor_4  g18927(new_n21231, new_n21213, new_n21276_1);
nor_5  g18928(new_n21276_1, new_n2798, new_n21277);
xor_4  g18929(new_n21276_1, new_n2798, new_n21278);
not_10 g18930(new_n21278, new_n21279);
xor_4  g18931(new_n21229, new_n21217, new_n21280);
nor_5  g18932(new_n21280, new_n2802, new_n21281);
xor_4  g18933(new_n21280, new_n2802, new_n21282);
not_10 g18934(new_n21282, new_n21283);
xor_4  g18935(new_n21227, new_n21220, new_n21284);
or_5   g18936(new_n21284, new_n2807, new_n21285);
xor_4  g18937(new_n21284, new_n2807, new_n21286);
not_10 g18938(new_n21286, new_n21287_1);
xor_4  g18939(new_n21221, n5060, new_n21288);
xor_4  g18940(new_n21288, new_n21225_1, new_n21289);
nand_5 g18941(new_n21289, new_n2811, new_n21290);
xor_4  g18942(new_n21224, n15332, new_n21291);
nor_5  g18943(new_n21291, new_n2813, new_n21292);
xor_4  g18944(new_n21289, new_n2811, new_n21293);
not_10 g18945(new_n21293, new_n21294);
or_5   g18946(new_n21294, new_n21292, new_n21295);
and_5  g18947(new_n21295, new_n21290, new_n21296);
or_5   g18948(new_n21296, new_n21287_1, new_n21297);
and_5  g18949(new_n21297, new_n21285, new_n21298_1);
nor_5  g18950(new_n21298_1, new_n21283, new_n21299);
nor_5  g18951(new_n21299, new_n21281, new_n21300);
nor_5  g18952(new_n21300, new_n21279, new_n21301);
nor_5  g18953(new_n21301, new_n21277, new_n21302_1);
nor_5  g18954(new_n21302_1, new_n21275, new_n21303);
nor_5  g18955(new_n21303, new_n21273, new_n21304);
nor_5  g18956(new_n21304, new_n21270, new_n21305);
nor_5  g18957(new_n21305, new_n21268, new_n21306);
nor_5  g18958(new_n21306, new_n21266, new_n21307);
nor_5  g18959(new_n21307, new_n21264, new_n21308);
xor_4  g18960(new_n21261, new_n2776, new_n21309);
not_10 g18961(new_n21309, new_n21310);
nor_5  g18962(new_n21310, new_n21308, new_n21311);
nor_5  g18963(new_n21311, new_n21262, new_n21312);
nor_5  g18964(new_n21312, new_n21260, new_n21313);
nor_5  g18965(new_n21313, new_n21258, new_n21314);
nor_5  g18966(new_n21314, new_n21256, new_n21315);
or_5   g18967(new_n21315, new_n21254_1, new_n21316);
xnor_4 g18968(new_n21316, new_n21250, n7277);
xor_4  g18969(new_n13655, new_n13647, n7280);
xnor_4 g18970(new_n5813, new_n5782_1, n7298);
xor_4  g18971(new_n19788, new_n19775, n7308);
xor_4  g18972(new_n20018, new_n7294, new_n21321);
nand_5 g18973(new_n20020, new_n7312, new_n21322);
not_10 g18974(new_n7312, new_n21323);
xor_4  g18975(new_n20020, new_n21323, new_n21324);
nand_5 g18976(new_n15255_1, new_n7316, new_n21325);
or_5   g18977(new_n15282, new_n15257, new_n21326);
and_5  g18978(new_n21326, new_n21325, new_n21327);
or_5   g18979(new_n21327, new_n21324, new_n21328);
and_5  g18980(new_n21328, new_n21322, new_n21329);
xor_4  g18981(new_n21329, new_n21321, new_n21330);
not_10 g18982(new_n21330, new_n21331);
xor_4  g18983(new_n21331, new_n20045, new_n21332);
xor_4  g18984(new_n21327, new_n21324, new_n21333);
nor_5  g18985(new_n21333, new_n20051, new_n21334);
not_10 g18986(new_n21334, new_n21335);
and_5  g18987(new_n19391, new_n15283, new_n21336);
and_5  g18988(new_n19422, new_n19392, new_n21337);
nor_5  g18989(new_n21337, new_n21336, new_n21338);
xor_4  g18990(new_n21333, new_n20051, new_n21339);
and_5  g18991(new_n21339, new_n21338, new_n21340);
not_10 g18992(new_n21340, new_n21341);
and_5  g18993(new_n21341, new_n21335, new_n21342);
xor_4  g18994(new_n21342, new_n21332, n7313);
xnor_4 g18995(new_n3712, new_n3686, n7346);
xor_4  g18996(new_n21009, new_n14300, new_n21345);
nor_5  g18997(new_n21009, new_n14303, new_n21346);
xor_4  g18998(new_n21009, new_n14303, new_n21347);
not_10 g18999(new_n21347, new_n21348);
and_5  g19000(new_n14309, new_n11521, new_n21349_1);
xnor_4 g19001(new_n14309, new_n11520, new_n21350);
not_10 g19002(new_n21350, new_n21351);
and_5  g19003(new_n14315, new_n11526, new_n21352);
xnor_4 g19004(new_n14315, new_n11525, new_n21353);
not_10 g19005(new_n21353, new_n21354);
nor_5  g19006(new_n14320, new_n11530, new_n21355);
not_10 g19007(new_n21355, new_n21356);
and_5  g19008(new_n6593, new_n6463, new_n21357);
and_5  g19009(new_n6627, new_n6594, new_n21358);
nor_5  g19010(new_n21358, new_n21357, new_n21359);
xor_4  g19011(new_n14320, new_n11530, new_n21360);
and_5  g19012(new_n21360, new_n21359, new_n21361);
not_10 g19013(new_n21361, new_n21362);
and_5  g19014(new_n21362, new_n21356, new_n21363);
nor_5  g19015(new_n21363, new_n21354, new_n21364);
nor_5  g19016(new_n21364, new_n21352, new_n21365_1);
nor_5  g19017(new_n21365_1, new_n21351, new_n21366);
nor_5  g19018(new_n21366, new_n21349_1, new_n21367_1);
nor_5  g19019(new_n21367_1, new_n21348, new_n21368);
nor_5  g19020(new_n21368, new_n21346, new_n21369);
xor_4  g19021(new_n21369, new_n21345, n7349);
xnor_4 g19022(new_n21312, new_n21260, n7363);
and_5  g19023(new_n4301, n16544, new_n21372);
not_10 g19024(new_n21372, new_n21373);
nor_5  g19025(new_n19994, new_n19991, new_n21374);
not_10 g19026(new_n21374, new_n21375);
and_5  g19027(new_n21375, new_n21373, new_n21376);
xor_4  g19028(new_n21376, new_n10389, new_n21377);
not_10 g19029(new_n21377, new_n21378);
nor_5  g19030(new_n19995, new_n10393, new_n21379);
nor_5  g19031(new_n20000, new_n19997, new_n21380);
nor_5  g19032(new_n21380, new_n21379, new_n21381);
xnor_4 g19033(new_n21381, new_n21378, n7390);
xor_4  g19034(new_n9263, new_n9261_1, n7403);
xor_4  g19035(new_n9456, new_n9413, n7408);
xnor_4 g19036(new_n20338, new_n20316, n7432);
nor_5  g19037(new_n18242, new_n15734, new_n21386);
nor_5  g19038(new_n18254_1, new_n18243, new_n21387);
or_5   g19039(new_n21387, new_n21386, n7475);
xor_4  g19040(new_n5231, new_n5229, n7477);
xnor_4 g19041(new_n9077, new_n9049, n7507);
or_5   g19042(new_n12195, new_n10538, new_n21391);
xor_4  g19043(new_n12195, n23895, new_n21392);
nand_5 g19044(new_n6877, n17351, new_n21393);
or_5   g19045(new_n6922, new_n6878, new_n21394);
and_5  g19046(new_n21394, new_n21393, new_n21395);
or_5   g19047(new_n21395, new_n21392, new_n21396_1);
and_5  g19048(new_n21396_1, new_n21391, new_n21397);
xor_4  g19049(new_n21397, new_n12241, new_n21398_1);
xnor_4 g19050(new_n21398_1, new_n17563, new_n21399_1);
not_10 g19051(new_n21399_1, new_n21400);
xor_4  g19052(new_n21395, new_n21392, new_n21401);
nor_5  g19053(new_n21401, new_n17569, new_n21402);
xnor_4 g19054(new_n21401, new_n17568, new_n21403);
not_10 g19055(new_n21403, new_n21404_1);
nor_5  g19056(new_n6923, new_n17572, new_n21405);
nor_5  g19057(new_n6993, new_n6925, new_n21406);
nor_5  g19058(new_n21406, new_n21405, new_n21407);
nor_5  g19059(new_n21407, new_n21404_1, new_n21408);
nor_5  g19060(new_n21408, new_n21402, new_n21409);
xnor_4 g19061(new_n21409, new_n21400, n7514);
xnor_4 g19062(new_n11062, new_n11033, n7558);
xnor_4 g19063(new_n12290, new_n12289, n7572);
xor_4  g19064(new_n6305, new_n4041, new_n21413);
or_5   g19065(new_n6306, new_n10513, new_n21414);
or_5   g19066(new_n20369, new_n20360, new_n21415);
and_5  g19067(new_n21415, new_n21414, new_n21416);
xor_4  g19068(new_n21416, new_n21413, new_n21417);
xor_4  g19069(new_n21417, new_n9908, new_n21418);
not_10 g19070(new_n21418, new_n21419);
nor_5  g19071(new_n20370, new_n9915, new_n21420);
nor_5  g19072(new_n20386, new_n20372, new_n21421);
nor_5  g19073(new_n21421, new_n21420, new_n21422);
xnor_4 g19074(new_n21422, new_n21419, n7575);
xor_4  g19075(new_n21145, new_n9852, new_n21424);
not_10 g19076(new_n21424, new_n21425);
nand_5 g19077(new_n21149, new_n9895, new_n21426);
xnor_4 g19078(new_n21149, new_n9895, new_n21427);
nand_5 g19079(new_n11085, new_n9899, new_n21428);
nand_5 g19080(new_n11117, new_n11086, new_n21429);
and_5  g19081(new_n21429, new_n21428, new_n21430);
or_5   g19082(new_n21430, new_n21427, new_n21431);
and_5  g19083(new_n21431, new_n21426, new_n21432);
xor_4  g19084(new_n21432, new_n21425, new_n21433);
xnor_4 g19085(new_n21433, new_n11722, new_n21434);
xor_4  g19086(new_n21430, new_n21427, new_n21435);
nand_5 g19087(new_n21435, new_n11729, new_n21436);
xor_4  g19088(new_n21435, new_n11729, new_n21437);
and_5  g19089(new_n11129, new_n11119, new_n21438);
not_10 g19090(new_n11165, new_n21439);
and_5  g19091(new_n21439, new_n11130, new_n21440);
nor_5  g19092(new_n21440, new_n21438, new_n21441);
nand_5 g19093(new_n21441, new_n21437, new_n21442);
and_5  g19094(new_n21442, new_n21436, new_n21443);
xor_4  g19095(new_n21443, new_n21434, n7585);
xor_4  g19096(new_n20860, new_n7832, new_n21445);
not_10 g19097(new_n21445, new_n21446_1);
nor_5  g19098(new_n20863, new_n7837, new_n21447);
xor_4  g19099(new_n20863, new_n7837, new_n21448);
not_10 g19100(new_n21448, new_n21449);
and_5  g19101(new_n20869_1, new_n7843, new_n21450);
xnor_4 g19102(new_n20869_1, new_n7842, new_n21451);
not_10 g19103(new_n21451, new_n21452);
nor_5  g19104(new_n20873, new_n7849, new_n21453);
xor_4  g19105(new_n20873, new_n7849, new_n21454);
not_10 g19106(new_n21454, new_n21455);
nor_5  g19107(new_n18336, new_n7854, new_n21456);
xor_4  g19108(new_n18336, new_n7854, new_n21457);
not_10 g19109(new_n21457, new_n21458);
nor_5  g19110(new_n18339, new_n7859, new_n21459);
xor_4  g19111(new_n18339, new_n7859, new_n21460);
not_10 g19112(new_n21460, new_n21461);
nor_5  g19113(new_n18344, new_n7864, new_n21462);
xor_4  g19114(new_n18344, new_n7864, new_n21463);
not_10 g19115(new_n7872, new_n21464);
nor_5  g19116(new_n18348, new_n21464, new_n21465);
xnor_4 g19117(new_n18348, new_n7872, new_n21466);
not_10 g19118(new_n21466, new_n21467);
nor_5  g19119(new_n18356, new_n7883, new_n21468);
not_10 g19120(new_n21468, new_n21469);
and_5  g19121(new_n21469, new_n7879, new_n21470);
xnor_4 g19122(new_n21468, new_n7879, new_n21471_1);
and_5  g19123(new_n21471_1, new_n18363, new_n21472_1);
nor_5  g19124(new_n21472_1, new_n21470, new_n21473);
nor_5  g19125(new_n21473, new_n21467, new_n21474);
nor_5  g19126(new_n21474, new_n21465, new_n21475);
not_10 g19127(new_n21475, new_n21476);
and_5  g19128(new_n21476, new_n21463, new_n21477);
nor_5  g19129(new_n21477, new_n21462, new_n21478);
nor_5  g19130(new_n21478, new_n21461, new_n21479);
nor_5  g19131(new_n21479, new_n21459, new_n21480);
nor_5  g19132(new_n21480, new_n21458, new_n21481);
nor_5  g19133(new_n21481, new_n21456, new_n21482);
nor_5  g19134(new_n21482, new_n21455, new_n21483);
nor_5  g19135(new_n21483, new_n21453, new_n21484);
nor_5  g19136(new_n21484, new_n21452, new_n21485);
nor_5  g19137(new_n21485, new_n21450, new_n21486);
nor_5  g19138(new_n21486, new_n21449, new_n21487);
nor_5  g19139(new_n21487, new_n21447, new_n21488);
xnor_4 g19140(new_n21488, new_n21446_1, n7588);
and_5  g19141(new_n6712, new_n2354, new_n21490);
and_5  g19142(new_n21490, new_n2350, new_n21491);
and_5  g19143(new_n21491, new_n11403_1, new_n21492);
and_5  g19144(new_n21492, new_n11400, new_n21493);
xor_4  g19145(new_n21493, new_n11982, new_n21494);
xor_4  g19146(new_n21494, new_n16340, new_n21495);
xor_4  g19147(new_n21492, new_n11400, new_n21496);
or_5   g19148(new_n21496, n11455, new_n21497);
xor_4  g19149(new_n21496, new_n16272, new_n21498);
xor_4  g19150(new_n21491, new_n11403_1, new_n21499);
or_5   g19151(new_n21499, n3945, new_n21500);
xor_4  g19152(new_n21499, new_n16275_1, new_n21501);
xor_4  g19153(new_n21490, new_n2350, new_n21502);
or_5   g19154(new_n21502, n5255, new_n21503);
xor_4  g19155(new_n21502, new_n16278, new_n21504);
or_5   g19156(new_n6713, n21649, new_n21505);
xor_4  g19157(new_n6713, new_n5179, new_n21506);
or_5   g19158(new_n6730, n18274, new_n21507);
nor_5  g19159(new_n6745, n3828, new_n21508);
xor_4  g19160(new_n6745, new_n5187, new_n21509);
or_5   g19161(new_n6740, n23842, new_n21510);
nand_5 g19162(n21654, n2387, new_n21511);
xor_4  g19163(new_n6740, n23842, new_n21512);
nand_5 g19164(new_n21512, new_n21511, new_n21513);
and_5  g19165(new_n21513, new_n21510, new_n21514);
nor_5  g19166(new_n21514, new_n21509, new_n21515);
or_5   g19167(new_n21515, new_n21508, new_n21516);
xor_4  g19168(new_n6730, n18274, new_n21517);
nand_5 g19169(new_n21517, new_n21516, new_n21518);
and_5  g19170(new_n21518, new_n21507, new_n21519);
or_5   g19171(new_n21519, new_n21506, new_n21520);
and_5  g19172(new_n21520, new_n21505, new_n21521);
or_5   g19173(new_n21521, new_n21504, new_n21522);
and_5  g19174(new_n21522, new_n21503, new_n21523);
or_5   g19175(new_n21523, new_n21501, new_n21524);
and_5  g19176(new_n21524, new_n21500, new_n21525_1);
or_5   g19177(new_n21525_1, new_n21498, new_n21526);
and_5  g19178(new_n21526, new_n21497, new_n21527);
xor_4  g19179(new_n21527, new_n21495, new_n21528);
xnor_4 g19180(new_n21528, new_n14666, new_n21529);
xor_4  g19181(new_n21525_1, new_n21498, new_n21530);
nand_5 g19182(new_n21530, new_n14709, new_n21531);
xor_4  g19183(new_n21530, new_n14709, new_n21532);
xor_4  g19184(new_n21523, new_n21501, new_n21533);
nor_5  g19185(new_n21533, new_n14712, new_n21534);
xnor_4 g19186(new_n21533, new_n14712, new_n21535);
xor_4  g19187(new_n21521, new_n21504, new_n21536);
or_5   g19188(new_n21536, new_n14717, new_n21537);
xor_4  g19189(new_n21519, new_n21506, new_n21538_1);
nor_5  g19190(new_n21538_1, new_n14721, new_n21539);
xor_4  g19191(new_n21517, new_n21516, new_n21540);
nor_5  g19192(new_n21540, new_n14725, new_n21541);
xor_4  g19193(new_n21540, new_n14724, new_n21542);
xnor_4 g19194(new_n21514, new_n21509, new_n21543);
nand_5 g19195(new_n21543, new_n14729, new_n21544);
xor_4  g19196(new_n21543, new_n14729, new_n21545);
or_5   g19197(new_n21512, new_n14732, new_n21546);
xor_4  g19198(new_n21512, new_n21511, new_n21547);
nor_5  g19199(new_n21547, new_n14734_1, new_n21548);
xor_4  g19200(n21654, n2387, new_n21549_1);
and_5  g19201(new_n21549_1, new_n14738, new_n21550);
or_5   g19202(new_n21550, new_n21548, new_n21551);
and_5  g19203(new_n21551, new_n21546, new_n21552);
nand_5 g19204(new_n21552, new_n21545, new_n21553);
and_5  g19205(new_n21553, new_n21544, new_n21554);
nor_5  g19206(new_n21554, new_n21542, new_n21555);
or_5   g19207(new_n21555, new_n21541, new_n21556);
xor_4  g19208(new_n21538_1, new_n14721, new_n21557);
and_5  g19209(new_n21557, new_n21556, new_n21558);
or_5   g19210(new_n21558, new_n21539, new_n21559);
xor_4  g19211(new_n21536, new_n14717, new_n21560);
nand_5 g19212(new_n21560, new_n21559, new_n21561);
and_5  g19213(new_n21561, new_n21537, new_n21562);
nor_5  g19214(new_n21562, new_n21535, new_n21563);
nor_5  g19215(new_n21563, new_n21534, new_n21564);
nand_5 g19216(new_n21564, new_n21532, new_n21565);
and_5  g19217(new_n21565, new_n21531, new_n21566);
xor_4  g19218(new_n21566, new_n21529, n7598);
xnor_4 g19219(new_n18252, new_n18248, n7607);
xnor_4 g19220(new_n5038, new_n5011_1, n7610);
xnor_4 g19221(new_n3378, new_n3366_1, n7616);
not_10 g19222(new_n16000, new_n21571);
xnor_4 g19223(n10514, n6105, new_n21572);
or_5   g19224(n18649, n3795, new_n21573);
xnor_4 g19225(n18649, n3795, new_n21574);
or_5   g19226(n25464, n6218, new_n21575);
xnor_4 g19227(n25464, n6218, new_n21576);
or_5   g19228(n20470, n4590, new_n21577);
xnor_4 g19229(n20470, n4590, new_n21578);
or_5   g19230(n26752, n21222, new_n21579);
xnor_4 g19231(n26752, n21222, new_n21580);
or_5   g19232(n9832, n6513, new_n21581);
xor_4  g19233(n9832, n6513, new_n21582);
nand_5 g19234(n3918, n1558, new_n21583);
or_5   g19235(n3918, n1558, new_n21584);
nor_5  g19236(n21749, n919, new_n21585);
nor_5  g19237(new_n16781, new_n16776, new_n21586);
nor_5  g19238(new_n21586, new_n21585, new_n21587);
nand_5 g19239(new_n21587, new_n21584, new_n21588);
and_5  g19240(new_n21588, new_n21583, new_n21589);
nand_5 g19241(new_n21589, new_n21582, new_n21590);
and_5  g19242(new_n21590, new_n21581, new_n21591);
or_5   g19243(new_n21591, new_n21580, new_n21592);
and_5  g19244(new_n21592, new_n21579, new_n21593);
or_5   g19245(new_n21593, new_n21578, new_n21594);
and_5  g19246(new_n21594, new_n21577, new_n21595);
or_5   g19247(new_n21595, new_n21576, new_n21596);
and_5  g19248(new_n21596, new_n21575, new_n21597);
or_5   g19249(new_n21597, new_n21574, new_n21598);
and_5  g19250(new_n21598, new_n21573, new_n21599_1);
xor_4  g19251(new_n21599_1, new_n21572, new_n21600);
nand_5 g19252(new_n21600, n9872, new_n21601);
xor_4  g19253(new_n21600, new_n21194, new_n21602);
xor_4  g19254(new_n21597, new_n21574, new_n21603);
nand_5 g19255(new_n21603, n5842, new_n21604);
xor_4  g19256(new_n21603, new_n21198, new_n21605);
xor_4  g19257(new_n21595, new_n21576, new_n21606);
nand_5 g19258(new_n21606, n6379, new_n21607);
xor_4  g19259(new_n21606, new_n21202, new_n21608);
xor_4  g19260(new_n21593, new_n21578, new_n21609);
nand_5 g19261(new_n21609, n2102, new_n21610);
xor_4  g19262(new_n21609, new_n21206, new_n21611);
xor_4  g19263(new_n21591, new_n21580, new_n21612);
nand_5 g19264(new_n21612, n17954, new_n21613);
xnor_4 g19265(new_n21612, n17954, new_n21614);
xor_4  g19266(new_n21589, new_n21582, new_n21615_1);
nand_5 g19267(new_n21615_1, n8256, new_n21616);
xor_4  g19268(new_n21615_1, new_n21212, new_n21617);
xor_4  g19269(n3918, n1558, new_n21618);
xor_4  g19270(new_n21618, new_n21587, new_n21619);
or_5   g19271(new_n21619, new_n21216, new_n21620);
xor_4  g19272(new_n21619, n24150, new_n21621);
nand_5 g19273(new_n16782, n19584, new_n21622);
nand_5 g19274(new_n16791, new_n16783, new_n21623);
and_5  g19275(new_n21623, new_n21622, new_n21624);
or_5   g19276(new_n21624, new_n21621, new_n21625);
and_5  g19277(new_n21625, new_n21620, new_n21626);
or_5   g19278(new_n21626, new_n21617, new_n21627);
and_5  g19279(new_n21627, new_n21616, new_n21628_1);
or_5   g19280(new_n21628_1, new_n21614, new_n21629);
and_5  g19281(new_n21629, new_n21613, new_n21630);
or_5   g19282(new_n21630, new_n21611, new_n21631);
and_5  g19283(new_n21631, new_n21610, new_n21632);
or_5   g19284(new_n21632, new_n21608, new_n21633);
and_5  g19285(new_n21633, new_n21607, new_n21634);
or_5   g19286(new_n21634, new_n21605, new_n21635);
and_5  g19287(new_n21635, new_n21604, new_n21636);
or_5   g19288(new_n21636, new_n21602, new_n21637_1);
and_5  g19289(new_n21637_1, new_n21601, new_n21638);
or_5   g19290(n10514, n6105, new_n21639);
or_5   g19291(new_n21599_1, new_n21572, new_n21640);
and_5  g19292(new_n21640, new_n21639, new_n21641);
nor_5  g19293(new_n21641, new_n21638, new_n21642);
xnor_4 g19294(new_n21642, new_n21571, new_n21643);
xor_4  g19295(new_n21641, new_n21638, new_n21644);
and_5  g19296(new_n21644, new_n15868, new_n21645_1);
xnor_4 g19297(new_n21644, new_n15869_1, new_n21646);
not_10 g19298(new_n15920, new_n21647);
xor_4  g19299(new_n21636, new_n21602, new_n21648);
and_5  g19300(new_n21648, new_n21647, new_n21649_1);
xnor_4 g19301(new_n21648, new_n15920, new_n21650);
xor_4  g19302(new_n21634, new_n21605, new_n21651);
and_5  g19303(new_n21651, new_n15927, new_n21652);
xor_4  g19304(new_n21651, new_n15927, new_n21653);
not_10 g19305(new_n21653, new_n21654_1);
xor_4  g19306(new_n21632, new_n21608, new_n21655);
nand_5 g19307(new_n21655, new_n15933, new_n21656);
xor_4  g19308(new_n21655, new_n15933, new_n21657);
xor_4  g19309(new_n21630, new_n21611, new_n21658);
nand_5 g19310(new_n21658, new_n15939, new_n21659);
xor_4  g19311(new_n21658, new_n15939, new_n21660);
xor_4  g19312(new_n21628_1, new_n21614, new_n21661);
not_10 g19313(new_n21661, new_n21662);
or_5   g19314(new_n21662, new_n15943, new_n21663);
xor_4  g19315(new_n21662, new_n15943, new_n21664);
xor_4  g19316(new_n21626, new_n21617, new_n21665_1);
nand_5 g19317(new_n21665_1, new_n15950, new_n21666);
xor_4  g19318(new_n21665_1, new_n15950, new_n21667);
xor_4  g19319(new_n21624, new_n21621, new_n21668);
nand_5 g19320(new_n21668, new_n15953, new_n21669);
xor_4  g19321(new_n21668, new_n15953, new_n21670);
not_10 g19322(new_n21670, new_n21671);
nand_5 g19323(new_n16792, new_n15970, new_n21672);
nand_5 g19324(new_n16800, new_n16793, new_n21673);
and_5  g19325(new_n21673, new_n21672, new_n21674_1);
or_5   g19326(new_n21674_1, new_n21671, new_n21675);
nand_5 g19327(new_n21675, new_n21669, new_n21676);
nand_5 g19328(new_n21676, new_n21667, new_n21677);
nand_5 g19329(new_n21677, new_n21666, new_n21678);
nand_5 g19330(new_n21678, new_n21664, new_n21679);
nand_5 g19331(new_n21679, new_n21663, new_n21680_1);
nand_5 g19332(new_n21680_1, new_n21660, new_n21681);
nand_5 g19333(new_n21681, new_n21659, new_n21682);
nand_5 g19334(new_n21682, new_n21657, new_n21683);
and_5  g19335(new_n21683, new_n21656, new_n21684);
nor_5  g19336(new_n21684, new_n21654_1, new_n21685_1);
nor_5  g19337(new_n21685_1, new_n21652, new_n21686);
not_10 g19338(new_n21686, new_n21687_1);
and_5  g19339(new_n21687_1, new_n21650, new_n21688);
nor_5  g19340(new_n21688, new_n21649_1, new_n21689);
not_10 g19341(new_n21689, new_n21690);
and_5  g19342(new_n21690, new_n21646, new_n21691);
nor_5  g19343(new_n21691, new_n21645_1, new_n21692);
xor_4  g19344(new_n21692, new_n21643, n7630);
or_5   g19345(new_n19135, new_n19106, new_n21694);
not_10 g19346(new_n19136, new_n21695);
or_5   g19347(new_n19145, new_n21695, new_n21696);
and_5  g19348(new_n21696, new_n21694, n7643);
xnor_4 g19349(new_n12425, new_n12397_1, n7647);
xnor_4 g19350(new_n10246, new_n10207, n7679);
xnor_4 g19351(new_n20556, new_n20531, n7686);
xor_4  g19352(new_n18602, new_n18578_1, new_n21701);
xor_4  g19353(new_n21701, new_n18620, n7698);
xor_4  g19354(new_n19792_1, new_n19769, n7708);
xor_4  g19355(new_n18592, n3324, new_n21704);
not_10 g19356(n17911, new_n21705);
or_5   g19357(new_n2913, new_n21705, new_n21706);
xor_4  g19358(new_n2913, new_n21705, new_n21707);
nand_5 g19359(new_n2953, new_n19296, new_n21708);
xor_4  g19360(new_n2953, n21997, new_n21709);
nand_5 g19361(new_n2958, new_n8652, new_n21710);
nand_5 g19362(new_n8679, new_n8653, new_n21711);
and_5  g19363(new_n21711, new_n21710, new_n21712);
or_5   g19364(new_n21712, new_n21709, new_n21713);
and_5  g19365(new_n21713, new_n21708, new_n21714);
nand_5 g19366(new_n21714, new_n21707, new_n21715);
and_5  g19367(new_n21715, new_n21706, new_n21716);
xor_4  g19368(new_n21716, new_n21704, new_n21717_1);
not_10 g19369(new_n21717_1, new_n21718);
xor_4  g19370(new_n6070, new_n4919, new_n21719_1);
nand_5 g19371(new_n6074, new_n4923, new_n21720);
nand_5 g19372(new_n16548, new_n16540, new_n21721);
and_5  g19373(new_n21721, new_n21720, new_n21722);
xor_4  g19374(new_n21722, new_n21719_1, new_n21723);
not_10 g19375(new_n21723, new_n21724);
xor_4  g19376(new_n21724, new_n21718, new_n21725);
xor_4  g19377(new_n21714, new_n21707, new_n21726);
nor_5  g19378(new_n21726, new_n16549, new_n21727);
xor_4  g19379(new_n21726, new_n16549, new_n21728);
not_10 g19380(new_n21728, new_n21729);
xor_4  g19381(new_n21712, new_n21709, new_n21730);
and_5  g19382(new_n21730, new_n16551, new_n21731);
xor_4  g19383(new_n21730, new_n16551, new_n21732);
not_10 g19384(new_n21732, new_n21733);
and_5  g19385(new_n8680, new_n8651, new_n21734);
nor_5  g19386(new_n8728, new_n8682, new_n21735_1);
nor_5  g19387(new_n21735_1, new_n21734, new_n21736);
nor_5  g19388(new_n21736, new_n21733, new_n21737);
nor_5  g19389(new_n21737, new_n21731, new_n21738);
nor_5  g19390(new_n21738, new_n21729, new_n21739);
nor_5  g19391(new_n21739, new_n21727, new_n21740);
not_10 g19392(new_n21740, new_n21741);
xnor_4 g19393(new_n21741, new_n21725, n7780);
or_5   g19394(new_n2592, new_n5537, new_n21743);
xor_4  g19395(new_n2592, new_n5537, new_n21744);
not_10 g19396(new_n21744, new_n21745);
or_5   g19397(new_n2596, new_n9811, new_n21746);
or_5   g19398(new_n9851, new_n9813, new_n21747);
and_5  g19399(new_n21747, new_n21746, new_n21748);
or_5   g19400(new_n21748, new_n21745, new_n21749_1);
and_5  g19401(new_n21749_1, new_n21743, new_n21750_1);
xnor_4 g19402(new_n21750_1, new_n14945, new_n21751);
not_10 g19403(new_n21751, new_n21752);
and_5  g19404(new_n17656, new_n2709, new_n21753_1);
xor_4  g19405(new_n17656, new_n2710, new_n21754);
nand_5 g19406(new_n9858, new_n2713, new_n21755);
or_5   g19407(new_n9892, new_n9859, new_n21756);
and_5  g19408(new_n21756, new_n21755, new_n21757);
nor_5  g19409(new_n21757, new_n21754, new_n21758);
nor_5  g19410(new_n21758, new_n21753_1, new_n21759);
not_10 g19411(new_n21759, new_n21760);
and_5  g19412(new_n17655, new_n4301, new_n21761);
xor_4  g19413(new_n21761, new_n10338, new_n21762);
xor_4  g19414(new_n21762, new_n21760, new_n21763);
xnor_4 g19415(new_n21763, new_n21752, new_n21764);
xor_4  g19416(new_n21748, new_n21745, new_n21765_1);
xor_4  g19417(new_n21757, new_n21754, new_n21766);
nor_5  g19418(new_n21766, new_n21765_1, new_n21767);
xor_4  g19419(new_n21766, new_n21765_1, new_n21768);
not_10 g19420(new_n21768, new_n21769);
nor_5  g19421(new_n9893, new_n9852, new_n21770);
not_10 g19422(new_n21770, new_n21771);
and_5  g19423(new_n9945, new_n9894, new_n21772);
not_10 g19424(new_n21772, new_n21773);
and_5  g19425(new_n21773, new_n21771, new_n21774);
nor_5  g19426(new_n21774, new_n21769, new_n21775);
nor_5  g19427(new_n21775, new_n21767, new_n21776);
not_10 g19428(new_n21776, new_n21777);
xnor_4 g19429(new_n21777, new_n21764, n7794);
xnor_4 g19430(new_n17839, new_n17834, n7811);
xor_4  g19431(new_n17781, new_n17776, n7830);
xnor_4 g19432(new_n21484, new_n21452, n7834);
xnor_4 g19433(new_n11158, new_n11144, n7884);
xor_4  g19434(new_n3056, new_n18219, n7937);
xnor_4 g19435(new_n3071, new_n3016, n7943);
xor_4  g19436(new_n9939, new_n9907, n7950);
xnor_4 g19437(new_n20048, new_n15816_1, new_n21786);
and_5  g19438(new_n20053, new_n15818, new_n21787);
nor_5  g19439(new_n20055, new_n15822, new_n21788);
xnor_4 g19440(new_n20055, new_n15821, new_n21789);
not_10 g19441(new_n21789, new_n21790);
and_5  g19442(new_n15567, new_n15521, new_n21791);
nor_5  g19443(new_n15613, new_n15569, new_n21792);
nor_5  g19444(new_n21792, new_n21791, new_n21793);
nor_5  g19445(new_n21793, new_n21790, new_n21794);
nor_5  g19446(new_n21794, new_n21788, new_n21795);
xor_4  g19447(new_n20053, new_n15818, new_n21796);
not_10 g19448(new_n21796, new_n21797);
nor_5  g19449(new_n21797, new_n21795, new_n21798);
nor_5  g19450(new_n21798, new_n21787, new_n21799);
xor_4  g19451(new_n21799, new_n21786, n7959);
xnor_4 g19452(new_n17843, new_n17827, n7968);
xnor_4 g19453(new_n18856, new_n18854, n7992);
xor_4  g19454(new_n13159, n9554, new_n21803);
nand_5 g19455(new_n13162, n26408, new_n21804);
xor_4  g19456(new_n13162, n26408, new_n21805);
nand_5 g19457(new_n10760, new_n7910, new_n21806);
nand_5 g19458(new_n17813, new_n17802, new_n21807);
and_5  g19459(new_n21807, new_n21806, new_n21808);
nand_5 g19460(new_n21808, new_n21805, new_n21809);
and_5  g19461(new_n21809, new_n21804, new_n21810);
xor_4  g19462(new_n21810, new_n21803, new_n21811);
xor_4  g19463(new_n21811, new_n19023, new_n21812);
not_10 g19464(new_n21812, new_n21813);
xor_4  g19465(new_n21808, new_n21805, new_n21814);
and_5  g19466(new_n21814, new_n19028, new_n21815);
xor_4  g19467(new_n21814, new_n19028, new_n21816);
not_10 g19468(new_n21816, new_n21817);
not_10 g19469(new_n17814, new_n21818);
and_5  g19470(new_n19033_1, new_n21818, new_n21819);
not_10 g19471(new_n21819, new_n21820_1);
xor_4  g19472(new_n19033_1, new_n21818, new_n21821);
and_5  g19473(new_n19039, new_n17817, new_n21822);
xor_4  g19474(new_n19039, new_n17817, new_n21823);
not_10 g19475(new_n21823, new_n21824);
and_5  g19476(new_n19047, new_n17821, new_n21825);
xor_4  g19477(new_n19047, new_n17821, new_n21826);
not_10 g19478(new_n21826, new_n21827);
and_5  g19479(new_n13258, new_n13247, new_n21828);
nor_5  g19480(new_n13265, new_n13260, new_n21829);
nor_5  g19481(new_n21829, new_n21828, new_n21830);
nor_5  g19482(new_n21830, new_n21827, new_n21831);
nor_5  g19483(new_n21831, new_n21825, new_n21832_1);
nor_5  g19484(new_n21832_1, new_n21824, new_n21833);
nor_5  g19485(new_n21833, new_n21822, new_n21834);
not_10 g19486(new_n21834, new_n21835);
and_5  g19487(new_n21835, new_n21821, new_n21836);
not_10 g19488(new_n21836, new_n21837);
and_5  g19489(new_n21837, new_n21820_1, new_n21838);
nor_5  g19490(new_n21838, new_n21817, new_n21839_1);
nor_5  g19491(new_n21839_1, new_n21815, new_n21840);
xnor_4 g19492(new_n21840, new_n21813, n7999);
xnor_4 g19493(new_n18480, new_n18466, n8027);
not_10 g19494(new_n14945, new_n21843);
nor_5  g19495(new_n21750_1, new_n21843, new_n21844);
nand_5 g19496(new_n6278, n8614, new_n21845);
xor_4  g19497(new_n6278, new_n5480, new_n21846);
nand_5 g19498(new_n6285, n15182, new_n21847);
or_5   g19499(new_n6292, n27037, new_n21848);
xor_4  g19500(new_n6292, new_n10512, new_n21849);
or_5   g19501(new_n6296, n8964, new_n21850);
xor_4  g19502(new_n6296, n8964, new_n21851);
nand_5 g19503(new_n6300, n20151, new_n21852);
and_5  g19504(new_n6305, n7693, new_n21853);
nor_5  g19505(new_n21416, new_n21413, new_n21854);
or_5   g19506(new_n21854, new_n21853, new_n21855);
xor_4  g19507(new_n6300, n20151, new_n21856);
nand_5 g19508(new_n21856, new_n21855, new_n21857);
and_5  g19509(new_n21857, new_n21852, new_n21858);
nand_5 g19510(new_n21858, new_n21851, new_n21859);
and_5  g19511(new_n21859, new_n21850, new_n21860);
or_5   g19512(new_n21860, new_n21849, new_n21861);
and_5  g19513(new_n21861, new_n21848, new_n21862);
xor_4  g19514(new_n6285, n15182, new_n21863);
nand_5 g19515(new_n21863, new_n21862, new_n21864);
and_5  g19516(new_n21864, new_n21847, new_n21865);
or_5   g19517(new_n21865, new_n21846, new_n21866);
and_5  g19518(new_n21866, new_n21845, new_n21867);
nor_5  g19519(new_n21867, new_n6235, new_n21868);
not_10 g19520(new_n21868, new_n21869);
and_5  g19521(new_n21869, new_n21844, new_n21870);
not_10 g19522(new_n21844, new_n21871);
and_5  g19523(new_n21868, new_n21871, new_n21872);
xor_4  g19524(new_n21867, new_n6235, new_n21873);
nor_5  g19525(new_n21873, new_n21752, new_n21874_1);
xnor_4 g19526(new_n21873, new_n21751, new_n21875);
not_10 g19527(new_n21875, new_n21876);
xnor_4 g19528(new_n21865, new_n21846, new_n21877);
and_5  g19529(new_n21877, new_n21765_1, new_n21878);
xor_4  g19530(new_n21877, new_n21765_1, new_n21879);
not_10 g19531(new_n21879, new_n21880);
xnor_4 g19532(new_n21863, new_n21862, new_n21881);
and_5  g19533(new_n21881, new_n9852, new_n21882);
xor_4  g19534(new_n21881, new_n9852, new_n21883);
not_10 g19535(new_n21883, new_n21884);
xor_4  g19536(new_n21860, new_n21849, new_n21885);
and_5  g19537(new_n21885, new_n9895, new_n21886);
xor_4  g19538(new_n21885, new_n9895, new_n21887);
not_10 g19539(new_n21887, new_n21888);
xor_4  g19540(new_n21858, new_n21851, new_n21889);
and_5  g19541(new_n21889, new_n9899, new_n21890);
xor_4  g19542(new_n21889, new_n9899, new_n21891);
not_10 g19543(new_n21891, new_n21892);
xor_4  g19544(new_n21856, new_n21855, new_n21893);
nor_5  g19545(new_n21893, new_n9904, new_n21894);
xor_4  g19546(new_n21893, new_n9904, new_n21895);
not_10 g19547(new_n21895, new_n21896);
nor_5  g19548(new_n21417, new_n9908, new_n21897);
nor_5  g19549(new_n21422, new_n21419, new_n21898_1);
nor_5  g19550(new_n21898_1, new_n21897, new_n21899);
nor_5  g19551(new_n21899, new_n21896, new_n21900);
nor_5  g19552(new_n21900, new_n21894, new_n21901);
nor_5  g19553(new_n21901, new_n21892, new_n21902);
nor_5  g19554(new_n21902, new_n21890, new_n21903);
nor_5  g19555(new_n21903, new_n21888, new_n21904);
nor_5  g19556(new_n21904, new_n21886, new_n21905_1);
nor_5  g19557(new_n21905_1, new_n21884, new_n21906);
nor_5  g19558(new_n21906, new_n21882, new_n21907);
nor_5  g19559(new_n21907, new_n21880, new_n21908);
nor_5  g19560(new_n21908, new_n21878, new_n21909);
nor_5  g19561(new_n21909, new_n21876, new_n21910);
nor_5  g19562(new_n21910, new_n21874_1, new_n21911);
nor_5  g19563(new_n21911, new_n21872, new_n21912);
or_5   g19564(new_n21912, new_n21870, n8031);
nand_5 g19565(new_n17656, n22626, new_n21914);
not_10 g19566(new_n21761, new_n21915_1);
or_5   g19567(new_n17656, n22626, new_n21916);
nand_5 g19568(new_n17665, new_n21916, new_n21917);
and_5  g19569(new_n21917, new_n21915_1, new_n21918);
and_5  g19570(new_n21918, new_n21914, new_n21919);
and_5  g19571(new_n21919, new_n20217, new_n21920);
xnor_4 g19572(new_n21919, new_n20217, new_n21921);
or_5   g19573(new_n17667, new_n17654, new_n21922);
nand_5 g19574(new_n17696, new_n17668, new_n21923);
and_5  g19575(new_n21923, new_n21922, new_n21924);
nor_5  g19576(new_n21924, new_n21921, new_n21925);
nor_5  g19577(new_n21925, new_n21920, new_n21926);
nor_5  g19578(new_n17706, n9554, new_n21927);
not_10 g19579(new_n17738_1, new_n21928);
nor_5  g19580(new_n21928, new_n21927, new_n21929);
not_10 g19581(new_n21929, new_n21930);
and_5  g19582(new_n17706, n9554, new_n21931);
nor_5  g19583(new_n21931, new_n20504, new_n21932);
and_5  g19584(new_n21932, new_n21930, new_n21933);
not_10 g19585(new_n21933, new_n21934_1);
nand_5 g19586(new_n21934_1, new_n21926, new_n21935);
xor_4  g19587(new_n21933, new_n21926, new_n21936);
xor_4  g19588(new_n21924, new_n21921, new_n21937);
or_5   g19589(new_n21937, new_n21934_1, new_n21938);
xor_4  g19590(new_n21937, new_n21933, new_n21939);
or_5   g19591(new_n17739, new_n17697, new_n21940);
nand_5 g19592(new_n17800, new_n17740, new_n21941);
and_5  g19593(new_n21941, new_n21940, new_n21942);
or_5   g19594(new_n21942, new_n21939, new_n21943_1);
and_5  g19595(new_n21943_1, new_n21938, new_n21944);
or_5   g19596(new_n21944, new_n21936, new_n21945);
and_5  g19597(new_n21945, new_n21935, n8042);
and_5  g19598(new_n10169, new_n10079, new_n21947);
nor_5  g19599(new_n10261_1, new_n10171, new_n21948);
or_5   g19600(new_n21948, new_n21947, n8095);
and_5  g19601(n23166, new_n9291, new_n21950);
not_10 g19602(new_n21950, new_n21951);
xor_4  g19603(n23166, n4306, new_n21952);
or_5   g19604(new_n9309, n3279, new_n21953);
xor_4  g19605(n10577, n3279, new_n21954);
or_5   g19606(n13914, new_n9312, new_n21955);
xor_4  g19607(n13914, n6381, new_n21956);
or_5   g19608(n14702, new_n9315, new_n21957_1);
or_5   g19609(new_n19953, new_n19942, new_n21958);
and_5  g19610(new_n21958, new_n21957_1, new_n21959);
or_5   g19611(new_n21959, new_n21956, new_n21960_1);
and_5  g19612(new_n21960_1, new_n21955, new_n21961);
or_5   g19613(new_n21961, new_n21954, new_n21962);
and_5  g19614(new_n21962, new_n21953, new_n21963);
nor_5  g19615(new_n21963, new_n21952, new_n21964);
not_10 g19616(new_n21964, new_n21965);
and_5  g19617(new_n21965, new_n21951, new_n21966);
xor_4  g19618(new_n21966, new_n9140, new_n21967);
xor_4  g19619(new_n21963, new_n21952, new_n21968);
nor_5  g19620(new_n21968, new_n9202, new_n21969);
xor_4  g19621(new_n21968, new_n9202, new_n21970);
not_10 g19622(new_n21970, new_n21971);
xor_4  g19623(new_n21961, new_n21954, new_n21972);
nor_5  g19624(new_n21972, new_n9208, new_n21973);
not_10 g19625(new_n21973, new_n21974);
xor_4  g19626(new_n21972, new_n9208, new_n21975);
xor_4  g19627(new_n21959, new_n21956, new_n21976_1);
nor_5  g19628(new_n21976_1, new_n9214, new_n21977);
not_10 g19629(new_n21977, new_n21978);
xor_4  g19630(new_n21976_1, new_n9214, new_n21979);
and_5  g19631(new_n19954, new_n9220_1, new_n21980);
and_5  g19632(new_n19968_1, new_n19955, new_n21981_1);
nor_5  g19633(new_n21981_1, new_n21980, new_n21982);
and_5  g19634(new_n21982, new_n21979, new_n21983);
not_10 g19635(new_n21983, new_n21984);
and_5  g19636(new_n21984, new_n21978, new_n21985);
not_10 g19637(new_n21985, new_n21986_1);
and_5  g19638(new_n21986_1, new_n21975, new_n21987);
not_10 g19639(new_n21987, new_n21988);
and_5  g19640(new_n21988, new_n21974, new_n21989);
nor_5  g19641(new_n21989, new_n21971, new_n21990);
nor_5  g19642(new_n21990, new_n21969, new_n21991);
not_10 g19643(new_n21991, new_n21992);
xnor_4 g19644(new_n21992, new_n21967, n8103);
xnor_4 g19645(new_n19291, new_n19273, n8109);
and_5  g19646(new_n19755, new_n19739, new_n21995);
nor_5  g19647(new_n19798_1, new_n19757, new_n21996);
or_5   g19648(new_n21996, new_n21995, n8127);
xor_4  g19649(new_n17179, new_n17174, n8130);
and_5  g19650(new_n3409, n4319, new_n21999);
xor_4  g19651(n8856, n4319, new_n22000);
or_5   g19652(new_n11982, n14130, new_n22001);
xor_4  g19653(n23463, n14130, new_n22002);
or_5   g19654(n16482, new_n11400, new_n22003);
xor_4  g19655(n16482, n13074, new_n22004);
or_5   g19656(new_n11403_1, n9942, new_n22005);
not_10 g19657(new_n2349, new_n22006);
or_5   g19658(new_n2382, new_n22006, new_n22007);
and_5  g19659(new_n22007, new_n22005, new_n22008);
or_5   g19660(new_n22008, new_n22004, new_n22009);
and_5  g19661(new_n22009, new_n22003, new_n22010);
or_5   g19662(new_n22010, new_n22002, new_n22011);
and_5  g19663(new_n22011, new_n22001, new_n22012);
nor_5  g19664(new_n22012, new_n22000, new_n22013);
nor_5  g19665(new_n22013, new_n21999, new_n22014);
xor_4  g19666(new_n22014, new_n7644, new_n22015);
nor_5  g19667(new_n22014, new_n7647_1, new_n22016_1);
xor_4  g19668(new_n22014, new_n7647_1, new_n22017);
not_10 g19669(new_n22017, new_n22018);
xor_4  g19670(new_n22012, new_n22000, new_n22019);
nor_5  g19671(new_n22019, new_n7653, new_n22020);
xor_4  g19672(new_n22019, new_n7653, new_n22021);
xor_4  g19673(new_n22010, new_n22002, new_n22022);
nor_5  g19674(new_n22022, new_n7658, new_n22023);
xor_4  g19675(new_n22022, new_n7658, new_n22024);
xor_4  g19676(new_n22008, new_n22004, new_n22025);
and_5  g19677(new_n22025, new_n7663, new_n22026);
xnor_4 g19678(new_n22025, new_n7663, new_n22027_1);
or_5   g19679(new_n2501, new_n2383, new_n22028);
nand_5 g19680(new_n2544, new_n2502, new_n22029);
and_5  g19681(new_n22029, new_n22028, new_n22030);
nor_5  g19682(new_n22030, new_n22027_1, new_n22031);
nor_5  g19683(new_n22031, new_n22026, new_n22032);
and_5  g19684(new_n22032, new_n22024, new_n22033);
nor_5  g19685(new_n22033, new_n22023, new_n22034);
not_10 g19686(new_n22034, new_n22035);
and_5  g19687(new_n22035, new_n22021, new_n22036);
nor_5  g19688(new_n22036, new_n22020, new_n22037);
nor_5  g19689(new_n22037, new_n22018, new_n22038);
nor_5  g19690(new_n22038, new_n22016_1, new_n22039);
xor_4  g19691(new_n22039, new_n22015, n8135);
xnor_4 g19692(new_n7696, new_n2533_1, n8139);
not_10 g19693(n26660, new_n22042);
and_5  g19694(new_n18628, new_n10855, new_n22043_1);
and_5  g19695(new_n22043_1, new_n22042, new_n22044);
xor_4  g19696(new_n22044, new_n10834_1, new_n22045);
xor_4  g19697(new_n22045, new_n2960, new_n22046);
xor_4  g19698(new_n22043_1, new_n22042, new_n22047);
nand_5 g19699(new_n22047, new_n2965, new_n22048);
xor_4  g19700(new_n22047, new_n2966, new_n22049);
nand_5 g19701(new_n18629, new_n2971_1, new_n22050_1);
nand_5 g19702(new_n18646, new_n18630, new_n22051);
and_5  g19703(new_n22051, new_n22050_1, new_n22052);
or_5   g19704(new_n22052, new_n22049, new_n22053);
and_5  g19705(new_n22053, new_n22048, new_n22054);
xor_4  g19706(new_n22054, new_n22046, new_n22055);
xor_4  g19707(new_n22055, new_n6934, new_n22056);
not_10 g19708(new_n22056, new_n22057);
xor_4  g19709(new_n22052, new_n22049, new_n22058);
nor_5  g19710(new_n22058, new_n6940, new_n22059);
xor_4  g19711(new_n22058, new_n6940, new_n22060);
not_10 g19712(new_n22060, new_n22061);
and_5  g19713(new_n18647, new_n6944, new_n22062);
nor_5  g19714(new_n18669, new_n18649_1, new_n22063_1);
nor_5  g19715(new_n22063_1, new_n22062, new_n22064);
nor_5  g19716(new_n22064, new_n22061, new_n22065);
nor_5  g19717(new_n22065, new_n22059, new_n22066);
xnor_4 g19718(new_n22066, new_n22057, n8148);
xor_4  g19719(new_n18007, new_n18006, n8149);
xnor_4 g19720(new_n3928, new_n3911, n8159);
xor_4  g19721(new_n11922, new_n11921, n8179);
xor_4  g19722(new_n15219, new_n15214, n8215);
xnor_4 g19723(new_n19289, new_n19277, n8267);
xnor_4 g19724(new_n20381, new_n20380, n8276);
not_10 g19725(new_n17510, new_n22074);
not_10 g19726(n14440, new_n22075);
and_5  g19727(new_n22044, new_n10834_1, new_n22076_1);
and_5  g19728(new_n22076_1, new_n16163, new_n22077);
and_5  g19729(new_n22077, new_n22075, new_n22078);
xor_4  g19730(new_n22078, new_n7728, new_n22079);
nor_5  g19731(new_n22079, new_n15402, new_n22080);
not_10 g19732(new_n22080, new_n22081);
xnor_4 g19733(new_n22079, new_n15402, new_n22082);
xor_4  g19734(new_n22077, new_n22075, new_n22083);
or_5   g19735(new_n22083, new_n2951, new_n22084);
xnor_4 g19736(new_n22083, new_n15418, new_n22085);
xor_4  g19737(new_n22076_1, new_n16163, new_n22086);
nand_5 g19738(new_n22086, new_n2954, new_n22087);
and_5  g19739(new_n22045, new_n2959, new_n22088);
nor_5  g19740(new_n22054, new_n22046, new_n22089);
or_5   g19741(new_n22089, new_n22088, new_n22090_1);
xnor_4 g19742(new_n22086, new_n2955, new_n22091);
nand_5 g19743(new_n22091, new_n22090_1, new_n22092);
and_5  g19744(new_n22092, new_n22087, new_n22093);
nand_5 g19745(new_n22093, new_n22085, new_n22094);
and_5  g19746(new_n22094, new_n22084, new_n22095);
nor_5  g19747(new_n22095, new_n22082, new_n22096);
not_10 g19748(new_n22096, new_n22097);
and_5  g19749(new_n22097, new_n22081, new_n22098);
and_5  g19750(new_n22078, new_n7728, new_n22099);
xor_4  g19751(new_n22099, new_n15427, new_n22100);
xor_4  g19752(new_n22100, new_n22098, new_n22101);
nor_5  g19753(new_n22101, new_n17563, new_n22102);
xnor_4 g19754(new_n22101, new_n17564, new_n22103);
xor_4  g19755(new_n22095, new_n22082, new_n22104);
and_5  g19756(new_n22104, new_n17569, new_n22105);
xnor_4 g19757(new_n22104, new_n17568, new_n22106);
xor_4  g19758(new_n22093, new_n22085, new_n22107_1);
and_5  g19759(new_n22107_1, new_n17572, new_n22108);
xor_4  g19760(new_n22091, new_n22090_1, new_n22109);
nor_5  g19761(new_n22109, new_n6928, new_n22110);
xor_4  g19762(new_n22109, new_n6928, new_n22111);
not_10 g19763(new_n22111, new_n22112);
nor_5  g19764(new_n22055, new_n6934, new_n22113_1);
nor_5  g19765(new_n22066, new_n22057, new_n22114);
nor_5  g19766(new_n22114, new_n22113_1, new_n22115);
nor_5  g19767(new_n22115, new_n22112, new_n22116);
or_5   g19768(new_n22116, new_n22110, new_n22117);
xnor_4 g19769(new_n22107_1, new_n6847, new_n22118);
and_5  g19770(new_n22118, new_n22117, new_n22119);
nor_5  g19771(new_n22119, new_n22108, new_n22120);
not_10 g19772(new_n22120, new_n22121);
and_5  g19773(new_n22121, new_n22106, new_n22122);
nor_5  g19774(new_n22122, new_n22105, new_n22123);
not_10 g19775(new_n22123, new_n22124_1);
and_5  g19776(new_n22124_1, new_n22103, new_n22125);
nor_5  g19777(new_n22125, new_n22102, new_n22126_1);
not_10 g19778(new_n22126_1, new_n22127);
or_5   g19779(new_n22127, new_n22074, new_n22128);
not_10 g19780(new_n22098, new_n22129);
not_10 g19781(new_n22099, new_n22130_1);
and_5  g19782(new_n22130_1, new_n15427, new_n22131);
and_5  g19783(new_n22131, new_n22129, new_n22132);
and_5  g19784(new_n22127, new_n22074, new_n22133);
nor_5  g19785(new_n22130_1, new_n15427, new_n22134);
nand_5 g19786(new_n22134, new_n22098, new_n22135);
and_5  g19787(new_n22135, new_n22133, new_n22136);
or_5   g19788(new_n22136, new_n22132, new_n22137);
and_5  g19789(new_n22137, new_n22128, n8288);
xor_4  g19790(new_n11456, new_n7467, n8306);
xor_4  g19791(new_n8042_1, new_n7995, n8320);
xnor_4 g19792(new_n12757, new_n12736, n8321);
xor_4  g19793(new_n16744, new_n16730, n8339);
xor_4  g19794(new_n9278, new_n9217_1, n8376);
xor_4  g19795(new_n19616, new_n10432_1, n8408);
xor_4  g19796(new_n14738, new_n14737, n8417);
xnor_4 g19797(new_n13210, new_n13191, n8432);
nand_5 g19798(new_n10337, new_n10336, new_n22147);
and_5  g19799(new_n22147, new_n10335, new_n22148);
nor_5  g19800(new_n10388_1, new_n10339, new_n22149);
nor_5  g19801(new_n22149, new_n22148, new_n22150_1);
nor_5  g19802(new_n22150_1, new_n10315, new_n22151);
nor_5  g19803(new_n10389, new_n10314, new_n22152);
nor_5  g19804(new_n10465, new_n10391, new_n22153);
nor_5  g19805(new_n22153, new_n22152, new_n22154);
or_5   g19806(new_n22154, new_n22151, new_n22155);
and_5  g19807(new_n22150_1, new_n10315, new_n22156);
or_5   g19808(new_n22156, new_n22153, new_n22157_1);
and_5  g19809(new_n22157_1, new_n22155, n8453);
xor_4  g19810(new_n16010, new_n16008, n8480);
xnor_4 g19811(new_n16911_1, new_n16886, n8489);
xor_4  g19812(new_n22034, new_n22021, n8505);
xnor_4 g19813(new_n20066, new_n20050, n8510);
xor_4  g19814(new_n12416, new_n17996, n8519);
xnor_4 g19815(new_n9931, new_n9929, n8535);
xor_4  g19816(new_n19784, new_n19781, n8550);
xnor_4 g19817(new_n20972, new_n20964, n8563);
xnor_4 g19818(new_n13653, new_n13651, n8594);
xnor_4 g19819(new_n6977, new_n6953, n8608);
xor_4  g19820(new_n4580, new_n4579, n8620);
xor_4  g19821(new_n7500, new_n7429, n8637);
xor_4  g19822(new_n17582, new_n17581, n8662);
xnor_4 g19823(new_n19338, new_n19329, n8716);
xor_4  g19824(new_n7999_1, new_n7997, new_n22173_1);
xor_4  g19825(new_n22173_1, new_n8040, n8744);
or_5   g19826(new_n13159, new_n7908, new_n22175);
or_5   g19827(new_n21810, new_n21803, new_n22176);
and_5  g19828(new_n22176, new_n22175, new_n22177);
xnor_4 g19829(new_n22177, new_n15732, new_n22178);
or_5   g19830(new_n6070, new_n4919, new_n22179);
nand_5 g19831(new_n21722, new_n21719_1, new_n22180);
and_5  g19832(new_n22180, new_n22179, new_n22181);
xnor_4 g19833(new_n22181, new_n18241_1, new_n22182);
xnor_4 g19834(new_n22182, new_n22178, new_n22183);
not_10 g19835(new_n22183, new_n22184);
and_5  g19836(new_n21811, new_n21724, new_n22185);
not_10 g19837(new_n22185, new_n22186);
xnor_4 g19838(new_n21811, new_n21723, new_n22187);
nor_5  g19839(new_n21814, new_n16549, new_n22188);
xor_4  g19840(new_n21814, new_n16549, new_n22189);
or_5   g19841(new_n17814, new_n16551, new_n22190);
or_5   g19842(new_n17849, new_n17816, new_n22191);
and_5  g19843(new_n22191, new_n22190, new_n22192);
and_5  g19844(new_n22192, new_n22189, new_n22193);
nor_5  g19845(new_n22193, new_n22188, new_n22194);
and_5  g19846(new_n22194, new_n22187, new_n22195);
not_10 g19847(new_n22195, new_n22196);
and_5  g19848(new_n22196, new_n22186, new_n22197);
xnor_4 g19849(new_n22197, new_n22184, n8803);
and_5  g19850(new_n20819, new_n11979, new_n22199);
or_5   g19851(new_n20820, new_n9141, new_n22200);
or_5   g19852(new_n20839, new_n20821, new_n22201_1);
and_5  g19853(new_n22201_1, new_n22200, new_n22202);
xor_4  g19854(new_n22202, new_n22199, new_n22203);
or_5   g19855(n16544, n4319, new_n22204);
or_5   g19856(new_n16240, new_n16221, new_n22205);
and_5  g19857(new_n22205, new_n22204, new_n22206);
xor_4  g19858(new_n22206, new_n22203, new_n22207);
or_5   g19859(new_n20840, new_n16241, new_n22208);
or_5   g19860(new_n20859, new_n20841, new_n22209);
and_5  g19861(new_n22209, new_n22208, new_n22210);
xnor_4 g19862(new_n22210, new_n22207, new_n22211);
not_10 g19863(new_n22211, new_n22212);
xnor_4 g19864(new_n22212, new_n7829, new_n22213_1);
nor_5  g19865(new_n20860, new_n7832, new_n22214);
nor_5  g19866(new_n21488, new_n21446_1, new_n22215);
nor_5  g19867(new_n22215, new_n22214, new_n22216);
xor_4  g19868(new_n22216, new_n22213_1, n8809);
not_10 g19869(new_n18241_1, new_n22218);
nor_5  g19870(new_n22181, new_n22218, new_n22219);
not_10 g19871(new_n18586, new_n22220);
or_5   g19872(new_n18592, n3324, new_n22221);
nand_5 g19873(new_n21716, new_n21704, new_n22222);
and_5  g19874(new_n22222, new_n22221, new_n22223);
and_5  g19875(new_n22223, new_n22220, new_n22224);
xor_4  g19876(new_n22224, new_n22219, new_n22225);
not_10 g19877(new_n22182, new_n22226);
xnor_4 g19878(new_n22223, new_n18586, new_n22227);
nor_5  g19879(new_n22227, new_n22226, new_n22228);
xnor_4 g19880(new_n22227, new_n22182, new_n22229);
not_10 g19881(new_n22229, new_n22230);
nor_5  g19882(new_n21724, new_n21718, new_n22231);
and_5  g19883(new_n21741, new_n21725, new_n22232);
nor_5  g19884(new_n22232, new_n22231, new_n22233);
nor_5  g19885(new_n22233, new_n22230, new_n22234);
nor_5  g19886(new_n22234, new_n22228, new_n22235);
xnor_4 g19887(new_n22235, new_n22225, n8821);
xnor_4 g19888(new_n15971, new_n15969, n8824);
xor_4  g19889(new_n18185, new_n18184, n8849);
xnor_4 g19890(new_n14136_1, new_n14127, n8861);
xnor_4 g19891(n22442, n8856, new_n22240);
not_10 g19892(new_n22240, new_n22241);
or_5   g19893(n14130, new_n8414, new_n22242);
or_5   g19894(new_n20607, new_n20584, new_n22243);
and_5  g19895(new_n22243, new_n22242, new_n22244);
xor_4  g19896(new_n22244, new_n22241, new_n22245);
xnor_4 g19897(n3324, n2272, new_n22246);
or_5   g19898(n25331, n17911, new_n22247);
or_5   g19899(new_n20576, new_n20573, new_n22248);
and_5  g19900(new_n22248, new_n22247, new_n22249);
xor_4  g19901(new_n22249, new_n22246, new_n22250);
xnor_4 g19902(new_n22250, new_n7586, new_n22251);
or_5   g19903(new_n20577, new_n7577, new_n22252);
nand_5 g19904(new_n20580, new_n20579, new_n22253_1);
nand_5 g19905(new_n22253_1, new_n20578, new_n22254);
and_5  g19906(new_n22254, new_n22252, new_n22255);
xor_4  g19907(new_n22255, new_n22251, new_n22256);
xnor_4 g19908(new_n22256, new_n22245, new_n22257);
nand_5 g19909(new_n20608, new_n20582_1, new_n22258);
nand_5 g19910(new_n20640, new_n20609_1, new_n22259);
and_5  g19911(new_n22259, new_n22258, new_n22260);
xor_4  g19912(new_n22260, new_n22257, n8862);
xor_4  g19913(new_n14017, new_n14016, n8884);
xor_4  g19914(new_n19520, new_n18675, n8909);
xor_4  g19915(new_n11948, new_n11892, n8911);
xnor_4 g19916(new_n11395, new_n11393, n8971);
xnor_4 g19917(new_n21907, new_n21880, n8982);
xnor_4 g19918(new_n5468, new_n5452, n8993);
xor_4  g19919(new_n14746_1, new_n14745, n9012);
nor_5  g19920(new_n20730, new_n20727, new_n22269);
not_10 g19921(new_n22269, new_n22270_1);
nor_5  g19922(new_n20735, new_n4447, new_n22271);
and_5  g19923(new_n22271, new_n20734, new_n22272);
xnor_4 g19924(new_n22272, new_n22270_1, new_n22273);
not_10 g19925(new_n20737, new_n22274_1);
nor_5  g19926(new_n22274_1, new_n20731, new_n22275);
nor_5  g19927(new_n20792, new_n20739, new_n22276);
nor_5  g19928(new_n22276, new_n22275, new_n22277);
xor_4  g19929(new_n22277, new_n22273, n9032);
xor_4  g19930(new_n16481_1, new_n16480, n9042);
xor_4  g19931(new_n17790, new_n17760, n9046);
xnor_4 g19932(new_n8338, new_n8278, n9047);
xnor_4 g19933(new_n15670, new_n15668, n9104);
nor_5  g19934(new_n21121, new_n21113, new_n22283_1);
nor_5  g19935(new_n22283_1, new_n15999, new_n22284);
and_5  g19936(new_n21121, new_n21113, new_n22285);
nor_5  g19937(new_n22285, new_n15816_1, new_n22286);
nor_5  g19938(new_n22286, new_n22284, new_n22287);
xor_4  g19939(new_n22287, new_n20011, new_n22288);
nor_5  g19940(new_n21123_1, new_n20011, new_n22289);
nor_5  g19941(new_n21134_1, new_n21125, new_n22290_1);
nor_5  g19942(new_n22290_1, new_n22289, new_n22291);
xor_4  g19943(new_n22291, new_n22288, n9129);
xnor_4 g19944(new_n19716, new_n19680_1, n9146);
xnor_4 g19945(new_n17996, new_n6736_1, n9164);
xor_4  g19946(new_n13123, new_n13121, n9166);
xor_4  g19947(new_n18605, new_n18578_1, new_n22296);
xor_4  g19948(new_n22296, new_n18617, n9182);
xnor_4 g19949(new_n7211, new_n7174, n9191);
xnor_4 g19950(new_n11955, new_n11883, n9217);
xor_4  g19951(new_n16649, new_n16648, n9220);
xnor_4 g19952(new_n19706, new_n19698, n9261);
xor_4  g19953(n22626, n3324, new_n22302);
or_5   g19954(new_n21705, n14440, new_n22303);
or_5   g19955(new_n19315_1, new_n19295, new_n22304);
and_5  g19956(new_n22304, new_n22303, new_n22305);
xor_4  g19957(new_n22305, new_n22302, new_n22306);
and_5  g19958(new_n22306, new_n18609, new_n22307);
not_10 g19959(new_n22307, new_n22308);
xnor_4 g19960(new_n22306, new_n18609, new_n22309_1);
nand_5 g19961(new_n19316, new_n3009, new_n22310);
nand_5 g19962(new_n19344, new_n19317, new_n22311_1);
and_5  g19963(new_n22311_1, new_n22310, new_n22312);
nor_5  g19964(new_n22312, new_n22309_1, new_n22313);
not_10 g19965(new_n22313, new_n22314);
and_5  g19966(new_n22314, new_n22308, new_n22315);
not_10 g19967(n3324, new_n22316);
or_5   g19968(n22626, new_n22316, new_n22317_1);
or_5   g19969(new_n22305, new_n22302, new_n22318);
and_5  g19970(new_n22318, new_n22317_1, new_n22319);
xnor_4 g19971(new_n22319, new_n18605, new_n22320);
xnor_4 g19972(new_n22320, new_n22315, n9287);
xor_4  g19973(new_n14570_1, new_n14559, n9308);
xnor_4 g19974(new_n5042, new_n4999, n9344);
xnor_4 g19975(new_n3710_1, new_n3691, n9364);
not_10 g19976(new_n22315, new_n22325);
nor_5  g19977(new_n22319, new_n18605, new_n22326);
and_5  g19978(new_n22326, new_n22325, new_n22327);
and_5  g19979(new_n22327, new_n18602, new_n22328);
not_10 g19980(new_n18602, new_n22329);
and_5  g19981(new_n22319, new_n18605, new_n22330);
and_5  g19982(new_n22330, new_n22315, new_n22331);
and_5  g19983(new_n22331, new_n22329, new_n22332_1);
or_5   g19984(new_n22332_1, new_n22328, n9371);
xor_4  g19985(new_n10433, new_n10432_1, n9382);
xor_4  g19986(new_n21944, new_n21936, n9403);
xnor_4 g19987(new_n13130, new_n13102, n9419);
xnor_4 g19988(new_n21682, new_n21657, n9423);
xor_4  g19989(new_n19340, new_n19325, n9430);
xor_4  g19990(n25120, n23272, new_n22339);
nand_5 g19991(new_n18901_1, n8363, new_n22340);
xor_4  g19992(n11481, n8363, new_n22341_1);
nand_5 g19993(new_n4360, n14680, new_n22342);
or_5   g19994(new_n16160, new_n16157, new_n22343);
and_5  g19995(new_n22343, new_n22342, new_n22344);
or_5   g19996(new_n22344, new_n22341_1, new_n22345);
and_5  g19997(new_n22345, new_n22340, new_n22346);
xor_4  g19998(new_n22346, new_n22339, new_n22347);
xor_4  g19999(new_n22347, new_n17667, new_n22348);
xor_4  g20000(new_n22344, new_n22341_1, new_n22349);
nand_5 g20001(new_n22349, new_n17693, new_n22350);
xnor_4 g20002(new_n22349, new_n17693, new_n22351);
or_5   g20003(new_n16168, new_n16162, new_n22352);
or_5   g20004(new_n16172, new_n16169, new_n22353_1);
and_5  g20005(new_n22353_1, new_n22352, new_n22354);
or_5   g20006(new_n22354, new_n22351, new_n22355);
and_5  g20007(new_n22355, new_n22350, new_n22356);
xnor_4 g20008(new_n22356, new_n22348, new_n22357);
not_10 g20009(new_n22357, new_n22358_1);
xor_4  g20010(new_n22358_1, new_n17739, new_n22359_1);
xor_4  g20011(new_n22354, new_n22351, new_n22360);
nor_5  g20012(new_n22360, new_n17742, new_n22361);
xor_4  g20013(new_n22360, new_n17742, new_n22362);
nor_5  g20014(new_n17748, new_n16173, new_n22363);
xnor_4 g20015(new_n17747, new_n16173, new_n22364);
nor_5  g20016(new_n17755, new_n10879, new_n22365);
xnor_4 g20017(new_n17754, new_n10879, new_n22366);
and_5  g20018(new_n17762, new_n10882, new_n22367);
xor_4  g20019(new_n17762, new_n10882, new_n22368);
nor_5  g20020(new_n17766, new_n10885, new_n22369);
nor_5  g20021(new_n17772, new_n10887, new_n22370);
nor_5  g20022(new_n15395, new_n15383, new_n22371);
or_5   g20023(new_n22371, new_n22370, new_n22372);
xor_4  g20024(new_n17766, new_n10885, new_n22373);
and_5  g20025(new_n22373, new_n22372, new_n22374);
nor_5  g20026(new_n22374, new_n22369, new_n22375);
and_5  g20027(new_n22375, new_n22368, new_n22376);
nor_5  g20028(new_n22376, new_n22367, new_n22377);
not_10 g20029(new_n22377, new_n22378);
and_5  g20030(new_n22378, new_n22366, new_n22379_1);
nor_5  g20031(new_n22379_1, new_n22365, new_n22380);
not_10 g20032(new_n22380, new_n22381);
and_5  g20033(new_n22381, new_n22364, new_n22382);
nor_5  g20034(new_n22382, new_n22363, new_n22383);
not_10 g20035(new_n22383, new_n22384);
and_5  g20036(new_n22384, new_n22362, new_n22385);
nor_5  g20037(new_n22385, new_n22361, new_n22386);
xor_4  g20038(new_n22386, new_n22359_1, n9435);
xnor_4 g20039(new_n16593, new_n16560, n9451);
xor_4  g20040(n12657, n10763, new_n22389);
or_5   g20041(n17077, new_n17115, new_n22390);
or_5   g20042(new_n19853, new_n19845, new_n22391);
and_5  g20043(new_n22391, new_n22390, new_n22392);
xor_4  g20044(new_n22392, new_n22389, new_n22393);
xnor_4 g20045(new_n22393, new_n20583, new_n22394);
nor_5  g20046(new_n19874, new_n19854, new_n22395);
not_10 g20047(new_n22395, new_n22396);
and_5  g20048(new_n19885, new_n19875, new_n22397);
not_10 g20049(new_n22397, new_n22398);
and_5  g20050(new_n22398, new_n22396, new_n22399);
xor_4  g20051(new_n22399, new_n22394, n9458);
or_5   g20052(n12507, new_n20890, new_n22401);
xor_4  g20053(n12507, n11220, new_n22402);
or_5   g20054(new_n18572_1, n15077, new_n22403);
or_5   g20055(new_n15306, new_n15284, new_n22404);
and_5  g20056(new_n22404, new_n22403, new_n22405);
or_5   g20057(new_n22405, new_n22402, new_n22406);
and_5  g20058(new_n22406, new_n22401, new_n22407);
xor_4  g20059(new_n22407, new_n21331, new_n22408);
xor_4  g20060(new_n22405, new_n22402, new_n22409);
nor_5  g20061(new_n22409, new_n21333, new_n22410);
xor_4  g20062(new_n22409, new_n21333, new_n22411);
not_10 g20063(new_n22411, new_n22412);
nor_5  g20064(new_n15307_1, new_n15283, new_n22413);
nor_5  g20065(new_n15353_1, new_n15309, new_n22414);
nor_5  g20066(new_n22414, new_n22413, new_n22415);
nor_5  g20067(new_n22415, new_n22412, new_n22416);
nor_5  g20068(new_n22416, new_n22410, new_n22417);
xor_4  g20069(new_n22417, new_n22408, n9459);
xnor_4 g20070(new_n15611, new_n15609, n9508);
xor_4  g20071(new_n13134, new_n13090, n9552);
xnor_4 g20072(new_n4583, new_n4581, n9556);
xnor_4 g20073(new_n11367, new_n8998, n9558);
xor_4  g20074(new_n21549_1, new_n14738, n9616);
xnor_4 g20075(new_n8724, new_n8693, n9622);
xor_4  g20076(new_n17105, new_n17088, n9626);
xnor_4 g20077(new_n4589, new_n4571, n9633);
or_5   g20078(new_n7779, n23272, new_n22427);
or_5   g20079(new_n22346, new_n22339, new_n22428);
and_5  g20080(new_n22428, new_n22427, new_n22429);
and_5  g20081(new_n22429, new_n21919, new_n22430);
xor_4  g20082(new_n22429, new_n21919, new_n22431);
nand_5 g20083(new_n22347, new_n17667, new_n22432);
not_10 g20084(new_n22348, new_n22433_1);
or_5   g20085(new_n22356, new_n22433_1, new_n22434);
and_5  g20086(new_n22434, new_n22432, new_n22435);
and_5  g20087(new_n22435, new_n22431, new_n22436);
nor_5  g20088(new_n22436, new_n22430, new_n22437);
nand_5 g20089(new_n22437, new_n5736, new_n22438);
xor_4  g20090(new_n22437, new_n5590, new_n22439);
xor_4  g20091(new_n22435, new_n22431, new_n22440);
or_5   g20092(new_n22440, new_n5736, new_n22441);
xnor_4 g20093(new_n22440, new_n5590, new_n22442_1);
nor_5  g20094(new_n22357, new_n5591, new_n22443);
and_5  g20095(new_n22360, new_n5661, new_n22444_1);
xnor_4 g20096(new_n22360, new_n5661, new_n22445);
nand_5 g20097(new_n16173, new_n5667, new_n22446);
or_5   g20098(new_n16177, new_n16174, new_n22447);
and_5  g20099(new_n22447, new_n22446, new_n22448);
nor_5  g20100(new_n22448, new_n22445, new_n22449);
nor_5  g20101(new_n22449, new_n22444_1, new_n22450);
xnor_4 g20102(new_n22358_1, new_n5591, new_n22451);
and_5  g20103(new_n22451, new_n22450, new_n22452);
nor_5  g20104(new_n22452, new_n22443, new_n22453);
nand_5 g20105(new_n22453, new_n22442_1, new_n22454);
and_5  g20106(new_n22454, new_n22441, new_n22455);
or_5   g20107(new_n22455, new_n22439, new_n22456);
and_5  g20108(new_n22456, new_n22438, n9635);
xnor_4 g20109(new_n20095, new_n20090, n9648);
xor_4  g20110(new_n5024_1, new_n5023, n9689);
xnor_4 g20111(new_n11060, new_n11037, n9695);
xor_4  g20112(new_n7718, new_n7660, n9699);
xnor_4 g20113(new_n17195, new_n15118_1, new_n22462);
nor_5  g20114(new_n16612, new_n15118_1, new_n22463);
and_5  g20115(new_n16656_1, new_n16613, new_n22464);
nor_5  g20116(new_n22464, new_n22463, new_n22465);
xor_4  g20117(new_n22465, new_n22462, n9726);
xor_4  g20118(new_n13665, new_n10233, n9753);
xnor_4 g20119(new_n3380, new_n3360, n9761);
xnor_4 g20120(new_n10250_1, new_n10195, n9763);
xnor_4 g20121(new_n14014, new_n14012, n9767);
xor_4  g20122(new_n14188, new_n13915, n9771);
xor_4  g20123(new_n22030, new_n22027_1, n9778);
xnor_4 g20124(new_n16383, new_n16374, n9783);
xnor_4 g20125(new_n6765, new_n6763, n9803);
not_10 g20126(n4319, new_n22475);
and_5  g20127(new_n21493, new_n11982, new_n22476);
and_5  g20128(new_n22476, new_n22475, new_n22477);
xor_4  g20129(new_n22476, new_n22475, new_n22478);
and_5  g20130(new_n22478, new_n18547, new_n22479);
nor_5  g20131(new_n22478, new_n18547, new_n22480);
and_5  g20132(new_n21494, new_n18552, new_n22481);
not_10 g20133(new_n22481, new_n22482);
nor_5  g20134(new_n21494, new_n18552, new_n22483);
and_5  g20135(new_n21496, new_n17255, new_n22484_1);
nor_5  g20136(new_n21496, new_n17255, new_n22485);
nor_5  g20137(new_n21499, new_n17259, new_n22486);
nand_5 g20138(new_n21502, new_n17264, new_n22487);
xnor_4 g20139(new_n21502, new_n17264, new_n22488);
nand_5 g20140(new_n6728, new_n6713, new_n22489_1);
or_5   g20141(new_n6752, new_n6729_1, new_n22490);
and_5  g20142(new_n22490, new_n22489_1, new_n22491);
or_5   g20143(new_n22491, new_n22488, new_n22492_1);
and_5  g20144(new_n22492_1, new_n22487, new_n22493);
xor_4  g20145(new_n21499, new_n17259, new_n22494_1);
and_5  g20146(new_n22494_1, new_n22493, new_n22495);
or_5   g20147(new_n22495, new_n22486, new_n22496);
or_5   g20148(new_n22496, new_n22485, new_n22497);
not_10 g20149(new_n22497, new_n22498);
nor_5  g20150(new_n22498, new_n22484_1, new_n22499);
or_5   g20151(new_n22499, new_n22483, new_n22500);
and_5  g20152(new_n22500, new_n22482, new_n22501);
or_5   g20153(new_n22501, new_n22480, new_n22502);
not_10 g20154(new_n22502, new_n22503);
nor_5  g20155(new_n22503, new_n22479, new_n22504);
xor_4  g20156(new_n22504, new_n18545, new_n22505);
xor_4  g20157(new_n22505, new_n22477, new_n22506);
not_10 g20158(new_n22506, new_n22507);
or_5   g20159(new_n22507, new_n3315, new_n22508);
xor_4  g20160(new_n22507, new_n3315, new_n22509);
xor_4  g20161(new_n22478, new_n18548, new_n22510);
xor_4  g20162(new_n22510, new_n22501, new_n22511);
or_5   g20163(new_n22511, new_n3324_1, new_n22512);
xnor_4 g20164(new_n22511, new_n3322, new_n22513);
not_10 g20165(new_n22513, new_n22514);
xor_4  g20166(new_n21494, new_n18553, new_n22515);
xor_4  g20167(new_n22515, new_n22499, new_n22516);
or_5   g20168(new_n22516, new_n3330, new_n22517);
xnor_4 g20169(new_n22516, new_n3328, new_n22518);
not_10 g20170(new_n22518, new_n22519);
xnor_4 g20171(new_n21496, new_n17255, new_n22520);
xor_4  g20172(new_n22520, new_n22496, new_n22521);
or_5   g20173(new_n22521, new_n3336, new_n22522);
xnor_4 g20174(new_n22521, new_n3334, new_n22523);
not_10 g20175(new_n22523, new_n22524);
xor_4  g20176(new_n22494_1, new_n22493, new_n22525);
nand_5 g20177(new_n22525, new_n3340_1, new_n22526);
xor_4  g20178(new_n22525, new_n3340_1, new_n22527);
not_10 g20179(new_n22527, new_n22528);
xor_4  g20180(new_n22491, new_n22488, new_n22529);
or_5   g20181(new_n22529, new_n3347, new_n22530);
xnor_4 g20182(new_n22529, new_n3345, new_n22531);
not_10 g20183(new_n22531, new_n22532);
or_5   g20184(new_n6753, new_n3353, new_n22533_1);
not_10 g20185(new_n6754, new_n22534);
or_5   g20186(new_n6773_1, new_n22534, new_n22535);
and_5  g20187(new_n22535, new_n22533_1, new_n22536);
or_5   g20188(new_n22536, new_n22532, new_n22537);
and_5  g20189(new_n22537, new_n22530, new_n22538);
or_5   g20190(new_n22538, new_n22528, new_n22539);
and_5  g20191(new_n22539, new_n22526, new_n22540);
or_5   g20192(new_n22540, new_n22524, new_n22541);
and_5  g20193(new_n22541, new_n22522, new_n22542);
or_5   g20194(new_n22542, new_n22519, new_n22543);
and_5  g20195(new_n22543, new_n22517, new_n22544);
or_5   g20196(new_n22544, new_n22514, new_n22545);
nand_5 g20197(new_n22545, new_n22512, new_n22546);
nand_5 g20198(new_n22546, new_n22509, new_n22547);
and_5  g20199(new_n22547, new_n22508, new_n22548);
and_5  g20200(new_n22504, new_n18545, new_n22549);
xor_4  g20201(new_n22477, new_n18502, new_n22550);
nand_5 g20202(new_n22550, new_n22549, new_n22551);
or_5   g20203(new_n22550, new_n22504, new_n22552);
and_5  g20204(new_n22552, new_n22551, new_n22553);
and_5  g20205(new_n22553, new_n22548, new_n22554_1);
nor_5  g20206(new_n22477, new_n18502, new_n22555);
and_5  g20207(new_n22555, new_n22504, new_n22556);
xor_4  g20208(new_n22556, new_n22554_1, n9833);
and_5  g20209(new_n17934, new_n8802, new_n22558);
and_5  g20210(new_n22558, new_n8798, new_n22559);
and_5  g20211(new_n22559, new_n18520, new_n22560);
nor_5  g20212(new_n22560, new_n18540, new_n22561);
xor_4  g20213(new_n22559, new_n18520, new_n22562);
nand_5 g20214(new_n22562, new_n18518, new_n22563);
xor_4  g20215(new_n22562, new_n18518, new_n22564);
not_10 g20216(new_n22564, new_n22565);
xor_4  g20217(new_n22558, new_n8798, new_n22566);
nand_5 g20218(new_n22566, new_n18523, new_n22567);
xnor_4 g20219(new_n22566, new_n18523, new_n22568);
nand_5 g20220(new_n17935, new_n17224, new_n22569);
nand_5 g20221(new_n17964, new_n17936, new_n22570);
and_5  g20222(new_n22570, new_n22569, new_n22571);
or_5   g20223(new_n22571, new_n22568, new_n22572);
and_5  g20224(new_n22572, new_n22567, new_n22573);
or_5   g20225(new_n22573, new_n22565, new_n22574);
and_5  g20226(new_n22574, new_n22563, new_n22575);
nand_5 g20227(new_n22575, new_n22561, new_n22576);
and_5  g20228(new_n17966, new_n8961, new_n22577);
and_5  g20229(new_n22577, new_n8954, new_n22578);
and_5  g20230(new_n22578, new_n8893, new_n22579);
xor_4  g20231(new_n22579, new_n16603, new_n22580);
xor_4  g20232(new_n22578, new_n8893, new_n22581);
nor_5  g20233(new_n22581, new_n13310, new_n22582);
not_10 g20234(new_n22582, new_n22583);
xor_4  g20235(new_n22577, new_n8954, new_n22584_1);
nor_5  g20236(new_n22584_1, new_n5337_1, new_n22585);
xor_4  g20237(new_n22584_1, new_n5337_1, new_n22586);
nand_5 g20238(new_n17967, new_n5377, new_n22587);
nand_5 g20239(new_n17972, new_n17968_1, new_n22588_1);
and_5  g20240(new_n22588_1, new_n22587, new_n22589_1);
and_5  g20241(new_n22589_1, new_n22586, new_n22590);
or_5   g20242(new_n22590, new_n22585, new_n22591_1);
xor_4  g20243(new_n22581, new_n13310, new_n22592);
and_5  g20244(new_n22592, new_n22591_1, new_n22593);
not_10 g20245(new_n22593, new_n22594);
and_5  g20246(new_n22594, new_n22583, new_n22595);
xnor_4 g20247(new_n22595, new_n22580, new_n22596);
xor_4  g20248(new_n22560, new_n18540, new_n22597_1);
xor_4  g20249(new_n22597_1, new_n22575, new_n22598);
nor_5  g20250(new_n22598, new_n22596, new_n22599);
xor_4  g20251(new_n22598, new_n22596, new_n22600);
not_10 g20252(new_n22600, new_n22601);
xor_4  g20253(new_n22573, new_n22565, new_n22602);
not_10 g20254(new_n22602, new_n22603);
xor_4  g20255(new_n22592, new_n22591_1, new_n22604);
and_5  g20256(new_n22604, new_n22603, new_n22605);
xor_4  g20257(new_n22604, new_n22603, new_n22606);
xor_4  g20258(new_n22589_1, new_n22586, new_n22607);
not_10 g20259(new_n22607, new_n22608);
xor_4  g20260(new_n22571, new_n22568, new_n22609);
nor_5  g20261(new_n22609, new_n22608, new_n22610);
xor_4  g20262(new_n22609, new_n22608, new_n22611);
not_10 g20263(new_n22611, new_n22612);
nor_5  g20264(new_n17973, new_n17965, new_n22613);
nor_5  g20265(new_n18014, new_n17975, new_n22614);
nor_5  g20266(new_n22614, new_n22613, new_n22615);
nor_5  g20267(new_n22615, new_n22612, new_n22616);
nor_5  g20268(new_n22616, new_n22610, new_n22617);
not_10 g20269(new_n22617, new_n22618);
and_5  g20270(new_n22618, new_n22606, new_n22619_1);
nor_5  g20271(new_n22619_1, new_n22605, new_n22620_1);
nor_5  g20272(new_n22620_1, new_n22601, new_n22621);
nor_5  g20273(new_n22621, new_n22599, new_n22622);
nor_5  g20274(new_n22622, new_n22576, new_n22623_1);
xnor_4 g20275(new_n22622, new_n22576, new_n22624);
nor_5  g20276(new_n22579, new_n16603, new_n22625);
not_10 g20277(new_n22595, new_n22626_1);
and_5  g20278(new_n22626_1, new_n22625, new_n22627);
and_5  g20279(new_n22627, new_n22624, new_n22628);
or_5   g20280(new_n22628, new_n22623_1, n9838);
xnor_4 g20281(new_n20250_1, new_n20246, n9867);
nor_5  g20282(new_n19808, new_n5653, new_n22631_1);
and_5  g20283(new_n19812, new_n19809, new_n22632);
nor_5  g20284(new_n22632, new_n22631_1, new_n22633);
nor_5  g20285(new_n22633, new_n21072, new_n22634);
xor_4  g20286(new_n22633, new_n21072, new_n22635);
or_5   g20287(new_n22635, new_n8269, new_n22636);
or_5   g20288(new_n19813, new_n8277, new_n22637);
or_5   g20289(new_n19818, new_n19815, new_n22638);
and_5  g20290(new_n22638, new_n22637, new_n22639);
xor_4  g20291(new_n22635, new_n8269, new_n22640);
not_10 g20292(new_n22640, new_n22641);
or_5   g20293(new_n22641, new_n22639, new_n22642);
and_5  g20294(new_n22642, new_n22636, new_n22643);
or_5   g20295(new_n22643, new_n22634, new_n22644);
and_5  g20296(new_n22644, new_n8163, n9890);
xor_4  g20297(new_n18562, new_n18551, n9917);
xnor_4 g20298(new_n21363, new_n21354, n9919);
xnor_4 g20299(new_n18738, new_n18723, n9938);
xnor_4 g20300(new_n18364, new_n18363, n9946);
xnor_4 g20301(n21784, n3740, new_n22650);
or_5   g20302(n5521, n2858, new_n22651);
xnor_4 g20303(n5521, n2858, new_n22652);
or_5   g20304(n11926, n2659, new_n22653);
xnor_4 g20305(n11926, n2659, new_n22654);
or_5   g20306(n24327, n4325, new_n22655);
xor_4  g20307(n24327, n4325, new_n22656);
nand_5 g20308(n22198, n5337, new_n22657);
or_5   g20309(n22198, n5337, new_n22658);
nor_5  g20310(n20826, n626, new_n22659);
nor_5  g20311(new_n13284, new_n13281, new_n22660_1);
nor_5  g20312(new_n22660_1, new_n22659, new_n22661);
nand_5 g20313(new_n22661, new_n22658, new_n22662);
and_5  g20314(new_n22662, new_n22657, new_n22663);
nand_5 g20315(new_n22663, new_n22656, new_n22664);
and_5  g20316(new_n22664, new_n22655, new_n22665);
or_5   g20317(new_n22665, new_n22654, new_n22666);
and_5  g20318(new_n22666, new_n22653, new_n22667);
or_5   g20319(new_n22667, new_n22652, new_n22668);
and_5  g20320(new_n22668, new_n22651, new_n22669);
xor_4  g20321(new_n22669, new_n22650, new_n22670);
xor_4  g20322(new_n22670, new_n4857, new_n22671);
xor_4  g20323(new_n22667, new_n22652, new_n22672);
nand_5 g20324(new_n22672, new_n4862, new_n22673);
xnor_4 g20325(new_n22672, new_n4862, new_n22674);
xor_4  g20326(new_n22665, new_n22654, new_n22675);
nand_5 g20327(new_n22675, new_n4866, new_n22676);
xor_4  g20328(new_n22663, new_n22656, new_n22677);
and_5  g20329(new_n22677, new_n4870, new_n22678);
xnor_4 g20330(new_n22677, new_n4870, new_n22679);
xor_4  g20331(n22198, n5337, new_n22680);
xor_4  g20332(new_n22680, new_n22661, new_n22681);
or_5   g20333(new_n22681, new_n4873, new_n22682);
or_5   g20334(new_n13285_1, new_n13280, new_n22683);
nand_5 g20335(new_n13286, new_n4876, new_n22684);
and_5  g20336(new_n22684, new_n22683, new_n22685);
xor_4  g20337(new_n22681, new_n4873, new_n22686);
nand_5 g20338(new_n22686, new_n22685, new_n22687);
and_5  g20339(new_n22687, new_n22682, new_n22688);
nor_5  g20340(new_n22688, new_n22679, new_n22689);
or_5   g20341(new_n22689, new_n22678, new_n22690);
xor_4  g20342(new_n22675, new_n4866, new_n22691);
nand_5 g20343(new_n22691, new_n22690, new_n22692);
and_5  g20344(new_n22692, new_n22676, new_n22693);
or_5   g20345(new_n22693, new_n22674, new_n22694);
and_5  g20346(new_n22694, new_n22673, new_n22695);
xor_4  g20347(new_n22695, new_n22671, new_n22696);
xnor_4 g20348(new_n22696, new_n17856, new_n22697_1);
xor_4  g20349(new_n22693, new_n22674, new_n22698);
nand_5 g20350(new_n22698, new_n17160, new_n22699);
xor_4  g20351(new_n22698, new_n17160, new_n22700);
not_10 g20352(new_n22700, new_n22701);
xor_4  g20353(new_n22691, new_n22690, new_n22702);
nand_5 g20354(new_n22702, new_n17162, new_n22703);
xor_4  g20355(new_n22702, new_n17162, new_n22704);
not_10 g20356(new_n22704, new_n22705);
xor_4  g20357(new_n22688, new_n22679, new_n22706);
nand_5 g20358(new_n22706, new_n3767, new_n22707);
xor_4  g20359(new_n22706, new_n3767, new_n22708);
xor_4  g20360(new_n22686, new_n22685, new_n22709);
or_5   g20361(new_n22709, new_n3770, new_n22710);
and_5  g20362(new_n13287, new_n3774, new_n22711);
nor_5  g20363(new_n13296, new_n13288, new_n22712);
or_5   g20364(new_n22712, new_n22711, new_n22713);
xor_4  g20365(new_n22709, new_n3770, new_n22714_1);
nand_5 g20366(new_n22714_1, new_n22713, new_n22715);
and_5  g20367(new_n22715, new_n22710, new_n22716);
nand_5 g20368(new_n22716, new_n22708, new_n22717);
and_5  g20369(new_n22717, new_n22707, new_n22718);
or_5   g20370(new_n22718, new_n22705, new_n22719);
and_5  g20371(new_n22719, new_n22703, new_n22720);
or_5   g20372(new_n22720, new_n22701, new_n22721);
and_5  g20373(new_n22721, new_n22699, new_n22722);
xor_4  g20374(new_n22722, new_n22697_1, n9968);
or_5   g20375(new_n21018, new_n14243, new_n22724);
xor_4  g20376(new_n21018, new_n14243, new_n22725);
nor_5  g20377(new_n21025, new_n14243, new_n22726);
xor_4  g20378(new_n21025, new_n14243, new_n22727);
and_5  g20379(new_n11545, new_n11481_1, new_n22728);
and_5  g20380(new_n11592, new_n11546, new_n22729);
nor_5  g20381(new_n22729, new_n22728, new_n22730);
and_5  g20382(new_n22730, new_n22727, new_n22731);
nor_5  g20383(new_n22731, new_n22726, new_n22732);
nand_5 g20384(new_n22732, new_n22725, new_n22733);
and_5  g20385(new_n22733, new_n22724, n10009);
xnor_4 g20386(new_n21774, new_n21769, n10010);
not_10 g20387(new_n15186, new_n22736);
and_5  g20388(new_n15118_1, new_n11259, new_n22737);
and_5  g20389(new_n15148, new_n15119, new_n22738);
nor_5  g20390(new_n22738, new_n22737, new_n22739);
nand_5 g20391(new_n22739, new_n22736, new_n22740);
xor_4  g20392(new_n22739, new_n15186, new_n22741);
or_5   g20393(new_n22736, new_n15149, new_n22742);
nand_5 g20394(new_n15233, new_n15187, new_n22743);
and_5  g20395(new_n22743, new_n22742, new_n22744);
or_5   g20396(new_n22744, new_n22741, new_n22745);
and_5  g20397(new_n22745, new_n22740, n10019);
xor_4  g20398(new_n15014, new_n14953, n10021);
xor_4  g20399(new_n9804, new_n9796, n10055);
xnor_4 g20400(new_n10902, new_n10884, n10101);
xnor_4 g20401(new_n4598, new_n4551, n10111);
nor_5  g20402(n16544, new_n22316, new_n22751);
not_10 g20403(new_n22751, new_n22752);
xor_4  g20404(n16544, n3324, new_n22753);
or_5   g20405(new_n21705, n6814, new_n22754);
xor_4  g20406(n17911, n6814, new_n22755);
or_5   g20407(new_n19296, n19701, new_n22756);
xor_4  g20408(n21997, n19701, new_n22757);
or_5   g20409(new_n8652, n23529, new_n22758);
xor_4  g20410(n25119, n23529, new_n22759);
or_5   g20411(n24620, new_n8654, new_n22760);
xor_4  g20412(n24620, n1163, new_n22761_1);
or_5   g20413(new_n8656_1, n5211, new_n22762);
or_5   g20414(n18537, new_n9162, new_n22763);
and_5  g20415(n12956, new_n8660, new_n22764_1);
nor_5  g20416(new_n9695_1, new_n9684, new_n22765);
nor_5  g20417(new_n22765, new_n22764_1, new_n22766);
nand_5 g20418(new_n22766, new_n22763, new_n22767);
and_5  g20419(new_n22767, new_n22762, new_n22768);
or_5   g20420(new_n22768, new_n22761_1, new_n22769);
and_5  g20421(new_n22769, new_n22760, new_n22770);
or_5   g20422(new_n22770, new_n22759, new_n22771);
and_5  g20423(new_n22771, new_n22758, new_n22772);
or_5   g20424(new_n22772, new_n22757, new_n22773);
and_5  g20425(new_n22773, new_n22756, new_n22774);
or_5   g20426(new_n22774, new_n22755, new_n22775);
and_5  g20427(new_n22775, new_n22754, new_n22776);
nor_5  g20428(new_n22776, new_n22753, new_n22777);
not_10 g20429(new_n22777, new_n22778);
and_5  g20430(new_n22778, new_n22752, new_n22779_1);
xor_4  g20431(new_n22779_1, new_n21926, new_n22780);
not_10 g20432(new_n22779_1, new_n22781);
or_5   g20433(new_n22781, new_n21937, new_n22782);
and_5  g20434(new_n22781, new_n21937, new_n22783);
not_10 g20435(new_n22783, new_n22784);
xor_4  g20436(new_n22776, new_n22753, new_n22785);
nor_5  g20437(new_n22785, new_n17698, new_n22786);
xor_4  g20438(new_n22785, new_n17698, new_n22787_1);
xor_4  g20439(new_n22774, new_n22755, new_n22788);
nor_5  g20440(new_n22788, new_n17743, new_n22789);
xor_4  g20441(new_n22788, new_n17743, new_n22790);
xor_4  g20442(new_n22772, new_n22757, new_n22791);
nor_5  g20443(new_n22791, new_n17750, new_n22792);
xor_4  g20444(new_n22791, new_n17750, new_n22793_1);
xor_4  g20445(new_n22770, new_n22759, new_n22794);
nor_5  g20446(new_n22794, new_n17757, new_n22795);
xor_4  g20447(new_n22794, new_n17757, new_n22796);
xor_4  g20448(new_n22768, new_n22761_1, new_n22797);
nor_5  g20449(new_n22797, new_n17764, new_n22798);
xnor_4 g20450(n18537, n5211, new_n22799);
xor_4  g20451(new_n22799, new_n22766, new_n22800);
and_5  g20452(new_n22800, new_n17768, new_n22801);
xnor_4 g20453(new_n22800, new_n17768, new_n22802);
or_5   g20454(new_n9696, new_n9683, new_n22803);
nand_5 g20455(new_n9717, new_n9697, new_n22804);
and_5  g20456(new_n22804, new_n22803, new_n22805);
nor_5  g20457(new_n22805, new_n22802, new_n22806);
nor_5  g20458(new_n22806, new_n22801, new_n22807);
xor_4  g20459(new_n22797, new_n17764, new_n22808);
and_5  g20460(new_n22808, new_n22807, new_n22809);
nor_5  g20461(new_n22809, new_n22798, new_n22810);
not_10 g20462(new_n22810, new_n22811);
and_5  g20463(new_n22811, new_n22796, new_n22812);
nor_5  g20464(new_n22812, new_n22795, new_n22813);
not_10 g20465(new_n22813, new_n22814);
and_5  g20466(new_n22814, new_n22793_1, new_n22815);
nor_5  g20467(new_n22815, new_n22792, new_n22816);
not_10 g20468(new_n22816, new_n22817);
and_5  g20469(new_n22817, new_n22790, new_n22818);
nor_5  g20470(new_n22818, new_n22789, new_n22819_1);
not_10 g20471(new_n22819_1, new_n22820);
and_5  g20472(new_n22820, new_n22787_1, new_n22821);
nor_5  g20473(new_n22821, new_n22786, new_n22822);
nand_5 g20474(new_n22822, new_n22784, new_n22823);
and_5  g20475(new_n22823, new_n22782, new_n22824);
xor_4  g20476(new_n22824, new_n22780, n10165);
xnor_4 g20477(new_n13372, new_n13371, n10236);
xnor_4 g20478(new_n14878, new_n14856, n10239);
xor_4  g20479(new_n6445, new_n6398, n10244);
xnor_4 g20480(new_n18667, new_n18653_1, n10261);
xor_4  g20481(new_n16217_1, new_n16203, n10262);
xor_4  g20482(new_n17416, new_n17415, n10287);
not_10 g20483(new_n15732, new_n22832);
nor_5  g20484(new_n22177, new_n22832, new_n22833);
xor_4  g20485(new_n22219, new_n22833, new_n22834);
and_5  g20486(new_n22226, new_n22178, new_n22835);
nor_5  g20487(new_n22197, new_n22184, new_n22836);
nor_5  g20488(new_n22836, new_n22835, new_n22837);
xnor_4 g20489(new_n22837, new_n22834, n10295);
xor_4  g20490(new_n15338, new_n15332_1, n10321);
xnor_4 g20491(new_n14880, new_n14853, n10326);
xor_4  g20492(new_n2819, new_n2809_1, n10327);
xnor_4 g20493(new_n21025, new_n21005, new_n22842);
xor_4  g20494(new_n22842, new_n21022, n10330);
xor_4  g20495(new_n21686, new_n21650, n10340);
xnor_4 g20496(new_n17413, new_n17411, new_n22845);
xor_4  g20497(new_n22845, new_n17417, n10345);
not_10 g20498(new_n4913_1, new_n22847);
and_5  g20499(new_n4916, new_n22847, new_n22848);
not_10 g20500(new_n22848, new_n22849);
nand_5 g20501(new_n19755, new_n22849, new_n22850);
nor_5  g20502(new_n19760, new_n4918, new_n22851);
xor_4  g20503(new_n19760, new_n4918, new_n22852);
not_10 g20504(new_n22852, new_n22853);
and_5  g20505(new_n19766, new_n4920, new_n22854);
xor_4  g20506(new_n19766, new_n4920, new_n22855);
not_10 g20507(new_n22855, new_n22856);
and_5  g20508(new_n19772, new_n4924, new_n22857);
xor_4  g20509(new_n19772, new_n4924, new_n22858_1);
not_10 g20510(new_n22858_1, new_n22859);
and_5  g20511(new_n19778, new_n4928, new_n22860);
xor_4  g20512(new_n19778, new_n4928, new_n22861);
not_10 g20513(new_n22861, new_n22862);
and_5  g20514(new_n20524, new_n4932, new_n22863);
xnor_4 g20515(new_n9589, new_n4932, new_n22864);
not_10 g20516(new_n22864, new_n22865);
and_5  g20517(new_n20528, new_n4936, new_n22866);
xnor_4 g20518(new_n9593, new_n4936, new_n22867);
not_10 g20519(new_n22867, new_n22868);
and_5  g20520(new_n20532, new_n4940, new_n22869);
xnor_4 g20521(new_n9598_1, new_n4940, new_n22870_1);
not_10 g20522(new_n22870_1, new_n22871_1);
and_5  g20523(new_n20536, new_n4944, new_n22872);
xnor_4 g20524(new_n9603, new_n4944, new_n22873);
not_10 g20525(new_n22873, new_n22874);
and_5  g20526(new_n9610, new_n4947_1, new_n22875);
xor_4  g20527(new_n9610, new_n4947_1, new_n22876);
and_5  g20528(new_n9616_1, new_n4953, new_n22877);
and_5  g20529(new_n22877, new_n9612, new_n22878);
not_10 g20530(new_n4950, new_n22879_1);
xnor_4 g20531(new_n22877, new_n9619, new_n22880);
and_5  g20532(new_n22880, new_n22879_1, new_n22881);
nor_5  g20533(new_n22881, new_n22878, new_n22882);
not_10 g20534(new_n22882, new_n22883);
and_5  g20535(new_n22883, new_n22876, new_n22884);
nor_5  g20536(new_n22884, new_n22875, new_n22885);
nor_5  g20537(new_n22885, new_n22874, new_n22886);
nor_5  g20538(new_n22886, new_n22872, new_n22887);
nor_5  g20539(new_n22887, new_n22871_1, new_n22888);
nor_5  g20540(new_n22888, new_n22869, new_n22889);
nor_5  g20541(new_n22889, new_n22868, new_n22890);
nor_5  g20542(new_n22890, new_n22866, new_n22891_1);
nor_5  g20543(new_n22891_1, new_n22865, new_n22892);
nor_5  g20544(new_n22892, new_n22863, new_n22893);
nor_5  g20545(new_n22893, new_n22862, new_n22894);
nor_5  g20546(new_n22894, new_n22860, new_n22895);
nor_5  g20547(new_n22895, new_n22859, new_n22896);
nor_5  g20548(new_n22896, new_n22857, new_n22897_1);
nor_5  g20549(new_n22897_1, new_n22856, new_n22898);
nor_5  g20550(new_n22898, new_n22854, new_n22899);
nor_5  g20551(new_n22899, new_n22853, new_n22900);
nor_5  g20552(new_n22900, new_n22851, new_n22901);
xnor_4 g20553(new_n19756_1, new_n22849, new_n22902);
nand_5 g20554(new_n22902, new_n22901, new_n22903_1);
and_5  g20555(new_n22903_1, new_n22850, n10356);
xor_4  g20556(new_n20336, new_n20335, n10385);
and_5  g20557(new_n20569, new_n19756_1, new_n22906);
or_5   g20558(new_n20569, new_n19756_1, new_n22907_1);
and_5  g20559(new_n22907_1, new_n20509, new_n22908);
nor_5  g20560(new_n22908, new_n22906, new_n22909);
nor_5  g20561(new_n22909, new_n20507, n10387);
xnor_4 g20562(new_n20780, new_n20763, n10388);
xor_4  g20563(new_n15985, new_n15934, n10390);
xor_4  g20564(new_n9706, new_n9705, n10404);
xnor_4 g20565(new_n16381, new_n16378, n10409);
xor_4  g20566(new_n16579, new_n8711, n10420);
xor_4  g20567(new_n18658, new_n6967_1, n10432);
xor_4  g20568(new_n21765_1, new_n21141, new_n22917);
not_10 g20569(new_n22917, new_n22918_1);
nand_5 g20570(new_n21145, new_n9852, new_n22919);
or_5   g20571(new_n21432, new_n21425, new_n22920);
and_5  g20572(new_n22920, new_n22919, new_n22921);
xor_4  g20573(new_n22921, new_n22918_1, new_n22922);
xor_4  g20574(new_n22922, new_n11716, new_n22923);
nand_5 g20575(new_n21433, new_n11722, new_n22924);
or_5   g20576(new_n21443, new_n21434, new_n22925);
and_5  g20577(new_n22925, new_n22924, new_n22926);
xor_4  g20578(new_n22926, new_n22923, n10484);
xnor_4 g20579(new_n11580_1, new_n11564_1, n10489);
xnor_4 g20580(new_n13811, new_n3638, n10525);
xor_4  g20581(new_n17990, new_n12404, new_n22930);
xor_4  g20582(new_n22930, new_n18001, n10540);
xor_4  g20583(new_n16489, new_n16463, n10561);
xor_4  g20584(new_n15991, new_n15922_1, n10564);
xor_4  g20585(new_n10233, new_n10231, n10588);
xnor_4 g20586(new_n10235, new_n10234, n10595);
xor_4  g20587(new_n21554, new_n21542, n10617);
xnor_4 g20588(new_n12769, new_n12700, n10628);
xnor_4 g20589(new_n10854, new_n5779, new_n22938);
not_10 g20590(new_n22938, new_n22939_1);
and_5  g20591(new_n10861, new_n5783, new_n22940);
xnor_4 g20592(new_n10861, new_n5784, new_n22941);
and_5  g20593(new_n10864, new_n5789, new_n22942);
not_10 g20594(new_n22942, new_n22943);
xor_4  g20595(new_n10864, new_n5789, new_n22944);
nor_5  g20596(new_n5829, new_n5795, new_n22945);
nor_5  g20597(new_n22945, new_n5839, new_n22946);
xnor_4 g20598(new_n22945, new_n5838, new_n22947);
and_5  g20599(new_n22947, new_n5803, new_n22948);
nor_5  g20600(new_n22948, new_n22946, new_n22949);
not_10 g20601(new_n22949, new_n22950);
and_5  g20602(new_n22950, new_n22944, new_n22951);
not_10 g20603(new_n22951, new_n22952);
and_5  g20604(new_n22952, new_n22943, new_n22953);
not_10 g20605(new_n22953, new_n22954);
and_5  g20606(new_n22954, new_n22941, new_n22955);
nor_5  g20607(new_n22955, new_n22940, new_n22956);
xnor_4 g20608(new_n22956, new_n22939_1, n10647);
and_5  g20609(new_n8478, new_n8472, new_n22958);
not_10 g20610(new_n22958, new_n22959);
nand_5 g20611(new_n3600, new_n3583, new_n22960);
nor_5  g20612(new_n3659, new_n3601, new_n22961);
nor_5  g20613(new_n22961, new_n20233, new_n22962);
and_5  g20614(new_n22962, new_n22960, new_n22963);
and_5  g20615(new_n22963, new_n13778, new_n22964);
xor_4  g20616(new_n22964, new_n22959, new_n22965);
not_10 g20617(new_n8479, new_n22966);
xnor_4 g20618(new_n22963, new_n13777, new_n22967);
nor_5  g20619(new_n22967, new_n22966, new_n22968);
or_5   g20620(new_n3660, new_n3530, new_n22969);
nand_5 g20621(new_n3722, new_n3661, new_n22970);
and_5  g20622(new_n22970, new_n22969, new_n22971);
xnor_4 g20623(new_n22967, new_n8479, new_n22972);
and_5  g20624(new_n22972, new_n22971, new_n22973);
nor_5  g20625(new_n22973, new_n22968, new_n22974);
xor_4  g20626(new_n22974, new_n22965, n10653);
xor_4  g20627(new_n9249, new_n9247, n10692);
xor_4  g20628(new_n15067, new_n15066, n10694);
xnor_4 g20629(new_n20638, new_n20612, n10701);
xnor_4 g20630(new_n6175, new_n6157, n10756);
not_10 g20631(n5101, new_n22980);
and_5  g20632(n6659, new_n22980, new_n22981);
not_10 g20633(new_n22981, new_n22982);
nor_5  g20634(new_n16343, new_n16339, new_n22983);
not_10 g20635(new_n22983, new_n22984);
and_5  g20636(new_n22984, new_n22982, new_n22985);
not_10 g20637(new_n22985, new_n22986);
nand_5 g20638(new_n16344, new_n16338, new_n22987);
nor_5  g20639(new_n16344, new_n16338, new_n22988);
nand_5 g20640(new_n16298, new_n16300, new_n22989);
or_5   g20641(new_n16298, new_n16300, new_n22990);
nand_5 g20642(new_n19675, new_n22990, new_n22991);
and_5  g20643(new_n22991, new_n22989, new_n22992);
or_5   g20644(new_n22992, new_n22988, new_n22993);
and_5  g20645(new_n22993, new_n22987, new_n22994);
and_5  g20646(new_n22994, new_n22986, new_n22995);
xor_4  g20647(new_n22995, new_n3399, new_n22996);
xnor_4 g20648(new_n22994, new_n22985, new_n22997);
and_5  g20649(new_n22997, new_n3316_1, new_n22998_1);
xnor_4 g20650(new_n22997, new_n3316_1, new_n22999);
xnor_4 g20651(new_n22992, new_n16345, new_n23000);
or_5   g20652(new_n23000, new_n3201, new_n23001);
xor_4  g20653(new_n23000, new_n3201, new_n23002);
or_5   g20654(new_n19676, new_n3208_1, new_n23003);
or_5   g20655(new_n19718, new_n19677, new_n23004);
and_5  g20656(new_n23004, new_n23003, new_n23005);
nand_5 g20657(new_n23005, new_n23002, new_n23006_1);
and_5  g20658(new_n23006_1, new_n23001, new_n23007_1);
nor_5  g20659(new_n23007_1, new_n22999, new_n23008);
nor_5  g20660(new_n23008, new_n22998_1, new_n23009_1);
xor_4  g20661(new_n23009_1, new_n22996, n10775);
xnor_4 g20662(new_n21473, new_n21467, n10780);
xnor_4 g20663(n17095, n1689, new_n23012);
or_5   g20664(n22591, n22274, new_n23013);
and_5  g20665(n26167, n24129, new_n23014_1);
xnor_4 g20666(n22591, n22274, new_n23015);
or_5   g20667(new_n23015, new_n23014_1, new_n23016);
and_5  g20668(new_n23016, new_n23013, new_n23017);
xor_4  g20669(new_n23017, new_n23012, new_n23018);
xor_4  g20670(new_n23018, new_n21164, new_n23019);
nor_5  g20671(new_n9091, new_n9090_1, new_n23020);
or_5   g20672(new_n23020, n7769, new_n23021);
xnor_4 g20673(new_n23015, new_n23014_1, new_n23022);
xor_4  g20674(new_n23020, n7769, new_n23023);
nand_5 g20675(new_n23023, new_n23022, new_n23024);
and_5  g20676(new_n23024, new_n23021, new_n23025);
xor_4  g20677(new_n23025, new_n23019, new_n23026);
xnor_4 g20678(new_n23026, new_n18846, new_n23027);
xor_4  g20679(new_n23023, new_n23022, new_n23028);
nand_5 g20680(new_n23028, new_n18850, new_n23029);
nor_5  g20681(new_n9092, new_n9089, new_n23030);
xor_4  g20682(new_n23028, new_n18850, new_n23031);
nand_5 g20683(new_n23031, new_n23030, new_n23032);
and_5  g20684(new_n23032, new_n23029, new_n23033);
xor_4  g20685(new_n23033, new_n23027, n10817);
nand_5 g20686(new_n22206, new_n22203, new_n23035_1);
nand_5 g20687(new_n22202, new_n22199, new_n23036);
nor_5  g20688(new_n22206, new_n22203, new_n23037);
or_5   g20689(new_n22210, new_n23037, new_n23038);
and_5  g20690(new_n23038, new_n23036, new_n23039_1);
and_5  g20691(new_n23039_1, new_n23035_1, new_n23040);
or_5   g20692(new_n23040, new_n7829, new_n23041);
nor_5  g20693(new_n22211, new_n7829, new_n23042);
not_10 g20694(new_n22216, new_n23043);
and_5  g20695(new_n23043, new_n22213_1, new_n23044);
nor_5  g20696(new_n23044, new_n23042, new_n23045);
xor_4  g20697(new_n23040, new_n7829, new_n23046);
nand_5 g20698(new_n23046, new_n23045, new_n23047_1);
and_5  g20699(new_n23047_1, new_n23041, n10834);
xor_4  g20700(new_n22455, new_n22439, n10851);
xor_4  g20701(new_n21985, new_n21975, n10874);
xor_4  g20702(new_n22643, new_n22634, new_n23051);
xor_4  g20703(new_n23051, new_n8163, n10924);
or_5   g20704(new_n11334, new_n11328, new_n23053);
nand_5 g20705(new_n11397, new_n11335, new_n23054);
and_5  g20706(new_n23054, new_n23053, n10943);
xor_4  g20707(new_n12177, new_n12131_1, n10961);
xnor_4 g20708(new_n10804, new_n10794, n11005);
xnor_4 g20709(new_n21738, new_n21729, n11023);
nor_5  g20710(new_n18506, new_n7312, new_n23059);
xor_4  g20711(new_n18506, new_n21323, new_n23060);
or_5   g20712(new_n18508, new_n7316, new_n23061);
xor_4  g20713(new_n18508, new_n7316, new_n23062);
nand_5 g20714(new_n17210, new_n7321, new_n23063);
xnor_4 g20715(new_n17210, new_n7321, new_n23064);
nand_5 g20716(new_n12358, new_n7326, new_n23065_1);
or_5   g20717(new_n12384_1, new_n12359, new_n23066_1);
and_5  g20718(new_n23066_1, new_n23065_1, new_n23067_1);
or_5   g20719(new_n23067_1, new_n23064, new_n23068_1);
and_5  g20720(new_n23068_1, new_n23063, new_n23069);
nand_5 g20721(new_n23069, new_n23062, new_n23070);
and_5  g20722(new_n23070, new_n23061, new_n23071);
nor_5  g20723(new_n23071, new_n23060, new_n23072);
nor_5  g20724(new_n23072, new_n23059, new_n23073);
nor_5  g20725(new_n23073, new_n7294, new_n23074);
and_5  g20726(new_n23074, new_n18535, new_n23075);
not_10 g20727(new_n23075, new_n23076);
not_10 g20728(new_n22596, new_n23077);
xor_4  g20729(new_n23073, new_n7294, new_n23078);
xor_4  g20730(new_n23078, new_n18534, new_n23079);
and_5  g20731(new_n23079, new_n23077, new_n23080);
xor_4  g20732(new_n23079, new_n23077, new_n23081);
not_10 g20733(new_n23081, new_n23082);
xor_4  g20734(new_n23071, new_n23060, new_n23083);
and_5  g20735(new_n23083, new_n22604, new_n23084);
xor_4  g20736(new_n23083, new_n22604, new_n23085);
not_10 g20737(new_n23085, new_n23086);
xor_4  g20738(new_n23069, new_n23062, new_n23087);
and_5  g20739(new_n23087, new_n22607, new_n23088);
not_10 g20740(new_n23088, new_n23089);
xnor_4 g20741(new_n23087, new_n22608, new_n23090);
xor_4  g20742(new_n23067_1, new_n23064, new_n23091);
nor_5  g20743(new_n23091, new_n17973, new_n23092);
xor_4  g20744(new_n23091, new_n17973, new_n23093);
not_10 g20745(new_n23093, new_n23094);
nor_5  g20746(new_n12385, new_n12355, new_n23095);
nor_5  g20747(new_n12430, new_n12387, new_n23096);
nor_5  g20748(new_n23096, new_n23095, new_n23097);
nor_5  g20749(new_n23097, new_n23094, new_n23098);
nor_5  g20750(new_n23098, new_n23092, new_n23099);
not_10 g20751(new_n23099, new_n23100);
and_5  g20752(new_n23100, new_n23090, new_n23101);
not_10 g20753(new_n23101, new_n23102);
and_5  g20754(new_n23102, new_n23089, new_n23103);
nor_5  g20755(new_n23103, new_n23086, new_n23104);
nor_5  g20756(new_n23104, new_n23084, new_n23105);
nor_5  g20757(new_n23105, new_n23082, new_n23106);
nor_5  g20758(new_n23106, new_n23080, new_n23107);
nor_5  g20759(new_n23107, new_n23076, new_n23108);
not_10 g20760(new_n22627, new_n23109);
xor_4  g20761(new_n23107, new_n23076, new_n23110);
nor_5  g20762(new_n23110, new_n23109, new_n23111);
or_5   g20763(new_n23111, new_n23108, n11025);
xor_4  g20764(new_n16836, new_n8798, new_n23113);
not_10 g20765(new_n23113, new_n23114);
or_5   g20766(new_n16839, new_n8802, new_n23115);
xor_4  g20767(new_n16839, new_n8802, new_n23116);
not_10 g20768(new_n23116, new_n23117);
or_5   g20769(new_n16842, new_n8806_1, new_n23118);
xor_4  g20770(new_n16842, new_n8806_1, new_n23119);
not_10 g20771(new_n23119, new_n23120_1);
or_5   g20772(new_n16845, new_n8810, new_n23121);
or_5   g20773(new_n19546, new_n19543, new_n23122);
and_5  g20774(new_n23122, new_n23121, new_n23123);
or_5   g20775(new_n23123, new_n23120_1, new_n23124);
and_5  g20776(new_n23124, new_n23118, new_n23125);
or_5   g20777(new_n23125, new_n23117, new_n23126);
and_5  g20778(new_n23126, new_n23115, new_n23127);
xor_4  g20779(new_n23127, new_n23114, new_n23128);
not_10 g20780(n3795, new_n23129);
not_10 g20781(n25464, new_n23130);
not_10 g20782(n4590, new_n23131);
and_5  g20783(new_n19549, new_n19548, new_n23132);
and_5  g20784(new_n23132, new_n23131, new_n23133);
and_5  g20785(new_n23133, new_n23130, new_n23134);
xor_4  g20786(new_n23134, new_n23129, new_n23135);
xor_4  g20787(new_n23135, new_n8958, new_n23136);
xor_4  g20788(new_n23133, new_n23130, new_n23137);
or_5   g20789(new_n23137, new_n8960, new_n23138);
xor_4  g20790(new_n23137, new_n8965, new_n23139);
xor_4  g20791(new_n23132, new_n23131, new_n23140);
or_5   g20792(new_n23140, new_n8967, new_n23141);
xor_4  g20793(new_n23140, new_n8968, new_n23142);
or_5   g20794(new_n19550, new_n8972, new_n23143);
or_5   g20795(new_n19555, new_n19551, new_n23144);
and_5  g20796(new_n23144, new_n23143, new_n23145);
or_5   g20797(new_n23145, new_n23142, new_n23146_1);
and_5  g20798(new_n23146_1, new_n23141, new_n23147);
or_5   g20799(new_n23147, new_n23139, new_n23148);
and_5  g20800(new_n23148, new_n23138, new_n23149);
xor_4  g20801(new_n23149, new_n23136, new_n23150);
xnor_4 g20802(new_n23150, new_n23128, new_n23151);
xor_4  g20803(new_n23125, new_n23117, new_n23152);
xnor_4 g20804(new_n23147, new_n23139, new_n23153);
nor_5  g20805(new_n23153, new_n23152, new_n23154);
xor_4  g20806(new_n23147, new_n23139, new_n23155);
xnor_4 g20807(new_n23155, new_n23152, new_n23156);
not_10 g20808(new_n23156, new_n23157);
xor_4  g20809(new_n23123, new_n23120_1, new_n23158);
xnor_4 g20810(new_n23145, new_n23142, new_n23159);
nor_5  g20811(new_n23159, new_n23158, new_n23160_1);
xor_4  g20812(new_n23145, new_n23142, new_n23161);
xnor_4 g20813(new_n23161, new_n23158, new_n23162);
not_10 g20814(new_n23162, new_n23163);
xnor_4 g20815(new_n19555, new_n19551, new_n23164);
nor_5  g20816(new_n23164, new_n19547, new_n23165);
nor_5  g20817(new_n19561, new_n19558, new_n23166_1);
nor_5  g20818(new_n23166_1, new_n23165, new_n23167);
nor_5  g20819(new_n23167, new_n23163, new_n23168);
nor_5  g20820(new_n23168, new_n23160_1, new_n23169);
nor_5  g20821(new_n23169, new_n23157, new_n23170);
or_5   g20822(new_n23170, new_n23154, new_n23171);
xnor_4 g20823(new_n23171, new_n23151, n11063);
xnor_4 g20824(new_n20777, new_n20767, n11078);
xnor_4 g20825(new_n21476, new_n21463, n11080);
xnor_4 g20826(new_n14138, new_n14121_1, n11094);
xnor_4 g20827(new_n22808, new_n22807, n11101);
xnor_4 g20828(new_n21547, new_n14732, new_n23177);
xor_4  g20829(new_n23177, new_n21550, n11103);
xnor_4 g20830(new_n6625, new_n6598, n11120);
xor_4  g20831(new_n5031_1, new_n5027, n11127);
xor_4  g20832(new_n15344, new_n15342, n11132);
xnor_4 g20833(new_n11389, new_n11345, n11134);
xnor_4 g20834(new_n3706, new_n3705, n11138);
xnor_4 g20835(new_n10699, new_n10687, n11182);
xor_4  g20836(new_n14148_1, new_n14103, n11234);
xor_4  g20837(new_n22178, new_n19019, new_n23186);
and_5  g20838(new_n21811, new_n19023, new_n23187);
nor_5  g20839(new_n21840, new_n21813, new_n23188);
nor_5  g20840(new_n23188, new_n23187, new_n23189);
xor_4  g20841(new_n23189, new_n23186, n11245);
xor_4  g20842(new_n8793, new_n8779, n11261);
xnor_4 g20843(new_n23169, new_n23157, n11275);
nand_5 g20844(new_n13839, new_n13770, n11290);
xnor_4 g20845(new_n9620, new_n9618, n11313);
xor_4  g20846(new_n17189, new_n16612, new_n23195);
xor_4  g20847(new_n23195, new_n17202_1, n11325);
xnor_4 g20848(new_n14196, new_n14195, n11326);
xor_4  g20849(new_n17426, new_n17396, n11330);
xnor_4 g20850(new_n11382, new_n11357, n11347);
xnor_4 g20851(new_n22883, new_n22876, n11348);
xnor_4 g20852(new_n15461, new_n15450, n11352);
and_5  g20853(n22442, new_n22316, new_n23202);
xor_4  g20854(n22442, n3324, new_n23203);
or_5   g20855(n17911, new_n8414, new_n23204);
and_5  g20856(new_n19296, n5400, new_n23205);
nor_5  g20857(new_n17632, new_n17624, new_n23206);
or_5   g20858(new_n23206, new_n23205, new_n23207);
xnor_4 g20859(n17911, n468, new_n23208);
nand_5 g20860(new_n23208, new_n23207, new_n23209);
and_5  g20861(new_n23209, new_n23204, new_n23210);
nor_5  g20862(new_n23210, new_n23203, new_n23211);
nor_5  g20863(new_n23211, new_n23202, new_n23212);
not_10 g20864(new_n23212, new_n23213);
and_5  g20865(new_n18164, new_n18158, new_n23214);
nor_5  g20866(new_n23214, new_n7778, new_n23215);
nor_5  g20867(new_n18164, new_n18158, new_n23216);
not_10 g20868(new_n23216, new_n23217);
and_5  g20869(new_n23217, new_n7778, new_n23218);
nor_5  g20870(new_n23218, new_n23215, new_n23219);
xor_4  g20871(new_n23219, new_n23213, new_n23220);
or_5   g20872(new_n23213, new_n18166, new_n23221);
and_5  g20873(new_n23213, new_n18166, new_n23222);
not_10 g20874(new_n23222, new_n23223);
xor_4  g20875(new_n23210, new_n23203, new_n23224);
nor_5  g20876(new_n23224, new_n18168, new_n23225);
not_10 g20877(new_n23225, new_n23226);
xor_4  g20878(new_n23224, new_n18168, new_n23227);
xor_4  g20879(new_n23208, new_n23207, new_n23228);
and_5  g20880(new_n23228, new_n18170, new_n23229);
xnor_4 g20881(new_n23228, new_n18170, new_n23230);
nand_5 g20882(new_n17633, new_n17623, new_n23231);
or_5   g20883(new_n17644, new_n17634, new_n23232);
and_5  g20884(new_n23232, new_n23231, new_n23233);
nor_5  g20885(new_n23233, new_n23230, new_n23234);
nor_5  g20886(new_n23234, new_n23229, new_n23235);
and_5  g20887(new_n23235, new_n23227, new_n23236);
not_10 g20888(new_n23236, new_n23237);
and_5  g20889(new_n23237, new_n23226, new_n23238_1);
nand_5 g20890(new_n23238_1, new_n23223, new_n23239);
and_5  g20891(new_n23239, new_n23221, new_n23240);
xor_4  g20892(new_n23240, new_n23220, n11375);
xor_4  g20893(new_n12802, new_n7198, n11379);
or_5   g20894(new_n12189, n2570, new_n23243);
or_5   g20895(new_n16833, new_n16804, new_n23244);
and_5  g20896(new_n23244, new_n23243, new_n23245);
xor_4  g20897(new_n23245, new_n12241, new_n23246);
or_5   g20898(new_n16834_1, new_n12194, new_n23247_1);
or_5   g20899(new_n16868, new_n16835, new_n23248_1);
and_5  g20900(new_n23248_1, new_n23247_1, new_n23249);
xor_4  g20901(new_n23249, new_n23246, new_n23250_1);
xnor_4 g20902(new_n23250_1, new_n6380, new_n23251);
and_5  g20903(new_n16869, new_n16803, new_n23252);
nor_5  g20904(new_n16917, new_n16871, new_n23253);
nor_5  g20905(new_n23253, new_n23252, new_n23254);
xnor_4 g20906(new_n23254, new_n23251, n11386);
xnor_4 g20907(new_n19708, new_n19694, n11391);
xnor_4 g20908(new_n21797, new_n21795, n11398);
xor_4  g20909(new_n13120, new_n13119, n11403);
xnor_4 g20910(new_n12520, new_n12514, n11419);
xnor_4 g20911(new_n19531_1, new_n19515_1, n11439);
xnor_4 g20912(n7569, n2570, new_n23261);
or_5   g20913(n19033, n17037, new_n23262);
xnor_4 g20914(n19033, n17037, new_n23263);
or_5   g20915(n5386, n655, new_n23264);
xnor_4 g20916(n5386, n655, new_n23265);
or_5   g20917(n26191, n18145, new_n23266);
xnor_4 g20918(n26191, n18145, new_n23267);
or_5   g20919(n26512, n10712, new_n23268);
xnor_4 g20920(n26512, n10712, new_n23269);
or_5   g20921(n25126, n19575, new_n23270_1);
xor_4  g20922(n25126, n19575, new_n23271);
nand_5 g20923(n19608, n15378, new_n23272_1);
or_5   g20924(n19608, n15378, new_n23273);
nor_5  g20925(n17095, n1689, new_n23274);
nor_5  g20926(new_n23017, new_n23012, new_n23275);
nor_5  g20927(new_n23275, new_n23274, new_n23276);
nand_5 g20928(new_n23276, new_n23273, new_n23277);
and_5  g20929(new_n23277, new_n23272_1, new_n23278);
nand_5 g20930(new_n23278, new_n23271, new_n23279);
and_5  g20931(new_n23279, new_n23270_1, new_n23280);
or_5   g20932(new_n23280, new_n23269, new_n23281);
and_5  g20933(new_n23281, new_n23268, new_n23282);
or_5   g20934(new_n23282, new_n23267, new_n23283);
and_5  g20935(new_n23283, new_n23266, new_n23284);
or_5   g20936(new_n23284, new_n23265, new_n23285);
and_5  g20937(new_n23285, new_n23264, new_n23286);
or_5   g20938(new_n23286, new_n23263, new_n23287);
and_5  g20939(new_n23287, new_n23262, new_n23288);
xor_4  g20940(new_n23288, new_n23261, new_n23289_1);
nor_5  g20941(new_n23289_1, n10514, new_n23290);
not_10 g20942(new_n23290, new_n23291);
xor_4  g20943(new_n23289_1, n10514, new_n23292);
xor_4  g20944(new_n23286, new_n23263, new_n23293);
nand_5 g20945(new_n23293, n18649, new_n23294);
xor_4  g20946(new_n23293, new_n21144, new_n23295);
xor_4  g20947(new_n23284, new_n23265, new_n23296);
nand_5 g20948(new_n23296, n6218, new_n23297);
xor_4  g20949(new_n23296, new_n21148, new_n23298);
xor_4  g20950(new_n23282, new_n23267, new_n23299);
nand_5 g20951(new_n23299, n20470, new_n23300);
xor_4  g20952(new_n23299, new_n21152, new_n23301);
xor_4  g20953(new_n23280, new_n23269, new_n23302);
nand_5 g20954(new_n23302, n21222, new_n23303);
xor_4  g20955(new_n23302, new_n21155, new_n23304_1);
xor_4  g20956(new_n23278, new_n23271, new_n23305_1);
nand_5 g20957(new_n23305_1, n9832, new_n23306);
xor_4  g20958(new_n23305_1, n9832, new_n23307);
xor_4  g20959(n19608, n15378, new_n23308);
xor_4  g20960(new_n23308, new_n23276, new_n23309);
nand_5 g20961(new_n23309, new_n21161, new_n23310);
xor_4  g20962(new_n23309, n1558, new_n23311);
or_5   g20963(new_n23018, n21749, new_n23312);
or_5   g20964(new_n23025, new_n23019, new_n23313);
and_5  g20965(new_n23313, new_n23312, new_n23314);
or_5   g20966(new_n23314, new_n23311, new_n23315);
and_5  g20967(new_n23315, new_n23310, new_n23316);
nand_5 g20968(new_n23316, new_n23307, new_n23317);
and_5  g20969(new_n23317, new_n23306, new_n23318);
or_5   g20970(new_n23318, new_n23304_1, new_n23319);
and_5  g20971(new_n23319, new_n23303, new_n23320);
or_5   g20972(new_n23320, new_n23301, new_n23321);
and_5  g20973(new_n23321, new_n23300, new_n23322);
or_5   g20974(new_n23322, new_n23298, new_n23323);
and_5  g20975(new_n23323, new_n23297, new_n23324);
or_5   g20976(new_n23324, new_n23295, new_n23325);
and_5  g20977(new_n23325, new_n23294, new_n23326);
and_5  g20978(new_n23326, new_n23292, new_n23327);
not_10 g20979(new_n23327, new_n23328);
and_5  g20980(new_n23328, new_n23291, new_n23329);
or_5   g20981(n7569, n2570, new_n23330);
or_5   g20982(new_n23288, new_n23261, new_n23331);
and_5  g20983(new_n23331, new_n23330, new_n23332);
xnor_4 g20984(new_n23332, new_n23329, new_n23333_1);
and_5  g20985(new_n23134, new_n23129, new_n23334);
and_5  g20986(new_n23334, new_n12546_1, new_n23335);
xor_4  g20987(new_n23335, new_n11334, new_n23336);
xor_4  g20988(new_n23334, new_n12546_1, new_n23337);
nor_5  g20989(new_n23337, new_n8891, new_n23338);
not_10 g20990(new_n23338, new_n23339);
xnor_4 g20991(new_n23337, new_n8892, new_n23340);
not_10 g20992(new_n23340, new_n23341_1);
or_5   g20993(new_n23135, new_n8953, new_n23342_1);
or_5   g20994(new_n23149, new_n23136, new_n23343);
and_5  g20995(new_n23343, new_n23342_1, new_n23344);
nor_5  g20996(new_n23344, new_n23341_1, new_n23345);
not_10 g20997(new_n23345, new_n23346);
and_5  g20998(new_n23346, new_n23339, new_n23347);
xor_4  g20999(new_n23347, new_n23336, new_n23348);
xor_4  g21000(new_n23348, new_n23333_1, new_n23349);
xor_4  g21001(new_n23326, new_n23292, new_n23350);
not_10 g21002(new_n23350, new_n23351);
xnor_4 g21003(new_n23344, new_n23340, new_n23352);
and_5  g21004(new_n23352, new_n23351, new_n23353);
xor_4  g21005(new_n23352, new_n23351, new_n23354);
xor_4  g21006(new_n23324, new_n23295, new_n23355_1);
and_5  g21007(new_n23355_1, new_n23150, new_n23356);
xor_4  g21008(new_n23355_1, new_n23150, new_n23357);
not_10 g21009(new_n23357, new_n23358);
xor_4  g21010(new_n23322, new_n23298, new_n23359);
nand_5 g21011(new_n23359, new_n23155, new_n23360);
xor_4  g21012(new_n23359, new_n23155, new_n23361);
not_10 g21013(new_n23361, new_n23362);
xor_4  g21014(new_n23320, new_n23301, new_n23363);
nand_5 g21015(new_n23363, new_n23161, new_n23364);
xor_4  g21016(new_n23363, new_n23161, new_n23365);
not_10 g21017(new_n23365, new_n23366);
xor_4  g21018(new_n23318, new_n23304_1, new_n23367);
nand_5 g21019(new_n23367, new_n19556, new_n23368);
xor_4  g21020(new_n23367, new_n19556, new_n23369_1);
not_10 g21021(new_n23369_1, new_n23370);
xor_4  g21022(new_n23316, new_n23307, new_n23371_1);
nand_5 g21023(new_n23371_1, new_n18816, new_n23372);
xnor_4 g21024(new_n23371_1, new_n18817, new_n23373);
xor_4  g21025(new_n23314, new_n23311, new_n23374);
or_5   g21026(new_n23374, new_n18840, new_n23375);
and_5  g21027(new_n23026, new_n18846, new_n23376);
nor_5  g21028(new_n23033, new_n23027, new_n23377);
or_5   g21029(new_n23377, new_n23376, new_n23378);
xnor_4 g21030(new_n23374, new_n18839, new_n23379);
not_10 g21031(new_n23379, new_n23380);
or_5   g21032(new_n23380, new_n23378, new_n23381);
nand_5 g21033(new_n23381, new_n23375, new_n23382);
nand_5 g21034(new_n23382, new_n23373, new_n23383);
and_5  g21035(new_n23383, new_n23372, new_n23384);
or_5   g21036(new_n23384, new_n23370, new_n23385);
and_5  g21037(new_n23385, new_n23368, new_n23386);
or_5   g21038(new_n23386, new_n23366, new_n23387);
and_5  g21039(new_n23387, new_n23364, new_n23388);
or_5   g21040(new_n23388, new_n23362, new_n23389);
and_5  g21041(new_n23389, new_n23360, new_n23390);
nor_5  g21042(new_n23390, new_n23358, new_n23391);
nor_5  g21043(new_n23391, new_n23356, new_n23392);
not_10 g21044(new_n23392, new_n23393);
and_5  g21045(new_n23393, new_n23354, new_n23394);
nor_5  g21046(new_n23394, new_n23353, new_n23395);
xor_4  g21047(new_n23395, new_n23349, n11462);
xnor_4 g21048(new_n20784, new_n20755, n11470);
xor_4  g21049(new_n15795, new_n15779, n11472);
xor_4  g21050(new_n19357_1, new_n7371, new_n23399);
xor_4  g21051(new_n23399, new_n19379, n11496);
xnor_4 g21052(new_n20560, new_n20523, n11506);
xnor_4 g21053(new_n22349, new_n5755, new_n23402);
not_10 g21054(new_n23402, new_n23403);
and_5  g21055(new_n16162, new_n5761, new_n23404);
xnor_4 g21056(new_n16161, new_n5761, new_n23405);
not_10 g21057(new_n23405, new_n23406);
and_5  g21058(new_n10833, new_n5767, new_n23407);
xnor_4 g21059(new_n10832, new_n5767, new_n23408);
not_10 g21060(new_n23408, new_n23409);
xnor_4 g21061(new_n10829, new_n10828, new_n23410);
and_5  g21062(new_n23410, new_n5773, new_n23411);
xnor_4 g21063(new_n10851_1, new_n5773, new_n23412);
not_10 g21064(new_n23412, new_n23413);
and_5  g21065(new_n10859, new_n5779, new_n23414_1);
nor_5  g21066(new_n22956, new_n22939_1, new_n23415);
nor_5  g21067(new_n23415, new_n23414_1, new_n23416);
nor_5  g21068(new_n23416, new_n23413, new_n23417);
nor_5  g21069(new_n23417, new_n23411, new_n23418);
nor_5  g21070(new_n23418, new_n23409, new_n23419);
nor_5  g21071(new_n23419, new_n23407, new_n23420);
nor_5  g21072(new_n23420, new_n23406, new_n23421);
nor_5  g21073(new_n23421, new_n23404, new_n23422);
xnor_4 g21074(new_n23422, new_n23403, n11515);
xnor_4 g21075(new_n21486, new_n21449, n11538);
xor_4  g21076(new_n19142, new_n19141_1, n11548);
xnor_4 g21077(new_n19409, new_n19404, n11564);
and_5  g21078(n22442, new_n3409, new_n23427);
not_10 g21079(new_n23427, new_n23428);
nor_5  g21080(new_n22244, new_n22241, new_n23429_1);
not_10 g21081(new_n23429_1, new_n23430_1);
and_5  g21082(new_n23430_1, new_n23428, new_n23431);
not_10 g21083(new_n23431, new_n23432);
or_5   g21084(n3324, n2272, new_n23433_1);
or_5   g21085(new_n22249, new_n22246, new_n23434_1);
and_5  g21086(new_n23434_1, new_n23433_1, new_n23435);
nor_5  g21087(new_n23435, new_n7590, new_n23436);
not_10 g21088(new_n23436, new_n23437);
or_5   g21089(new_n22250, new_n7586, new_n23438);
or_5   g21090(new_n22255, new_n22251, new_n23439);
and_5  g21091(new_n23439, new_n23438, new_n23440);
xor_4  g21092(new_n23435, new_n7590, new_n23441);
and_5  g21093(new_n23441, new_n23440, new_n23442);
not_10 g21094(new_n23442, new_n23443);
and_5  g21095(new_n23443, new_n23437, new_n23444);
xor_4  g21096(new_n23444, new_n23432, new_n23445);
xor_4  g21097(new_n23441, new_n23440, new_n23446);
and_5  g21098(new_n23446, new_n23432, new_n23447);
xor_4  g21099(new_n23446, new_n23432, new_n23448);
and_5  g21100(new_n22256, new_n22245, new_n23449);
nor_5  g21101(new_n22260, new_n22257, new_n23450_1);
nor_5  g21102(new_n23450_1, new_n23449, new_n23451);
and_5  g21103(new_n23451, new_n23448, new_n23452);
nor_5  g21104(new_n23452, new_n23447, new_n23453);
xor_4  g21105(new_n23453, new_n23445, n11591);
or_5   g21106(new_n8468, new_n8462, new_n23455);
and_5  g21107(new_n8479, new_n8469, new_n23456);
or_5   g21108(new_n8479, new_n8469, new_n23457);
and_5  g21109(new_n8538, new_n23457, new_n23458);
not_10 g21110(new_n23458, new_n23459);
nand_5 g21111(new_n23459, new_n22959, new_n23460);
nor_5  g21112(new_n23460, new_n23456, new_n23461);
and_5  g21113(new_n23461, new_n23455, n11607);
xor_4  g21114(new_n19073, new_n19043, n11647);
xor_4  g21115(new_n23233, new_n23230, n11674);
xor_4  g21116(new_n20035, new_n15816_1, new_n23465);
or_5   g21117(new_n20048, new_n15999, new_n23466);
nand_5 g21118(new_n21799, new_n21786, new_n23467);
and_5  g21119(new_n23467, new_n23466, new_n23468);
xor_4  g21120(new_n23468, new_n23465, n11682);
xor_4  g21121(new_n22453, new_n22442_1, n11710);
xnor_4 g21122(new_n14142, new_n14113, n11712);
xor_4  g21123(new_n22120, new_n22106, n11724);
xnor_4 g21124(new_n18475, new_n18473, n11741);
xor_4  g21125(new_n18220, new_n3048, n11770);
xnor_4 g21126(new_n8522, new_n8521, n11771);
xnor_4 g21127(new_n19254, new_n19220_1, n11818);
xor_4  g21128(new_n22949, new_n22944, n11837);
and_5  g21129(new_n16500, new_n3533, new_n23478);
xor_4  g21130(new_n23478, new_n20241, new_n23479);
and_5  g21131(new_n23479, new_n5965, new_n23480_1);
not_10 g21132(new_n23480_1, new_n23481);
xor_4  g21133(new_n23479, new_n5966, new_n23482);
nand_5 g21134(new_n16501, new_n5970, new_n23483);
nand_5 g21135(new_n16537, new_n16502_1, new_n23484);
and_5  g21136(new_n23484, new_n23483, new_n23485);
nor_5  g21137(new_n23485, new_n23482, new_n23486);
not_10 g21138(new_n23486, new_n23487);
and_5  g21139(new_n23487, new_n23481, new_n23488);
and_5  g21140(new_n23478, new_n20241, new_n23489);
xor_4  g21141(new_n23489, new_n13717, new_n23490);
xor_4  g21142(new_n23490, new_n23488, new_n23491);
xnor_4 g21143(new_n23491, new_n22226, new_n23492);
xor_4  g21144(new_n23485, new_n23482, new_n23493_1);
nor_5  g21145(new_n23493_1, new_n21723, new_n23494);
xor_4  g21146(new_n23493_1, new_n21723, new_n23495);
not_10 g21147(new_n23495, new_n23496);
and_5  g21148(new_n16549, new_n16539, new_n23497);
not_10 g21149(new_n23497, new_n23498);
not_10 g21150(new_n16597, new_n23499);
and_5  g21151(new_n23499, new_n16550, new_n23500);
not_10 g21152(new_n23500, new_n23501);
and_5  g21153(new_n23501, new_n23498, new_n23502);
nor_5  g21154(new_n23502, new_n23496, new_n23503);
nor_5  g21155(new_n23503, new_n23494, new_n23504);
not_10 g21156(new_n23504, new_n23505);
xnor_4 g21157(new_n23505, new_n23492, n11842);
xnor_4 g21158(new_n16122, new_n16102, n11843);
xnor_4 g21159(new_n18860, new_n18843_1, n11905);
xnor_4 g21160(new_n11574, new_n11567, n11965);
xnor_4 g21161(new_n18734, new_n18731, n12000);
xor_4  g21162(new_n16674_1, new_n16671, n12003);
xor_4  g21163(new_n17271, new_n17270, n12011);
xnor_4 g21164(new_n17785, new_n17771, n12072);
xor_4  g21165(new_n10900, new_n10899, n12131);
xor_4  g21166(new_n16651, new_n16617_1, n12146);
xnor_4 g21167(new_n16905_1, new_n16899, n12157);
xnor_4 g21168(new_n10461, new_n10401, n12158);
xor_4  g21169(new_n22542, new_n22518, n12179);
xnor_4 g21170(new_n6449, new_n6393, n12192);
xnor_4 g21171(new_n22885, new_n22874, n12223);
xor_4  g21172(new_n10457, new_n10406, n12225);
xor_4  g21173(new_n22953, new_n22941, n12228);
xnor_4 g21174(new_n13650, new_n7246, n12235);
xor_4  g21175(new_n9266, new_n9235, n12302);
xnor_4 g21176(new_n17049, new_n17017, n12304);
xor_4  g21177(n19196, n1742, new_n23526);
or_5   g21178(new_n16811, n4858, new_n23527);
xor_4  g21179(n23586, n4858, new_n23528);
or_5   g21180(new_n16814, n8244, new_n23529_1);
xor_4  g21181(n21226, n8244, new_n23530);
or_5   g21182(n9493, new_n12210, new_n23531);
or_5   g21183(n20036, new_n6529, new_n23532);
or_5   g21184(new_n19975, new_n19970, new_n23533);
and_5  g21185(new_n23533, new_n23532, new_n23534);
xnor_4 g21186(n9493, n4426, new_n23535);
nand_5 g21187(new_n23535, new_n23534, new_n23536);
and_5  g21188(new_n23536, new_n23531, new_n23537);
or_5   g21189(new_n23537, new_n23530, new_n23538);
and_5  g21190(new_n23538, new_n23529_1, new_n23539);
or_5   g21191(new_n23539, new_n23528, new_n23540);
and_5  g21192(new_n23540, new_n23527, new_n23541_1);
xor_4  g21193(new_n23541_1, new_n23526, new_n23542);
xor_4  g21194(new_n23542, new_n19929, new_n23543);
not_10 g21195(new_n23543, new_n23544);
xor_4  g21196(new_n23539, new_n23528, new_n23545);
nor_5  g21197(new_n23545, new_n18456, new_n23546_1);
xor_4  g21198(new_n23545, new_n18456, new_n23547);
not_10 g21199(new_n23547, new_n23548);
xor_4  g21200(new_n23537, new_n23530, new_n23549);
nor_5  g21201(new_n23549, new_n18460, new_n23550_1);
xor_4  g21202(new_n23549, new_n18460, new_n23551);
xor_4  g21203(new_n23535, new_n23534, new_n23552);
nor_5  g21204(new_n23552, new_n18464, new_n23553);
xor_4  g21205(new_n23552, new_n18464, new_n23554);
nor_5  g21206(new_n19976, new_n18467_1, new_n23555);
nor_5  g21207(new_n19986, new_n19978, new_n23556);
nor_5  g21208(new_n23556, new_n23555, new_n23557);
not_10 g21209(new_n23557, new_n23558);
and_5  g21210(new_n23558, new_n23554, new_n23559);
nor_5  g21211(new_n23559, new_n23553, new_n23560);
not_10 g21212(new_n23560, new_n23561);
and_5  g21213(new_n23561, new_n23551, new_n23562);
nor_5  g21214(new_n23562, new_n23550_1, new_n23563);
nor_5  g21215(new_n23563, new_n23548, new_n23564);
nor_5  g21216(new_n23564, new_n23546_1, new_n23565);
xnor_4 g21217(new_n23565, new_n23544, n12324);
xnor_4 g21218(new_n21793, new_n21790, n12325);
xor_4  g21219(new_n10701_1, new_n10681, n12329);
xor_4  g21220(new_n8791, new_n8789, n12330);
xnor_4 g21221(new_n5819, new_n5764, n12346);
xor_4  g21222(new_n7707, new_n7679_1, n12349);
xnor_4 g21223(new_n19704, new_n19702, n12364);
nand_5 g21224(new_n22428, new_n22427, new_n23573);
nand_5 g21225(new_n23573, new_n5740, new_n23574);
xnor_4 g21226(new_n22429, new_n5740, new_n23575);
and_5  g21227(new_n23573, new_n9973, new_n23576);
xnor_4 g21228(new_n22429, new_n9973, new_n23577);
xnor_4 g21229(new_n22346, new_n22339, new_n23578);
and_5  g21230(new_n23578, new_n5749, new_n23579);
xnor_4 g21231(new_n22347, new_n5749, new_n23580);
not_10 g21232(new_n23580, new_n23581);
xnor_4 g21233(new_n22344, new_n22341_1, new_n23582);
and_5  g21234(new_n23582, new_n5755, new_n23583);
nor_5  g21235(new_n23422, new_n23403, new_n23584);
nor_5  g21236(new_n23584, new_n23583, new_n23585_1);
nor_5  g21237(new_n23585_1, new_n23581, new_n23586_1);
nor_5  g21238(new_n23586_1, new_n23579, new_n23587);
not_10 g21239(new_n23587, new_n23588_1);
and_5  g21240(new_n23588_1, new_n23577, new_n23589);
nor_5  g21241(new_n23589, new_n23576, new_n23590);
nand_5 g21242(new_n23590, new_n23575, new_n23591);
and_5  g21243(new_n23591, new_n23574, n12383);
xor_4  g21244(new_n8712, new_n8711, n12397);
xor_4  g21245(new_n17419, new_n17409, n12408);
nand_5 g21246(new_n20035, new_n15999, new_n23595);
or_5   g21247(new_n23468, new_n23465, new_n23596);
and_5  g21248(new_n23596, new_n23595, n12449);
xnor_4 g21249(new_n21564, new_n21532, n12461);
nor_5  g21250(new_n21397, new_n12241, new_n23599);
not_10 g21251(new_n23599, new_n23600);
and_5  g21252(new_n23600, new_n17510, new_n23601);
nor_5  g21253(new_n23600, new_n17510, new_n23602);
nor_5  g21254(new_n21398_1, new_n17564, new_n23603);
nor_5  g21255(new_n21409, new_n21400, new_n23604);
nor_5  g21256(new_n23604, new_n23603, new_n23605);
nor_5  g21257(new_n23605, new_n23602, new_n23606);
or_5   g21258(new_n23606, new_n23601, n12462);
xor_4  g21259(new_n22553, new_n22548, n12467);
nor_5  g21260(new_n16241, n3324, new_n23609);
nor_5  g21261(new_n16268, new_n16243_1, new_n23610);
nor_5  g21262(new_n23610, new_n23609, new_n23611);
not_10 g21263(new_n23611, new_n23612);
or_5   g21264(new_n23612, new_n22206, new_n23613);
or_5   g21265(new_n16345, new_n16337, new_n23614);
or_5   g21266(new_n16344, n13419, new_n23615);
and_5  g21267(new_n23615, new_n23614, new_n23616);
and_5  g21268(new_n23616, new_n22985, new_n23617);
xor_4  g21269(new_n23612, new_n22206, new_n23618);
xor_4  g21270(new_n23616, new_n22985, new_n23619_1);
or_5   g21271(new_n23619_1, new_n23618, new_n23620);
xor_4  g21272(new_n23619_1, new_n23618, new_n23621);
nor_5  g21273(new_n16346, new_n16269, new_n23622);
and_5  g21274(new_n16393, new_n16347, new_n23623);
nor_5  g21275(new_n23623, new_n23622, new_n23624_1);
nand_5 g21276(new_n23624_1, new_n23621, new_n23625);
and_5  g21277(new_n23625, new_n23620, new_n23626);
xor_4  g21278(new_n23626, new_n23617, new_n23627);
xor_4  g21279(new_n23627, new_n23613, n12469);
xnor_4 g21280(new_n11163, new_n11136, n12515);
and_5  g21281(n10250, new_n14262, new_n23630);
not_10 g21282(new_n23630, new_n23631);
xor_4  g21283(n10250, n5140, new_n23632);
or_5   g21284(new_n12199, n6204, new_n23633);
xor_4  g21285(n7674, n6204, new_n23634);
or_5   g21286(new_n12202, n3349, new_n23635);
xor_4  g21287(n6397, n3349, new_n23636);
or_5   g21288(new_n12205, n1742, new_n23637_1);
or_5   g21289(new_n23541_1, new_n23526, new_n23638);
and_5  g21290(new_n23638, new_n23637_1, new_n23639);
or_5   g21291(new_n23639, new_n23636, new_n23640);
and_5  g21292(new_n23640, new_n23635, new_n23641);
or_5   g21293(new_n23641, new_n23634, new_n23642);
and_5  g21294(new_n23642, new_n23633, new_n23643);
nor_5  g21295(new_n23643, new_n23632, new_n23644);
not_10 g21296(new_n23644, new_n23645);
and_5  g21297(new_n23645, new_n23631, new_n23646);
not_10 g21298(new_n23646, new_n23647);
xor_4  g21299(new_n23647, new_n22287, new_n23648);
and_5  g21300(new_n23646, new_n21123_1, new_n23649);
nor_5  g21301(new_n23646, new_n21123_1, new_n23650);
not_10 g21302(new_n23650, new_n23651);
xor_4  g21303(new_n23643, new_n23632, new_n23652);
nor_5  g21304(new_n23652, new_n21126, new_n23653);
xor_4  g21305(new_n23652, new_n21126, new_n23654);
not_10 g21306(new_n23654, new_n23655);
xor_4  g21307(new_n23641, new_n23634, new_n23656);
nor_5  g21308(new_n23656, new_n19922_1, new_n23657_1);
xor_4  g21309(new_n23656, new_n19922_1, new_n23658);
not_10 g21310(new_n23658, new_n23659);
xor_4  g21311(new_n23639, new_n23636, new_n23660);
nor_5  g21312(new_n23660, new_n19926, new_n23661);
xor_4  g21313(new_n23660, new_n19926, new_n23662);
nor_5  g21314(new_n23542, new_n19929, new_n23663_1);
nor_5  g21315(new_n23565, new_n23544, new_n23664);
nor_5  g21316(new_n23664, new_n23663_1, new_n23665);
not_10 g21317(new_n23665, new_n23666);
and_5  g21318(new_n23666, new_n23662, new_n23667);
nor_5  g21319(new_n23667, new_n23661, new_n23668);
nor_5  g21320(new_n23668, new_n23659, new_n23669_1);
nor_5  g21321(new_n23669_1, new_n23657_1, new_n23670);
nor_5  g21322(new_n23670, new_n23655, new_n23671);
nor_5  g21323(new_n23671, new_n23653, new_n23672);
and_5  g21324(new_n23672, new_n23651, new_n23673);
nor_5  g21325(new_n23673, new_n23649, new_n23674);
xor_4  g21326(new_n23674, new_n23648, n12516);
xor_4  g21327(new_n7476, new_n7464, n12540);
xnor_4 g21328(new_n11929, new_n11927, n12545);
xnor_4 g21329(new_n20782, new_n20759, n12552);
xnor_4 g21330(new_n8328, new_n8304, n12566);
xnor_4 g21331(new_n13609, new_n13590, n12569);
xnor_4 g21332(new_n6453, new_n6383_1, n12607);
xnor_4 g21333(new_n10259, new_n10177, n12620);
xnor_4 g21334(new_n3716, new_n3676, n12621);
xnor_4 g21335(new_n18661, new_n18659, n12654);
xor_4  g21336(new_n19979, new_n15365, n12665);
xnor_4 g21337(new_n17459, new_n17450_1, n12670);
xor_4  g21338(new_n7690, new_n2528, n12707);
xnor_4 g21339(new_n7201, new_n7191, n12725);
xnor_4 g21340(new_n16391, new_n16353, n12727);
xor_4  g21341(new_n9937, new_n9912, n12740);
xor_4  g21342(new_n21096, new_n21095_1, n12742);
xor_4  g21343(new_n21291, new_n2813, n12746);
xor_4  g21344(new_n9441, new_n9440, n12756);
xnor_4 g21345(new_n7218, new_n7157, n12783);
xor_4  g21346(new_n23646, new_n21123_1, new_n23695);
xor_4  g21347(new_n23695, new_n23672, n12801);
xor_4  g21348(new_n18114, new_n18107, n12812);
xnor_4 g21349(new_n16595, new_n16555, n12816);
or_5   g21350(new_n17654, n6659, new_n23699);
or_5   g21351(new_n18712, new_n18693_1, new_n23700);
and_5  g21352(new_n23700, new_n23699, new_n23701);
and_5  g21353(new_n23701, new_n20217, new_n23702);
xor_4  g21354(new_n23701, new_n20217, new_n23703);
or_5   g21355(new_n23703, new_n23618, new_n23704);
xor_4  g21356(new_n23703, new_n23618, new_n23705);
not_10 g21357(new_n23705, new_n23706);
nand_5 g21358(new_n18713, new_n16269, new_n23707);
or_5   g21359(new_n18742, new_n18715, new_n23708);
and_5  g21360(new_n23708, new_n23707, new_n23709);
or_5   g21361(new_n23709, new_n23706, new_n23710);
and_5  g21362(new_n23710, new_n23704, new_n23711);
or_5   g21363(new_n23711, new_n23702, new_n23712);
and_5  g21364(new_n23712, new_n23613, n12843);
xnor_4 g21365(new_n21339, new_n21338, n12864);
not_10 g21366(new_n19134, new_n23715);
or_5   g21367(new_n22670, new_n4857, new_n23716);
nand_5 g21368(new_n22695, new_n22671, new_n23717_1);
and_5  g21369(new_n23717_1, new_n23716, new_n23718);
nor_5  g21370(n21784, n3740, new_n23719_1);
nor_5  g21371(new_n22669, new_n22650, new_n23720);
or_5   g21372(new_n23720, new_n23719_1, new_n23721);
xor_4  g21373(new_n23721, new_n4916, new_n23722);
xor_4  g21374(new_n23722, new_n23718, new_n23723);
nor_5  g21375(new_n23723, new_n23715, new_n23724);
and_5  g21376(new_n22696, new_n17857, new_n23725);
and_5  g21377(new_n22722, new_n22697_1, new_n23726);
or_5   g21378(new_n23726, new_n23725, new_n23727);
xnor_4 g21379(new_n23723, new_n19134, new_n23728);
and_5  g21380(new_n23728, new_n23727, new_n23729);
nor_5  g21381(new_n23729, new_n23724, new_n23730);
or_5   g21382(new_n23721, new_n4916, new_n23731);
and_5  g21383(new_n23721, new_n4916, new_n23732);
or_5   g21384(new_n23732, new_n23718, new_n23733);
and_5  g21385(new_n23733, new_n23731, new_n23734);
and_5  g21386(new_n23734, new_n23730, n12865);
xnor_4 g21387(new_n13212, new_n13187, n12870);
xnor_4 g21388(new_n21300, new_n21279, n12873);
and_5  g21389(new_n22833, new_n18935, new_n23738);
xor_4  g21390(new_n22833, new_n18934, new_n23739);
and_5  g21391(new_n22178, new_n19019, new_n23740);
not_10 g21392(new_n23189, new_n23741);
and_5  g21393(new_n23741, new_n23186, new_n23742);
nor_5  g21394(new_n23742, new_n23740, new_n23743);
nor_5  g21395(new_n23743, new_n23739, new_n23744);
or_5   g21396(new_n23744, new_n23738, n12904);
xor_4  g21397(new_n10706, new_n10705, n12941);
xnor_4 g21398(new_n11446, new_n11438, n12942);
xnor_4 g21399(new_n5899, new_n3787, new_n23748_1);
xor_4  g21400(new_n23748_1, new_n5904_1, n12978);
xnor_4 g21401(new_n9952, new_n8024, n12980);
xor_4  g21402(new_n6612_1, new_n4720, n12985);
xnor_4 g21403(new_n14882, new_n14849_1, n12987);
and_5  g21404(new_n20890, n2160, new_n23753);
not_10 g21405(new_n23753, new_n23754);
nor_5  g21406(new_n17128, new_n17111, new_n23755_1);
not_10 g21407(new_n23755_1, new_n23756);
and_5  g21408(new_n23756, new_n23754, new_n23757);
xor_4  g21409(new_n23757, new_n15149, new_n23758);
and_5  g21410(new_n17129, new_n15188, new_n23759);
and_5  g21411(new_n17150, new_n17130_1, new_n23760);
nor_5  g21412(new_n23760, new_n23759, new_n23761);
xor_4  g21413(new_n23761, new_n23758, n12992);
nor_5  g21414(new_n22478, n6659, new_n23763);
nor_5  g21415(new_n21494, n23250, new_n23764);
nor_5  g21416(new_n21527, new_n21495, new_n23765);
nor_5  g21417(new_n23765, new_n23764, new_n23766);
and_5  g21418(new_n22478, n6659, new_n23767);
nor_5  g21419(new_n23767, new_n23766, new_n23768);
nor_5  g21420(new_n23768, new_n23763, new_n23769);
nor_5  g21421(new_n23769, new_n22477, new_n23770);
not_10 g21422(new_n23770, new_n23771);
xnor_4 g21423(new_n23771, new_n20226, new_n23772);
xnor_4 g21424(new_n22478, n6659, new_n23773);
xor_4  g21425(new_n23773, new_n23766, new_n23774);
nor_5  g21426(new_n23774, new_n20245, new_n23775_1);
nor_5  g21427(new_n21528, new_n14665, new_n23776);
and_5  g21428(new_n21566, new_n21529, new_n23777);
or_5   g21429(new_n23777, new_n23776, new_n23778);
xor_4  g21430(new_n23774, new_n20245, new_n23779);
and_5  g21431(new_n23779, new_n23778, new_n23780);
nor_5  g21432(new_n23780, new_n23775_1, new_n23781);
xor_4  g21433(new_n23781, new_n23772, n13005);
xor_4  g21434(new_n20327, new_n16990, n13043);
xnor_4 g21435(new_n18196, new_n18194, n13048);
xor_4  g21436(new_n15749_1, new_n15748, n13054);
xnor_4 g21437(new_n18366, new_n18354, n13082);
xnor_4 g21438(new_n7209, new_n7180, n13096);
xnor_4 g21439(new_n18368, new_n18347, n13116);
xor_4  g21440(new_n20342, new_n20308, n13122);
xnor_4 g21441(new_n6431_1, new_n6430, n13141);
xor_4  g21442(new_n20177, new_n20170, n13144);
xnor_4 g21443(new_n20788_1, new_n20747, n13168);
xnor_4 g21444(new_n21480, new_n21458, n13198);
xnor_4 g21445(new_n14876, new_n14860, n13199);
xnor_4 g21446(new_n14996, new_n14981, n13204);
xnor_4 g21447(new_n10448, new_n10421, n13209);
xnor_4 g21448(new_n19966, new_n19958, n13270);
xnor_4 g21449(new_n13491, new_n13466, n13273);
xor_4  g21450(new_n22544, new_n22513, n13285);
xnor_4 g21451(new_n21905_1, new_n21884, n13338);
xnor_4 g21452(new_n8036, new_n8012, n13407);
xnor_4 g21453(new_n5458, new_n4259, new_n23802);
xor_4  g21454(new_n23802, new_n16634, n13409);
xnor_4 g21455(new_n5472_1, new_n5442, n13456);
and_5  g21456(new_n21871, new_n21251, new_n23805);
and_5  g21457(new_n21765_1, new_n21141, new_n23806);
nor_5  g21458(new_n22921, new_n22918_1, new_n23807);
nor_5  g21459(new_n23807, new_n23806, new_n23808);
not_10 g21460(new_n23808, new_n23809);
nor_5  g21461(new_n21752, new_n21139, new_n23810);
nor_5  g21462(new_n23810, new_n23809, new_n23811);
and_5  g21463(new_n23811, new_n23805, new_n23812);
xor_4  g21464(new_n21752, new_n21251, new_n23813);
xor_4  g21465(new_n23813, new_n23809, new_n23814);
and_5  g21466(new_n23814, new_n11614, new_n23815);
xor_4  g21467(new_n23814, new_n11614, new_n23816);
nand_5 g21468(new_n22922, new_n11715, new_n23817);
or_5   g21469(new_n22926, new_n22923, new_n23818);
and_5  g21470(new_n23818, new_n23817, new_n23819);
and_5  g21471(new_n23819, new_n23816, new_n23820);
or_5   g21472(new_n23820, new_n23815, new_n23821);
xor_4  g21473(new_n21871, new_n21251, new_n23822);
and_5  g21474(new_n23822, new_n23808, new_n23823);
nor_5  g21475(new_n23822, new_n23811, new_n23824);
nor_5  g21476(new_n23824, new_n23823, new_n23825);
not_10 g21477(new_n23825, new_n23826);
and_5  g21478(new_n23826, new_n23821, new_n23827);
or_5   g21479(new_n23827, new_n23812, n13457);
xnor_4 g21480(new_n12462_1, new_n12452, n13477);
xor_4  g21481(new_n12818, new_n12816_1, n13484);
xnor_4 g21482(new_n20980, new_n20948, n13486);
xor_4  g21483(new_n22440, new_n21933, new_n23832);
or_5   g21484(new_n22358_1, new_n17739, new_n23833);
nand_5 g21485(new_n22386, new_n22359_1, new_n23834);
and_5  g21486(new_n23834, new_n23833, new_n23835);
xor_4  g21487(new_n23835, new_n23832, n13487);
xnor_4 g21488(new_n5236, new_n5214, n13500);
xor_4  g21489(new_n4587, new_n4585, n13501);
xor_4  g21490(new_n6438, new_n6414, n13506);
xnor_4 g21491(new_n6172, new_n6163, n13548);
xnor_4 g21492(new_n23386, new_n23366, n13551);
xnor_4 g21493(new_n5036, new_n5017, n13602);
xnor_4 g21494(new_n17841, new_n17831, n13626);
xor_4  g21495(new_n8323, new_n8314, n13683);
xnor_4 g21496(new_n20562, new_n20520, n13710);
xor_4  g21497(new_n20181, new_n20164, n13722);
xor_4  g21498(new_n14507, new_n14444, new_n23847);
xor_4  g21499(new_n23847, new_n14594, n13754);
xor_4  g21500(new_n2825, new_n2794, n13764);
xnor_4 g21501(new_n14735, new_n14732, new_n23850);
xor_4  g21502(new_n23850, new_n14739, n13798);
xnor_4 g21503(new_n17845, new_n17824, n13835);
xnor_4 g21504(new_n16215_1, new_n16214, n13850);
xor_4  g21505(new_n18356, new_n7883, n13922);
xor_4  g21506(new_n19937, new_n19928, n13923);
xnor_4 g21507(new_n11935, new_n11933, n14004);
xor_4  g21508(new_n12181, new_n12124, n14036);
xnor_4 g21509(new_n21989, new_n21971, n14059);
xor_4  g21510(new_n17642, new_n17638_1, n14081);
xor_4  g21511(new_n19373, new_n19367_1, n14095);
xor_4  g21512(new_n6760, new_n3367, n14107);
xnor_4 g21513(new_n9079, new_n9043, n14121);
xor_4  g21514(new_n12416, new_n12415, n14126);
xor_4  g21515(new_n20187_1, new_n20158, n14136);
not_10 g21516(new_n23757, new_n23865);
nor_5  g21517(new_n23865, new_n15149, new_n23866);
and_5  g21518(new_n23865, new_n15149, new_n23867);
nor_5  g21519(new_n23761, new_n23867, new_n23868);
nor_5  g21520(new_n23868, new_n23866, new_n23869);
xor_4  g21521(new_n23757, new_n22739, new_n23870);
xor_4  g21522(new_n23870, new_n23869, n14147);
xor_4  g21523(new_n21689, new_n21646, n14174);
xnor_4 g21524(new_n16913, new_n16881, n14190);
xnor_4 g21525(new_n5470, new_n5448, n14211);
xnor_4 g21526(new_n17098, new_n17095_1, n14222);
xor_4  g21527(new_n13833, new_n13783_1, n14267);
xor_4  g21528(new_n5806, new_n5794, n14271);
xnor_4 g21529(new_n9623, new_n9611, n14277);
xnor_4 g21530(new_n8517, new_n8515, n14294);
xnor_4 g21531(new_n23393, new_n23354, n14310);
xnor_4 g21532(new_n23416, new_n23413, n14326);
xnor_4 g21533(new_n12765, new_n12712, n14342);
xnor_4 g21534(new_n18858_1, new_n18849, n14353);
not_10 g21535(new_n21966, new_n23884);
nor_5  g21536(new_n23884, new_n11965_1, new_n23885);
nor_5  g21537(new_n21966, new_n9140, new_n23886);
and_5  g21538(new_n21992, new_n21967, new_n23887);
nor_5  g21539(new_n23887, new_n23886, new_n23888_1);
or_5   g21540(new_n23888_1, new_n23885, new_n23889);
and_5  g21541(new_n23884, new_n11965_1, new_n23890);
or_5   g21542(new_n23890, new_n23887, new_n23891);
and_5  g21543(new_n23891, new_n23889, n14364);
xor_4  g21544(new_n22448, new_n22445, n14375);
xnor_4 g21545(new_n22893, new_n22862, n14412);
not_10 g21546(new_n11878, new_n23895_1);
nor_5  g21547(new_n18060, new_n6273, new_n23896);
not_10 g21548(new_n23896, new_n23897);
nor_5  g21549(new_n18086, new_n23897, new_n23898);
xnor_4 g21550(new_n23898, new_n23895_1, new_n23899_1);
nor_5  g21551(new_n18087, new_n11879, new_n23900);
not_10 g21552(new_n18088, new_n23901);
nor_5  g21553(new_n18126, new_n23901, new_n23902);
nor_5  g21554(new_n23902, new_n23900, new_n23903_1);
xor_4  g21555(new_n23903_1, new_n23899_1, n14414);
xor_4  g21556(new_n15965, new_n15964, n14457);
xnor_4 g21557(new_n5040, new_n5005, n14464);
xnor_4 g21558(new_n11161, new_n11140, n14471);
nor_5  g21559(new_n20217, new_n8478, new_n23908);
not_10 g21560(new_n20218, new_n23909);
nor_5  g21561(new_n20225, new_n23909, new_n23910);
nor_5  g21562(new_n23910, new_n23908, new_n23911);
xor_4  g21563(new_n23911, new_n23771, new_n23912_1);
nor_5  g21564(new_n23771, new_n20226, new_n23913_1);
and_5  g21565(new_n23771, new_n20226, new_n23914);
nor_5  g21566(new_n23781, new_n23914, new_n23915);
nor_5  g21567(new_n23915, new_n23913_1, new_n23916);
xor_4  g21568(new_n23916, new_n23912_1, n14475);
xor_4  g21569(new_n12752, new_n12751, n14541);
not_10 g21570(new_n22219, new_n23919);
nor_5  g21571(new_n22224, new_n23919, new_n23920);
nor_5  g21572(new_n22235, new_n22225, new_n23921);
or_5   g21573(new_n23921, new_n23920, n14546);
xor_4  g21574(new_n11371, new_n11370, n14547);
xnor_4 g21575(new_n13128, new_n13108, n14593);
xnor_4 g21576(new_n9627, new_n9601, n14636);
xnor_4 g21577(new_n23563, new_n23548, n14701);
xnor_4 g21578(new_n12523, new_n12511, n14734);
xnor_4 g21579(new_n7216, new_n7163, n14746);
xnor_4 g21580(new_n9928, new_n9926_1, n14763);
xor_4  g21581(new_n23099, new_n23090, n14772);
xnor_4 g21582(new_n22451, new_n22450, n14801);
xnor_4 g21583(new_n22037, new_n22018, n14819);
xnor_4 g21584(new_n15008, new_n14965, n14827);
xnor_4 g21585(new_n21407, new_n21404_1, n14839);
xnor_4 g21586(new_n17837, new_n17836, n14849);
nor_5  g21587(new_n21249, new_n14946, new_n23936);
and_5  g21588(new_n21316, new_n21250, new_n23937);
nor_5  g21589(new_n23937, new_n23936, new_n23938);
nor_5  g21590(new_n23938, new_n21246, n14891);
xor_4  g21591(new_n6574, new_n4749, n14931);
nand_5 g21592(new_n23898, new_n23895_1, new_n23941);
nor_5  g21593(new_n23903_1, new_n23941, new_n23942_1);
nor_5  g21594(new_n23898, new_n23895_1, new_n23943);
and_5  g21595(new_n23903_1, new_n23943, new_n23944);
or_5   g21596(new_n23944, new_n23942_1, n14944);
xor_4  g21597(new_n18853, new_n9089, n14977);
xnor_4 g21598(new_n13137_1, new_n13085, n14989);
xnor_4 g21599(new_n11054, new_n11044_1, n15002);
xnor_4 g21600(new_n22947, new_n5803, n15004);
xor_4  g21601(new_n9274, new_n9223, n15011);
xor_4  g21602(new_n23005, new_n23002, n15019);
and_5  g21603(new_n15733, new_n15724, new_n23952);
nor_5  g21604(new_n15756, new_n15735, new_n23953);
or_5   g21605(new_n23953, new_n23952, n15031);
xor_4  g21606(new_n18357, new_n18356, n15033);
xor_4  g21607(new_n12288, new_n7246, n15052);
xnor_4 g21608(new_n20097, new_n20086_1, n15082);
xnor_4 g21609(new_n8326, new_n8309_1, n15094);
xor_4  g21610(new_n11996, new_n11993, n15118);
xnor_4 g21611(new_n23743, new_n23739, n15128);
xnor_4 g21612(new_n19258, new_n19212, n15139);
xnor_4 g21613(new_n17195, new_n17189, new_n23962);
xor_4  g21614(new_n23962, new_n17204, n15145);
xnor_4 g21615(new_n15231, new_n15193, n15165);
xor_4  g21616(new_n15667, new_n5100, n15176);
xor_4  g21617(new_n20775, new_n20774_1, n15180);
xnor_4 g21618(new_n16653, new_n16615, n15205);
xor_4  g21619(new_n5463, new_n16633, n15230);
xor_4  g21620(new_n17455, new_n17454, n15255);
xnor_4 g21621(new_n9941, new_n9903, n15275);
xnor_4 g21622(new_n14337, new_n14332, n15300);
nor_5  g21623(new_n23489, new_n13717, new_n23972);
and_5  g21624(new_n23972, new_n23488, new_n23973);
and_5  g21625(new_n23489, new_n13717, new_n23974_1);
not_10 g21626(new_n23974_1, new_n23975);
nor_5  g21627(new_n23975, new_n23488, new_n23976);
nor_5  g21628(new_n23976, new_n23973, new_n23977);
xor_4  g21629(new_n23977, new_n22219, new_n23978);
nor_5  g21630(new_n23491, new_n22182, new_n23979);
and_5  g21631(new_n23505, new_n23492, new_n23980);
nor_5  g21632(new_n23980, new_n23979, new_n23981);
xor_4  g21633(new_n23981, new_n23978, n15307);
xnor_4 g21634(new_n20564, new_n20517, n15327);
xnor_4 g21635(new_n20550, new_n20542, n15345);
xnor_4 g21636(new_n13125, new_n13115, n15353);
xor_4  g21637(new_n23590, new_n23575, n15366);
xnor_4 g21638(new_n23734, new_n23730, n15382);
xnor_4 g21639(new_n9448, new_n9429, n15407);
xor_4  g21640(new_n15362, new_n13916, n15428);
not_10 g21641(new_n23329, new_n23990);
nor_5  g21642(new_n23332, new_n23990, new_n23991);
not_10 g21643(new_n23991, new_n23992);
and_5  g21644(new_n23348, new_n23333_1, new_n23993);
not_10 g21645(new_n23395, new_n23994);
and_5  g21646(new_n23994, new_n23349, new_n23995);
nor_5  g21647(new_n23995, new_n23993, new_n23996);
not_10 g21648(new_n23996, new_n23997);
nand_5 g21649(new_n23997, new_n23992, new_n23998);
nor_5  g21650(new_n23335, new_n11334, new_n23999);
not_10 g21651(new_n23347, new_n24000);
and_5  g21652(new_n24000, new_n23999, new_n24001);
not_10 g21653(new_n24001, new_n24002_1);
nor_5  g21654(new_n24002_1, new_n23991, new_n24003);
or_5   g21655(new_n24003, new_n23995, new_n24004_1);
and_5  g21656(new_n24004_1, new_n23998, n15435);
or_5   g21657(new_n22964, new_n22959, new_n24006);
nor_5  g21658(new_n22974, new_n24006, new_n24007);
and_5  g21659(new_n22964, new_n22959, new_n24008);
and_5  g21660(new_n22974, new_n24008, new_n24009);
or_5   g21661(new_n24009, new_n24007, n15438);
xnor_4 g21662(new_n23388, new_n23362, n15465);
xor_4  g21663(new_n8711, new_n6700, n15467);
xnor_4 g21664(new_n8046, new_n7983, n15470);
xnor_4 g21665(new_n15012, new_n14957, n15477);
xnor_4 g21666(new_n23668, new_n23659, n15481);
xor_4  g21667(new_n15457, new_n15454, n15496);
xor_4  g21668(new_n12427, new_n12392, n15501);
xor_4  g21669(new_n19377, new_n19362, n15555);
xnor_4 g21670(new_n21838, new_n21817, n15558);
and_5  g21671(new_n23919, new_n22833, new_n24020);
nor_5  g21672(new_n22837, new_n22834, new_n24021);
or_5   g21673(new_n24021, new_n24020, n15559);
or_5   g21674(n23895, new_n22980, new_n24023);
or_5   g21675(new_n20814, new_n20795_1, new_n24024);
and_5  g21676(new_n24024, new_n24023, new_n24025);
nand_5 g21677(new_n24025, new_n23040, new_n24026);
and_5  g21678(new_n20860, new_n20815, new_n24027);
and_5  g21679(new_n20884, new_n20861, new_n24028);
nor_5  g21680(new_n24028, new_n24027, new_n24029);
nor_5  g21681(new_n24025, new_n22211, new_n24030);
nor_5  g21682(new_n24030, new_n24029, new_n24031);
not_10 g21683(new_n24031, new_n24032_1);
or_5   g21684(new_n24032_1, new_n23040, new_n24033);
nand_5 g21685(new_n24025, new_n22212, new_n24034);
nand_5 g21686(new_n24034, new_n24032_1, new_n24035);
and_5  g21687(new_n24035, new_n24033, new_n24036);
and_5  g21688(new_n24036, new_n24026, n15570);
xnor_4 g21689(new_n12771, new_n12694, n15573);
xnor_4 g21690(new_n11953, new_n11951, n15588);
xnor_4 g21691(new_n22032, new_n22024, n15590);
xnor_4 g21692(new_n22618, new_n22606, n15598);
xnor_4 g21693(new_n9629, new_n9596, n15614);
xnor_4 g21694(new_n23105, new_n23082, n15662);
xnor_4 g21695(new_n3384, new_n3348, n15716);
xnor_4 g21696(new_n14884, new_n14846, n15749);
xnor_4 g21697(new_n19287, new_n19281, n15762);
xnor_4 g21698(new_n9963, new_n8024, n15793);
xnor_4 g21699(new_n22887, new_n22871_1, n15812);
xnor_4 g21700(new_n12767, new_n12706, n15815);
xnor_4 g21701(new_n8513, new_n8511, n15816);
xnor_4 g21702(new_n12295, new_n12280, n15831);
xnor_4 g21703(new_n9802, new_n9801, n15846);
xnor_4 g21704(new_n8575, new_n8574, n15859);
not_10 g21705(new_n8207, new_n24054);
and_5  g21706(new_n8208, n23272, new_n24055);
and_5  g21707(new_n20434, new_n20419, new_n24056);
nor_5  g21708(new_n24056, new_n24055, new_n24057);
nor_5  g21709(new_n24057, new_n24054, new_n24058);
xor_4  g21710(new_n24058, new_n22272, new_n24059);
xor_4  g21711(new_n24057, new_n24054, new_n24060);
or_5   g21712(new_n24060, new_n22274_1, new_n24061);
or_5   g21713(new_n20435, new_n20417, new_n24062);
nand_5 g21714(new_n20460, new_n20436_1, new_n24063);
and_5  g21715(new_n24063, new_n24062, new_n24064);
xnor_4 g21716(new_n24060, new_n20737, new_n24065);
not_10 g21717(new_n24065, new_n24066);
or_5   g21718(new_n24066, new_n24064, new_n24067);
and_5  g21719(new_n24067, new_n24061, new_n24068);
xor_4  g21720(new_n24068, new_n24059, n15869);
xnor_4 g21721(new_n19420, new_n19395, n15885);
nor_5  g21722(new_n21642, new_n21571, new_n24071);
and_5  g21723(new_n21692, new_n24071, new_n24072);
and_5  g21724(new_n21691, new_n21642, new_n24073);
or_5   g21725(new_n24073, new_n24072, n15889);
xnor_4 g21726(new_n19407, new_n14195, n15917);
xor_4  g21727(new_n14188, new_n14187, n15922);
xor_4  g21728(new_n7193, new_n7192, n15947);
and_5  g21729(new_n20018, new_n7294, new_n24078);
and_5  g21730(new_n21329, new_n21321, new_n24079);
nor_5  g21731(new_n24079, new_n24078, new_n24080);
xnor_4 g21732(new_n24080, new_n20045, new_n24081);
nor_5  g21733(new_n21331, new_n20045, new_n24082);
not_10 g21734(new_n21342, new_n24083);
and_5  g21735(new_n24083, new_n21332, new_n24084);
nor_5  g21736(new_n24084, new_n24082, new_n24085_1);
xor_4  g21737(new_n24085_1, new_n24081, n15956);
xor_4  g21738(new_n13936, new_n13933, n15958);
nor_5  g21739(new_n17492, new_n12486, new_n24088);
not_10 g21740(new_n12490, new_n24089);
and_5  g21741(new_n17492, new_n24089, new_n24090);
or_5   g21742(new_n24090, new_n24088, new_n24091);
not_10 g21743(new_n17484, new_n24092_1);
nor_5  g21744(new_n24092_1, new_n12486, new_n24093_1);
nor_5  g21745(new_n17487, new_n24093_1, new_n24094);
and_5  g21746(new_n24094, new_n24091, n15986);
xnor_4 g21747(new_n23502, new_n23496, n16013);
nor_5  g21748(new_n22407, new_n21331, new_n24097_1);
and_5  g21749(new_n22407, new_n21331, new_n24098);
nor_5  g21750(new_n22417, new_n24098, new_n24099);
nor_5  g21751(new_n24099, new_n24097_1, new_n24100);
xnor_4 g21752(new_n24080, new_n22407, new_n24101);
xor_4  g21753(new_n24101, new_n24100, n16060);
or_5   g21754(new_n16834_1, new_n18520, new_n24103);
xor_4  g21755(new_n16834_1, n25972, new_n24104);
or_5   g21756(new_n16836, new_n8798, new_n24105_1);
or_5   g21757(new_n23127, new_n23114, new_n24106);
and_5  g21758(new_n24106, new_n24105_1, new_n24107);
or_5   g21759(new_n24107, new_n24104, new_n24108);
and_5  g21760(new_n24108, new_n24103, new_n24109);
nor_5  g21761(new_n24109, new_n23245, new_n24110);
not_10 g21762(new_n23348, new_n24111);
xor_4  g21763(new_n24109, new_n23245, new_n24112);
nor_5  g21764(new_n24112, new_n24111, new_n24113);
xnor_4 g21765(new_n24112, new_n23348, new_n24114);
not_10 g21766(new_n23352, new_n24115);
xor_4  g21767(new_n24107, new_n24104, new_n24116);
nor_5  g21768(new_n24116, new_n24115, new_n24117);
xnor_4 g21769(new_n24116, new_n23352, new_n24118);
xnor_4 g21770(new_n23149, new_n23136, new_n24119_1);
nor_5  g21771(new_n24119_1, new_n23128, new_n24120);
and_5  g21772(new_n23171, new_n23151, new_n24121);
or_5   g21773(new_n24121, new_n24120, new_n24122);
and_5  g21774(new_n24122, new_n24118, new_n24123);
or_5   g21775(new_n24123, new_n24117, new_n24124);
and_5  g21776(new_n24124, new_n24114, new_n24125);
nor_5  g21777(new_n24125, new_n24113, new_n24126);
xor_4  g21778(new_n24126, new_n24110, new_n24127);
xor_4  g21779(new_n24127, new_n24002_1, n16062);
xnor_4 g21780(new_n23588_1, new_n23577, n16068);
xnor_4 g21781(new_n23819, new_n23816, n16080);
and_5  g21782(new_n23250_1, new_n6380, new_n24131);
nor_5  g21783(new_n23254, new_n23251, new_n24132);
or_5   g21784(new_n24132, new_n24131, new_n24133_1);
nor_5  g21785(new_n23245, new_n12246, new_n24134);
not_10 g21786(new_n24134, new_n24135);
nor_5  g21787(new_n23249, new_n23246, new_n24136);
not_10 g21788(new_n24136, new_n24137);
and_5  g21789(new_n24137, new_n24135, new_n24138);
xor_4  g21790(new_n24138, new_n24133_1, n16098);
xnor_4 g21791(new_n18049, new_n18041, n16110);
xnor_4 g21792(new_n15607, new_n15577, n16142);
xnor_4 g21793(new_n17043, new_n17029, n16185);
xnor_4 g21794(new_n12814, new_n12791, n16196);
xnor_4 g21795(new_n21360, new_n21359, n16206);
xor_4  g21796(new_n21441, new_n21437, n16215);
xnor_4 g21797(new_n19529, new_n19519, n16218);
xor_4  g21798(new_n3921, new_n3920, n16219);
xnor_4 g21799(new_n6970, new_n6969, n16230);
xor_4  g21800(new_n8572, new_n8564, n16243);
xnor_4 g21801(new_n17783, new_n17774, n16275);
xor_4  g21802(new_n10452, new_n10450, n16279);
nor_5  g21803(new_n20927, new_n20085, new_n24152);
nor_5  g21804(new_n20990, new_n20928, new_n24153);
or_5   g21805(new_n24153, new_n24152, n16322);
xor_4  g21806(new_n17794, new_n17753, n16327);
xnor_4 g21807(new_n21832_1, new_n21824, n16350);
xor_4  g21808(new_n6702, new_n6700, n16367);
xor_4  g21809(new_n19634, new_n19632, n16379);
xnor_4 g21810(new_n20554, new_n20535, n16398);
xnor_4 g21811(new_n13923_1, new_n13922_1, n16406);
xnor_4 g21812(new_n22620_1, new_n22601, n16407);
xnor_4 g21813(new_n24124, new_n24114, n16419);
xnor_4 g21814(new_n8532, new_n8486, n16424);
xor_4  g21815(new_n14303, new_n14237, new_n24164);
xor_4  g21816(new_n24164, new_n14351, n16428);
xnor_4 g21817(new_n12315_1, new_n12245, n16433);
xnor_4 g21818(new_n12311, new_n12255, n16440);
xor_4  g21819(new_n18051, new_n18037, n16445);
xnor_4 g21820(new_n14589, new_n14520, n16460);
xnor_4 g21821(new_n20456, new_n20446, n16481);
or_5   g21822(new_n15186, new_n11328, new_n24171);
nor_5  g21823(new_n15186, new_n11336, new_n24172_1);
nor_5  g21824(new_n21054, new_n21036, new_n24173);
nor_5  g21825(new_n24173, new_n24172_1, new_n24174);
xor_4  g21826(new_n15186, new_n11328, new_n24175);
nand_5 g21827(new_n24175, new_n24174, new_n24176);
and_5  g21828(new_n24176, new_n24171, n16493);
xnor_4 g21829(new_n4765, new_n4737, n16506);
xnor_4 g21830(new_n13203, new_n13202, n16516);
xor_4  g21831(new_n22714_1, new_n22713, n16517);
xnor_4 g21832(new_n16114, new_n16112, n16527);
xnor_4 g21833(new_n11045, new_n9387, n16554);
xor_4  g21834(new_n6168, new_n6167, n16583);
xor_4  g21835(new_n22150_1, new_n10314, new_n24184);
xor_4  g21836(new_n24184, new_n22154, n16584);
xnor_4 g21837(new_n19712, new_n19686, n16589);
xor_4  g21838(new_n20064, new_n20063, n16596);
xnor_4 g21839(new_n22899, new_n22853, n16617);
xnor_4 g21840(new_n7713, new_n7670_1, n16630);
xor_4  g21841(new_n22880, new_n4950, n16640);
xor_4  g21842(new_n2528, new_n2526, n16656);
xor_4  g21843(new_n6989, new_n6931, n16674);
xor_4  g21844(new_n14585, new_n14526, n16682);
xor_4  g21845(new_n22813, new_n22793_1, n16684);
xnor_4 g21846(new_n10802, new_n10798, n16688);
xnor_4 g21847(new_n6434, new_n6424, n16733);
xor_4  g21848(new_n8032, new_n8031_1, n16798);
xnor_4 g21849(new_n17146, new_n17145, n16834);
xnor_4 g21850(new_n3069, new_n3022, n16837);
xnor_4 g21851(new_n22415, new_n22412, n16841);
xnor_4 g21852(new_n5103, new_n5102, n16885);
xor_4  g21853(new_n8340, new_n8272, n16905);
nor_5  g21854(new_n22331, new_n22327, new_n24203);
xor_4  g21855(new_n24203, new_n22329, n16951);
xor_4  g21856(new_n16638, new_n16628, n16954);
xor_4  g21857(new_n8510_1, new_n8509, n16989);
xnor_4 g21858(new_n19637, new_n19602_1, n17006);
xnor_4 g21859(new_n13813, new_n13812, n17068);
xnor_4 g21860(new_n15596, new_n15595, n17070);
xnor_4 g21861(new_n20986_1, new_n20936_1, n17075);
xnor_4 g21862(new_n17421_1, new_n17405, n17084);
xor_4  g21863(new_n4756, new_n4754, n17104);
xnor_4 g21864(new_n13611, new_n13585, n17106);
xor_4  g21865(new_n9933, new_n9922, n17119);
xnor_4 g21866(new_n13496, new_n13454, n17130);
xnor_4 g21867(new_n23384, new_n23370, n17138);
xnor_4 g21868(new_n22716, new_n22708, n17163);
xor_4  g21869(new_n20636, new_n20635, n17168);
xnor_4 g21870(new_n11744, new_n11735, n17202);
xor_4  g21871(new_n19883, new_n19881, n17219);
xor_4  g21872(new_n19075, new_n19037, n17232);
xnor_4 g21873(new_n15706, new_n15702, n17236);
xor_4  g21874(new_n10711, new_n10710_1, n17243);
xnor_4 g21875(new_n11377, new_n11363, n17263);
nand_5 g21876(new_n20046, new_n20035, new_n24225);
nand_5 g21877(new_n20068, new_n20047, new_n24226);
and_5  g21878(new_n24226, new_n24225, n17285);
xor_4  g21879(new_n11941, new_n11906, n17320);
xor_4  g21880(new_n2829, new_n2784, n17337);
xor_4  g21881(new_n22538, new_n22527, n17344);
xnor_4 g21882(new_n22546, new_n22509, n17359);
xor_4  g21883(new_n14564, new_n13666, n17387);
xor_4  g21884(new_n5101_1, new_n5100, n17391);
xnor_4 g21885(new_n19630, new_n19608_1, n17392);
xor_4  g21886(new_n22816, new_n22790, n17421);
xor_4  g21887(new_n12459, new_n16004, n17432);
xnor_4 g21888(new_n21680_1, new_n21660, n17436);
xor_4  g21889(new_n7192, new_n4719, n17440);
xor_4  g21890(new_n8607, new_n6167, n17450);
and_5  g21891(new_n19384, new_n7417, new_n24240);
nor_5  g21892(new_n7417, new_n7371, new_n24241);
and_5  g21893(new_n7417, new_n7371, new_n24242);
nor_5  g21894(new_n7506, new_n24242, new_n24243);
nor_5  g21895(new_n24243, new_n24241, new_n24244);
or_5   g21896(new_n24244, new_n24240, new_n24245);
nor_5  g21897(new_n19384, new_n7417, new_n24246);
or_5   g21898(new_n24246, new_n24243, new_n24247);
and_5  g21899(new_n24247, new_n24245, n17461);
xor_4  g21900(new_n23779, new_n23778, n17466);
xor_4  g21901(new_n13830, new_n13786, n17493);
xor_4  g21902(new_n22192, new_n22189, n17500);
xnor_4 g21903(new_n23097, new_n23094, n17524);
xnor_4 g21904(new_n5817, new_n5770, n17529);
xor_4  g21905(new_n15388, new_n5849, new_n24254);
xor_4  g21906(new_n24254, new_n15391, n17557);
xnor_4 g21907(new_n17051, new_n17013, n17583);
xnor_4 g21908(new_n14575_1, new_n14549, n17592);
xnor_4 g21909(new_n8519_1, new_n8504, n17638);
xnor_4 g21910(new_n20458, new_n20441_1, n17687);
xnor_4 g21911(new_n14146, new_n14107_1, n17721);
xor_4  g21912(new_n22383, new_n22362, n17735);
nor_5  g21913(new_n21915_1, new_n10338, new_n24262);
and_5  g21914(new_n24262, new_n21760, new_n24263);
and_5  g21915(new_n21915_1, new_n10338, new_n24264);
and_5  g21916(new_n24264, new_n21759, new_n24265);
nor_5  g21917(new_n24265, new_n24263, new_n24266);
nand_5 g21918(new_n24266, new_n21844, new_n24267);
or_5   g21919(new_n24266, new_n21844, new_n24268);
nor_5  g21920(new_n21763, new_n21751, new_n24269);
and_5  g21921(new_n21777, new_n21764, new_n24270);
nor_5  g21922(new_n24270, new_n24269, new_n24271);
and_5  g21923(new_n24271, new_n24268, new_n24272);
nor_5  g21924(new_n24272, new_n24263, new_n24273);
and_5  g21925(new_n24273, new_n24267, n17738);
xor_4  g21926(new_n15790, new_n15787, n17746);
xnor_4 g21927(new_n23558, new_n23554, n17749);
xnor_4 g21928(new_n19250, new_n19228_1, n17820);
xnor_4 g21929(new_n14572, new_n14555, n17855);
nor_5  g21930(new_n4916, new_n22847, new_n24279);
and_5  g21931(new_n4974, new_n24279, new_n24280);
nor_5  g21932(new_n4974, new_n22849, new_n24281);
or_5   g21933(new_n24281, new_n24280, new_n24282);
nand_5 g21934(new_n4975, new_n4815, new_n24283);
nand_5 g21935(new_n5050, new_n4976, new_n24284);
and_5  g21936(new_n24284, new_n24283, new_n24285);
nor_5  g21937(new_n24285, new_n24282, new_n24286);
nor_5  g21938(new_n24286, new_n24280, n17877);
xnor_4 g21939(new_n15996, new_n15994, n17889);
and_5  g21940(new_n23444, new_n23431, new_n24289_1);
or_5   g21941(new_n23453, new_n24289_1, new_n24290);
nor_5  g21942(new_n23444, new_n23431, new_n24291);
or_5   g21943(new_n23452, new_n24291, new_n24292);
and_5  g21944(new_n24292, new_n24290, n17912);
xor_4  g21945(new_n22805, new_n22802, n17927);
xnor_4 g21946(new_n22891_1, new_n22865, n17931);
xnor_4 g21947(new_n8027_1, new_n8026, n17948);
xor_4  g21948(new_n16212, new_n16209, n17956);
or_5   g21949(new_n13148, new_n12915, new_n24298);
not_10 g21950(new_n13063, new_n24299);
nor_5  g21951(new_n24299, new_n12915, new_n24300);
or_5   g21952(new_n13147, new_n24300, new_n24301);
and_5  g21953(new_n24301, new_n24298, n17963);
and_5  g21954(new_n3408, n6659, new_n24303);
not_10 g21955(new_n24303, new_n24304);
nor_5  g21956(new_n18031, new_n18016, new_n24305);
not_10 g21957(new_n24305, new_n24306);
and_5  g21958(new_n24306, new_n24304, new_n24307_1);
not_10 g21959(new_n24307_1, new_n24308);
nor_5  g21960(new_n24308, new_n13448, new_n24309);
nor_5  g21961(new_n24307_1, new_n13452, new_n24310);
xor_4  g21962(new_n24307_1, new_n13452, new_n24311);
nor_5  g21963(new_n18032, new_n13457_1, new_n24312);
and_5  g21964(new_n18053, new_n18033, new_n24313);
nor_5  g21965(new_n24313, new_n24312, new_n24314);
and_5  g21966(new_n24314, new_n24311, new_n24315);
nor_5  g21967(new_n24315, new_n24310, new_n24316);
or_5   g21968(new_n24316, new_n24309, new_n24317);
and_5  g21969(new_n24308, new_n13448, new_n24318);
or_5   g21970(new_n24318, new_n24315, new_n24319_1);
and_5  g21971(new_n24319_1, new_n24317, n17976);
xor_4  g21972(new_n7213, new_n7168, n17998);
xnor_4 g21973(new_n14989_1, new_n2813, n18025);
xnor_4 g21974(new_n21310, new_n21308, n18043);
xnor_4 g21975(new_n22730, new_n22727, n18045);
xnor_4 g21976(new_n3926, new_n3916, n18059);
xnor_4 g21977(new_n20984, new_n20940, n18061);
xnor_4 g21978(new_n3392, new_n3325, n18071);
xnor_4 g21979(new_n10256, new_n10183, n18143);
xnor_4 g21980(new_n22194, new_n22187, n18152);
xor_4  g21981(new_n7699, new_n7689, n18193);
xnor_4 g21982(new_n11987, new_n11978, new_n24331);
xor_4  g21983(new_n24331, new_n12000_1, n18232);
xor_4  g21984(new_n17423, new_n17400, n18238);
xnor_4 g21985(new_n19063, new_n19060, n18241);
xnor_4 g21986(new_n21676, new_n21667, n18254);
xor_4  g21987(new_n22380, new_n22364, n18288);
xnor_4 g21988(new_n12540_1, new_n12492, n18301);
xor_4  g21989(new_n22718, new_n22704, n18304);
xnor_4 g21990(new_n13837, new_n13780, n18310);
xnor_4 g21991(new_n6704, new_n6703, n18311);
xnor_4 g21992(new_n18192, new_n18173, n18323);
xnor_4 g21993(new_n5474, new_n5437, n18332);
xor_4  g21994(new_n22902, new_n22901, n18343);
xnor_4 g21995(new_n19964, new_n19961, n18350);
xnor_4 g21996(new_n18665, new_n18663, n18362);
xnor_4 g21997(new_n5046_1, new_n4987, n18377);
xor_4  g21998(new_n4108, new_n4083, n18405);
xor_4  g21999(new_n17274, new_n17261, n18414);
xor_4  g22000(new_n15076, new_n15065, n18418);
xnor_4 g22001(new_n8334, new_n8288_1, n18437);
xnor_4 g22002(new_n20790, new_n20743, n18439);
xnor_4 g22003(new_n11444, new_n11443, n18445);
xor_4  g22004(new_n6985_1, new_n6937, n18467);
xor_4  g22005(new_n19083, new_n19022, n18482);
xnor_4 g22006(new_n19418, new_n19397, n18509);
xnor_4 g22007(new_n14378, new_n9255, n18513);
xor_4  g22008(new_n15605, new_n15603, n18515);
xor_4  g22009(new_n16487, new_n16467, n18572);
and_5  g22010(new_n24126, new_n24110, new_n24359);
or_5   g22011(new_n24359, new_n24002_1, new_n24360);
nor_5  g22012(new_n24126, new_n24110, new_n24361);
or_5   g22013(new_n24361, new_n24001, new_n24362);
and_5  g22014(new_n24362, new_n24360, n18574);
xnor_4 g22015(new_n21830, new_n21827, n18576);
xnor_4 g22016(new_n23235, new_n23227, n18582);
xnor_4 g22017(new_n20552, new_n20539, n18583);
xnor_4 g22018(new_n20969, new_n20968, n18610);
xor_4  g22019(new_n22744, new_n22741, n18635);
xor_4  g22020(new_n6770, new_n6769, n18653);
xnor_4 g22021(new_n3720, new_n3666, n18679);
xnor_4 g22022(new_n21098, new_n21090, n18693);
xnor_4 g22023(new_n3067_1, new_n3028, n18708);
xnor_4 g22024(new_n23600, new_n22074, new_n24373_1);
xor_4  g22025(new_n24373_1, new_n23605, n18721);
xnor_4 g22026(new_n19256, new_n19216, n18725);
xnor_4 g22027(new_n21482, new_n21455, n18751);
xnor_4 g22028(new_n17045, new_n17025, n18780);
xnor_4 g22029(new_n20197, new_n20149_1, n18782);
not_10 g22030(new_n7644, new_n24379);
and_5  g22031(new_n24379, new_n7558_1, new_n24380);
or_5   g22032(new_n7726, new_n24380, new_n24381);
nor_5  g22033(new_n24379, new_n7558_1, new_n24382);
or_5   g22034(new_n7725, new_n24382, new_n24383);
and_5  g22035(new_n24383, new_n24381, n18802);
xor_4  g22036(new_n11156, new_n11155, n18830);
xor_4  g22037(new_n13235, new_n13229, n18831);
xnor_4 g22038(new_n12293, new_n12284, n18843);
xnor_4 g22039(new_n3063, new_n3039, n18858);
xnor_4 g22040(new_n10242, new_n10219, n18859);
xnor_4 g22041(new_n17798, new_n17746_1, n18864);
xnor_4 g22042(new_n4608, new_n4532, n18865);
xnor_4 g22043(new_n22118, new_n22117, n18886);
xnor_4 g22044(new_n17041, new_n17039, n18887);
xnor_4 g22045(new_n9081, new_n9037, n18919);
xnor_4 g22046(new_n12755, new_n12743, n18940);
xor_4  g22047(new_n23728, new_n23727, n18945);
xnor_4 g22048(new_n23420, new_n23406, n18970);
xor_4  g22049(new_n24092_1, new_n12490, new_n24398);
xor_4  g22050(new_n24398, new_n17492, n18977);
xnor_4 g22051(new_n15708, new_n15698, n18982);
xor_4  g22052(new_n21560, new_n21559, n18999);
xnor_4 g22053(new_n5823, new_n5752_1, n19044);
xor_4  g22054(new_n15393, new_n15386, n19125);
xnor_4 g22055(new_n5821, new_n5758, n19141);
xor_4  g22056(new_n17906, new_n14516, new_n24405);
not_10 g22057(new_n24405, new_n24406_1);
nor_5  g22058(new_n17910, new_n14523, new_n24407);
xor_4  g22059(new_n17910, new_n14523, new_n24408);
not_10 g22060(new_n24408, new_n24409);
and_5  g22061(new_n17913, new_n14527, new_n24410);
nor_5  g22062(new_n19293, new_n19269, new_n24411);
nor_5  g22063(new_n24411, new_n24410, new_n24412);
nor_5  g22064(new_n24412, new_n24409, new_n24413);
nor_5  g22065(new_n24413, new_n24407, new_n24414);
xnor_4 g22066(new_n24414, new_n24406_1, n19164);
xnor_4 g22067(new_n8527, new_n8526_1, n19174);
xnor_4 g22068(new_n21736, new_n21733, n19176);
xor_4  g22069(new_n22720, new_n22700, n19202);
xnor_4 g22070(new_n20880, new_n20871, n19220);
xor_4  g22071(new_n8044, new_n7989, n19221);
xnor_4 g22072(new_n11578, new_n11576, n19223);
xor_4  g22073(new_n17779, new_n17778, n19224);
xnor_4 g22074(new_n16152, new_n16140, n19233);
xnor_4 g22075(new_n13218, new_n13177, n19244);
xnor_4 g22076(new_n9083, new_n9031, n19314);
xnor_4 g22077(new_n11058, new_n11056_1, n19315);
xor_4  g22078(new_n13824, new_n13792, n19323);
xor_4  g22079(new_n22536, new_n22531, n19333);
and_5  g22080(new_n17902, new_n17899, new_n24429);
or_5   g22081(new_n24429, new_n10170, new_n24430);
and_5  g22082(new_n17903, new_n10176, new_n24431_1);
nor_5  g22083(new_n17926, new_n17905, new_n24432);
nor_5  g22084(new_n24432, new_n24431_1, new_n24433);
xor_4  g22085(new_n24429, new_n10170, new_n24434);
nand_5 g22086(new_n24434, new_n24433, new_n24435);
and_5  g22087(new_n24435, new_n24430, n19348);
xnor_4 g22088(new_n17441, new_n17374, n19354);
xnor_4 g22089(new_n11385, new_n11353, n19367);
xor_4  g22090(new_n19796, new_n19762, n19385);
xor_4  g22091(new_n17560, new_n17510, new_n24440);
xor_4  g22092(new_n24440, new_n17594, n19389);
xnor_4 g22093(new_n16915, new_n16876, n19401);
xor_4  g22094(new_n23007_1, new_n22999, n19414);
xnor_4 g22095(new_n19984, new_n18475, n19424);
xnor_4 g22096(new_n22124_1, new_n22103, n19450);
not_10 g22097(new_n14444, new_n24446);
and_5  g22098(new_n24429, new_n24446, new_n24447);
xor_4  g22099(new_n24429, new_n14444, new_n24448);
and_5  g22100(new_n17903, new_n14514, new_n24449);
xor_4  g22101(new_n17903, new_n14514, new_n24450);
and_5  g22102(new_n17906, new_n14516, new_n24451);
nor_5  g22103(new_n24414, new_n24406_1, new_n24452);
nor_5  g22104(new_n24452, new_n24451, new_n24453);
not_10 g22105(new_n24453, new_n24454);
and_5  g22106(new_n24454, new_n24450, new_n24455);
nor_5  g22107(new_n24455, new_n24449, new_n24456);
nor_5  g22108(new_n24456, new_n24448, new_n24457);
or_5   g22109(new_n24457, new_n24447, n19458);
xor_4  g22110(new_n15792, new_n15784, n19467);
xnor_4 g22111(new_n8336, new_n8283, n19496);
xor_4  g22112(new_n15752, new_n15743_1, n19523);
xnor_4 g22113(new_n4596, new_n4556, n19570);
xnor_4 g22114(new_n12421, new_n12410, n19602);
xnor_4 g22115(new_n12804, new_n12799, n19617);
xnor_4 g22116(new_n14144, new_n14110, n19623);
xor_4  g22117(new_n23046, new_n23045, n19641);
xnor_4 g22118(new_n22820, new_n22787_1, n19648);
xor_4  g22119(new_n16485, new_n16471, n19664);
xnor_4 g22120(new_n20633, new_n20617, n19736);
or_5   g22121(new_n23009_1, new_n22995, new_n24470);
nor_5  g22122(new_n22995, new_n3399, new_n24471);
or_5   g22123(new_n23008, new_n24471, new_n24472_1);
and_5  g22124(new_n24472_1, new_n24470, n19749);
xor_4  g22125(new_n15463, new_n15446, n19756);
xor_4  g22126(new_n12419, new_n12417, n19767);
xor_4  g22127(new_n3317, new_n3315, new_n24476_1);
xor_4  g22128(new_n24476_1, new_n3394, n19780);
xnor_4 g22129(new_n23624_1, new_n23621, n19792);
xnor_4 g22130(new_n21298_1, new_n21283, n19798);
xor_4  g22131(new_n17143, new_n17140, n19873);
or_5   g22132(new_n19123, new_n19097, new_n24481);
nor_5  g22133(new_n19107_1, new_n19097, new_n24482);
or_5   g22134(new_n19122, new_n24482, new_n24483_1);
and_5  g22135(new_n24483_1, new_n24481, n19909);
xor_4  g22136(new_n20631, new_n20621, n19916);
xnor_4 g22137(new_n21302_1, new_n21275, n19923);
xor_4  g22138(new_n19639, new_n19599, n19930);
xnor_4 g22139(new_n6455, new_n6343, n19968);
xnor_4 g22140(new_n20179_1, new_n20167, n19988);
not_10 g22141(new_n21376, new_n24490);
nor_5  g22142(new_n22150_1, new_n24490, new_n24491);
nor_5  g22143(new_n21376, new_n10389, new_n24492);
nor_5  g22144(new_n21381, new_n21378, new_n24493);
nor_5  g22145(new_n24493, new_n24492, new_n24494);
or_5   g22146(new_n24494, new_n24491, new_n24495);
and_5  g22147(new_n22150_1, new_n24490, new_n24496);
or_5   g22148(new_n24496, new_n24493, new_n24497);
and_5  g22149(new_n24497, new_n24495, n20004);
xnor_4 g22150(new_n21478, new_n21461, n20017);
xor_4  g22151(new_n19077, new_n19032, n20033);
xnor_4 g22152(new_n14343, new_n14341, n20061);
xnor_4 g22153(new_n18615, new_n18612, n20069);
and_5  g22154(new_n14946, new_n14937, new_n24503);
nor_5  g22155(new_n15017, new_n14948, new_n24504);
or_5   g22156(new_n24504, new_n24503, n20086);
xnor_4 g22157(new_n20061_1, new_n20057, n20096);
xor_4  g22158(new_n13815, new_n13806, n20103);
xor_4  g22159(new_n11945, new_n11899, n20126);
xnor_4 g22160(new_n21909, new_n21876, n20149);
xor_4  g22161(new_n12307, new_n12259, n20187);
xnor_4 g22162(new_n18012, new_n17979, n20279);
nand_5 g22163(new_n23219, new_n23212, new_n24512_1);
and_5  g22164(new_n23223, new_n24512_1, new_n24513);
not_10 g22165(new_n23219, new_n24514);
nand_5 g22166(new_n23238_1, new_n24514, new_n24515);
or_5   g22167(new_n23238_1, new_n18166, new_n24516);
and_5  g22168(new_n24516, new_n24515, new_n24517);
and_5  g22169(new_n24517, new_n24513, n20287);
xnor_4 g22170(new_n21132, new_n21129, n20301);
or_5   g22171(new_n8342, new_n8268, new_n24520);
and_5  g22172(new_n24520, new_n8163, n20330);
xor_4  g22173(new_n12301, new_n12267, n20333);
and_5  g22174(new_n10648, new_n10510, new_n24523);
and_5  g22175(new_n10718, new_n24523, new_n24524);
or_5   g22176(new_n10648, new_n10510, new_n24525);
nor_5  g22177(new_n10718, new_n24525, new_n24526);
or_5   g22178(new_n24526, new_n24524, n20355);
xor_4  g22179(new_n8565, new_n5224, n20366);
xor_4  g22180(new_n19833, new_n19827, n20388);
xnor_4 g22181(new_n22889, new_n22868, n20402);
xnor_4 g22182(new_n15977, new_n15951, n20403);
xor_4  g22183(new_n3048, new_n3046, n20424);
xnor_4 g22184(new_n20974, new_n20960, n20436);
xor_4  g22185(new_n8321_1, new_n8320_1, n20441);
xnor_4 g22186(new_n7724, new_n7650, n20445);
xnor_4 g22187(new_n5048, new_n4981, n20450);
xor_4  g22188(new_n17056, new_n6702, n20490);
xor_4  g22189(new_n20878, new_n20875, n20495);
and_5  g22190(new_n16001, new_n16000, new_n24539);
and_5  g22191(new_n24539, new_n15998, new_n24540);
or_5   g22192(new_n16001, new_n16000, new_n24541);
nor_5  g22193(new_n24541, new_n15998, new_n24542);
or_5   g22194(new_n24542, new_n24540, n20515);
or_5   g22195(new_n23626, new_n23617, new_n24544);
and_5  g22196(new_n24544, new_n23613, n20533);
xnor_4 g22197(new_n18477, new_n18470, n20582);
xor_4  g22198(new_n20340, new_n20312, n20590);
xnor_4 g22199(new_n3376, new_n3374, n20602);
xnor_4 g22200(new_n17037_1, new_n17035_1, n20609);
xnor_4 g22201(new_n6619, new_n6610, n20623);
xor_4  g22202(new_n21314, new_n21255, n20629);
xnor_4 g22203(new_n14339, new_n14329, n20661);
xnor_4 g22204(new_n8611, new_n8609, n20673);
xnor_4 g22205(new_n21306, new_n21266, n20678);
or_5   g22206(new_n15433, new_n12188, new_n24555);
nand_5 g22207(new_n15472, new_n24555, new_n24556);
and_5  g22208(new_n15433, new_n12188, new_n24557);
nor_5  g22209(new_n24557, new_n15429, new_n24558_1);
and_5  g22210(new_n24558_1, new_n24556, n20680);
xnor_4 g22211(new_n6429, new_n4156, n20685);
xor_4  g22212(new_n24307_1, new_n13448, new_n24561);
xor_4  g22213(new_n24561, new_n24316, n20691);
xnor_4 g22214(new_n16483, new_n16475, n20696);
xnor_4 g22215(new_n23382, new_n23373, n20704);
xor_4  g22216(new_n22373, new_n22372, n20705);
xor_4  g22217(new_n10252, new_n10189, n20709);
xnor_4 g22218(new_n15351, new_n15314, n20713);
xnor_4 g22219(new_n8785, new_n8784, n20722);
nor_5  g22220(new_n23911, new_n20238, new_n24569);
and_5  g22221(new_n20238, new_n20226, new_n24570);
nor_5  g22222(new_n20238, new_n20226, new_n24571);
nor_5  g22223(new_n20252, new_n24571, new_n24572);
nor_5  g22224(new_n24572, new_n24570, new_n24573);
or_5   g22225(new_n24573, new_n24569, new_n24574);
and_5  g22226(new_n23911, new_n20238, new_n24575);
or_5   g22227(new_n24575, new_n24572, new_n24576_1);
and_5  g22228(new_n24576_1, new_n24574, n20723);
xor_4  g22229(new_n23213, new_n18166, new_n24578);
xor_4  g22230(new_n24578, new_n23238_1, n20748);
xor_4  g22231(new_n5466, new_n5456, n20761);
xnor_4 g22232(new_n20982, new_n20944, n20774);
xnor_4 g22233(new_n24456, new_n24448, n20788);
nor_5  g22234(new_n23757, new_n22739, new_n24583);
or_5   g22235(new_n24583, new_n23869, new_n24584);
and_5  g22236(new_n23757, new_n22739, new_n24585);
or_5   g22237(new_n24585, new_n23868, new_n24586);
and_5  g22238(new_n24586, new_n24584, n20795);
xor_4  g22239(new_n21018, new_n21005, new_n24588);
nand_5 g22240(new_n21025, new_n21005, new_n24589);
nand_5 g22241(new_n24589, new_n21022, new_n24590);
and_5  g22242(new_n24590, new_n21026, new_n24591);
xor_4  g22243(new_n24591, new_n24588, n20803);
xor_4  g22244(new_n24285, new_n24282, n20869);
xnor_4 g22245(new_n23561, new_n23551, n20879);
xnor_4 g22246(new_n6441, new_n6409, n20915);
xor_4  g22247(n19282, n2160, new_n24596);
or_5   g22248(n12657, new_n17112, new_n24597);
or_5   g22249(new_n22392, new_n22389, new_n24598);
and_5  g22250(new_n24598, new_n24597, new_n24599);
xor_4  g22251(new_n24599, new_n24596, new_n24600);
nor_5  g22252(new_n24600, new_n22256, new_n24601);
nor_5  g22253(new_n22393, new_n20582_1, new_n24602_1);
not_10 g22254(new_n24602_1, new_n24603);
not_10 g22255(new_n22399, new_n24604_1);
and_5  g22256(new_n24604_1, new_n22394, new_n24605);
not_10 g22257(new_n24605, new_n24606);
and_5  g22258(new_n24606, new_n24603, new_n24607);
xor_4  g22259(new_n24600, new_n22256, new_n24608);
not_10 g22260(new_n24608, new_n24609);
nor_5  g22261(new_n24609, new_n24607, new_n24610);
nor_5  g22262(new_n24610, new_n24601, new_n24611);
nand_5 g22263(new_n7295, n2160, new_n24612);
or_5   g22264(new_n24599, new_n24596, new_n24613);
and_5  g22265(new_n24613, new_n24612, new_n24614);
and_5  g22266(new_n24614, new_n23446, new_n24615);
not_10 g22267(new_n24615, new_n24616);
nor_5  g22268(new_n24616, new_n24611, new_n24617);
and_5  g22269(new_n24617, new_n23444, new_n24618_1);
nor_5  g22270(new_n24614, new_n23446, new_n24619);
and_5  g22271(new_n24619, new_n24611, new_n24620_1);
not_10 g22272(new_n24620_1, new_n24621);
nor_5  g22273(new_n24621, new_n23444, new_n24622);
or_5   g22274(new_n24622, new_n24618_1, n20935);
xor_4  g22275(new_n22810, new_n22796, n20936);
xnor_4 g22276(new_n17471, new_n17469, n21008);
xor_4  g22277(new_n20193, new_n20152, n21017);
nand_5 g22278(new_n23977, new_n22219, new_n24627);
or_5   g22279(new_n23977, new_n22219, new_n24628);
and_5  g22280(new_n23981, new_n24628, new_n24629_1);
nor_5  g22281(new_n24629_1, new_n23976, new_n24630);
and_5  g22282(new_n24630, new_n24627, n21034);
xor_4  g22283(new_n22972, new_n22971, n21046);
xnor_4 g22284(new_n8722, new_n8698, n21062);
xor_4  g22285(new_n23711, new_n23702, new_n24634);
xor_4  g22286(new_n24634, new_n23613, n21093);
xor_4  g22287(new_n9969, new_n8020, n21094);
xnor_4 g22288(new_n15228, new_n15198, n21123);
xor_4  g22289(new_n19527, new_n18687, n21154);
xnor_4 g22290(new_n16124, new_n16098_1, n21157);
xnor_4 g22291(new_n21901, new_n21892, n21168);
xor_4  g22292(new_n7467, new_n7465, n21173);
xnor_4 g22293(new_n4592, new_n4566, n21176);
xnor_4 g22294(new_n14872, new_n14866, n21182);
or_5   g22295(new_n22781, new_n21926, new_n24644);
nand_5 g22296(new_n22822, new_n21926, new_n24645);
and_5  g22297(new_n24645, new_n24644, new_n24646);
or_5   g22298(new_n22822, new_n21937, new_n24647);
and_5  g22299(new_n24647, new_n22784, new_n24648);
and_5  g22300(new_n24648, new_n24646, n21193);
xnor_4 g22301(new_n9713, new_n9712, n21203);
xor_4  g22302(new_n17034, new_n2547_1, n21225);
xnor_4 g22303(new_n20566, new_n20514, n21238);
xnor_4 g22304(new_n14345_1, new_n14323_1, n21254);
xnor_4 g22305(new_n20786, new_n20751, n21298);
xor_4  g22306(new_n20545, new_n9616_1, n21302);
xnor_4 g22307(new_n20629_1, new_n20625, n21349);
xnor_4 g22308(new_n16642, new_n16640_1, n21365);
xnor_4 g22309(new_n15754, new_n15740, n21367);
xor_4  g22310(new_n12173, new_n12136, n21396);
xor_4  g22311(new_n7721_1, new_n7655, n21399);
xor_4  g22312(new_n3403, new_n3397, n21404);
xnor_4 g22313(new_n8613, new_n8602, n21446);
xnor_4 g22314(new_n11998, new_n11990, n21472);
xor_4  g22315(new_n7496, new_n7435, n21525);
xnor_4 g22316(new_n17847, new_n17820_1, n21549);
xnor_4 g22317(new_n20454, new_n20451, n21615);
nand_5 g22318(new_n24514, new_n13931, new_n24667);
xor_4  g22319(new_n24514, new_n7975, new_n24668);
or_5   g22320(new_n18166, new_n13931, new_n24669);
nand_5 g22321(new_n18198, new_n18167, new_n24670);
and_5  g22322(new_n24670, new_n24669, new_n24671);
or_5   g22323(new_n24671, new_n24668, new_n24672);
and_5  g22324(new_n24672, new_n24667, n21628);
nand_5 g22325(new_n22437, new_n21934_1, new_n24674);
xor_4  g22326(new_n22437, new_n21933, new_n24675);
or_5   g22327(new_n22440, new_n21934_1, new_n24676);
or_5   g22328(new_n23835, new_n23832, new_n24677);
and_5  g22329(new_n24677, new_n24676, new_n24678);
or_5   g22330(new_n24678, new_n24675, new_n24679);
and_5  g22331(new_n24679, new_n24674, n21637);
xnor_4 g22332(new_n22375, new_n22368, n21645);
xor_4  g22333(new_n12453, new_n6612_1, n21665);
xnor_4 g22334(new_n15470_1, new_n15438_1, n21680);
xnor_4 g22335(new_n22897_1, new_n22856, n21685);
xnor_4 g22336(new_n19252, new_n19224_1, n21717);
xnor_4 g22337(new_n17457, new_n17452, n21719);
xnor_4 g22338(new_n19243, new_n19240, n21750);
xnor_4 g22339(new_n22641, new_n22639, n21765);
xnor_4 g22340(new_n24609, new_n24607, n21800);
xor_4  g22341(new_n4289, new_n4288, new_n24690);
xor_4  g22342(new_n24690, new_n4293, n21820);
xor_4  g22343(new_n20184, new_n20161, n21874);
xor_4  g22344(new_n13817, new_n13802, n21943);
xnor_4 g22345(new_n16646, new_n16622, n21960);
xor_4  g22346(new_n7199, new_n7198, n21976);
xnor_4 g22347(new_n11588, new_n11556, n21986);
xnor_4 g22348(new_n11387, new_n11349, n22016);
xnor_4 g22349(new_n19246, new_n19236, n22027);
xnor_4 g22350(new_n13607, new_n13597, n22050);
xnor_4 g22351(new_n4158, new_n4156, n22063);
xnor_4 g22352(new_n21899, new_n21896, n22076);
or_5   g22353(new_n21009, new_n14300, new_n24702);
nand_5 g22354(new_n21369, new_n21345, new_n24703);
and_5  g22355(new_n24703, new_n24702, n22090);
xnor_4 g22356(new_n23418, new_n23409, n22107);
xnor_4 g22357(new_n18370, new_n18342, n22113);
nor_5  g22358(new_n14299, new_n14237, new_n24707);
or_5   g22359(new_n14353_1, new_n24707, new_n24708);
and_5  g22360(new_n14299, new_n14237, new_n24709);
or_5   g22361(new_n14352, new_n24709, new_n24710);
and_5  g22362(new_n24710, new_n24708, n22124);
nand_5 g22363(new_n24080, new_n20046, new_n24712);
nand_5 g22364(new_n24085_1, new_n24081, new_n24713);
and_5  g22365(new_n24713, new_n24712, n22126);
nor_5  g22366(new_n24620_1, new_n24617, new_n24715_1);
xor_4  g22367(new_n24715_1, new_n23444, n22130);
xor_4  g22368(new_n18560, new_n18559, n22144);
xor_4  g22369(new_n23825, new_n23821, n22150);
xnor_4 g22370(new_n20384, new_n20376, n22157);
xnor_4 g22371(new_n24412, new_n24409, n22213);
xnor_4 g22372(new_n10697, new_n10696, n22283);
xor_4  g22373(new_n21047, new_n21046_1, n22311);
xnor_4 g22374(new_n9085, new_n9025, n22317);
xor_4  g22375(new_n18120, new_n18097, n22341);
not_10 g22376(new_n18868, new_n24725);
not_10 g22377(new_n7228, new_n24726);
and_5  g22378(new_n7241, new_n24726, new_n24727);
and_5  g22379(new_n24727, new_n7222, new_n24728);
nor_5  g22380(new_n7241, new_n24726, new_n24729);
not_10 g22381(new_n24729, new_n24730);
nor_5  g22382(new_n24730, new_n7222, new_n24731);
nor_5  g22383(new_n24731, new_n24728, new_n24732_1);
xor_4  g22384(new_n24732_1, new_n24725, n22353);
xor_4  g22385(new_n18117, new_n18102, n22444);
xor_4  g22386(new_n10439, new_n10438, n22467);
xor_4  g22387(new_n9064, new_n9062, n22484);
xor_4  g22388(new_n4604, new_n4539, n22489);
xnor_4 g22389(new_n8535_1, new_n8483, n22494);
xnor_4 g22390(new_n10703, new_n10677, n22533);
xor_4  g22391(new_n23379, new_n23378, n22584);
or_5   g22392(new_n18566, new_n18541, new_n24741);
and_5  g22393(new_n24741, new_n18502, n22589);
xor_4  g22394(new_n24453, new_n24450, n22620);
xor_4  g22395(new_n8608_1, new_n8606, n22623);
xnor_4 g22396(new_n17589, new_n17571, n22697);
xnor_4 g22397(new_n9075, new_n9054, n22714);
xnor_4 g22398(new_n12313, new_n12250, n22761);
xnor_4 g22399(new_n19710, new_n19690, n22779);
xnor_4 g22400(new_n23390, new_n23358, n22787);
xor_4  g22401(new_n2542, new_n2508, n22819);
xor_4  g22402(new_n9439, new_n4580, n22858);
xor_4  g22403(new_n21966, new_n11965_1, new_n24752);
xor_4  g22404(new_n24752, new_n23888_1, n22870);
xor_4  g22405(new_n9935, new_n9917_1, n22891);
xor_4  g22406(new_n20333_1, new_n20321, n22897);
xnor_4 g22407(new_n10463, new_n10396, n22903);
xnor_4 g22408(new_n14886, new_n14842, n22907);
xor_4  g22409(new_n7206, new_n7204, n22910);
xnor_4 g22410(new_n12779, new_n12773, n22914);
xor_4  g22411(new_n5829, new_n5795, n22939);
xnor_4 g22412(new_n19838, new_n18744, new_n24761);
xor_4  g22413(new_n24761, new_n19836, n22998);
xnor_4 g22414(new_n9071, new_n9070, n23006);
xnor_4 g22415(new_n13237, new_n13227, n23007);
xnor_4 g22416(new_n18760, new_n18757, n23009);
xnor_4 g22417(new_n17439, new_n17380, n23014);
xor_4  g22418(new_n24678, new_n24675, n23047);
xnor_4 g22419(new_n18190, new_n18176, n23058);
and_5  g22420(new_n19265, new_n19260, n23066);
and_5  g22421(new_n19151, new_n10509, new_n24770);
nor_5  g22422(new_n24770, new_n19153, new_n24771);
xor_4  g22423(new_n24771, new_n19148, n23067);
xor_4  g22424(new_n16636, new_n16630_1, n23238);
xnor_4 g22425(new_n17924, new_n17909, n23247);
xor_4  g22426(new_n15598_1, new_n15592, n23248);
xor_4  g22427(new_n18003, new_n17989, n23270);
xnor_4 g22428(new_n23451, new_n23448, n23289);
xnor_4 g22429(new_n5476, new_n5432, n23305);
xnor_4 g22430(new_n21674_1, new_n21671, n23341);
xor_4  g22431(new_n9615, new_n4953, n23342);
and_5  g22432(new_n22014, new_n24379, new_n24781);
or_5   g22433(new_n22039, new_n24781, new_n24782);
nor_5  g22434(new_n22014, new_n24379, new_n24783);
or_5   g22435(new_n22038, new_n24783, new_n24784_1);
and_5  g22436(new_n24784_1, new_n24782, n23355);
xnor_4 g22437(new_n19935, new_n19932, n23371);
xnor_4 g22438(new_n15983, new_n15940, n23401);
xor_4  g22439(new_n13604, new_n13602_1, n23414);
xnor_4 g22440(new_n18009, new_n17983, n23429);
or_5   g22441(new_n22277, new_n22269, new_n24790);
and_5  g22442(new_n22272, new_n22270_1, new_n24791);
or_5   g22443(new_n24791, new_n22276, new_n24792);
and_5  g22444(new_n24792, new_n24790, n23433);
xor_4  g22445(new_n19069, new_n19053, n23434);
and_5  g22446(new_n24080, new_n22407, new_n24795);
or_5   g22447(new_n24795, new_n24100, new_n24796);
nor_5  g22448(new_n24080, new_n22407, new_n24797);
or_5   g22449(new_n24797, new_n24099, new_n24798);
and_5  g22450(new_n24798, new_n24796, n23450);
xor_4  g22451(new_n17435, new_n17384, n23471);
xor_4  g22452(new_n21684, new_n21653, n23480);
xor_4  g22453(new_n18402, new_n18397, n23546);
xnor_4 g22454(new_n21296, new_n21287_1, n23550);
xor_4  g22455(new_n7484, new_n7453, n23585);
xor_4  g22456(new_n20331, new_n20324, n23588);
xor_4  g22457(new_n21557, new_n21556, n23619);
xor_4  g22458(new_n3059, new_n3045, n23624);
xnor_4 g22459(new_n12159, new_n12151, n23628);
xor_4  g22460(new_n22540, new_n22523, n23637);
xnor_4 g22461(new_n23167, new_n23163, n23663);
xor_4  g22462(new_n12161_1, new_n12148, n23669);
xnor_4 g22463(new_n13493, new_n13460_1, n23684);
xnor_4 g22464(new_n19623_1, new_n19615, n23690);
xnor_4 g22465(new_n22895, new_n22859, n23714);
not_10 g22466(new_n24138, new_n24815);
and_5  g22467(new_n24815, new_n24133_1, n23719);
xnor_4 g22468(new_n21982, new_n21979, n23748);
xor_4  g22469(new_n11151, new_n7244, n23856);
xor_4  g22470(new_n7481, new_n7479, n23883);
xor_4  g22471(new_n14867, new_n5866, new_n24820);
xor_4  g22472(new_n24820, new_n14869, n23888);
xnor_4 g22473(new_n3382, new_n3354, n23899);
xor_4  g22474(new_n15390, new_n9706, n23903);
xnor_4 g22475(new_n13216, new_n13180, n23924);
xor_4  g22476(new_n17102, new_n17100, n23935);
xnor_4 g22477(new_n13489, new_n13472, n23942);
xnor_4 g22478(new_n18228, new_n18218, n23954);
xor_4  g22479(new_n19342, new_n19320, n23958);
xor_4  g22480(new_n23031, new_n23030, n23986);
xor_4  g22481(new_n17473, new_n17467, n24002);
xnor_4 g22482(new_n13374, new_n13367_1, n24039);
xor_4  g22483(new_n24065, new_n24064, n24052);
xnor_4 g22484(new_n20976, new_n20956, n24092);
xnor_4 g22485(new_n16120, new_n16118, n24096);
xnor_4 g22486(new_n12531, new_n12499, n24097);
xor_4  g22487(new_n12169, new_n12140, n24105);
xnor_4 g22488(new_n18740, new_n18719, n24119);
xnor_4 g22489(new_n15467_1, new_n15442, n24133);
xnor_4 g22490(new_n20558, new_n20527, n24141);
xnor_4 g22491(new_n21869, new_n21871, new_n24840_1);
xor_4  g22492(new_n24840_1, new_n21911, n24145);
xnor_4 g22493(new_n22615, new_n22612, n24146);
xor_4  g22494(new_n13139, new_n13079, n24155);
xnor_4 g22495(new_n24314, new_n24311, n24160);
xnor_4 g22496(new_n9454, new_n9417, n24167);
nor_5  g22497(new_n21105, new_n21100, n24172);
xnor_4 g22498(new_n14874, new_n14863, n24177);
xor_4  g22499(new_n24175, new_n24174, n24228);
xor_4  g22500(new_n18123, new_n18092, n24258);
or_5   g22501(new_n18868, new_n7228, new_n24850);
and_5  g22502(new_n24731, new_n24725, new_n24851);
or_5   g22503(new_n24851, new_n24728, new_n24852);
and_5  g22504(new_n24852, new_n24850, n24260);
xnor_4 g22505(new_n19714, new_n19683, n24289);
xnor_4 g22506(new_n4759, new_n4746, n24297);
xor_4  g22507(new_n12157_1, new_n3917, n24307);
xnor_4 g22508(new_n2536, new_n2525, n24342);
xnor_4 g22509(new_n16644, new_n16625, n24345);
xnor_4 g22510(new_n9715, new_n9704, n24347);
xnor_4 g22511(new_n5044, new_n4993, n24373);
xor_4  g22512(new_n18676, new_n18675, n24406);
xor_4  g22513(new_n14198, new_n14186, n24415);
xnor_4 g22514(new_n11051, new_n11050, n24421);
xnor_4 g22515(new_n14021, new_n13997, n24431);
xnor_4 g22516(new_n12299, new_n12271, n24472);
nor_5  g22517(new_n23459, new_n22959, new_n24866);
nor_5  g22518(new_n24866, new_n23461, new_n24867);
xor_4  g22519(new_n24867, new_n23455, n24476);
xnor_4 g22520(new_n10455, new_n10412, n24483);
xor_4  g22521(new_n13916, new_n13915, n24501);
xor_4  g22522(new_n18785, new_n18779, n24512);
xnor_4 g22523(new_n4763, new_n4761, n24558);
xor_4  g22524(new_n2814, new_n2813, n24576);
xnor_4 g22525(new_n2817, new_n2815, n24579);
xnor_4 g22526(new_n21052, new_n21039, n24602);
xnor_4 g22527(new_n14748, new_n14719, n24604);
xnor_4 g22528(new_n23585_1, new_n23581, n24626);
xor_4  g22529(new_n22627, new_n22624, n24629);
xor_4  g22530(new_n22377, new_n22366, n24636);
xnor_4 g22531(new_n22115, new_n22112, n24715);
xnor_4 g22532(new_n20988, new_n20932, n24723);
xor_4  g22533(new_n17368, new_n17323, new_n24882);
xor_4  g22534(new_n24882, new_n17443, n24749);
xnor_4 g22535(new_n20978, new_n20952, n24758);
xor_4  g22536(new_n23665, new_n23662, n24784);
xnor_4 g22537(new_n16798_1, new_n16797, n24807);
xor_4  g22538(new_n9964, new_n9963, n24826);
xor_4  g22539(new_n7715, new_n7665, n24840);
xor_4  g22540(new_n10238, new_n10225, n24841);
xor_4  g22541(new_n5234, new_n5220, n24853);
xnor_4 g22542(new_n3065, new_n3034, n24857);
xnor_4 g22543(new_n6436, new_n6420, n24887);
xor_4  g22544(new_n9443, new_n9436, n24934);
xor_4  g22545(new_n7504, new_n7422, n24998);
xnor_4 g22546(new_n11931, new_n11916, n25006);
xnor_4 g22547(new_n21365_1, new_n21351, n25032);
xnor_4 g22548(new_n16748, new_n16727, n25062);
xor_4  g22549(new_n20141, new_n17323, new_n24898);
xor_4  g22550(new_n24898, new_n20201, n25083);
xor_4  g22551(new_n13484_1, new_n13481, n25097);
xnor_4 g22552(new_n18395, new_n18392, n25133);
xnor_4 g22553(new_n19071, new_n19049, n25155);
xnor_4 g22554(new_n24614, new_n23446, new_n24903);
xor_4  g22555(new_n24903, new_n24611, n25181);
xnor_4 g22556(new_n21367_1, new_n21348, n25200);
not_10 g22557(new_n22132, new_n24906);
and_5  g22558(new_n22135, new_n24906, new_n24907);
xor_4  g22559(new_n22126_1, new_n17510, new_n24908);
xor_4  g22560(new_n24908, new_n24907, n25209);
xnor_4 g22561(new_n15674, new_n15672, n25215);
xor_4  g22562(new_n18873, new_n18870, n25244);
xnor_4 g22563(new_n18483_1, new_n18462, n25254);
xor_4  g22564(new_n21562, new_n21535, n25256);
nand_5 g22565(new_n24025, new_n22211, new_n24914);
nand_5 g22566(new_n24914, new_n24032_1, new_n24915);
xor_4  g22567(new_n24025, new_n23040, new_n24916);
xor_4  g22568(new_n24916, new_n24915, n25293);
xor_4  g22569(new_n21552, new_n21545, n25328);
xor_4  g22570(new_n11367, new_n4291, n25332);
and_5  g22571(new_n23647, new_n22287, new_n24920);
or_5   g22572(new_n23674, new_n24920, new_n24921);
nor_5  g22573(new_n23647, new_n22287, new_n24922);
or_5   g22574(new_n23673, new_n24922, new_n24923);
and_5  g22575(new_n24923, new_n24921, n25337);
xor_4  g22576(new_n11737, new_n11133, new_n24925);
xor_4  g22577(new_n24925, new_n11742, n25356);
xor_4  g22578(new_n9258, new_n9246_1, n25362);
xor_4  g22579(new_n14998, new_n14977_1, n25412);
xor_4  g22580(new_n15967_1, new_n15966, n25460);
xor_4  g22581(new_n7488, new_n7447, n25468);
xnor_4 g22582(new_n15002_1, new_n14973, n25499);
xor_4  g22583(new_n20548, new_n20546, n25513);
xnor_4 g22584(new_n12529, new_n12502, n25518);
xor_4  g22585(new_n13827, new_n13789, n25532);
xor_4  g22586(new_n20882, new_n20865, n25539);
xor_4  g22587(new_n17585, new_n17575, n25550);
xnor_4 g22588(new_n21678, new_n21664, n25611);
xnor_4 g22589(new_n5460, new_n5458, new_n24938);
xor_4  g22590(new_n24938, new_n5464, n25614);
xnor_4 g22591(new_n13214, new_n13184, n25619);
and_5  g22592(new_n23911, new_n23771, new_n24941);
or_5   g22593(new_n23916, new_n24941, new_n24942);
nor_5  g22594(new_n23911, new_n23771, new_n24943);
or_5   g22595(new_n23915, new_n24943, new_n24944);
and_5  g22596(new_n24944, new_n24942, n25665);
xnor_4 g22597(new_n9450, new_n9425, n25706);
xor_4  g22598(new_n23911, new_n20237, new_n24947);
xor_4  g22599(new_n24947, new_n24573, n25719);
xor_4  g22600(new_n9943, new_n9898, n25756);
not_10 g22601(new_n13407_1, new_n24950);
nor_5  g22602(new_n13448, new_n24950, new_n24951);
or_5   g22603(new_n13498, new_n24951, new_n24952);
and_5  g22604(new_n13448, new_n24950, new_n24953);
or_5   g22605(new_n13497, new_n24953, new_n24954);
and_5  g22606(new_n24954, new_n24952, n25758);
xor_4  g22607(new_n15390, new_n5831, n25773);
xnor_4 g22608(new_n21471_1, new_n18363, n25784);
xnor_4 g22609(new_n8524, new_n8499, n25792);
xor_4  g22610(new_n6981, new_n6943, n25816);
xnor_4 g22611(new_n6443, new_n6403, n25826);
xor_4  g22612(new_n12745, new_n12744, n25839);
xnor_4 g22613(new_n14583, new_n14531, n25840);
xnor_4 g22614(new_n8330, new_n8298, n25873);
xor_4  g22615(new_n24671, new_n24668, n25934);
xnor_4 g22616(new_n21903, new_n21888, n25938);
xnor_4 g22617(new_n22233, new_n22230, n25985);
xor_4  g22618(new_n14373, new_n9249, n25994);
nor_5  g22619(new_n19016, new_n18935, new_n24968);
and_5  g22620(new_n19087, new_n19017, new_n24969);
or_5   g22621(new_n24969, new_n24968, n26084);
xnor_4 g22622(new_n23670, new_n23655, n26096);
nor_5  g22623(new_n11957, new_n11878, new_n24972);
and_5  g22624(new_n24972, new_n11854, n26111);
xor_4  g22625(new_n11937, new_n11910, n26113);
xor_4  g22626(new_n20998, new_n20994, n26156);
xor_4  g22627(new_n17787, new_n17765, n26159);
xnor_4 g22628(new_n3718, new_n3671, n26179);
xor_4  g22629(new_n14565, new_n14564, n26220);
xnor_4 g22630(new_n23709, new_n23706, n26229);
xnor_4 g22631(new_n13132, new_n13096_1, n26237);
xnor_4 g22632(new_n16385, new_n16370, n26250);
xor_4  g22633(new_n21942, new_n21939, n26274);
xnor_4 g22634(new_n16389, new_n16359, n26287);
xor_4  g22635(new_n22150_1, new_n21376, new_n24984);
xor_4  g22636(new_n24984, new_n24494, n26317);
and_5  g22637(new_n19384, new_n19357_1, new_n24986);
or_5   g22638(new_n24986, new_n19381, new_n24987);
nor_5  g22639(new_n19384, new_n19357_1, new_n24988);
or_5   g22640(new_n24988, new_n19380, new_n24989);
and_5  g22641(new_n24989, new_n24987, n26353);
xnor_4 g22642(new_n21049, new_n21042, n26375);
or_5   g22643(new_n24058, new_n22272, new_n24992);
not_10 g22644(new_n24059, new_n24993);
or_5   g22645(new_n24068, new_n24993, new_n24994);
and_5  g22646(new_n24994, new_n24992, n26396);
xor_4  g22647(new_n5463, new_n5462, n26429);
xnor_4 g22648(new_n15079, new_n15061, n26431);
xnor_4 g22649(new_n7220, new_n7151, n26439);
xnor_4 g22650(new_n21294, new_n21292, n26492);
xnor_4 g22651(new_n10446, new_n10444, n26515);
xnor_4 g22652(new_n2540, new_n2514, n26538);
xnor_4 g22653(new_n15600, new_n15588_1, n26590);
xor_4  g22654(new_n20174, new_n17416, n26598);
xor_4  g22655(new_n24025, new_n22212, new_n25004);
xor_4  g22656(new_n25004, new_n24029, n26605);
xnor_4 g22657(new_n24002_1, new_n23992, new_n25006_1);
xor_4  g22658(new_n25006_1, new_n23997, n26656);
xnor_4 g22659(new_n11925, new_n11923, n26674);
xnor_4 g22660(new_n9807, new_n9791, n26675);
xnor_4 g22661(new_n21304, new_n21270, n26681);
nor_5  g22662(new_n5740, new_n5536, new_n25011);
or_5   g22663(new_n5827, new_n25011, new_n25012);
and_5  g22664(new_n5740, new_n5536, new_n25013);
or_5   g22665(new_n5826, new_n25013, new_n25014);
and_5  g22666(new_n25014, new_n25012, n26696);
xor_4  g22667(new_n15347, new_n15320, n26698);
xor_4  g22668(new_n16111, new_n5856, n26707);
xor_4  g22669(new_n24434, new_n24433, n26719);
xnor_4 g22670(new_n9445_1, new_n9433, n26727);
or_5   g22671(new_n22287, new_n20011, new_n25020);
nand_5 g22672(new_n22291, new_n22288, new_n25021);
and_5  g22673(new_n25021, new_n25020, n26729);
xor_4  g22674(new_n22312, new_n22309_1, n26745);
xnor_4 g22675(new_n8038, new_n8006_1, n26775);
xor_4  g22676(new_n10806, new_n10788, n26780);
xor_4  g22677(new_n22732, new_n22725, n26794);
xnor_4 g22678(new_n3390_1, new_n3331, n26795);
xnor_4 g22679(new_n11068, new_n11021, n26801);
xnor_4 g22680(new_n11450, new_n11432, n26815);
xnor_4 g22681(new_n24122, new_n24118, n26847);
xnor_4 g22682(new_n19384, new_n7417, new_n25031);
xor_4  g22683(new_n25031, new_n24244, n26900);
xor_4  g22684(new_n19534, new_n19533, n26902);
xor_4  g22685(new_n18047, new_n18044, n26905);
xnor_4 g22686(new_n8332, new_n8293, n26921);
xnor_4 g22687(new_n23103, new_n23086, n26923);
xnor_4 g22688(new_n11153, new_n11152, n26929);
xor_4  g22689(new_n13145, new_n13069, n26930);
xnor_4 g22690(new_n16387, new_n16365, n26943);
xor_4  g22691(new_n15004_1, new_n14969, n26970);
xor_4  g22692(new_n21834, new_n21821, n27004);
xnor_4 g22693(new_n10715, new_n10654, n27011);
xnor_4 g22694(new_n20199, new_n20145, n27019);
xnor_4 g22695(new_n5033, new_n5022, n27031);
xor_4  g22696(new_n22781, new_n21937, new_n25045);
xor_4  g22697(new_n25045, new_n22822, n27051);
xor_4  g22698(new_n17918, new_n17915, n27072);
xnor_4 g22699(new_n15989, new_n15928, n27079);
xnor_4 g22700(new_n15066, new_n4291, n27096);
xor_4  g22701(new_n14741, new_n14731, n27110);
xnor_4 g22702(new_n14134, new_n14131, n27112);
xor_4  g22703(new_n23110, new_n23109, n27130);
xor_4  g22704(new_n16742, new_n16733_1, n27145);
not_10 g22705(new_n15118_1, new_n25054);
nand_5 g22706(new_n17195, new_n25054, new_n25055);
nand_5 g22707(new_n22465, new_n22462, new_n25056);
and_5  g22708(new_n25056, new_n25055, n27158);
xnor_4 g22709(new_n22064, new_n22061, n27163);
xor_4  g22710(new_n24266, new_n21844, new_n25059);
xor_4  g22711(new_n25059, new_n24271, n27194);
endmodule


