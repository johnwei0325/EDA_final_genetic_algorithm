// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Thu Jun 27 02:53:54 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067_1, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095, new_n1096,
    new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269_1, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333_1, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355, new_n1356,
    new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471_1,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1, new_n2432,
    new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1, new_n2510,
    new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3263, new_n3264, new_n3265, new_n3266, new_n3267,
    new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1, new_n3273,
    new_n3274, new_n3275, new_n3276, new_n3277, new_n3278, new_n3279,
    new_n3280, new_n3281, new_n3282, new_n3283, new_n3284, new_n3285,
    new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290, new_n3291,
    new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297,
    new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303,
    new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309,
    new_n3310, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321,
    new_n3322, new_n3323, new_n3324, new_n3325, new_n3326, new_n3327,
    new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339_1,
    new_n3340, new_n3341, new_n3342_1, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986_1, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992_1, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005_1, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086_1, new_n4087, new_n4088_1, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094_1, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141_1, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155_1, new_n4156, new_n4157,
    new_n4158, new_n4159_1, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187_1,
    new_n4188, new_n4189_1, new_n4190_1, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203_1, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4211,
    new_n4212, new_n4213, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226_1, new_n4227, new_n4228, new_n4229,
    new_n4230_1, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300_1, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312_1, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326_1, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333_1, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370_1, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378_1, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397_1,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436_1, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4451, new_n4452, new_n4453, new_n4454, new_n4455,
    new_n4456, new_n4457, new_n4458, new_n4459, new_n4460, new_n4461,
    new_n4462, new_n4463, new_n4464, new_n4465, new_n4466, new_n4467,
    new_n4468, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473,
    new_n4474, new_n4475, new_n4476, new_n4477, new_n4478, new_n4479,
    new_n4480, new_n4481, new_n4482, new_n4483, new_n4484, new_n4485,
    new_n4486, new_n4487, new_n4488, new_n4489, new_n4490, new_n4491,
    new_n4492, new_n4493, new_n4494, new_n4495, new_n4496, new_n4497,
    new_n4498, new_n4499_1, new_n4500, new_n4501, new_n4502, new_n4503,
    new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509,
    new_n4510, new_n4511, new_n4512, new_n4513, new_n4514, new_n4515,
    new_n4516_1, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521,
    new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527,
    new_n4528, new_n4529, new_n4530, new_n4531, new_n4532, new_n4533,
    new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539,
    new_n4540, new_n4541, new_n4542, new_n4543, new_n4544, new_n4545,
    new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551,
    new_n4552, new_n4553_1, new_n4554, new_n4555, new_n4556, new_n4557,
    new_n4558, new_n4559, new_n4560, new_n4561, new_n4562, new_n4563,
    new_n4564, new_n4565, new_n4566, new_n4567, new_n4568, new_n4569,
    new_n4570, new_n4571, new_n4572, new_n4573, new_n4574, new_n4575,
    new_n4576, new_n4577, new_n4578, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599,
    new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605,
    new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611,
    new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617,
    new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623,
    new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634_1, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686_1, new_n4687, new_n4688, new_n4689_1,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733_1, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757_1, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805_1, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817_1, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826_1, new_n4827,
    new_n4828_1, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212_1, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314_1, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1,
    new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643, new_n5644,
    new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859, new_n5860_1,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934_1, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089_1,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254_1, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273_1, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294_1,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358_1, new_n6359_1, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429_1, new_n6430, new_n6431_1, new_n6434, new_n6435,
    new_n6436, new_n6437, new_n6438, new_n6439, new_n6440, new_n6441_1,
    new_n6442, new_n6443, new_n6444, new_n6445_1, new_n6446, new_n6447,
    new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453,
    new_n6454, new_n6455, new_n6456, new_n6457, new_n6458, new_n6459,
    new_n6460, new_n6461, new_n6462, new_n6463, new_n6464, new_n6465,
    new_n6466, new_n6467, new_n6468, new_n6469, new_n6470, new_n6471,
    new_n6472, new_n6473, new_n6474, new_n6475, new_n6476, new_n6477,
    new_n6478, new_n6479, new_n6480, new_n6481, new_n6482, new_n6483,
    new_n6484, new_n6485, new_n6486, new_n6487, new_n6488, new_n6489,
    new_n6490, new_n6491, new_n6492, new_n6493, new_n6494, new_n6495,
    new_n6496, new_n6497, new_n6498, new_n6499, new_n6500, new_n6501,
    new_n6502, new_n6503, new_n6504, new_n6505, new_n6506, new_n6507,
    new_n6508, new_n6509, new_n6510, new_n6511, new_n6512, new_n6513,
    new_n6514, new_n6515, new_n6516, new_n6517, new_n6518, new_n6519,
    new_n6520, new_n6521, new_n6522, new_n6523, new_n6524, new_n6525,
    new_n6526, new_n6527, new_n6528, new_n6529, new_n6530, new_n6531,
    new_n6532, new_n6533, new_n6534, new_n6535, new_n6536, new_n6537,
    new_n6538, new_n6539, new_n6540, new_n6541, new_n6542, new_n6543,
    new_n6544, new_n6545, new_n6546, new_n6547, new_n6548, new_n6549,
    new_n6550, new_n6551, new_n6552, new_n6553, new_n6554, new_n6555,
    new_n6556, new_n6557, new_n6558, new_n6559, new_n6560, new_n6561,
    new_n6562, new_n6563, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578_1, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604_1, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611_1, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645_1,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687_1,
    new_n6688, new_n6689_1, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703_1, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742_1, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770_1, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776_1, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797_1, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806_1, new_n6807,
    new_n6808, new_n6809_1, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822_1, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860_1, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877_1, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941,
    new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947,
    new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986_1, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013,
    new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019,
    new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025,
    new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031,
    new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159_1, new_n7160_1, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193_1,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265_1,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270_1, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294_1, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320_1, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523_1,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7635, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009,
    new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028_1, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100_1, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202_1, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303_1, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336_1, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384_1, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398_1, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8431, new_n8432, new_n8433_1, new_n8434, new_n8435, new_n8436,
    new_n8437, new_n8438, new_n8439, new_n8440, new_n8441, new_n8442,
    new_n8443, new_n8447, new_n8448, new_n8449, new_n8450, new_n8451,
    new_n8452, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595_1, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665_1, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717_1, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759_1, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819_1, new_n8820, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930,
    new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080_1,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111_1, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137_1, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189_1, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195_1, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241_1, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338,
    new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9344,
    new_n9345, new_n9346, new_n9347, new_n9348, new_n9349, new_n9350,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387_1, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400_1, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457_1, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571_1, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578_1, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583_1, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637_1, new_n9638, new_n9639, new_n9640_1, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706_1, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725_1,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756_1, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820_1, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920_1, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956_1, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022_1, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174_1, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217_1, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223_1, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278_1, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295, new_n10296, new_n10297,
    new_n10298, new_n10299, new_n10300, new_n10301, new_n10302, new_n10303,
    new_n10304, new_n10305, new_n10306, new_n10307, new_n10308, new_n10309,
    new_n10310, new_n10311, new_n10312, new_n10313, new_n10314, new_n10315,
    new_n10316, new_n10317, new_n10318, new_n10319, new_n10320, new_n10321,
    new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327_1, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391_1, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439_1, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451_1, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476_1,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510_1, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545_1, new_n10546,
    new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558,
    new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564,
    new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570,
    new_n10571, new_n10572, new_n10573, new_n10574, new_n10575, new_n10576,
    new_n10577, new_n10578, new_n10579, new_n10580, new_n10581, new_n10582,
    new_n10583, new_n10584, new_n10585, new_n10586, new_n10587, new_n10588,
    new_n10589_1, new_n10590, new_n10591, new_n10592, new_n10593,
    new_n10594, new_n10595, new_n10596, new_n10597, new_n10598, new_n10599,
    new_n10600, new_n10601, new_n10602, new_n10603, new_n10604, new_n10605,
    new_n10606, new_n10607, new_n10608, new_n10609, new_n10610, new_n10611,
    new_n10612, new_n10613, new_n10614, new_n10615, new_n10616, new_n10617,
    new_n10618, new_n10619, new_n10620, new_n10621, new_n10622, new_n10623,
    new_n10624, new_n10625, new_n10626, new_n10627, new_n10628, new_n10629,
    new_n10630, new_n10631, new_n10632, new_n10633, new_n10634, new_n10635,
    new_n10636, new_n10637, new_n10638, new_n10639, new_n10640, new_n10641,
    new_n10642, new_n10643, new_n10644_1, new_n10645, new_n10646,
    new_n10647, new_n10648, new_n10649, new_n10650, new_n10651, new_n10652,
    new_n10653, new_n10654, new_n10655, new_n10656, new_n10657, new_n10658,
    new_n10659, new_n10660, new_n10661, new_n10662, new_n10663, new_n10664,
    new_n10665, new_n10666, new_n10667, new_n10668, new_n10669, new_n10670,
    new_n10671, new_n10672, new_n10673, new_n10674, new_n10675, new_n10676,
    new_n10677, new_n10678_1, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685_1, new_n10686,
    new_n10687, new_n10688, new_n10689, new_n10690, new_n10691, new_n10692,
    new_n10693, new_n10694, new_n10695_1, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10701, new_n10702, new_n10703,
    new_n10704, new_n10705, new_n10706, new_n10707, new_n10708, new_n10709,
    new_n10710, new_n10711, new_n10712, new_n10713, new_n10714, new_n10715,
    new_n10716, new_n10717, new_n10718, new_n10719, new_n10720, new_n10721,
    new_n10722, new_n10723, new_n10724, new_n10725, new_n10726, new_n10727,
    new_n10728, new_n10729, new_n10730, new_n10731, new_n10732, new_n10733,
    new_n10734, new_n10735, new_n10736, new_n10737, new_n10738, new_n10739,
    new_n10740, new_n10741, new_n10742, new_n10743, new_n10744, new_n10745,
    new_n10746, new_n10747, new_n10748, new_n10749, new_n10750, new_n10751,
    new_n10752, new_n10753, new_n10754, new_n10755, new_n10756, new_n10757,
    new_n10758, new_n10759, new_n10760, new_n10761, new_n10762, new_n10763,
    new_n10764, new_n10765, new_n10766, new_n10767, new_n10768, new_n10769,
    new_n10770, new_n10771, new_n10772, new_n10773, new_n10774, new_n10775,
    new_n10776, new_n10777, new_n10778, new_n10779, new_n10780, new_n10781,
    new_n10782, new_n10783, new_n10784, new_n10785, new_n10786, new_n10787,
    new_n10788, new_n10789_1, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848_1, new_n10849, new_n10850, new_n10851_1,
    new_n10852, new_n10853, new_n10854, new_n10855, new_n10856, new_n10857,
    new_n10858, new_n10859, new_n10860, new_n10861, new_n10862, new_n10863,
    new_n10864, new_n10865, new_n10866, new_n10867, new_n10868, new_n10869,
    new_n10870, new_n10871, new_n10872, new_n10873, new_n10874, new_n10875,
    new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881,
    new_n10882, new_n10883, new_n10884, new_n10885, new_n10886, new_n10887,
    new_n10888, new_n10889, new_n10890, new_n10891, new_n10892, new_n10893,
    new_n10894, new_n10895, new_n10896, new_n10897, new_n10898_1,
    new_n10899, new_n10900, new_n10901, new_n10902, new_n10903, new_n10904,
    new_n10905, new_n10906, new_n10907, new_n10908, new_n10909, new_n10910,
    new_n10911, new_n10912, new_n10913_1, new_n10914, new_n10915,
    new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921,
    new_n10922, new_n10923, new_n10924, new_n10925, new_n10926, new_n10927,
    new_n10928_1, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944,
    new_n10945, new_n10946, new_n10947, new_n10948, new_n10949_1,
    new_n10950, new_n10951, new_n10952, new_n10953, new_n10954, new_n10955,
    new_n10956, new_n10957, new_n10958, new_n10959, new_n10960, new_n10961,
    new_n10962, new_n10963, new_n10964, new_n10965_1, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989,
    new_n10990_1, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023_1,
    new_n11024, new_n11025, new_n11026, new_n11027, new_n11028, new_n11029,
    new_n11030, new_n11031, new_n11032, new_n11033, new_n11034, new_n11035,
    new_n11036, new_n11037, new_n11038, new_n11039, new_n11040, new_n11041,
    new_n11042, new_n11043, new_n11044, new_n11045, new_n11046, new_n11047,
    new_n11048, new_n11049, new_n11050, new_n11051, new_n11052, new_n11053,
    new_n11054, new_n11055, new_n11056, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063, new_n11064, new_n11065,
    new_n11066, new_n11067, new_n11068, new_n11069, new_n11070, new_n11071,
    new_n11072, new_n11073, new_n11074, new_n11075, new_n11076, new_n11077,
    new_n11078, new_n11079, new_n11080, new_n11081, new_n11082, new_n11083,
    new_n11084, new_n11085, new_n11086, new_n11087, new_n11088, new_n11089,
    new_n11090, new_n11091, new_n11092, new_n11093, new_n11094, new_n11095,
    new_n11096, new_n11097, new_n11098, new_n11099, new_n11100, new_n11101,
    new_n11102, new_n11103, new_n11104, new_n11105, new_n11106, new_n11107,
    new_n11108, new_n11109, new_n11110, new_n11111, new_n11112, new_n11113,
    new_n11114, new_n11115, new_n11116, new_n11117, new_n11118, new_n11119,
    new_n11120, new_n11121, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127, new_n11128, new_n11129, new_n11130, new_n11131,
    new_n11132, new_n11133, new_n11134, new_n11135, new_n11136, new_n11137,
    new_n11138, new_n11139, new_n11140, new_n11141, new_n11142, new_n11143,
    new_n11144, new_n11145, new_n11146, new_n11147, new_n11148, new_n11149,
    new_n11150, new_n11151, new_n11152, new_n11153_1, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11181,
    new_n11182, new_n11183, new_n11184, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201, new_n11202, new_n11203, new_n11204, new_n11205,
    new_n11206, new_n11207, new_n11208, new_n11209, new_n11210, new_n11211,
    new_n11212, new_n11213, new_n11214, new_n11215, new_n11216_1,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221,
    new_n11222_1, new_n11223, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238,
    new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244,
    new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257_1, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11312, new_n11313, new_n11314, new_n11315,
    new_n11316, new_n11317, new_n11318, new_n11319, new_n11320, new_n11321,
    new_n11322, new_n11323, new_n11324, new_n11325, new_n11326_1,
    new_n11327, new_n11328, new_n11329, new_n11330, new_n11331, new_n11332,
    new_n11333, new_n11334, new_n11335, new_n11336, new_n11337, new_n11338,
    new_n11339, new_n11340, new_n11341, new_n11342, new_n11343, new_n11344,
    new_n11345, new_n11346, new_n11347, new_n11348, new_n11349, new_n11350,
    new_n11351, new_n11352, new_n11353, new_n11354, new_n11355, new_n11356,
    new_n11357, new_n11358, new_n11359, new_n11360, new_n11361, new_n11362,
    new_n11363, new_n11364, new_n11365, new_n11366, new_n11367, new_n11368,
    new_n11369, new_n11370, new_n11371, new_n11372, new_n11373, new_n11374,
    new_n11375, new_n11376, new_n11377, new_n11378, new_n11379, new_n11380,
    new_n11381, new_n11382, new_n11383, new_n11384, new_n11385, new_n11386,
    new_n11387, new_n11388, new_n11389, new_n11390, new_n11391, new_n11392,
    new_n11393, new_n11394, new_n11395, new_n11396, new_n11397, new_n11398,
    new_n11399, new_n11400, new_n11401, new_n11402, new_n11403, new_n11404,
    new_n11405, new_n11406, new_n11407_1, new_n11408, new_n11409,
    new_n11410, new_n11411, new_n11412, new_n11413, new_n11414, new_n11415,
    new_n11416, new_n11417, new_n11418, new_n11419, new_n11420, new_n11421,
    new_n11422, new_n11423_1, new_n11424, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444,
    new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450,
    new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462,
    new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468,
    new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478_1, new_n11479,
    new_n11480, new_n11481, new_n11482, new_n11483, new_n11484, new_n11485,
    new_n11486, new_n11487, new_n11488, new_n11489, new_n11490, new_n11491,
    new_n11492, new_n11493, new_n11494, new_n11495, new_n11496, new_n11497,
    new_n11498, new_n11499, new_n11500, new_n11501, new_n11502, new_n11503,
    new_n11504, new_n11505, new_n11506, new_n11507, new_n11508, new_n11509,
    new_n11510, new_n11511, new_n11512, new_n11513, new_n11514, new_n11515,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536_1, new_n11537, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11571, new_n11572, new_n11573, new_n11574,
    new_n11575, new_n11576, new_n11577, new_n11578, new_n11579, new_n11580,
    new_n11581, new_n11582, new_n11583, new_n11584, new_n11585, new_n11586,
    new_n11587, new_n11588, new_n11589, new_n11590, new_n11591, new_n11592,
    new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607, new_n11608, new_n11609, new_n11610,
    new_n11611, new_n11612, new_n11613, new_n11614, new_n11615, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652,
    new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658,
    new_n11659, new_n11660, new_n11661, new_n11662_1, new_n11663,
    new_n11664, new_n11665, new_n11666, new_n11667, new_n11668, new_n11669,
    new_n11670, new_n11671, new_n11672, new_n11673, new_n11674, new_n11675,
    new_n11676, new_n11677, new_n11678, new_n11679, new_n11680, new_n11681,
    new_n11682, new_n11683, new_n11684, new_n11685, new_n11686, new_n11687,
    new_n11688, new_n11689, new_n11690, new_n11691, new_n11692, new_n11693,
    new_n11694, new_n11695, new_n11696, new_n11697, new_n11698, new_n11699,
    new_n11700, new_n11701, new_n11702, new_n11703, new_n11704, new_n11705,
    new_n11706, new_n11707_1, new_n11708, new_n11709, new_n11710,
    new_n11711, new_n11712, new_n11713, new_n11714, new_n11715, new_n11716,
    new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722,
    new_n11723, new_n11724, new_n11725, new_n11726, new_n11727,
    new_n11728_1, new_n11729, new_n11730, new_n11731, new_n11732,
    new_n11733, new_n11734, new_n11735, new_n11736, new_n11737, new_n11738,
    new_n11739, new_n11740, new_n11741, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749, new_n11750,
    new_n11751, new_n11752, new_n11753, new_n11754, new_n11755_1,
    new_n11756, new_n11757_1, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780_1, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11790, new_n11791_1, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11817, new_n11818,
    new_n11819, new_n11820, new_n11821_1, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876_1,
    new_n11877_1, new_n11878, new_n11879, new_n11880, new_n11881,
    new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887,
    new_n11888, new_n11889, new_n11890, new_n11891, new_n11892_1,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917_1, new_n11918, new_n11919_1, new_n11920, new_n11921,
    new_n11922_1, new_n11923, new_n11924, new_n11925, new_n11926,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956,
    new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962,
    new_n11963, new_n11964, new_n11965, new_n11966, new_n11967_1,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999_1, new_n12000_1, new_n12001, new_n12002,
    new_n12003, new_n12004, new_n12005_1, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014_1, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020_1, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025_1, new_n12026, new_n12027, new_n12028,
    new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044_1, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069_1, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076_1, new_n12077, new_n12078,
    new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108,
    new_n12109, new_n12110, new_n12111_1, new_n12112, new_n12113,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121, new_n12122, new_n12123, new_n12124, new_n12125,
    new_n12126, new_n12127, new_n12128, new_n12129, new_n12130, new_n12131,
    new_n12132, new_n12133, new_n12134, new_n12135, new_n12136, new_n12137,
    new_n12138, new_n12139, new_n12140, new_n12141, new_n12142, new_n12143,
    new_n12144, new_n12145_1, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12209, new_n12210, new_n12211, new_n12212, new_n12213,
    new_n12214, new_n12215, new_n12216, new_n12217, new_n12218, new_n12219,
    new_n12220, new_n12221_1, new_n12222, new_n12223, new_n12224,
    new_n12225, new_n12226, new_n12227, new_n12228, new_n12229, new_n12230,
    new_n12231, new_n12232, new_n12233, new_n12234, new_n12235, new_n12236,
    new_n12237, new_n12238, new_n12239, new_n12240, new_n12241, new_n12242,
    new_n12243, new_n12244, new_n12245, new_n12246, new_n12247_1,
    new_n12248, new_n12249, new_n12250, new_n12251, new_n12252, new_n12253,
    new_n12254, new_n12255, new_n12256, new_n12257, new_n12258, new_n12259,
    new_n12260, new_n12261, new_n12262, new_n12263, new_n12264, new_n12265,
    new_n12266, new_n12267, new_n12268, new_n12269, new_n12270, new_n12271,
    new_n12272, new_n12273, new_n12274, new_n12275, new_n12276, new_n12277,
    new_n12278, new_n12279, new_n12280, new_n12281, new_n12282, new_n12283,
    new_n12284, new_n12285, new_n12286, new_n12287, new_n12288, new_n12289,
    new_n12290, new_n12291, new_n12292, new_n12293, new_n12294, new_n12295,
    new_n12296, new_n12297, new_n12298, new_n12299_1, new_n12300,
    new_n12301, new_n12302, new_n12303, new_n12304, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12322, new_n12323, new_n12324,
    new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336,
    new_n12337, new_n12338, new_n12339, new_n12340, new_n12341, new_n12342,
    new_n12343, new_n12344, new_n12345, new_n12346, new_n12347, new_n12348,
    new_n12349, new_n12350, new_n12351, new_n12352, new_n12353, new_n12354,
    new_n12355, new_n12356, new_n12357, new_n12358, new_n12359, new_n12360,
    new_n12361, new_n12362, new_n12363, new_n12364, new_n12365, new_n12366,
    new_n12367, new_n12368, new_n12369, new_n12370, new_n12371, new_n12372,
    new_n12373, new_n12374, new_n12375, new_n12376, new_n12377, new_n12378,
    new_n12379, new_n12380, new_n12381, new_n12382, new_n12383, new_n12384,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391_1, new_n12392, new_n12393, new_n12394, new_n12395,
    new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413,
    new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444_1, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489_1,
    new_n12490, new_n12491, new_n12492, new_n12493, new_n12494, new_n12495,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506, new_n12507,
    new_n12508, new_n12509, new_n12510, new_n12511_1, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540, new_n12541, new_n12542,
    new_n12543, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554,
    new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560,
    new_n12561, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591_1,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626, new_n12627,
    new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648_1, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702, new_n12703,
    new_n12704_1, new_n12705_1, new_n12706_1, new_n12707, new_n12708,
    new_n12709_1, new_n12710, new_n12711, new_n12712, new_n12713,
    new_n12714, new_n12715, new_n12716, new_n12717, new_n12718, new_n12719,
    new_n12720_1, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12740, new_n12741, new_n12742,
    new_n12743, new_n12744, new_n12745, new_n12746, new_n12747, new_n12748,
    new_n12749, new_n12750, new_n12751, new_n12752, new_n12753_1,
    new_n12754, new_n12755, new_n12756, new_n12757, new_n12758, new_n12759,
    new_n12760, new_n12761, new_n12762, new_n12763, new_n12764, new_n12765,
    new_n12766, new_n12767, new_n12768, new_n12769, new_n12770, new_n12771,
    new_n12772, new_n12773, new_n12774, new_n12775, new_n12776,
    new_n12777_1, new_n12778, new_n12779, new_n12780, new_n12781,
    new_n12782, new_n12783, new_n12784, new_n12785, new_n12786, new_n12787,
    new_n12788, new_n12789, new_n12790, new_n12791, new_n12792, new_n12793,
    new_n12794, new_n12795, new_n12796, new_n12797, new_n12798, new_n12799,
    new_n12800, new_n12801, new_n12802, new_n12803, new_n12804, new_n12805,
    new_n12806, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925_1,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947_1, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128,
    new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134,
    new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140,
    new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368,
    new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374,
    new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380,
    new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386,
    new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392,
    new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398,
    new_n13399, new_n13400, new_n13401, new_n13402, new_n13403, new_n13404,
    new_n13405, new_n13406, new_n13407, new_n13408, new_n13409, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422,
    new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458,
    new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464,
    new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470,
    new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476,
    new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482,
    new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488,
    new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500,
    new_n13501, new_n13502, new_n13503, new_n13504, new_n13505, new_n13506,
    new_n13507, new_n13508, new_n13509, new_n13510, new_n13511, new_n13512,
    new_n13513, new_n13515, new_n13517, new_n13518, new_n13519, new_n13520,
    new_n13521, new_n13522, new_n13523, new_n13524, new_n13525, new_n13526,
    new_n13527, new_n13528, new_n13529, new_n13530, new_n13531, new_n13532,
    new_n13533, new_n13534, new_n13535, new_n13536, new_n13537, new_n13538,
    new_n13539, new_n13540, new_n13541, new_n13542, new_n13543, new_n13544,
    new_n13545, new_n13546, new_n13547, new_n13548, new_n13549, new_n13550,
    new_n13551, new_n13552, new_n13553, new_n13554, new_n13555, new_n13556,
    new_n13557, new_n13558, new_n13559, new_n13560, new_n13561, new_n13562,
    new_n13563, new_n13564, new_n13565, new_n13566, new_n13567, new_n13568,
    new_n13569, new_n13570, new_n13571, new_n13572, new_n13573, new_n13574,
    new_n13575, new_n13576, new_n13577, new_n13578, new_n13579, new_n13580,
    new_n13581, new_n13582, new_n13583, new_n13584, new_n13585, new_n13586,
    new_n13587, new_n13588, new_n13589, new_n13590, new_n13591, new_n13592,
    new_n13593, new_n13594, new_n13595, new_n13596, new_n13597, new_n13598,
    new_n13599, new_n13600, new_n13601, new_n13602, new_n13603, new_n13604,
    new_n13605, new_n13606, new_n13607, new_n13608, new_n13609, new_n13610,
    new_n13611, new_n13612, new_n13613, new_n13614, new_n13615, new_n13616,
    new_n13617, new_n13618, new_n13619, new_n13620, new_n13621, new_n13622,
    new_n13623, new_n13624, new_n13625, new_n13626, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634,
    new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640,
    new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646,
    new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652,
    new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658,
    new_n13659, new_n13660, new_n13661, new_n13662, new_n13663, new_n13664,
    new_n13665, new_n13666, new_n13667, new_n13668, new_n13669, new_n13670,
    new_n13671, new_n13672, new_n13673, new_n13674, new_n13675, new_n13676,
    new_n13677, new_n13678, new_n13679, new_n13680, new_n13681, new_n13682,
    new_n13683, new_n13684, new_n13685, new_n13686, new_n13687, new_n13688,
    new_n13689, new_n13690, new_n13691, new_n13692, new_n13693, new_n13694,
    new_n13695, new_n13696, new_n13697, new_n13698, new_n13699, new_n13700,
    new_n13701, new_n13702, new_n13703, new_n13704, new_n13705, new_n13706,
    new_n13707, new_n13708, new_n13709, new_n13710, new_n13711, new_n13712,
    new_n13713, new_n13714, new_n13715, new_n13716, new_n13717, new_n13718,
    new_n13719, new_n13720, new_n13721, new_n13722, new_n13723, new_n13724,
    new_n13725, new_n13726, new_n13727, new_n13728, new_n13729, new_n13730,
    new_n13731, new_n13732, new_n13733, new_n13734, new_n13735, new_n13736,
    new_n13737, new_n13738, new_n13739, new_n13740, new_n13741, new_n13742,
    new_n13743, new_n13744, new_n13745, new_n13746, new_n13747, new_n13748,
    new_n13760, new_n13761, new_n13762, new_n13763, new_n13764, new_n13765,
    new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771,
    new_n13772, new_n13773, new_n13774, new_n13775, new_n13776, new_n13777,
    new_n13778, new_n13779, new_n13780, new_n13781, new_n13782, new_n13783,
    new_n13784, new_n13785, new_n13786, new_n13787, new_n13788, new_n13789,
    new_n13790, new_n13791, new_n13792, new_n13793, new_n13794, new_n13795,
    new_n13796, new_n13797, new_n13798, new_n13799, new_n13800, new_n13801,
    new_n13802, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807,
    new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813,
    new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819,
    new_n13820, new_n13821, new_n13822, new_n13823, new_n13824, new_n13825,
    new_n13826, new_n13827, new_n13828, new_n13829, new_n13830, new_n13831,
    new_n13832, new_n13833, new_n13834, new_n13835, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047,
    new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14053,
    new_n14054, new_n14055, new_n14056, new_n14059, new_n14064, new_n14071,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081, new_n14082, new_n14083,
    new_n14084, new_n14085, new_n14086, new_n14087, new_n14088, new_n14089,
    new_n14090, new_n14091, new_n14092, new_n14093, new_n14094, new_n14095,
    new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101,
    new_n14102, new_n14103, new_n14104, new_n14105, new_n14106, new_n14107,
    new_n14108, new_n14109, new_n14110, new_n14111, new_n14112, new_n14113,
    new_n14114, new_n14115, new_n14116, new_n14117, new_n14118, new_n14119,
    new_n14120, new_n14121, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126, new_n14127, new_n14128, new_n14129, new_n14130, new_n14131,
    new_n14132, new_n14133, new_n14134, new_n14135, new_n14136, new_n14137,
    new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143,
    new_n14144, new_n14145, new_n14146, new_n14147, new_n14148, new_n14149,
    new_n14150, new_n14151, new_n14152, new_n14153, new_n14154, new_n14155,
    new_n14156, new_n14157, new_n14158, new_n14159, new_n14160, new_n14161,
    new_n14162, new_n14163, new_n14164, new_n14165, new_n14166, new_n14167,
    new_n14168, new_n14169, new_n14170, new_n14171, new_n14172, new_n14173,
    new_n14174, new_n14175, new_n14176, new_n14177, new_n14178, new_n14179,
    new_n14180, new_n14181, new_n14182, new_n14183, new_n14184, new_n14185,
    new_n14186, new_n14187, new_n14188, new_n14189, new_n14190, new_n14191,
    new_n14192, new_n14193, new_n14194, new_n14195, new_n14196, new_n14197,
    new_n14198, new_n14199, new_n14200, new_n14201, new_n14202, new_n14203,
    new_n14204, new_n14205, new_n14206, new_n14207, new_n14208, new_n14209,
    new_n14210, new_n14211, new_n14212, new_n14213, new_n14214, new_n14215,
    new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221,
    new_n14222, new_n14223, new_n14224, new_n14225, new_n14226, new_n14227,
    new_n14228, new_n14229, new_n14230, new_n14231, new_n14232, new_n14233,
    new_n14234, new_n14235, new_n14236, new_n14237, new_n14238, new_n14239,
    new_n14240, new_n14241, new_n14242, new_n14243, new_n14244, new_n14245,
    new_n14246, new_n14247, new_n14248, new_n14249, new_n14250, new_n14251,
    new_n14252, new_n14253, new_n14254, new_n14255, new_n14256, new_n14257,
    new_n14258, new_n14259, new_n14260, new_n14261, new_n14262, new_n14263,
    new_n14264, new_n14265, new_n14266, new_n14267, new_n14268, new_n14269,
    new_n14270, new_n14271, new_n14272, new_n14273, new_n14274, new_n14275,
    new_n14276, new_n14277, new_n14278, new_n14279, new_n14280, new_n14281,
    new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287,
    new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293,
    new_n14294, new_n14295, new_n14296, new_n14297, new_n14298, new_n14299,
    new_n14300, new_n14301, new_n14302, new_n14303, new_n14304, new_n14305,
    new_n14306, new_n14307, new_n14308, new_n14309, new_n14319;
and_8  g00000(n6687, n6038, new_n377);
and_8  g00001(n8336, n7354, new_n378);
and_8  g00002(n11222, n8028, new_n379);
and_8  g00003(n12069, n1564, new_n380);
xor_4  g00004(new_n380, new_n379, new_n381_1);
xor_4  g00005(new_n381_1, new_n378, new_n382);
xor_4  g00006(new_n382, new_n377, n112);
and_8  g00007(n12720, n4312, new_n384);
and_8  g00008(n12025, n6038, new_n385);
and_8  g00009(n12705, n2509, new_n386);
xor_4  g00010(new_n386, new_n385, new_n387);
xor_4  g00011(new_n387, new_n384, new_n388);
and_8  g00012(n12705, n6038, new_n389);
and_8  g00013(n12720, n1097, new_n390);
or_8   g00014(new_n390, new_n389, new_n391);
and_8  g00015(n4312, n2509, new_n392);
xnor_4 g00016(new_n390, new_n389, new_n393);
or_8   g00017(new_n393, new_n392, new_n394);
and_8  g00018(new_n394, new_n391, new_n395);
xor_4  g00019(new_n395, new_n388, new_n396);
and_8  g00020(n2508, n1097, new_n397_1);
and_8  g00021(n5964, n2585, new_n398);
xor_4  g00022(new_n398, new_n397_1, new_n399);
xor_4  g00023(new_n399, new_n396, new_n400);
nand_5 g00024(n5964, n2508, new_n401);
xor_4  g00025(new_n393, new_n392, new_n402);
and_8  g00026(new_n402, new_n401, new_n403);
nor_6  g00027(new_n402, new_n401, new_n404);
or_8   g00028(new_n404, new_n403, new_n405_1);
and_8  g00029(n6038, n4312, new_n406);
and_8  g00030(n12720, n5964, new_n407);
or_8   g00031(new_n407, new_n406, new_n408);
nand_5 g00032(new_n407, new_n406, new_n409);
nand_5 g00033(n2509, n1097, new_n410);
nand_5 g00034(new_n410, new_n409, new_n411);
and_8  g00035(new_n411, new_n408, new_n412);
nor_6  g00036(new_n412, new_n405_1, new_n413);
nor_6  g00037(new_n413, new_n403, new_n414);
xor_4  g00038(new_n414, new_n400, new_n415);
and_8  g00039(n5305, n2585, new_n416);
and_8  g00040(new_n412, new_n405_1, new_n417);
or_8   g00041(new_n417, new_n413, new_n418);
or_8   g00042(new_n418, new_n416, new_n419);
not_8  g00043(new_n416, new_n420);
xor_4  g00044(new_n418, new_n420, new_n421);
and_8  g00045(n5305, n2508, new_n422);
and_8  g00046(n6038, n1097, new_n423);
and_8  g00047(n12720, n5305, new_n424);
and_8  g00048(new_n424, new_n423, new_n425);
or_8   g00049(new_n424, new_n423, new_n426);
and_8  g00050(n5964, n2509, new_n427);
and_8  g00051(new_n427, new_n426, new_n428);
or_8   g00052(new_n428, new_n425, new_n429);
and_8  g00053(new_n429, new_n422, new_n430);
xor_4  g00054(new_n429, new_n422, new_n431);
and_8  g00055(new_n409, new_n408, new_n432);
xnor_4 g00056(new_n432, new_n410, new_n433);
and_8  g00057(new_n433, new_n431, new_n434);
or_8   g00058(new_n434, new_n430, new_n435);
or_8   g00059(new_n435, new_n421, new_n436);
and_8  g00060(new_n436, new_n419, new_n437);
and_8  g00061(new_n437, new_n415, new_n438);
and_8  g00062(new_n387, new_n384, new_n439);
and_8  g00063(new_n395, new_n388, new_n440);
or_8   g00064(new_n440, new_n439, new_n441);
and_8  g00065(n5964, n4005, new_n442);
and_8  g00066(n2585, n1097, new_n443);
and_8  g00067(n12706, n5305, new_n444);
xnor_4 g00068(new_n444, new_n443, new_n445);
xor_4  g00069(new_n445, new_n442, new_n446);
xor_4  g00070(new_n446, new_n441, new_n447_1);
and_8  g00071(new_n386, new_n385, new_n448);
and_8  g00072(n4312, n2508, new_n449);
xnor_4 g00073(new_n449, new_n448, new_n450);
and_8  g00074(n12025, n2509, new_n451);
and_8  g00075(n12720, n12705, new_n452);
and_8  g00076(n11257, n6038, new_n453);
xnor_4 g00077(new_n453, new_n452, new_n454);
xor_4  g00078(new_n454, new_n451, new_n455);
xor_4  g00079(new_n455, new_n450, new_n456);
xor_4  g00080(new_n456, new_n447_1, new_n457);
nand_5 g00081(new_n399, new_n396, new_n458);
and_8  g00082(new_n398, new_n397_1, new_n459);
and_8  g00083(new_n414, new_n400, new_n460);
and_8  g00084(new_n460, new_n459, new_n461);
nor_6  g00085(new_n460, new_n459, new_n462);
or_8   g00086(new_n462, new_n461, new_n463);
and_8  g00087(new_n463, new_n458, new_n464);
xor_4  g00088(new_n464, new_n457, new_n465);
xor_4  g00089(new_n465, new_n438, new_n466);
and_8  g00090(n5305, n4005, new_n467);
xor_4  g00091(new_n437, new_n415, new_n468);
and_8  g00092(new_n468, new_n467, new_n469);
or_8   g00093(new_n468, new_n467, new_n470);
xnor_4 g00094(new_n433, new_n431, new_n471);
xor_4  g00095(new_n424, new_n423, new_n472);
and_8  g00096(n6038, n5964, new_n473);
and_8  g00097(n5305, n2509, new_n474);
nand_5 g00098(new_n474, new_n473, new_n475);
or_8   g00099(new_n475, new_n472, new_n476);
or_8   g00100(new_n476, new_n471, new_n477);
xor_4  g00101(new_n435, new_n421, new_n478);
or_8   g00102(new_n478, new_n477, new_n479);
not_8  g00103(new_n479, new_n480);
and_8  g00104(new_n480, new_n470, new_n481);
or_8   g00105(new_n481, new_n469, new_n482);
xor_4  g00106(new_n482, new_n466, new_n483);
and_8  g00107(n8759, n5105, new_n484);
and_8  g00108(n12299, n7354, new_n485);
and_8  g00109(n8759, n1209, new_n486);
or_8   g00110(new_n486, new_n485, new_n487);
and_8  g00111(new_n486, new_n485, new_n488);
and_8  g00112(n7500, n6776, new_n489);
or_8   g00113(new_n489, new_n488, new_n490);
and_8  g00114(new_n490, new_n487, new_n491);
xor_4  g00115(new_n491, new_n484, new_n492);
nand_5 g00116(n12299, n7500, new_n493);
and_8  g00117(n7436, n7354, new_n494);
and_8  g00118(n6776, n1209, new_n495);
xnor_4 g00119(new_n495, new_n494, new_n496);
xor_4  g00120(new_n496, new_n493, new_n497);
and_8  g00121(new_n497, new_n492, new_n498);
nor_6  g00122(new_n497, new_n492, new_n499);
or_8   g00123(new_n499, new_n498, new_n500);
and_8  g00124(n8759, n7354, new_n501);
not_8  g00125(new_n501, new_n502);
and_8  g00126(new_n502, new_n489, new_n503_1);
nor_6  g00127(new_n503_1, new_n487, new_n504);
or_8   g00128(new_n504, new_n488, new_n505);
nand_5 g00129(new_n505, new_n489, new_n506);
or_8   g00130(new_n506, new_n500, new_n507);
not_8  g00131(new_n507, new_n508);
nand_5 g00132(n8759, n4141, new_n509);
and_8  g00133(n6776, n5105, new_n510);
or_8   g00134(new_n495, new_n494, new_n511);
and_8  g00135(n12299, n7500, new_n512);
or_8   g00136(new_n496, new_n512, new_n513);
and_8  g00137(new_n513, new_n511, new_n514);
and_8  g00138(new_n514, new_n510, new_n515);
nor_6  g00139(new_n514, new_n510, new_n516);
or_8   g00140(new_n516, new_n515, new_n517);
and_8  g00141(n7500, n7436, new_n518);
and_8  g00142(n12299, n1209, new_n519);
and_8  g00143(n8276, n7354, new_n520);
xnor_4 g00144(new_n520, new_n519, new_n521_1);
xor_4  g00145(new_n521_1, new_n518, new_n522);
nor_6  g00146(new_n522, new_n517, new_n523);
and_8  g00147(new_n522, new_n517, new_n524);
or_8   g00148(new_n524, new_n523, new_n525);
or_8   g00149(new_n525, new_n509, new_n526);
not_8  g00150(new_n526, new_n527);
and_8  g00151(new_n525, new_n509, new_n528);
or_8   g00152(new_n528, new_n527, new_n529);
and_8  g00153(new_n491, new_n484, new_n530);
or_8   g00154(new_n498, new_n530, new_n531);
not_8  g00155(new_n531, new_n532);
xor_4  g00156(new_n532, new_n529, new_n533_1);
and_8  g00157(new_n533_1, new_n508, new_n534);
and_8  g00158(n8759, n4928, new_n535);
and_8  g00159(n7436, n1209, new_n536);
and_8  g00160(n8276, n7500, new_n537);
and_8  g00161(n9241, n7354, new_n538);
xor_4  g00162(new_n538, new_n537, new_n539);
xor_4  g00163(new_n539, new_n536, new_n540);
or_8   g00164(new_n520, new_n519, new_n541);
or_8   g00165(new_n521_1, new_n518, new_n542);
and_8  g00166(new_n542, new_n541, new_n543);
xor_4  g00167(new_n543, new_n540, new_n544);
and_8  g00168(n6776, n4141, new_n545);
and_8  g00169(n12299, n5105, new_n546);
xor_4  g00170(new_n546, new_n545, new_n547);
xor_4  g00171(new_n547, new_n544, new_n548);
or_8   g00172(new_n523, new_n515, new_n549);
and_8  g00173(new_n549, new_n548, new_n550);
nor_6  g00174(new_n549, new_n548, new_n551);
or_8   g00175(new_n551, new_n550, new_n552);
or_8   g00176(new_n532, new_n529, new_n553);
and_8  g00177(new_n553, new_n526, new_n554);
xor_4  g00178(new_n554, new_n552, new_n555);
and_8  g00179(new_n555, new_n535, new_n556);
not_8  g00180(new_n535, new_n557);
not_8  g00181(new_n552, new_n558);
xor_4  g00182(new_n554, new_n558, new_n559);
and_8  g00183(new_n559, new_n557, new_n560);
or_8   g00184(new_n560, new_n556, new_n561);
xor_4  g00185(new_n561, new_n534, new_n562);
xor_4  g00186(new_n533_1, new_n508, new_n563);
xor_4  g00187(new_n506, new_n500, new_n564);
and_8  g00188(n5331, n1564, new_n565);
and_8  g00189(n8028, n7965, new_n566);
xor_4  g00190(new_n566, new_n565, new_n567);
and_8  g00191(new_n567, new_n501, new_n568);
and_8  g00192(n7354, n6776, new_n569);
and_8  g00193(n8759, n7500, new_n570);
xor_4  g00194(new_n570, new_n569, new_n571);
nor_6  g00195(new_n571, new_n568, new_n572);
and_8  g00196(new_n566, new_n565, new_n573);
and_8  g00197(n5331, n1512, new_n574);
and_8  g00198(n8476, n1564, new_n575);
xor_4  g00199(new_n575, new_n574, new_n576);
xor_4  g00200(new_n576, new_n573, new_n577);
and_8  g00201(n8028, n7388, new_n578);
and_8  g00202(n10848, n7965, new_n579);
xor_4  g00203(new_n579, new_n578, new_n580);
nor_6  g00204(new_n580, new_n577, new_n581);
and_8  g00205(new_n580, new_n577, new_n582);
or_8   g00206(new_n582, new_n581, new_n583);
xor_4  g00207(new_n571, new_n568, new_n584);
and_8  g00208(new_n584, new_n583, new_n585);
or_8   g00209(new_n585, new_n572, new_n586);
not_8  g00210(new_n586, new_n587);
and_8  g00211(new_n503_1, new_n487, new_n588);
nor_6  g00212(new_n588, new_n505, new_n589);
or_8   g00213(new_n589, new_n587, new_n590);
not_8  g00214(n7388, new_n591);
not_8  g00215(n10848, new_n592);
or_8   g00216(new_n592, new_n591, new_n593);
or_8   g00217(new_n593, new_n566, new_n594);
and_8  g00218(n11892, n8028, new_n595);
and_8  g00219(n7965, n1980, new_n596);
nor_6  g00220(new_n596, new_n595, new_n597);
and_8  g00221(n11892, n1980, new_n598);
and_8  g00222(new_n598, new_n566, new_n599);
or_8   g00223(new_n599, new_n597, new_n600);
and_8  g00224(new_n600, new_n594, new_n601);
nor_6  g00225(new_n597, new_n594, new_n602);
or_8   g00226(new_n602, new_n601, new_n603);
and_8  g00227(n8476, n1512, new_n604);
not_8  g00228(new_n604, new_n605);
or_8   g00229(new_n605, new_n565, new_n606);
and_8  g00230(n2530, n1564, new_n607);
and_8  g00231(n5331, n533, new_n608);
or_8   g00232(new_n608, new_n607, new_n609);
not_8  g00233(new_n609, new_n610);
and_8  g00234(new_n610, new_n606, new_n611);
and_8  g00235(new_n608, new_n607, new_n612);
or_8   g00236(new_n612, new_n611, new_n613);
nor_6  g00237(new_n610, new_n606, new_n614);
or_8   g00238(new_n614, new_n613, new_n615_1);
xor_4  g00239(new_n615_1, new_n603, new_n616);
and_8  g00240(new_n576, new_n573, new_n617);
or_8   g00241(new_n582, new_n617, new_n618);
xor_4  g00242(new_n618, new_n616, new_n619);
xor_4  g00243(new_n589, new_n586, new_n620);
or_8   g00244(new_n620, new_n619, new_n621);
and_8  g00245(new_n621, new_n590, new_n622);
or_8   g00246(new_n622, new_n564, new_n623);
and_8  g00247(n5331, n2802, new_n624);
or_8   g00248(new_n612, new_n604, new_n625);
and_8  g00249(new_n625, new_n609, new_n626);
xor_4  g00250(new_n626, new_n624, new_n627);
and_8  g00251(n2530, n1512, new_n628);
and_8  g00252(n12648, n1564, new_n629);
and_8  g00253(n8476, n533, new_n630);
nor_6  g00254(new_n630, new_n629, new_n631);
and_8  g00255(new_n630, new_n629, new_n632);
or_8   g00256(new_n632, new_n631, new_n633);
and_8  g00257(new_n633, new_n628, new_n634);
nor_6  g00258(new_n633, new_n628, new_n635);
or_8   g00259(new_n635, new_n634, new_n636);
xor_4  g00260(new_n636, new_n627, new_n637);
and_8  g00261(new_n613, new_n604, new_n638);
xor_4  g00262(new_n638, new_n637, new_n639);
and_8  g00263(n7965, n7294, new_n640);
or_8   g00264(new_n596, new_n595, new_n641);
and_8  g00265(n10848, n7388, new_n642);
or_8   g00266(new_n599, new_n642, new_n643);
and_8  g00267(new_n643, new_n641, new_n644);
xor_4  g00268(new_n644, new_n640, new_n645);
and_8  g00269(n11892, n10848, new_n646);
and_8  g00270(n7388, n1980, new_n647);
and_8  g00271(n8028, n2393, new_n648);
xor_4  g00272(new_n648, new_n647, new_n649);
xor_4  g00273(new_n649, new_n646, new_n650);
and_8  g00274(new_n650, new_n645, new_n651);
nor_6  g00275(new_n650, new_n645, new_n652);
or_8   g00276(new_n652, new_n651, new_n653);
nand_5 g00277(new_n601, new_n642, new_n654);
nor_6  g00278(new_n654, new_n653, new_n655);
and_8  g00279(new_n654, new_n653, new_n656);
or_8   g00280(new_n656, new_n655, new_n657);
xor_4  g00281(new_n657, new_n639, new_n658_1);
nor_6  g00282(new_n615_1, new_n603, new_n659);
and_8  g00283(new_n618, new_n616, new_n660);
or_8   g00284(new_n660, new_n659, new_n661);
not_8  g00285(new_n661, new_n662);
xor_4  g00286(new_n662, new_n658_1, new_n663);
and_8  g00287(new_n506, new_n500, new_n664);
or_8   g00288(new_n664, new_n508, new_n665);
xor_4  g00289(new_n622, new_n665, new_n666);
or_8   g00290(new_n666, new_n663, new_n667);
and_8  g00291(new_n667, new_n623, new_n668);
or_8   g00292(new_n668, new_n563, new_n669);
and_8  g00293(new_n644, new_n640, new_n670);
or_8   g00294(new_n651, new_n670, new_n671_1);
and_8  g00295(n12704, n7965, new_n672);
and_8  g00296(n7388, n7294, new_n673);
or_8   g00297(new_n648, new_n647, new_n674);
and_8  g00298(new_n648, new_n647, new_n675);
or_8   g00299(new_n675, new_n646, new_n676);
and_8  g00300(new_n676, new_n674, new_n677);
xor_4  g00301(new_n677, new_n673, new_n678);
and_8  g00302(n10848, n2393, new_n679);
and_8  g00303(n8028, n5860, new_n680);
xor_4  g00304(new_n680, new_n598, new_n681);
xor_4  g00305(new_n681, new_n679, new_n682);
xor_4  g00306(new_n682, new_n678, new_n683);
or_8   g00307(new_n683, new_n672, new_n684);
not_8  g00308(new_n672, new_n685);
and_8  g00309(new_n682, new_n678, new_n686);
nor_6  g00310(new_n682, new_n678, new_n687);
or_8   g00311(new_n687, new_n686, new_n688);
or_8   g00312(new_n688, new_n685, new_n689);
and_8  g00313(new_n689, new_n684, new_n690);
xor_4  g00314(new_n690, new_n671_1, new_n691);
xor_4  g00315(new_n691, new_n655, new_n692);
nand_5 g00316(new_n638, new_n637, new_n693);
not_8  g00317(new_n693, new_n694);
not_8  g00318(n5331, new_n695);
not_8  g00319(n6806, new_n696);
or_8   g00320(new_n696, new_n695, new_n697);
and_8  g00321(n8476, n2802, new_n698);
nor_6  g00322(new_n635, new_n631, new_n699);
xor_4  g00323(new_n699, new_n698, new_n700);
not_8  g00324(n1512, new_n701);
not_8  g00325(n12648, new_n702);
or_8   g00326(new_n702, new_n701, new_n703);
and_8  g00327(n2530, n533, new_n704);
and_8  g00328(n10545, n1564, new_n705);
xnor_4 g00329(new_n705, new_n704, new_n706);
xor_4  g00330(new_n706, new_n703, new_n707);
and_8  g00331(new_n707, new_n700, new_n708);
or_8   g00332(new_n635, new_n631, new_n709);
xor_4  g00333(new_n709, new_n698, new_n710);
and_8  g00334(n12648, n1512, new_n711);
xor_4  g00335(new_n706, new_n711, new_n712);
and_8  g00336(new_n712, new_n710, new_n713);
or_8   g00337(new_n713, new_n708, new_n714);
nor_6  g00338(new_n714, new_n697, new_n715);
and_8  g00339(new_n714, new_n697, new_n716);
or_8   g00340(new_n716, new_n715, new_n717);
and_8  g00341(new_n626, new_n624, new_n718);
and_8  g00342(new_n636, new_n627, new_n719);
or_8   g00343(new_n719, new_n718, new_n720);
not_8  g00344(new_n720, new_n721);
or_8   g00345(new_n721, new_n717, new_n722);
xor_4  g00346(new_n714, new_n697, new_n723);
or_8   g00347(new_n720, new_n723, new_n724);
and_8  g00348(new_n724, new_n722, new_n725);
and_8  g00349(new_n725, new_n694, new_n726);
and_8  g00350(new_n720, new_n723, new_n727);
and_8  g00351(new_n721, new_n717, new_n728);
or_8   g00352(new_n728, new_n727, new_n729);
and_8  g00353(new_n729, new_n693, new_n730);
or_8   g00354(new_n730, new_n726, new_n731);
nor_6  g00355(new_n636, new_n627, new_n732);
or_8   g00356(new_n732, new_n719, new_n733);
xor_4  g00357(new_n638, new_n733, new_n734);
and_8  g00358(new_n657, new_n734, new_n735);
xor_4  g00359(new_n657, new_n734, new_n736);
and_8  g00360(new_n662, new_n736, new_n737);
or_8   g00361(new_n737, new_n735, new_n738);
or_8   g00362(new_n738, new_n731, new_n739);
or_8   g00363(new_n729, new_n693, new_n740);
or_8   g00364(new_n725, new_n694, new_n741);
and_8  g00365(new_n741, new_n740, new_n742);
not_8  g00366(new_n735, new_n743);
or_8   g00367(new_n661, new_n658_1, new_n744);
and_8  g00368(new_n744, new_n743, new_n745);
or_8   g00369(new_n745, new_n742, new_n746);
and_8  g00370(new_n746, new_n739, new_n747);
xor_4  g00371(new_n747, new_n692, new_n748);
xor_4  g00372(new_n533_1, new_n507, new_n749);
not_8  g00373(new_n623, new_n750);
xor_4  g00374(new_n662, new_n736, new_n751);
xor_4  g00375(new_n622, new_n564, new_n752);
and_8  g00376(new_n752, new_n751, new_n753_1);
or_8   g00377(new_n753_1, new_n750, new_n754);
and_8  g00378(new_n754, new_n749, new_n755);
and_8  g00379(new_n668, new_n563, new_n756);
or_8   g00380(new_n756, new_n755, new_n757);
or_8   g00381(new_n757, new_n748, new_n758);
and_8  g00382(new_n758, new_n669, new_n759);
xor_4  g00383(new_n759, new_n562, new_n760);
and_8  g00384(new_n738, new_n731, new_n761);
not_8  g00385(new_n692, new_n762);
and_8  g00386(new_n747, new_n762, new_n763);
nor_6  g00387(new_n763, new_n761, new_n764);
and_8  g00388(n5331, n5069, new_n765);
not_8  g00389(new_n765, new_n766);
and_8  g00390(n12648, n533, new_n767);
and_8  g00391(n10545, n1512, new_n768);
and_8  g00392(n7690, n1564, new_n769);
xor_4  g00393(new_n769, new_n768, new_n770);
xor_4  g00394(new_n770, new_n767, new_n771);
or_8   g00395(new_n705, new_n704, new_n772);
or_8   g00396(new_n706, new_n711, new_n773);
and_8  g00397(new_n773, new_n772, new_n774);
and_8  g00398(new_n774, new_n771, new_n775);
nor_6  g00399(new_n774, new_n771, new_n776);
or_8   g00400(new_n776, new_n775, new_n777);
and_8  g00401(n8476, n6806, new_n778);
and_8  g00402(n2802, n2530, new_n779);
xor_4  g00403(new_n779, new_n778, new_n780);
not_8  g00404(new_n780, new_n781);
or_8   g00405(new_n781, new_n777, new_n782);
xor_4  g00406(new_n774, new_n771, new_n783_1);
or_8   g00407(new_n780, new_n783_1, new_n784);
and_8  g00408(new_n784, new_n782, new_n785);
and_8  g00409(new_n699, new_n698, new_n786);
or_8   g00410(new_n708, new_n786, new_n787);
and_8  g00411(new_n787, new_n785, new_n788);
nor_6  g00412(new_n787, new_n785, new_n789);
or_8   g00413(new_n789, new_n788, new_n790);
not_8  g00414(new_n790, new_n791);
or_8   g00415(new_n727, new_n715, new_n792);
and_8  g00416(new_n792, new_n791, new_n793);
not_8  g00417(new_n715, new_n794);
and_8  g00418(new_n722, new_n794, new_n795);
and_8  g00419(new_n795, new_n790, new_n796);
or_8   g00420(new_n796, new_n793, new_n797);
or_8   g00421(new_n797, new_n766, new_n798);
or_8   g00422(new_n795, new_n790, new_n799);
or_8   g00423(new_n792, new_n791, new_n800);
and_8  g00424(new_n800, new_n799, new_n801);
or_8   g00425(new_n801, new_n765, new_n802);
and_8  g00426(new_n802, new_n798, new_n803);
xor_4  g00427(new_n803, new_n726, new_n804);
and_8  g00428(new_n804, new_n764, new_n805);
or_8   g00429(new_n763, new_n761, new_n806_1);
xor_4  g00430(new_n803, new_n740, new_n807);
and_8  g00431(new_n807, new_n806_1, new_n808);
or_8   g00432(new_n808, new_n805, new_n809);
nand_5 g00433(new_n691, new_n655, new_n810);
and_8  g00434(n7965, n5814, new_n811);
and_8  g00435(n2393, n1980, new_n812);
and_8  g00436(n8028, n3986, new_n813);
and_8  g00437(n10848, n5860, new_n814);
xor_4  g00438(new_n814, new_n813, new_n815);
xor_4  g00439(new_n815, new_n812, new_n816);
or_8   g00440(new_n680, new_n598, new_n817);
and_8  g00441(new_n680, new_n598, new_n818);
or_8   g00442(new_n818, new_n679, new_n819);
and_8  g00443(new_n819, new_n817, new_n820);
xor_4  g00444(new_n820, new_n816, new_n821);
and_8  g00445(n12704, n7388, new_n822);
and_8  g00446(n11892, n7294, new_n823);
xor_4  g00447(new_n823, new_n822, new_n824);
xor_4  g00448(new_n824, new_n821, new_n825);
and_8  g00449(new_n677, new_n673, new_n826);
or_8   g00450(new_n686, new_n826, new_n827);
xor_4  g00451(new_n827, new_n825, new_n828);
not_8  g00452(new_n684, new_n829);
not_8  g00453(new_n671_1, new_n830);
and_8  g00454(new_n689, new_n830, new_n831);
nor_6  g00455(new_n831, new_n829, new_n832);
xor_4  g00456(new_n832, new_n828, new_n833);
xor_4  g00457(new_n833, new_n811, new_n834);
or_8   g00458(new_n834, new_n810, new_n835);
not_8  g00459(new_n810, new_n836);
and_8  g00460(new_n833, new_n811, new_n837_1);
nor_6  g00461(new_n833, new_n811, new_n838);
or_8   g00462(new_n838, new_n837_1, new_n839);
or_8   g00463(new_n839, new_n836, new_n840);
and_8  g00464(new_n840, new_n835, new_n841);
xor_4  g00465(new_n841, new_n809, new_n842);
and_8  g00466(new_n842, new_n760, new_n843);
not_8  g00467(new_n534, new_n844_1);
xor_4  g00468(new_n561, new_n844_1, new_n845);
xor_4  g00469(new_n759, new_n845, new_n846);
or_8   g00470(new_n807, new_n806_1, new_n847);
or_8   g00471(new_n804, new_n764, new_n848);
and_8  g00472(new_n848, new_n847, new_n849);
xor_4  g00473(new_n841, new_n849, new_n850);
and_8  g00474(new_n850, new_n846, new_n851);
or_8   g00475(new_n851, new_n843, new_n852);
xor_4  g00476(new_n468, new_n467, new_n853);
xor_4  g00477(new_n853, new_n480, new_n854);
and_8  g00478(new_n854, new_n852, new_n855);
xnor_4 g00479(new_n478, new_n477, new_n856);
xor_4  g00480(new_n757, new_n748, new_n857);
nor_6  g00481(new_n857, new_n856, new_n858);
and_8  g00482(new_n857, new_n856, new_n859);
or_8   g00483(new_n859, new_n858, new_n860);
xnor_4 g00484(new_n476, new_n471, new_n861);
xor_4  g00485(new_n752, new_n751, new_n862);
nor_6  g00486(new_n862, new_n861, new_n863);
xor_4  g00487(new_n620, new_n619, new_n864);
not_8  g00488(new_n472, new_n865);
and_8  g00489(n6038, n5305, new_n866);
not_8  g00490(new_n866, new_n867);
nand_5 g00491(new_n867, new_n427, new_n868);
and_8  g00492(new_n868, new_n865, new_n869);
nand_5 g00493(new_n867, new_n428, new_n870);
not_8  g00494(new_n870, new_n871);
or_8   g00495(new_n871, new_n869, new_n872);
nand_5 g00496(new_n872, new_n864, new_n873);
xnor_4 g00497(new_n872, new_n864, new_n874);
xor_4  g00498(new_n567, new_n501, new_n875);
and_8  g00499(new_n875, new_n866, new_n876);
xor_4  g00500(new_n474, new_n473, new_n877);
or_8   g00501(new_n877, new_n876, new_n878);
xnor_4 g00502(new_n584, new_n583, new_n879);
xnor_4 g00503(new_n877, new_n876, new_n880);
or_8   g00504(new_n880, new_n879, new_n881);
and_8  g00505(new_n881, new_n878, new_n882);
or_8   g00506(new_n882, new_n874, new_n883);
and_8  g00507(new_n883, new_n873, new_n884);
xor_4  g00508(new_n862, new_n861, new_n885);
and_8  g00509(new_n885, new_n884, new_n886);
or_8   g00510(new_n886, new_n863, new_n887);
not_8  g00511(new_n887, new_n888);
nor_6  g00512(new_n888, new_n860, new_n889);
or_8   g00513(new_n889, new_n858, new_n890);
or_8   g00514(new_n850, new_n846, new_n891);
or_8   g00515(new_n842, new_n760, new_n892);
and_8  g00516(new_n892, new_n891, new_n893);
xor_4  g00517(new_n853, new_n479, new_n894);
or_8   g00518(new_n894, new_n893, new_n895);
or_8   g00519(new_n854, new_n852, new_n896);
and_8  g00520(new_n896, new_n895, new_n897);
and_8  g00521(new_n897, new_n890, new_n898);
or_8   g00522(new_n898, new_n855, new_n899);
or_8   g00523(new_n899, new_n483, new_n900);
not_8  g00524(new_n483, new_n901);
not_8  g00525(new_n858, new_n902);
or_8   g00526(new_n888, new_n860, new_n903);
and_8  g00527(new_n903, new_n902, new_n904);
and_8  g00528(new_n894, new_n893, new_n905);
or_8   g00529(new_n905, new_n855, new_n906);
or_8   g00530(new_n906, new_n904, new_n907);
and_8  g00531(new_n907, new_n895, new_n908);
or_8   g00532(new_n908, new_n901, new_n909);
and_8  g00533(new_n909, new_n900, new_n910);
or_8   g00534(new_n554, new_n552, new_n911_1);
nand_5 g00535(new_n539, new_n536, new_n912);
nand_5 g00536(new_n543, new_n540, new_n913);
and_8  g00537(new_n913, new_n912, new_n914);
and_8  g00538(n6776, n4928, new_n915);
and_8  g00539(n12299, n4141, new_n916);
and_8  g00540(n8759, n8236, new_n917);
xnor_4 g00541(new_n917, new_n916, new_n918);
xor_4  g00542(new_n918, new_n915, new_n919);
xor_4  g00543(new_n919, new_n914, new_n920);
and_8  g00544(new_n538, new_n537, new_n921);
and_8  g00545(n7436, n5105, new_n922);
xnor_4 g00546(new_n922, new_n921, new_n923);
and_8  g00547(n9241, n7500, new_n924);
and_8  g00548(n8276, n1209, new_n925);
and_8  g00549(n10510, n7354, new_n926);
xnor_4 g00550(new_n926, new_n925, new_n927);
xor_4  g00551(new_n927, new_n924, new_n928);
xor_4  g00552(new_n928, new_n923, new_n929);
xor_4  g00553(new_n929, new_n920, new_n930);
and_8  g00554(new_n547, new_n544, new_n931);
and_8  g00555(new_n546, new_n545, new_n932);
xor_4  g00556(new_n550, new_n932, new_n933);
or_8   g00557(new_n933, new_n931, new_n934);
and_8  g00558(new_n934, new_n930, new_n935);
not_8  g00559(new_n929, new_n936);
xor_4  g00560(new_n936, new_n920, new_n937);
nor_6  g00561(new_n933, new_n931, new_n938);
and_8  g00562(new_n938, new_n937, new_n939);
or_8   g00563(new_n939, new_n935, new_n940);
and_8  g00564(new_n940, new_n911_1, new_n941);
xor_4  g00565(new_n525, new_n509, new_n942);
and_8  g00566(new_n531, new_n942, new_n943);
or_8   g00567(new_n943, new_n527, new_n944);
and_8  g00568(new_n944, new_n558, new_n945);
or_8   g00569(new_n938, new_n937, new_n946);
or_8   g00570(new_n934, new_n930, new_n947);
and_8  g00571(new_n947, new_n946, new_n948);
and_8  g00572(new_n948, new_n945, new_n949);
or_8   g00573(new_n949, new_n941, new_n950);
or_8   g00574(new_n559, new_n557, new_n951);
or_8   g00575(new_n561, new_n844_1, new_n952);
and_8  g00576(new_n952, new_n951, new_n953);
xor_4  g00577(new_n953, new_n950, new_n954);
not_8  g00578(new_n954, new_n955);
and_8  g00579(new_n770, new_n767, new_n956);
nor_6  g00580(new_n775, new_n956, new_n957);
and_8  g00581(n8476, n5069, new_n958);
and_8  g00582(n6806, n2530, new_n959);
and_8  g00583(n12044, n5331, new_n960);
xnor_4 g00584(new_n960, new_n959, new_n961);
xor_4  g00585(new_n961, new_n958, new_n962);
xnor_4 g00586(new_n962, new_n957, new_n963);
and_8  g00587(new_n769, new_n768, new_n964);
and_8  g00588(n12648, n2802, new_n965);
xnor_4 g00589(new_n965, new_n964, new_n966);
and_8  g00590(n7690, n1512, new_n967);
and_8  g00591(n10545, n533, new_n968);
and_8  g00592(n3616, n1564, new_n969);
xnor_4 g00593(new_n969, new_n968, new_n970);
xor_4  g00594(new_n970, new_n967, new_n971);
xor_4  g00595(new_n971, new_n966, new_n972);
nor_6  g00596(new_n972, new_n963, new_n973);
and_8  g00597(new_n972, new_n963, new_n974);
or_8   g00598(new_n974, new_n973, new_n975);
not_8  g00599(new_n782, new_n976);
and_8  g00600(new_n779, new_n778, new_n977);
xor_4  g00601(new_n788, new_n977, new_n978);
or_8   g00602(new_n978, new_n976, new_n979);
and_8  g00603(new_n979, new_n975, new_n980);
nor_6  g00604(new_n979, new_n975, new_n981);
or_8   g00605(new_n981, new_n980, new_n982);
and_8  g00606(new_n982, new_n799, new_n983);
xor_4  g00607(new_n979, new_n975, new_n984);
and_8  g00608(new_n984, new_n793, new_n985);
nor_6  g00609(new_n985, new_n983, new_n986);
and_8  g00610(new_n797, new_n766, new_n987);
or_8   g00611(new_n987, new_n740, new_n988);
and_8  g00612(new_n988, new_n798, new_n989);
xor_4  g00613(new_n989, new_n986, new_n990);
and_8  g00614(new_n832, new_n828, new_n991);
and_8  g00615(new_n815, new_n812, new_n992_1);
and_8  g00616(new_n820, new_n816, new_n993);
nor_6  g00617(new_n993, new_n992_1, new_n994);
and_8  g00618(n7388, n5814, new_n995);
and_8  g00619(n12704, n11892, new_n996_1);
and_8  g00620(n7965, n4903, new_n997);
xnor_4 g00621(new_n997, new_n996_1, new_n998);
xor_4  g00622(new_n998, new_n995, new_n999);
xor_4  g00623(new_n999, new_n994, new_n1000);
and_8  g00624(new_n814, new_n813, new_n1001);
and_8  g00625(n7294, n2393, new_n1002);
xnor_4 g00626(new_n1002, new_n1001, new_n1003);
and_8  g00627(n10848, n3986, new_n1004);
and_8  g00628(n5860, n1980, new_n1005);
and_8  g00629(n8028, n5857, new_n1006);
xnor_4 g00630(new_n1006, new_n1005, new_n1007);
xor_4  g00631(new_n1007, new_n1004, new_n1008);
xor_4  g00632(new_n1008, new_n1003, new_n1009);
xor_4  g00633(new_n1009, new_n1000, new_n1010);
and_8  g00634(new_n824, new_n821, new_n1011);
and_8  g00635(new_n823, new_n822, new_n1012);
and_8  g00636(new_n827, new_n825, new_n1013);
xor_4  g00637(new_n1013, new_n1012, new_n1014);
or_8   g00638(new_n1014, new_n1011, new_n1015);
xor_4  g00639(new_n1015, new_n1010, new_n1016);
or_8   g00640(new_n1016, new_n991, new_n1017);
not_8  g00641(new_n991, new_n1018);
and_8  g00642(new_n1015, new_n1010, new_n1019);
nor_6  g00643(new_n1015, new_n1010, new_n1020_1);
or_8   g00644(new_n1020_1, new_n1019, new_n1021);
or_8   g00645(new_n1021, new_n1018, new_n1022);
and_8  g00646(new_n1022, new_n1017, new_n1023);
or_8   g00647(new_n833, new_n811, new_n1024);
or_8   g00648(new_n837_1, new_n836, new_n1025);
and_8  g00649(new_n1025, new_n1024, new_n1026);
nor_6  g00650(new_n1026, new_n1023, new_n1027);
and_8  g00651(new_n1026, new_n1023, new_n1028);
or_8   g00652(new_n1028, new_n1027, new_n1029);
or_8   g00653(new_n1029, new_n990, new_n1030);
or_8   g00654(new_n985, new_n983, new_n1031);
xor_4  g00655(new_n989, new_n1031, new_n1032);
xor_4  g00656(new_n1026, new_n1023, new_n1033);
or_8   g00657(new_n1033, new_n1032, new_n1034);
and_8  g00658(new_n1034, new_n1030, new_n1035);
or_8   g00659(new_n841, new_n808, new_n1036);
and_8  g00660(new_n1036, new_n847, new_n1037);
xor_4  g00661(new_n1037, new_n1035, new_n1038);
and_8  g00662(new_n1038, new_n955, new_n1039);
and_8  g00663(new_n1037, new_n1035, new_n1040);
nor_6  g00664(new_n1037, new_n1035, new_n1041);
or_8   g00665(new_n1041, new_n1040, new_n1042);
and_8  g00666(new_n1042, new_n954, new_n1043);
or_8   g00667(new_n1043, new_n1039, new_n1044);
nor_6  g00668(new_n759, new_n845, new_n1045);
or_8   g00669(new_n851, new_n1045, new_n1046);
or_8   g00670(new_n1046, new_n1044, new_n1047);
or_8   g00671(new_n1042, new_n954, new_n1048);
or_8   g00672(new_n1038, new_n955, new_n1049);
and_8  g00673(new_n1049, new_n1048, new_n1050);
not_8  g00674(new_n1046, new_n1051);
or_8   g00675(new_n1051, new_n1050, new_n1052);
and_8  g00676(new_n1052, new_n1047, new_n1053);
xor_4  g00677(new_n1053, new_n910, n226);
and_8  g00678(n5305, n4634, new_n1055);
and_8  g00679(n10223, n5305, new_n1056);
and_8  g00680(n7265, n1097, new_n1057);
or_8   g00681(new_n1057, new_n1056, new_n1058);
and_8  g00682(n7265, n5305, new_n1059);
and_8  g00683(n10223, n1097, new_n1060);
and_8  g00684(new_n1060, new_n1059, new_n1061);
and_8  g00685(n5964, n2879, new_n1062);
or_8   g00686(new_n1062, new_n1061, new_n1063);
and_8  g00687(new_n1063, new_n1058, new_n1064);
xor_4  g00688(new_n1064, new_n1055, new_n1065);
and_8  g00689(n2879, n1097, new_n1066);
and_8  g00690(n10223, n5964, new_n1067_1);
and_8  g00691(n7265, n4312, new_n1068);
xor_4  g00692(new_n1068, new_n1067_1, new_n1069);
xor_4  g00693(new_n1069, new_n1066, new_n1070);
xor_4  g00694(new_n1070, new_n1065, new_n1071);
not_8  g00695(new_n1059, new_n1072);
nand_5 g00696(new_n1062, new_n1072, new_n1073);
not_8  g00697(new_n1061, new_n1074);
nand_5 g00698(new_n1074, new_n1058, new_n1075);
nand_5 g00699(new_n1075, new_n1073, new_n1076);
not_8  g00700(new_n1076, new_n1077);
and_8  g00701(new_n1077, new_n1062, new_n1078);
xnor_4 g00702(new_n1078, new_n1071, new_n1079);
not_8  g00703(new_n1073, new_n1080);
and_8  g00704(new_n1080, new_n1058, new_n1081);
or_8   g00705(new_n1081, new_n1077, new_n1082);
and_8  g00706(n8759, n7946, new_n1083);
and_8  g00707(n5331, n2558, new_n1084);
and_8  g00708(n9763, n7965, new_n1085);
xor_4  g00709(new_n1085, new_n1084, new_n1086);
and_8  g00710(new_n1086, new_n1083, new_n1087);
and_8  g00711(n7946, n6776, new_n1088);
and_8  g00712(n8759, n2024, new_n1089);
xor_4  g00713(new_n1089, new_n1088, new_n1090);
nand_5 g00714(new_n1090, new_n1087, new_n1091);
and_8  g00715(new_n1085, new_n1084, new_n1092);
and_8  g00716(n9111, n7965, new_n1093);
and_8  g00717(n9763, n7388, new_n1094_1);
xor_4  g00718(new_n1094_1, new_n1093, new_n1095);
xor_4  g00719(new_n1095, new_n1092, new_n1096);
not_8  g00720(new_n1096, new_n1097_1);
and_8  g00721(n5331, n2498, new_n1098);
and_8  g00722(n8476, n2558, new_n1099);
xor_4  g00723(new_n1099, new_n1098, new_n1100);
xor_4  g00724(new_n1100, new_n1097_1, new_n1101);
xnor_4 g00725(new_n1090, new_n1087, new_n1102);
or_8   g00726(new_n1102, new_n1101, new_n1103);
and_8  g00727(new_n1103, new_n1091, new_n1104);
not_8  g00728(new_n1083, new_n1105);
and_8  g00729(n6776, n2024, new_n1106);
and_8  g00730(new_n1106, new_n1105, new_n1107);
and_8  g00731(n12299, n7946, new_n1108);
and_8  g00732(n9189, n8759, new_n1109);
xor_4  g00733(new_n1109, new_n1108, new_n1110);
or_8   g00734(new_n1110, new_n1107, new_n1111);
or_8   g00735(new_n1109, new_n1108, new_n1112);
nand_5 g00736(new_n1112, new_n1107, new_n1113);
and_8  g00737(new_n1113, new_n1111, new_n1114);
xor_4  g00738(new_n1114, new_n1104, new_n1115);
or_8   g00739(new_n1095, new_n1092, new_n1116);
or_8   g00740(new_n1100, new_n1097_1, new_n1117);
and_8  g00741(new_n1117, new_n1116, new_n1118);
not_8  g00742(n9111, new_n1119);
or_8   g00743(new_n1119, new_n591, new_n1120);
or_8   g00744(new_n1120, new_n1085, new_n1121);
and_8  g00745(n11892, n3342, new_n1122);
and_8  g00746(new_n1122, new_n1085, new_n1123);
and_8  g00747(n11892, n9763, new_n1124);
and_8  g00748(n7965, n3342, new_n1125);
nor_6  g00749(new_n1125, new_n1124, new_n1126);
or_8   g00750(new_n1126, new_n1123, new_n1127);
nand_5 g00751(new_n1127, new_n1121, new_n1128);
or_8   g00752(new_n1126, new_n1121, new_n1129);
and_8  g00753(new_n1129, new_n1128, new_n1130);
and_8  g00754(new_n1130, new_n1118, new_n1131);
nor_6  g00755(new_n1130, new_n1118, new_n1132);
or_8   g00756(new_n1132, new_n1131, new_n1133);
not_8  g00757(n2558, new_n1134);
or_8   g00758(new_n695, new_n1134, new_n1135);
and_8  g00759(n8476, n2498, new_n1136_1);
and_8  g00760(new_n1136_1, new_n1135, new_n1137);
and_8  g00761(n2558, n2530, new_n1138_1);
and_8  g00762(n5579, n5331, new_n1139);
nor_6  g00763(new_n1139, new_n1138_1, new_n1140);
nand_5 g00764(new_n1140, new_n1137, new_n1141);
and_8  g00765(n5579, n2530, new_n1142);
and_8  g00766(new_n1142, new_n1084, new_n1143);
or_8   g00767(new_n1143, new_n1140, new_n1144);
or_8   g00768(new_n1144, new_n1137, new_n1145);
and_8  g00769(new_n1145, new_n1141, new_n1146);
xor_4  g00770(new_n1146, new_n1133, new_n1147);
xor_4  g00771(new_n1147, new_n1115, new_n1148);
nor_6  g00772(new_n1148, new_n1082, new_n1149);
not_8  g00773(new_n1149, new_n1150);
xor_4  g00774(new_n1086, new_n1083, new_n1151);
and_8  g00775(new_n1151, new_n1059, new_n1152);
and_8  g00776(n7265, n5964, new_n1153);
and_8  g00777(n5305, n2879, new_n1154);
xor_4  g00778(new_n1154, new_n1153, new_n1155);
or_8   g00779(new_n1155, new_n1152, new_n1156);
xor_4  g00780(new_n1102, new_n1101, new_n1157);
xor_4  g00781(new_n1155, new_n1152, new_n1158);
not_8  g00782(new_n1158, new_n1159);
or_8   g00783(new_n1159, new_n1157, new_n1160);
nand_5 g00784(new_n1160, new_n1156, new_n1161);
and_8  g00785(new_n1148, new_n1082, new_n1162);
or_8   g00786(new_n1162, new_n1149, new_n1163);
or_8   g00787(new_n1163, new_n1161, new_n1164);
and_8  g00788(new_n1164, new_n1150, new_n1165);
nor_6  g00789(new_n1165, new_n1079, new_n1166);
and_8  g00790(new_n1165, new_n1079, new_n1167);
or_8   g00791(new_n1167, new_n1166, new_n1168);
and_8  g00792(n8759, n2522, new_n1169);
and_8  g00793(new_n1109, new_n1108, new_n1170);
or_8   g00794(new_n1170, new_n1106, new_n1171);
and_8  g00795(new_n1171, new_n1112, new_n1172);
xor_4  g00796(new_n1172, new_n1169, new_n1173);
and_8  g00797(n12299, n2024, new_n1174);
and_8  g00798(n7946, n7436, new_n1175);
and_8  g00799(n9189, n6776, new_n1176);
xor_4  g00800(new_n1176, new_n1175, new_n1177);
xor_4  g00801(new_n1177, new_n1174, new_n1178);
xnor_4 g00802(new_n1178, new_n1173, new_n1179);
nand_5 g00803(n6776, n2024, new_n1180);
or_8   g00804(new_n1111, new_n1180, new_n1181);
xor_4  g00805(new_n1181, new_n1179, new_n1182);
not_8  g00806(new_n1104, new_n1183);
or_8   g00807(new_n1114, new_n1183, new_n1184);
or_8   g00808(new_n1147, new_n1115, new_n1185);
and_8  g00809(new_n1185, new_n1184, new_n1186);
and_8  g00810(new_n1186, new_n1182, new_n1187);
nor_6  g00811(new_n1186, new_n1182, new_n1188);
or_8   g00812(new_n1188, new_n1187, new_n1189);
and_8  g00813(n5331, n521, new_n1190);
or_8   g00814(new_n1139, new_n1138_1, new_n1191);
or_8   g00815(new_n1143, new_n1136_1, new_n1192);
and_8  g00816(new_n1192, new_n1191, new_n1193);
xor_4  g00817(new_n1193, new_n1190, new_n1194);
and_8  g00818(n2530, n2498, new_n1195);
and_8  g00819(n12648, n2558, new_n1196);
and_8  g00820(n8476, n5579, new_n1197);
nor_6  g00821(new_n1197, new_n1196, new_n1198_1);
and_8  g00822(new_n1197, new_n1196, new_n1199_1);
or_8   g00823(new_n1199_1, new_n1198_1, new_n1200);
and_8  g00824(new_n1200, new_n1195, new_n1201);
nor_6  g00825(new_n1200, new_n1195, new_n1202);
or_8   g00826(new_n1202, new_n1201, new_n1203);
xor_4  g00827(new_n1203, new_n1194, new_n1204);
and_8  g00828(new_n1099, new_n1098, new_n1205);
and_8  g00829(new_n1144, new_n1205, new_n1206);
xor_4  g00830(new_n1206, new_n1204, new_n1207);
and_8  g00831(n7965, n806, new_n1208);
and_8  g00832(n9111, n7388, new_n1209_1);
or_8   g00833(new_n1125, new_n1124, new_n1210);
and_8  g00834(new_n1210, new_n1209_1, new_n1211);
or_8   g00835(new_n1211, new_n1123, new_n1212);
xor_4  g00836(new_n1212, new_n1208, new_n1213);
and_8  g00837(n11892, n9111, new_n1214);
and_8  g00838(n9763, n2393, new_n1215);
and_8  g00839(n7388, n3342, new_n1216);
nor_6  g00840(new_n1216, new_n1215, new_n1217);
and_8  g00841(new_n1216, new_n1215, new_n1218);
or_8   g00842(new_n1218, new_n1217, new_n1219);
and_8  g00843(new_n1219, new_n1214, new_n1220);
nor_6  g00844(new_n1219, new_n1214, new_n1221);
or_8   g00845(new_n1221, new_n1220, new_n1222);
and_8  g00846(new_n1222, new_n1213, new_n1223);
nor_6  g00847(new_n1222, new_n1213, new_n1224);
or_8   g00848(new_n1224, new_n1223, new_n1225);
or_8   g00849(new_n1128, new_n1120, new_n1226);
nor_6  g00850(new_n1226, new_n1225, new_n1227);
and_8  g00851(new_n1226, new_n1225, new_n1228);
or_8   g00852(new_n1228, new_n1227, new_n1229);
xor_4  g00853(new_n1229, new_n1207, new_n1230);
not_8  g00854(new_n1132, new_n1231);
not_8  g00855(new_n1146, new_n1232);
or_8   g00856(new_n1232, new_n1133, new_n1233);
and_8  g00857(new_n1233, new_n1231, new_n1234);
xor_4  g00858(new_n1234, new_n1230, new_n1235);
xor_4  g00859(new_n1235, new_n1189, new_n1236);
not_8  g00860(new_n1236, new_n1237);
xor_4  g00861(new_n1237, new_n1168, n381);
and_8  g00862(n7862, n6038, new_n1239);
and_8  g00863(n7354, n6877, new_n1240);
and_8  g00864(n4805, n1564, new_n1241);
and_8  g00865(n8028, n7236, new_n1242);
xor_4  g00866(new_n1242, new_n1241, new_n1243);
xor_4  g00867(new_n1243, new_n1240, new_n1244);
xor_4  g00868(new_n1244, new_n1239, n397);
and_8  g00869(n6687, n4370, new_n1246);
and_8  g00870(n11407, n4189, new_n1247);
and_8  g00871(n11877, n6687, new_n1248);
or_8   g00872(new_n1248, new_n1247, new_n1249);
and_8  g00873(new_n1248, new_n1247, new_n1250);
and_8  g00874(n5212, n2564, new_n1251);
or_8   g00875(new_n1251, new_n1250, new_n1252);
and_8  g00876(new_n1252, new_n1249, new_n1253);
xor_4  g00877(new_n1253, new_n1246, new_n1254);
and_8  g00878(n5212, n4189, new_n1255);
and_8  g00879(n11407, n6770, new_n1256);
and_8  g00880(n11877, n2564, new_n1257);
xnor_4 g00881(new_n1257, new_n1256, new_n1258);
xnor_4 g00882(new_n1258, new_n1255, new_n1259);
xor_4  g00883(new_n1259, new_n1254, new_n1260);
nand_5 g00884(n11407, n6687, new_n1261);
and_8  g00885(new_n1261, new_n1251, new_n1262);
nor_6  g00886(new_n1262, new_n1249, new_n1263);
or_8   g00887(new_n1263, new_n1250, new_n1264);
and_8  g00888(new_n1264, new_n1251, new_n1265);
xnor_4 g00889(new_n1265, new_n1260, new_n1266);
and_8  g00890(n12709, n8336, new_n1267);
and_8  g00891(n11222, n10990, new_n1268);
and_8  g00892(n12489, n12069, new_n1269_1);
xor_4  g00893(new_n1269_1, new_n1268, new_n1270);
and_8  g00894(new_n1270, new_n1267, new_n1271);
and_8  g00895(n11728, n8336, new_n1272);
and_8  g00896(n12709, n10928, new_n1273);
xor_4  g00897(new_n1273, new_n1272, new_n1274);
nor_6  g00898(new_n1274, new_n1271, new_n1275);
and_8  g00899(new_n1269_1, new_n1268, new_n1276);
and_8  g00900(n11222, n5760, new_n1277);
and_8  g00901(n11153, n10990, new_n1278);
xor_4  g00902(new_n1278, new_n1277, new_n1279);
xor_4  g00903(new_n1279, new_n1276, new_n1280);
and_8  g00904(n12069, n7159, new_n1281);
and_8  g00905(n12489, n12391, new_n1282);
xor_4  g00906(new_n1282, new_n1281, new_n1283);
xor_4  g00907(new_n1283, new_n1280, new_n1284);
xnor_4 g00908(new_n1274, new_n1271, new_n1285);
nor_6  g00909(new_n1285, new_n1284, new_n1286);
or_8   g00910(new_n1286, new_n1275, new_n1287);
not_8  g00911(new_n1287, new_n1288);
and_8  g00912(n11728, n10928, new_n1289);
not_8  g00913(new_n1289, new_n1290);
or_8   g00914(new_n1290, new_n1267, new_n1291);
and_8  g00915(n6986, n6429, new_n1292);
and_8  g00916(new_n1292, new_n1267, new_n1293);
nand_5 g00917(n12709, n6986, new_n1294);
nand_5 g00918(n8336, n6429, new_n1295);
and_8  g00919(new_n1295, new_n1294, new_n1296);
or_8   g00920(new_n1296, new_n1293, new_n1297);
nand_5 g00921(new_n1297, new_n1291, new_n1298);
or_8   g00922(new_n1296, new_n1291, new_n1299);
and_8  g00923(new_n1299, new_n1298, new_n1300);
xor_4  g00924(new_n1300, new_n1288, new_n1301);
and_8  g00925(n12391, n7159, new_n1302);
not_8  g00926(new_n1302, new_n1303);
or_8   g00927(new_n1303, new_n1269_1, new_n1304);
and_8  g00928(n12489, n7891, new_n1305);
and_8  g00929(n12777, n12069, new_n1306);
or_8   g00930(new_n1306, new_n1305, new_n1307);
not_8  g00931(new_n1307, new_n1308);
and_8  g00932(new_n1308, new_n1304, new_n1309);
and_8  g00933(new_n1306, new_n1305, new_n1310);
or_8   g00934(new_n1310, new_n1309, new_n1311);
nor_6  g00935(new_n1308, new_n1304, new_n1312);
or_8   g00936(new_n1312, new_n1311, new_n1313);
and_8  g00937(n11153, n5760, new_n1314);
not_8  g00938(new_n1314, new_n1315);
nor_6  g00939(new_n1315, new_n1268, new_n1316);
and_8  g00940(n10990, n5314, new_n1317);
and_8  g00941(n11222, n1478, new_n1318);
xor_4  g00942(new_n1318, new_n1317, new_n1319);
or_8   g00943(new_n1319, new_n1316, new_n1320);
not_8  g00944(new_n1320, new_n1321);
or_8   g00945(new_n1318, new_n1317, new_n1322);
and_8  g00946(new_n1322, new_n1316, new_n1323);
or_8   g00947(new_n1323, new_n1321, new_n1324);
nor_6  g00948(new_n1324, new_n1313, new_n1325);
and_8  g00949(new_n1324, new_n1313, new_n1326);
or_8   g00950(new_n1326, new_n1325, new_n1327);
and_8  g00951(new_n1279, new_n1276, new_n1328);
and_8  g00952(new_n1283, new_n1280, new_n1329);
or_8   g00953(new_n1329, new_n1328, new_n1330);
xor_4  g00954(new_n1330, new_n1327, new_n1331);
xor_4  g00955(new_n1331, new_n1301, new_n1332);
not_8  g00956(new_n1264, new_n1333_1);
nand_5 g00957(new_n1262, new_n1249, new_n1334);
and_8  g00958(new_n1334, new_n1333_1, new_n1335);
not_8  g00959(new_n1335, new_n1336);
nand_5 g00960(new_n1336, new_n1332, new_n1337);
xor_4  g00961(new_n1335, new_n1332, new_n1338);
not_8  g00962(new_n1261, new_n1339);
xor_4  g00963(new_n1270, new_n1267, new_n1340);
and_8  g00964(new_n1340, new_n1339, new_n1341);
and_8  g00965(n11407, n2564, new_n1342);
and_8  g00966(n6687, n5212, new_n1343);
xor_4  g00967(new_n1343, new_n1342, new_n1344);
or_8   g00968(new_n1344, new_n1341, new_n1345);
xnor_4 g00969(new_n1285, new_n1284, new_n1346);
xnor_4 g00970(new_n1344, new_n1341, new_n1347);
or_8   g00971(new_n1347, new_n1346, new_n1348);
and_8  g00972(new_n1348, new_n1345, new_n1349);
or_8   g00973(new_n1349, new_n1338, new_n1350);
and_8  g00974(new_n1350, new_n1337, new_n1351);
xor_4  g00975(new_n1351, new_n1266, new_n1352);
and_8  g00976(n8819, n8336, new_n1353_1);
and_8  g00977(n11728, n6986, new_n1354);
and_8  g00978(n10928, n6429, new_n1355);
and_8  g00979(n12709, n2226, new_n1356);
xor_4  g00980(new_n1356, new_n1355, new_n1357_1);
xor_4  g00981(new_n1357_1, new_n1354, new_n1358);
xor_4  g00982(new_n1358, new_n1353_1, new_n1359);
nor_6  g00983(new_n1296, new_n1290, new_n1360);
or_8   g00984(new_n1360, new_n1293, new_n1361);
xor_4  g00985(new_n1361, new_n1359, new_n1362);
not_8  g00986(new_n1298, new_n1363);
and_8  g00987(new_n1363, new_n1289, new_n1364);
xor_4  g00988(new_n1364, new_n1362, new_n1365);
and_8  g00989(n12069, n6254, new_n1366);
or_8   g00990(new_n1310, new_n1302, new_n1367);
and_8  g00991(new_n1367, new_n1307, new_n1368);
and_8  g00992(new_n1368, new_n1366, new_n1369);
nor_6  g00993(new_n1368, new_n1366, new_n1370);
or_8   g00994(new_n1370, new_n1369, new_n1371);
and_8  g00995(n12489, n7160, new_n1372);
and_8  g00996(n12777, n12391, new_n1373);
and_8  g00997(n7891, n7159, new_n1374);
nor_6  g00998(new_n1374, new_n1373, new_n1375);
and_8  g00999(new_n1374, new_n1373, new_n1376);
or_8   g01000(new_n1376, new_n1375, new_n1377);
xor_4  g01001(new_n1377, new_n1372, new_n1378);
xor_4  g01002(new_n1378, new_n1371, new_n1379);
and_8  g01003(new_n1311, new_n1302, new_n1380);
or_8   g01004(new_n1380, new_n1379, new_n1381);
nor_6  g01005(new_n1378, new_n1371, new_n1382);
and_8  g01006(new_n1378, new_n1371, new_n1383);
or_8   g01007(new_n1383, new_n1382, new_n1384);
nor_6  g01008(new_n1310, new_n1309, new_n1385);
or_8   g01009(new_n1385, new_n1303, new_n1386);
or_8   g01010(new_n1386, new_n1384, new_n1387);
and_8  g01011(new_n1387, new_n1381, new_n1388);
and_8  g01012(n11791, n11222, new_n1389);
and_8  g01013(new_n1318, new_n1317, new_n1390);
or_8   g01014(new_n1390, new_n1314, new_n1391);
and_8  g01015(new_n1391, new_n1322, new_n1392);
and_8  g01016(new_n1392, new_n1389, new_n1393);
nor_6  g01017(new_n1392, new_n1389, new_n1394);
or_8   g01018(new_n1394, new_n1393, new_n1395);
and_8  g01019(n5760, n5314, new_n1396);
and_8  g01020(n10990, n996, new_n1397);
and_8  g01021(n11153, n1478, new_n1398);
nor_6  g01022(new_n1398, new_n1397, new_n1399);
and_8  g01023(new_n1398, new_n1397, new_n1400);
or_8   g01024(new_n1400, new_n1399, new_n1401);
xor_4  g01025(new_n1401, new_n1396, new_n1402);
nor_6  g01026(new_n1402, new_n1395, new_n1403);
and_8  g01027(new_n1402, new_n1395, new_n1404);
or_8   g01028(new_n1404, new_n1403, new_n1405);
or_8   g01029(new_n1320, new_n1315, new_n1406);
or_8   g01030(new_n1406, new_n1405, new_n1407);
xor_4  g01031(new_n1402, new_n1395, new_n1408);
not_8  g01032(new_n1406, new_n1409);
or_8   g01033(new_n1409, new_n1408, new_n1410);
and_8  g01034(new_n1410, new_n1407, new_n1411);
and_8  g01035(new_n1411, new_n1388, new_n1412);
and_8  g01036(new_n1386, new_n1384, new_n1413);
and_8  g01037(new_n1380, new_n1379, new_n1414);
or_8   g01038(new_n1414, new_n1413, new_n1415);
and_8  g01039(new_n1409, new_n1408, new_n1416);
and_8  g01040(new_n1406, new_n1405, new_n1417);
or_8   g01041(new_n1417, new_n1416, new_n1418);
and_8  g01042(new_n1418, new_n1415, new_n1419);
or_8   g01043(new_n1419, new_n1412, new_n1420);
not_8  g01044(new_n1330, new_n1421);
nor_6  g01045(new_n1421, new_n1327, new_n1422);
or_8   g01046(new_n1422, new_n1325, new_n1423);
nor_6  g01047(new_n1423, new_n1420, new_n1424);
and_8  g01048(new_n1423, new_n1420, new_n1425);
or_8   g01049(new_n1425, new_n1424, new_n1426);
xor_4  g01050(new_n1426, new_n1365, new_n1427);
nor_6  g01051(new_n1300, new_n1288, new_n1428);
and_8  g01052(new_n1331, new_n1301, new_n1429);
or_8   g01053(new_n1429, new_n1428, new_n1430);
xor_4  g01054(new_n1430, new_n1427, new_n1431);
xor_4  g01055(new_n1431, new_n1352, n658);
and_8  g01056(n7862, n2585, new_n1433);
not_8  g01057(new_n1433, new_n1434);
and_8  g01058(n2508, n1333, new_n1435);
and_8  g01059(n11757, n6038, new_n1436);
and_8  g01060(n12720, n1333, new_n1437);
or_8   g01061(new_n1437, new_n1436, new_n1438);
and_8  g01062(new_n1437, new_n1436, new_n1439);
and_8  g01063(n3172, n2509, new_n1440);
or_8   g01064(new_n1440, new_n1439, new_n1441);
and_8  g01065(new_n1441, new_n1438, new_n1442);
xnor_4 g01066(new_n1442, new_n1435, new_n1443);
and_8  g01067(n11757, n2509, new_n1444);
and_8  g01068(n6038, n5240, new_n1445);
and_8  g01069(n12720, n3172, new_n1446);
xnor_4 g01070(new_n1446, new_n1445, new_n1447);
xor_4  g01071(new_n1447, new_n1444, new_n1448);
nor_6  g01072(new_n1448, new_n1443, new_n1449);
and_8  g01073(new_n1448, new_n1443, new_n1450);
or_8   g01074(new_n1450, new_n1449, new_n1451);
and_8  g01075(new_n1451, new_n1434, new_n1452);
xor_4  g01076(new_n1451, new_n1434, new_n1453);
and_8  g01077(n7862, n2508, new_n1454);
and_8  g01078(n2509, n1333, new_n1455);
and_8  g01079(n6038, n3172, new_n1456);
and_8  g01080(n12720, n7862, new_n1457);
or_8   g01081(new_n1457, new_n1456, new_n1458);
and_8  g01082(new_n1458, new_n1455, new_n1459);
and_8  g01083(new_n1457, new_n1456, new_n1460);
or_8   g01084(new_n1460, new_n1459, new_n1461);
and_8  g01085(new_n1461, new_n1454, new_n1462);
xor_4  g01086(new_n1461, new_n1454, new_n1463);
xor_4  g01087(new_n1437, new_n1436, new_n1464);
xor_4  g01088(new_n1464, new_n1440, new_n1465);
and_8  g01089(new_n1465, new_n1463, new_n1466);
or_8   g01090(new_n1466, new_n1462, new_n1467);
not_8  g01091(new_n1467, new_n1468);
and_8  g01092(new_n1468, new_n1453, new_n1469);
or_8   g01093(new_n1469, new_n1452, new_n1470);
and_8  g01094(n12720, n11757, new_n1471_1);
and_8  g01095(n5240, n2509, new_n1472);
and_8  g01096(n11821, n6038, new_n1473);
xor_4  g01097(new_n1473, new_n1472, new_n1474);
xor_4  g01098(new_n1474, new_n1471_1, new_n1475);
or_8   g01099(new_n1446, new_n1445, new_n1476);
or_8   g01100(new_n1447, new_n1444, new_n1477);
and_8  g01101(new_n1477, new_n1476, new_n1478_1);
xor_4  g01102(new_n1478_1, new_n1475, new_n1479);
and_8  g01103(new_n1442, new_n1435, new_n1480);
or_8   g01104(new_n1449, new_n1480, new_n1481);
and_8  g01105(n2585, n1333, new_n1482);
and_8  g01106(n3172, n2508, new_n1483);
xor_4  g01107(new_n1483, new_n1482, new_n1484);
or_8   g01108(new_n1484, new_n1481, new_n1485);
nor_6  g01109(new_n1449, new_n1480, new_n1486);
not_8  g01110(new_n1484, new_n1487);
or_8   g01111(new_n1487, new_n1486, new_n1488);
and_8  g01112(new_n1488, new_n1485, new_n1489);
and_8  g01113(new_n1489, new_n1479, new_n1490);
not_8  g01114(new_n1479, new_n1491);
and_8  g01115(new_n1487, new_n1486, new_n1492);
and_8  g01116(new_n1484, new_n1481, new_n1493);
or_8   g01117(new_n1493, new_n1492, new_n1494);
and_8  g01118(new_n1494, new_n1491, new_n1495);
or_8   g01119(new_n1495, new_n1490, new_n1496);
or_8   g01120(new_n1496, new_n1470, new_n1497);
and_8  g01121(new_n1483, new_n1482, new_n1498);
and_8  g01122(new_n1485, new_n1479, new_n1499);
xor_4  g01123(new_n1499, new_n1498, new_n1500);
nor_6  g01124(new_n1500, new_n1493, new_n1501);
and_8  g01125(new_n1473, new_n1472, new_n1502);
and_8  g01126(n11757, n2508, new_n1503);
xnor_4 g01127(new_n1503, new_n1502, new_n1504);
and_8  g01128(n11821, n2509, new_n1505);
and_8  g01129(n12720, n5240, new_n1506);
and_8  g01130(n9080, n6038, new_n1507);
xnor_4 g01131(new_n1507, new_n1506, new_n1508);
xor_4  g01132(new_n1508, new_n1505, new_n1509);
xnor_4 g01133(new_n1509, new_n1504, new_n1510_1);
and_8  g01134(new_n1474, new_n1471_1, new_n1511);
and_8  g01135(new_n1478_1, new_n1475, new_n1512_1);
or_8   g01136(new_n1512_1, new_n1511, new_n1513);
not_8  g01137(new_n1513, new_n1514);
and_8  g01138(n4005, n1333, new_n1515);
and_8  g01139(n3172, n2585, new_n1516);
and_8  g01140(n12706, n7862, new_n1517);
xnor_4 g01141(new_n1517, new_n1516, new_n1518);
xor_4  g01142(new_n1518, new_n1515, new_n1519);
xor_4  g01143(new_n1519, new_n1514, new_n1520);
xor_4  g01144(new_n1520, new_n1510_1, new_n1521);
or_8   g01145(new_n1521, new_n1501, new_n1522);
or_8   g01146(new_n1500, new_n1493, new_n1523_1);
not_8  g01147(new_n1521, new_n1524);
or_8   g01148(new_n1524, new_n1523_1, new_n1525);
and_8  g01149(new_n1525, new_n1522, new_n1526);
xor_4  g01150(new_n1526, new_n1497, new_n1527);
and_8  g01151(n7862, n4005, new_n1528);
not_8  g01152(new_n1452, new_n1529);
xor_4  g01153(new_n1451, new_n1433, new_n1530);
or_8   g01154(new_n1467, new_n1530, new_n1531);
and_8  g01155(new_n1531, new_n1529, new_n1532);
nor_6  g01156(new_n1495, new_n1490, new_n1533);
or_8   g01157(new_n1533, new_n1532, new_n1534);
and_8  g01158(new_n1534, new_n1497, new_n1535);
and_8  g01159(new_n1535, new_n1528, new_n1536);
not_8  g01160(new_n1536, new_n1537);
xnor_4 g01161(new_n1465, new_n1463, new_n1538);
xnor_4 g01162(new_n1457, new_n1456, new_n1539);
and_8  g01163(n6038, n1333, new_n1540);
and_8  g01164(n7862, n2509, new_n1541);
and_8  g01165(new_n1541, new_n1540, new_n1542);
and_8  g01166(new_n1542, new_n1539, new_n1543);
not_8  g01167(new_n1543, new_n1544);
or_8   g01168(new_n1544, new_n1538, new_n1545);
xor_4  g01169(new_n1467, new_n1530, new_n1546);
or_8   g01170(new_n1546, new_n1545, new_n1547);
nor_6  g01171(new_n1535, new_n1528, new_n1548);
or_8   g01172(new_n1548, new_n1536, new_n1549);
or_8   g01173(new_n1549, new_n1547, new_n1550);
and_8  g01174(new_n1550, new_n1537, new_n1551);
xor_4  g01175(new_n1551, new_n1527, new_n1552);
and_8  g01176(n6877, n5105, new_n1553);
and_8  g01177(n6877, n1209, new_n1554);
and_8  g01178(n7354, n2464, new_n1555);
and_8  g01179(new_n1555, new_n1554, new_n1556);
or_8   g01180(new_n1555, new_n1554, new_n1557);
and_8  g01181(n9400, n7500, new_n1558);
and_8  g01182(new_n1558, new_n1557, new_n1559);
or_8   g01183(new_n1559, new_n1556, new_n1560);
xor_4  g01184(new_n1560, new_n1553, new_n1561);
and_8  g01185(n7500, n2464, new_n1562);
and_8  g01186(n9400, n1209, new_n1563);
and_8  g01187(n11311, n7354, new_n1564_1);
xor_4  g01188(new_n1564_1, new_n1563, new_n1565);
xor_4  g01189(new_n1565, new_n1562, new_n1566);
xnor_4 g01190(new_n1566, new_n1561, new_n1567);
xnor_4 g01191(new_n1555, new_n1554, new_n1568);
and_8  g01192(n9400, n7354, new_n1569);
and_8  g01193(n7500, n6877, new_n1570);
and_8  g01194(new_n1570, new_n1569, new_n1571);
and_8  g01195(new_n1571, new_n1568, new_n1572);
not_8  g01196(new_n1572, new_n1573);
or_8   g01197(new_n1573, new_n1567, new_n1574);
nand_5 g01198(n11311, n7500, new_n1575);
and_8  g01199(n2464, n1209, new_n1576_1);
and_8  g01200(n7354, n4187, new_n1577);
xnor_4 g01201(new_n1577, new_n1576_1, new_n1578);
xor_4  g01202(new_n1578, new_n1575, new_n1579);
and_8  g01203(n9400, n5105, new_n1580);
or_8   g01204(new_n1564_1, new_n1563, new_n1581);
and_8  g01205(new_n1564_1, new_n1563, new_n1582);
or_8   g01206(new_n1582, new_n1562, new_n1583);
and_8  g01207(new_n1583, new_n1581, new_n1584);
xor_4  g01208(new_n1584, new_n1580, new_n1585);
xnor_4 g01209(new_n1585, new_n1579, new_n1586);
and_8  g01210(n6877, n4141, new_n1587);
and_8  g01211(new_n1560, new_n1553, new_n1588);
and_8  g01212(new_n1566, new_n1561, new_n1589);
or_8   g01213(new_n1589, new_n1588, new_n1590);
xor_4  g01214(new_n1590, new_n1587, new_n1591);
xor_4  g01215(new_n1591, new_n1586, new_n1592);
or_8   g01216(new_n1592, new_n1574, new_n1593);
and_8  g01217(n6877, n4928, new_n1594);
nor_6  g01218(new_n1590, new_n1587, new_n1595);
and_8  g01219(new_n1591, new_n1586, new_n1596);
or_8   g01220(new_n1596, new_n1595, new_n1597);
and_8  g01221(n11311, n1209, new_n1598);
and_8  g01222(n7500, n4187, new_n1599);
and_8  g01223(n7354, n4203, new_n1600);
xor_4  g01224(new_n1600, new_n1599, new_n1601);
xor_4  g01225(new_n1601, new_n1598, new_n1602);
or_8   g01226(new_n1577, new_n1576_1, new_n1603);
not_8  g01227(new_n1575, new_n1604);
or_8   g01228(new_n1578, new_n1604, new_n1605);
and_8  g01229(new_n1605, new_n1603, new_n1606);
xor_4  g01230(new_n1606, new_n1602, new_n1607);
not_8  g01231(new_n1607, new_n1608);
and_8  g01232(new_n1584, new_n1580, new_n1609);
and_8  g01233(new_n1585, new_n1579, new_n1610);
or_8   g01234(new_n1610, new_n1609, new_n1611);
and_8  g01235(n9400, n4141, new_n1612);
and_8  g01236(n5105, n2464, new_n1613);
xor_4  g01237(new_n1613, new_n1612, new_n1614);
or_8   g01238(new_n1614, new_n1611, new_n1615);
nor_6  g01239(new_n1610, new_n1609, new_n1616);
not_8  g01240(new_n1614, new_n1617);
or_8   g01241(new_n1617, new_n1616, new_n1618);
and_8  g01242(new_n1618, new_n1615, new_n1619);
xor_4  g01243(new_n1619, new_n1608, new_n1620);
or_8   g01244(new_n1620, new_n1597, new_n1621);
nor_6  g01245(new_n1596, new_n1595, new_n1622);
xor_4  g01246(new_n1619, new_n1607, new_n1623);
or_8   g01247(new_n1623, new_n1622, new_n1624);
and_8  g01248(new_n1624, new_n1621, new_n1625);
and_8  g01249(new_n1625, new_n1594, new_n1626);
nor_6  g01250(new_n1625, new_n1594, new_n1627);
or_8   g01251(new_n1627, new_n1626, new_n1628);
xor_4  g01252(new_n1628, new_n1593, new_n1629);
not_8  g01253(new_n1629, new_n1630);
and_8  g01254(n7294, n7236, new_n1631);
and_8  g01255(n10848, n3992, new_n1632);
and_8  g01256(n8384, n8028, new_n1633);
and_8  g01257(n7236, n1980, new_n1634);
or_8   g01258(new_n1634, new_n1633, new_n1635);
and_8  g01259(new_n1635, new_n1632, new_n1636);
and_8  g01260(new_n1634, new_n1633, new_n1637);
or_8   g01261(new_n1637, new_n1636, new_n1638);
xor_4  g01262(new_n1638, new_n1631, new_n1639);
and_8  g01263(n8028, n6358, new_n1640);
and_8  g01264(n10848, n8384, new_n1641);
and_8  g01265(n3992, n1980, new_n1642);
nor_6  g01266(new_n1642, new_n1641, new_n1643);
and_8  g01267(new_n1642, new_n1641, new_n1644);
or_8   g01268(new_n1644, new_n1643, new_n1645);
xnor_4 g01269(new_n1645, new_n1640, new_n1646);
and_8  g01270(new_n1646, new_n1639, new_n1647);
nor_6  g01271(new_n1646, new_n1639, new_n1648);
or_8   g01272(new_n1648, new_n1647, new_n1649);
xnor_4 g01273(new_n1634, new_n1633, new_n1650);
and_8  g01274(n10848, n7236, new_n1651);
and_8  g01275(n8028, n3992, new_n1652);
and_8  g01276(new_n1652, new_n1651, new_n1653);
nand_5 g01277(new_n1653, new_n1650, new_n1654);
or_8   g01278(new_n1654, new_n1649, new_n1655);
and_8  g01279(n10848, n6358, new_n1656);
not_8  g01280(new_n1656, new_n1657);
and_8  g01281(n8384, n1980, new_n1658_1);
and_8  g01282(n8028, n5198, new_n1659);
xnor_4 g01283(new_n1659, new_n1658_1, new_n1660);
xor_4  g01284(new_n1660, new_n1657, new_n1661);
not_8  g01285(new_n1661, new_n1662);
and_8  g01286(n7294, n3992, new_n1663);
or_8   g01287(new_n1642, new_n1641, new_n1664);
or_8   g01288(new_n1645, new_n1640, new_n1665);
and_8  g01289(new_n1665, new_n1664, new_n1666);
xor_4  g01290(new_n1666, new_n1663, new_n1667);
xor_4  g01291(new_n1667, new_n1662, new_n1668);
and_8  g01292(n12704, n7236, new_n1669);
and_8  g01293(new_n1638, new_n1631, new_n1670);
or_8   g01294(new_n1647, new_n1670, new_n1671);
xor_4  g01295(new_n1671, new_n1669, new_n1672);
xor_4  g01296(new_n1672, new_n1668, new_n1673);
or_8   g01297(new_n1673, new_n1655, new_n1674);
and_8  g01298(n7236, n5814, new_n1675);
not_8  g01299(new_n1675, new_n1676);
and_8  g01300(new_n1666, new_n1663, new_n1677);
and_8  g01301(new_n1667, new_n1661, new_n1678);
or_8   g01302(new_n1678, new_n1677, new_n1679);
and_8  g01303(n8384, n7294, new_n1680);
and_8  g01304(n12704, n3992, new_n1681);
xor_4  g01305(new_n1681, new_n1680, new_n1682);
and_8  g01306(new_n1682, new_n1679, new_n1683);
nor_6  g01307(new_n1682, new_n1679, new_n1684);
or_8   g01308(new_n1684, new_n1683, new_n1685);
and_8  g01309(n6358, n1980, new_n1686);
not_8  g01310(new_n1686, new_n1687);
or_8   g01311(new_n1659, new_n1658_1, new_n1688);
or_8   g01312(new_n1660, new_n1656, new_n1689);
and_8  g01313(new_n1689, new_n1688, new_n1690);
xor_4  g01314(new_n1690, new_n1687, new_n1691);
and_8  g01315(n10848, n5198, new_n1692);
and_8  g01316(n8028, n1471, new_n1693);
xor_4  g01317(new_n1693, new_n1692, new_n1694);
xor_4  g01318(new_n1694, new_n1691, new_n1695);
or_8   g01319(new_n1695, new_n1685, new_n1696);
xor_4  g01320(new_n1682, new_n1679, new_n1697);
not_8  g01321(new_n1694, new_n1698);
xor_4  g01322(new_n1698, new_n1691, new_n1699);
or_8   g01323(new_n1699, new_n1697, new_n1700);
and_8  g01324(new_n1700, new_n1696, new_n1701);
nor_6  g01325(new_n1671, new_n1669, new_n1702);
and_8  g01326(new_n1672, new_n1668, new_n1703);
nor_6  g01327(new_n1703, new_n1702, new_n1704);
and_8  g01328(new_n1704, new_n1701, new_n1705);
and_8  g01329(new_n1699, new_n1697, new_n1706);
and_8  g01330(new_n1695, new_n1685, new_n1707);
or_8   g01331(new_n1707, new_n1706, new_n1708);
or_8   g01332(new_n1703, new_n1702, new_n1709);
and_8  g01333(new_n1709, new_n1708, new_n1710);
or_8   g01334(new_n1710, new_n1705, new_n1711);
or_8   g01335(new_n1711, new_n1676, new_n1712);
or_8   g01336(new_n1709, new_n1708, new_n1713);
or_8   g01337(new_n1704, new_n1701, new_n1714);
and_8  g01338(new_n1714, new_n1713, new_n1715);
or_8   g01339(new_n1715, new_n1675, new_n1716);
and_8  g01340(new_n1716, new_n1712, new_n1717);
xor_4  g01341(new_n1717, new_n1674, new_n1718);
and_8  g01342(n4805, n2802, new_n1719);
and_8  g01343(n5283, n1564, new_n1720);
and_8  g01344(n4805, n533, new_n1721);
and_8  g01345(new_n1721, new_n1720, new_n1722);
or_8   g01346(new_n1721, new_n1720, new_n1723);
and_8  g01347(n11478, n1512, new_n1724);
and_8  g01348(new_n1724, new_n1723, new_n1725);
or_8   g01349(new_n1725, new_n1722, new_n1726);
xor_4  g01350(new_n1726, new_n1719, new_n1727);
and_8  g01351(n1564, n137, new_n1728);
and_8  g01352(n5283, n1512, new_n1729);
and_8  g01353(n11478, n533, new_n1730);
nor_6  g01354(new_n1730, new_n1729, new_n1731);
and_8  g01355(new_n1730, new_n1729, new_n1732);
or_8   g01356(new_n1732, new_n1731, new_n1733);
xnor_4 g01357(new_n1733, new_n1728, new_n1734);
and_8  g01358(new_n1734, new_n1727, new_n1735);
nor_6  g01359(new_n1734, new_n1727, new_n1736);
or_8   g01360(new_n1736, new_n1735, new_n1737);
xor_4  g01361(new_n1721, new_n1720, new_n1738);
and_8  g01362(n4805, n1512, new_n1739);
and_8  g01363(n11478, n1564, new_n1740);
nand_5 g01364(new_n1740, new_n1739, new_n1741);
or_8   g01365(new_n1741, new_n1738, new_n1742);
or_8   g01366(new_n1742, new_n1737, new_n1743);
and_8  g01367(n6806, n4805, new_n1744);
and_8  g01368(n11478, n2802, new_n1745);
or_8   g01369(new_n1730, new_n1729, new_n1746);
or_8   g01370(new_n1733, new_n1728, new_n1747);
and_8  g01371(new_n1747, new_n1746, new_n1748);
xor_4  g01372(new_n1748, new_n1745, new_n1749);
and_8  g01373(n1512, n137, new_n1750);
not_8  g01374(new_n1750, new_n1751);
and_8  g01375(n5283, n533, new_n1752);
and_8  g01376(n6294, n1564, new_n1753);
xor_4  g01377(new_n1753, new_n1752, new_n1754);
xor_4  g01378(new_n1754, new_n1751, new_n1755);
xor_4  g01379(new_n1755, new_n1749, new_n1756);
xor_4  g01380(new_n1756, new_n1744, new_n1757);
and_8  g01381(new_n1726, new_n1719, new_n1758);
or_8   g01382(new_n1735, new_n1758, new_n1759);
xor_4  g01383(new_n1759, new_n1757, new_n1760);
or_8   g01384(new_n1760, new_n1743, new_n1761);
and_8  g01385(n5069, n4805, new_n1762);
not_8  g01386(new_n1762, new_n1763);
and_8  g01387(n533, n137, new_n1764);
and_8  g01388(n6294, n1512, new_n1765);
and_8  g01389(n6797, n1564, new_n1766);
xor_4  g01390(new_n1766, new_n1765, new_n1767);
and_8  g01391(new_n1767, new_n1764, new_n1768);
nor_6  g01392(new_n1767, new_n1764, new_n1769);
or_8   g01393(new_n1769, new_n1768, new_n1770);
nor_6  g01394(new_n1753, new_n1752, new_n1771);
and_8  g01395(new_n1754, new_n1751, new_n1772);
or_8   g01396(new_n1772, new_n1771, new_n1773);
nor_6  g01397(new_n1773, new_n1770, new_n1774);
and_8  g01398(new_n1773, new_n1770, new_n1775);
or_8   g01399(new_n1775, new_n1774, new_n1776);
and_8  g01400(n11478, n6806, new_n1777);
and_8  g01401(n5283, n2802, new_n1778);
xor_4  g01402(new_n1778, new_n1777, new_n1779);
not_8  g01403(new_n1779, new_n1780);
or_8   g01404(new_n1780, new_n1776, new_n1781);
xor_4  g01405(new_n1773, new_n1770, new_n1782);
or_8   g01406(new_n1779, new_n1782, new_n1783);
and_8  g01407(new_n1783, new_n1781, new_n1784);
and_8  g01408(new_n1748, new_n1745, new_n1785);
not_8  g01409(new_n1755, new_n1786);
and_8  g01410(new_n1786, new_n1749, new_n1787);
or_8   g01411(new_n1787, new_n1785, new_n1788);
xor_4  g01412(new_n1788, new_n1784, new_n1789);
not_8  g01413(new_n1744, new_n1790);
and_8  g01414(new_n1756, new_n1790, new_n1791);
not_8  g01415(new_n1791, new_n1792);
or_8   g01416(new_n1759, new_n1757, new_n1793);
and_8  g01417(new_n1793, new_n1792, new_n1794);
and_8  g01418(new_n1794, new_n1789, new_n1795);
not_8  g01419(new_n1789, new_n1796);
xor_4  g01420(new_n1756, new_n1790, new_n1797);
not_8  g01421(new_n1759, new_n1798_1);
and_8  g01422(new_n1798_1, new_n1797, new_n1799);
or_8   g01423(new_n1799, new_n1791, new_n1800);
and_8  g01424(new_n1800, new_n1796, new_n1801);
or_8   g01425(new_n1801, new_n1795, new_n1802);
or_8   g01426(new_n1802, new_n1763, new_n1803);
or_8   g01427(new_n1800, new_n1796, new_n1804);
or_8   g01428(new_n1794, new_n1789, new_n1805);
and_8  g01429(new_n1805, new_n1804, new_n1806);
or_8   g01430(new_n1806, new_n1762, new_n1807);
and_8  g01431(new_n1807, new_n1803, new_n1808);
xor_4  g01432(new_n1808, new_n1761, new_n1809);
and_8  g01433(new_n1809, new_n1718, new_n1810);
not_8  g01434(new_n1674, new_n1811);
xor_4  g01435(new_n1717, new_n1811, new_n1812);
not_8  g01436(new_n1761, new_n1813);
xor_4  g01437(new_n1808, new_n1813, new_n1814);
and_8  g01438(new_n1814, new_n1812, new_n1815);
or_8   g01439(new_n1815, new_n1810, new_n1816);
xor_4  g01440(new_n1673, new_n1655, new_n1817);
xor_4  g01441(new_n1742, new_n1737, new_n1818);
xor_4  g01442(new_n1654, new_n1649, new_n1819);
or_8   g01443(new_n1819, new_n1818, new_n1820);
and_8  g01444(new_n1242, new_n1241, new_n1821);
xor_4  g01445(new_n1740, new_n1739, new_n1822);
or_8   g01446(new_n1822, new_n1821, new_n1823);
xnor_4 g01447(new_n1822, new_n1821, new_n1824);
xor_4  g01448(new_n1652, new_n1651, new_n1825);
or_8   g01449(new_n1825, new_n1824, new_n1826);
and_8  g01450(new_n1826, new_n1823, new_n1827);
not_8  g01451(new_n1241, new_n1828);
and_8  g01452(new_n1724, new_n1828, new_n1829);
or_8   g01453(new_n1829, new_n1738, new_n1830);
nand_5 g01454(new_n1725, new_n1828, new_n1831);
and_8  g01455(new_n1831, new_n1830, new_n1832);
or_8   g01456(new_n1832, new_n1827, new_n1833);
xnor_4 g01457(new_n1832, new_n1827, new_n1834);
not_8  g01458(new_n1242, new_n1835_1);
nand_5 g01459(new_n1632, new_n1835_1, new_n1836);
nand_5 g01460(new_n1836, new_n1650, new_n1837);
nand_5 g01461(new_n1636, new_n1835_1, new_n1838);
and_8  g01462(new_n1838, new_n1837, new_n1839);
or_8   g01463(new_n1839, new_n1834, new_n1840);
and_8  g01464(new_n1840, new_n1833, new_n1841);
not_8  g01465(new_n1820, new_n1842);
and_8  g01466(new_n1819, new_n1818, new_n1843);
or_8   g01467(new_n1843, new_n1842, new_n1844);
or_8   g01468(new_n1844, new_n1841, new_n1845);
and_8  g01469(new_n1845, new_n1820, new_n1846);
or_8   g01470(new_n1846, new_n1817, new_n1847_1);
xor_4  g01471(new_n1760, new_n1743, new_n1848);
nor_6  g01472(new_n1846, new_n1817, new_n1849);
and_8  g01473(new_n1846, new_n1817, new_n1850);
or_8   g01474(new_n1850, new_n1849, new_n1851);
or_8   g01475(new_n1851, new_n1848, new_n1852);
and_8  g01476(new_n1852, new_n1847_1, new_n1853);
or_8   g01477(new_n1853, new_n1816, new_n1854);
or_8   g01478(new_n1814, new_n1812, new_n1855);
or_8   g01479(new_n1809, new_n1718, new_n1856);
and_8  g01480(new_n1856, new_n1855, new_n1857);
not_8  g01481(new_n1848, new_n1858);
xor_4  g01482(new_n1846, new_n1817, new_n1859);
and_8  g01483(new_n1859, new_n1858, new_n1860);
or_8   g01484(new_n1860, new_n1849, new_n1861);
or_8   g01485(new_n1861, new_n1857, new_n1862);
and_8  g01486(new_n1862, new_n1854, new_n1863);
and_8  g01487(new_n1863, new_n1630, new_n1864);
and_8  g01488(new_n1861, new_n1857, new_n1865);
and_8  g01489(new_n1853, new_n1816, new_n1866);
or_8   g01490(new_n1866, new_n1865, new_n1867);
or_8   g01491(new_n1867, new_n1629, new_n1868);
or_8   g01492(new_n1863, new_n1630, new_n1869);
and_8  g01493(new_n1869, new_n1868, new_n1870);
xor_4  g01494(new_n1592, new_n1574, new_n1871);
not_8  g01495(new_n1871, new_n1872);
or_8   g01496(new_n1859, new_n1858, new_n1873);
and_8  g01497(new_n1873, new_n1852, new_n1874);
or_8   g01498(new_n1874, new_n1872, new_n1875);
and_8  g01499(new_n1851, new_n1848, new_n1876);
or_8   g01500(new_n1876, new_n1860, new_n1877);
and_8  g01501(new_n1877, new_n1871, new_n1878);
and_8  g01502(new_n1874, new_n1872, new_n1879);
or_8   g01503(new_n1879, new_n1878, new_n1880);
xor_4  g01504(new_n1572, new_n1567, new_n1881);
xor_4  g01505(new_n1844, new_n1841, new_n1882);
or_8   g01506(new_n1882, new_n1881, new_n1883);
not_8  g01507(new_n1883, new_n1884);
and_8  g01508(new_n1882, new_n1881, new_n1885);
or_8   g01509(new_n1885, new_n1884, new_n1886);
xor_4  g01510(new_n1839, new_n1834, new_n1887);
not_8  g01511(new_n1240, new_n1888);
and_8  g01512(new_n1558, new_n1888, new_n1889);
not_8  g01513(new_n1889, new_n1890);
or_8   g01514(new_n1890, new_n1557, new_n1891);
or_8   g01515(new_n1889, new_n1568, new_n1892);
and_8  g01516(new_n1892, new_n1891, new_n1893);
nor_6  g01517(new_n1893, new_n1887, new_n1894);
not_8  g01518(new_n1894, new_n1895);
and_8  g01519(new_n1893, new_n1887, new_n1896);
or_8   g01520(new_n1896, new_n1894, new_n1897);
xnor_4 g01521(new_n1825, new_n1824, new_n1898);
xor_4  g01522(new_n1570, new_n1569, new_n1899);
and_8  g01523(new_n1899, new_n1898, new_n1900);
nand_5 g01524(new_n1243, new_n1240, new_n1901);
not_8  g01525(new_n1901, new_n1902);
xor_4  g01526(new_n1899, new_n1898, new_n1903);
and_8  g01527(new_n1903, new_n1902, new_n1904);
or_8   g01528(new_n1904, new_n1900, new_n1905);
not_8  g01529(new_n1905, new_n1906_1);
or_8   g01530(new_n1906_1, new_n1897, new_n1907);
and_8  g01531(new_n1907, new_n1895, new_n1908);
or_8   g01532(new_n1908, new_n1886, new_n1909);
and_8  g01533(new_n1909, new_n1883, new_n1910);
or_8   g01534(new_n1910, new_n1880, new_n1911);
and_8  g01535(new_n1911, new_n1875, new_n1912);
and_8  g01536(new_n1912, new_n1870, new_n1913);
or_8   g01537(new_n1913, new_n1864, new_n1914);
and_8  g01538(new_n1601, new_n1598, new_n1915);
and_8  g01539(new_n1606, new_n1602, new_n1916);
or_8   g01540(new_n1916, new_n1915, new_n1917);
and_8  g01541(n9400, n4928, new_n1918);
and_8  g01542(n4141, n2464, new_n1919);
and_8  g01543(n8236, n6877, new_n1920);
xor_4  g01544(new_n1920, new_n1919, new_n1921);
xor_4  g01545(new_n1921, new_n1918, new_n1922);
xor_4  g01546(new_n1922, new_n1917, new_n1923);
and_8  g01547(new_n1600, new_n1599, new_n1924);
and_8  g01548(n11311, n5105, new_n1925);
xnor_4 g01549(new_n1925, new_n1924, new_n1926);
and_8  g01550(n7500, n4203, new_n1927);
and_8  g01551(n4187, n1209, new_n1928);
and_8  g01552(n12753, n7354, new_n1929);
xnor_4 g01553(new_n1929, new_n1928, new_n1930);
xor_4  g01554(new_n1930, new_n1927, new_n1931);
xor_4  g01555(new_n1931, new_n1926, new_n1932);
xor_4  g01556(new_n1932, new_n1923, new_n1933);
not_8  g01557(new_n1618, new_n1934);
and_8  g01558(new_n1613, new_n1612, new_n1935);
and_8  g01559(new_n1615, new_n1607, new_n1936);
xor_4  g01560(new_n1936, new_n1935, new_n1937);
or_8   g01561(new_n1937, new_n1934, new_n1938);
xor_4  g01562(new_n1938, new_n1933, new_n1939);
xor_4  g01563(new_n1939, new_n1621, new_n1940);
not_8  g01564(new_n1626, new_n1941);
or_8   g01565(new_n1628, new_n1593, new_n1942);
and_8  g01566(new_n1942, new_n1941, new_n1943);
xor_4  g01567(new_n1943, new_n1940, new_n1944);
or_8   g01568(new_n1690, new_n1686, new_n1945);
or_8   g01569(new_n1694, new_n1691, new_n1946);
and_8  g01570(new_n1946, new_n1945, new_n1947);
and_8  g01571(n5814, n3992, new_n1948);
and_8  g01572(n12704, n8384, new_n1949);
and_8  g01573(n7236, n4903, new_n1950);
xnor_4 g01574(new_n1950, new_n1949, new_n1951);
xor_4  g01575(new_n1951, new_n1948, new_n1952);
xor_4  g01576(new_n1952, new_n1947, new_n1953);
and_8  g01577(new_n1693, new_n1692, new_n1954);
and_8  g01578(n7294, n6358, new_n1955);
xnor_4 g01579(new_n1955, new_n1954, new_n1956);
nand_5 g01580(n10848, n1471, new_n1957);
and_8  g01581(n5198, n1980, new_n1958);
and_8  g01582(n8028, n7646, new_n1959);
xor_4  g01583(new_n1959, new_n1958, new_n1960);
xor_4  g01584(new_n1960, new_n1957, new_n1961);
xor_4  g01585(new_n1961, new_n1956, new_n1962);
or_8   g01586(new_n1962, new_n1953, new_n1963);
not_8  g01587(new_n1952, new_n1964);
xor_4  g01588(new_n1964, new_n1947, new_n1965);
not_8  g01589(new_n1962, new_n1966);
or_8   g01590(new_n1966, new_n1965, new_n1967);
and_8  g01591(new_n1967, new_n1963, new_n1968);
not_8  g01592(new_n1683, new_n1969);
nand_5 g01593(new_n1681, new_n1680, new_n1970);
not_8  g01594(new_n1970, new_n1971);
and_8  g01595(new_n1706, new_n1971, new_n1972);
and_8  g01596(new_n1696, new_n1970, new_n1973);
or_8   g01597(new_n1973, new_n1972, new_n1974);
and_8  g01598(new_n1974, new_n1969, new_n1975);
or_8   g01599(new_n1975, new_n1968, new_n1976);
and_8  g01600(new_n1966, new_n1965, new_n1977);
and_8  g01601(new_n1962, new_n1953, new_n1978);
or_8   g01602(new_n1978, new_n1977, new_n1979);
or_8   g01603(new_n1696, new_n1970, new_n1980_1);
or_8   g01604(new_n1706, new_n1971, new_n1981);
and_8  g01605(new_n1981, new_n1980_1, new_n1982);
or_8   g01606(new_n1982, new_n1683, new_n1983);
or_8   g01607(new_n1983, new_n1979, new_n1984);
and_8  g01608(new_n1984, new_n1976, new_n1985);
xor_4  g01609(new_n1985, new_n1705, new_n1986);
not_8  g01610(new_n1712, new_n1987);
and_8  g01611(new_n1717, new_n1811, new_n1988);
or_8   g01612(new_n1988, new_n1987, new_n1989);
and_8  g01613(new_n1989, new_n1986, new_n1990);
xor_4  g01614(new_n1985, new_n1713, new_n1991);
nor_6  g01615(new_n1988, new_n1987, new_n1992);
and_8  g01616(new_n1992, new_n1991, new_n1993);
or_8   g01617(new_n1993, new_n1990, new_n1994);
and_8  g01618(new_n1806, new_n1762, new_n1995);
and_8  g01619(new_n1802, new_n1763, new_n1996);
or_8   g01620(new_n1996, new_n1995, new_n1997);
or_8   g01621(new_n1997, new_n1761, new_n1998);
and_8  g01622(new_n1998, new_n1803, new_n1999);
nor_6  g01623(new_n1774, new_n1768, new_n2000);
and_8  g01624(n11478, n5069, new_n2001);
and_8  g01625(n6806, n5283, new_n2002);
and_8  g01626(n12044, n4805, new_n2003);
xnor_4 g01627(new_n2003, new_n2002, new_n2004);
xor_4  g01628(new_n2004, new_n2001, new_n2005);
and_8  g01629(new_n2005, new_n2000, new_n2006);
nor_6  g01630(new_n2005, new_n2000, new_n2007);
or_8   g01631(new_n2007, new_n2006, new_n2008);
and_8  g01632(new_n1766, new_n1765, new_n2009);
and_8  g01633(n2802, n137, new_n2010);
xnor_4 g01634(new_n2010, new_n2009, new_n2011);
and_8  g01635(n6797, n1512, new_n2012);
and_8  g01636(n6294, n533, new_n2013);
and_8  g01637(n3146, n1564, new_n2014);
xnor_4 g01638(new_n2014, new_n2013, new_n2015);
xor_4  g01639(new_n2015, new_n2012, new_n2016);
xor_4  g01640(new_n2016, new_n2011, new_n2017);
xor_4  g01641(new_n2017, new_n2008, new_n2018);
and_8  g01642(new_n1778, new_n1777, new_n2019);
and_8  g01643(new_n1788, new_n1784, new_n2020);
and_8  g01644(new_n2020, new_n2019, new_n2021);
nor_6  g01645(new_n2020, new_n2019, new_n2022);
or_8   g01646(new_n2022, new_n2021, new_n2023);
and_8  g01647(new_n2023, new_n1781, new_n2024_1);
nor_6  g01648(new_n2024_1, new_n2018, new_n2025);
and_8  g01649(new_n2024_1, new_n2018, new_n2026);
or_8   g01650(new_n2026, new_n2025, new_n2027);
xor_4  g01651(new_n2027, new_n1804, new_n2028);
xor_4  g01652(new_n2028, new_n1999, new_n2029);
and_8  g01653(new_n2029, new_n1994, new_n2030);
or_8   g01654(new_n1992, new_n1991, new_n2031);
or_8   g01655(new_n1989, new_n1986, new_n2032);
and_8  g01656(new_n2032, new_n2031, new_n2033);
and_8  g01657(new_n1808, new_n1813, new_n2034);
or_8   g01658(new_n2034, new_n1995, new_n2035);
xor_4  g01659(new_n2028, new_n2035, new_n2036);
and_8  g01660(new_n2036, new_n2033, new_n2037);
or_8   g01661(new_n2037, new_n2030, new_n2038);
and_8  g01662(new_n1854, new_n1855, new_n2039);
nor_6  g01663(new_n2039, new_n2038, new_n2040);
and_8  g01664(new_n2039, new_n2038, new_n2041);
or_8   g01665(new_n2041, new_n2040, new_n2042);
or_8   g01666(new_n2042, new_n1944, new_n2043);
not_8  g01667(new_n1944, new_n2044);
xor_4  g01668(new_n2039, new_n2038, new_n2045);
or_8   g01669(new_n2045, new_n2044, new_n2046);
and_8  g01670(new_n2046, new_n2043, new_n2047);
and_8  g01671(new_n2047, new_n1914, new_n2048);
nor_6  g01672(new_n1913, new_n1864, new_n2049);
and_8  g01673(new_n2045, new_n2044, new_n2050);
and_8  g01674(new_n2042, new_n1944, new_n2051);
or_8   g01675(new_n2051, new_n2050, new_n2052);
and_8  g01676(new_n2052, new_n2049, new_n2053);
or_8   g01677(new_n2053, new_n2048, new_n2054);
and_8  g01678(new_n2054, new_n1552, new_n2055);
not_8  g01679(new_n1552, new_n2056);
or_8   g01680(new_n2052, new_n2049, new_n2057);
or_8   g01681(new_n2047, new_n1914, new_n2058);
and_8  g01682(new_n2058, new_n2057, new_n2059);
or_8   g01683(new_n2059, new_n2056, new_n2060);
or_8   g01684(new_n2054, new_n1552, new_n2061);
and_8  g01685(new_n2061, new_n2060, new_n2062);
xor_4  g01686(new_n1549, new_n1547, new_n2063);
nor_6  g01687(new_n1912, new_n1870, new_n2064);
or_8   g01688(new_n2064, new_n1913, new_n2065);
and_8  g01689(new_n2065, new_n2063, new_n2066);
xor_4  g01690(new_n1546, new_n1545, new_n2067);
xor_4  g01691(new_n1910, new_n1880, new_n2068);
or_8   g01692(new_n2068, new_n2067, new_n2069);
not_8  g01693(new_n2067, new_n2070);
nor_6  g01694(new_n1910, new_n1880, new_n2071);
and_8  g01695(new_n1910, new_n1880, new_n2072);
or_8   g01696(new_n2072, new_n2071, new_n2073);
and_8  g01697(new_n2073, new_n2070, new_n2074);
and_8  g01698(new_n2068, new_n2067, new_n2075);
or_8   g01699(new_n2075, new_n2074, new_n2076);
xor_4  g01700(new_n1544, new_n1538, new_n2077);
xor_4  g01701(new_n1908, new_n1886, new_n2078);
nor_6  g01702(new_n2078, new_n2077, new_n2079);
not_8  g01703(new_n2079, new_n2080);
xor_4  g01704(new_n1905, new_n1897, new_n2081);
not_8  g01705(new_n2081, new_n2082);
not_8  g01706(new_n1239, new_n2083);
nand_5 g01707(new_n1455, new_n2083, new_n2084);
nand_5 g01708(new_n2084, new_n1539, new_n2085);
nand_5 g01709(new_n1459, new_n2083, new_n2086);
and_8  g01710(new_n2086, new_n2085, new_n2087_1);
or_8   g01711(new_n2087_1, new_n2082, new_n2088);
xor_4  g01712(new_n2087_1, new_n2081, new_n2089);
and_8  g01713(new_n1244, new_n1239, new_n2090);
xor_4  g01714(new_n1541, new_n1540, new_n2091);
or_8   g01715(new_n2091, new_n2090, new_n2092);
xor_4  g01716(new_n1903, new_n1902, new_n2093);
xnor_4 g01717(new_n2091, new_n2090, new_n2094);
or_8   g01718(new_n2094, new_n2093, new_n2095);
and_8  g01719(new_n2095, new_n2092, new_n2096_1);
or_8   g01720(new_n2096_1, new_n2089, new_n2097);
and_8  g01721(new_n2097, new_n2088, new_n2098);
and_8  g01722(new_n2078, new_n2077, new_n2099);
or_8   g01723(new_n2099, new_n2079, new_n2100);
or_8   g01724(new_n2100, new_n2098, new_n2101);
and_8  g01725(new_n2101, new_n2080, new_n2102);
or_8   g01726(new_n2102, new_n2076, new_n2103);
and_8  g01727(new_n2103, new_n2069, new_n2104);
not_8  g01728(new_n2063, new_n2105);
xor_4  g01729(new_n1912, new_n1870, new_n2106);
or_8   g01730(new_n2106, new_n2105, new_n2107);
or_8   g01731(new_n2065, new_n2063, new_n2108);
and_8  g01732(new_n2108, new_n2107, new_n2109);
and_8  g01733(new_n2109, new_n2104, new_n2110);
or_8   g01734(new_n2110, new_n2066, new_n2111);
and_8  g01735(new_n2111, new_n2062, new_n2112);
or_8   g01736(new_n2112, new_n2055, new_n2113);
or_8   g01737(new_n2048, new_n2050, new_n2114);
nor_6  g01738(new_n2040, new_n2030, new_n2115);
xor_4  g01739(new_n1521, new_n1523_1, new_n2116);
or_8   g01740(new_n2116, new_n1497, new_n2117);
not_8  g01741(new_n2117, new_n2118);
not_8  g01742(new_n1497, new_n2119);
xor_4  g01743(new_n1526, new_n2119, new_n2120);
not_8  g01744(new_n1547, new_n2121);
xor_4  g01745(new_n1535, new_n1528, new_n2122);
and_8  g01746(new_n2122, new_n2121, new_n2123);
or_8   g01747(new_n2123, new_n1536, new_n2124);
and_8  g01748(new_n2124, new_n2120, new_n2125);
or_8   g01749(new_n2125, new_n2118, new_n2126);
and_8  g01750(new_n1985, new_n1705, new_n2127);
or_8   g01751(new_n1990, new_n2127, new_n2128);
or_8   g01752(new_n2128, new_n2126, new_n2129);
or_8   g01753(new_n1551, new_n1527, new_n2130);
and_8  g01754(new_n2130, new_n2117, new_n2131_1);
nor_6  g01755(new_n1990, new_n2127, new_n2132);
or_8   g01756(new_n2132, new_n2131_1, new_n2133);
and_8  g01757(new_n2133, new_n2129, new_n2134);
and_8  g01758(new_n1976, new_n1980_1, new_n2135);
and_8  g01759(new_n2010, new_n2009, new_n2136);
nor_6  g01760(new_n2016, new_n2011, new_n2137);
or_8   g01761(new_n2137, new_n2136, new_n2138);
nand_5 g01762(n7862, n615, new_n2139);
and_8  g01763(n4903, n3992, new_n2140);
and_8  g01764(n6806, n137, new_n2141);
xor_4  g01765(new_n2141, new_n2140, new_n2142);
xnor_4 g01766(new_n2142, new_n2139, new_n2143);
xor_4  g01767(new_n2143, new_n2138, new_n2144);
and_8  g01768(n6797, n533, new_n2145);
and_8  g01769(n8384, n5814, new_n2146);
xor_4  g01770(new_n2146, new_n2145, new_n2147);
and_8  g01771(n12044, n11478, new_n2148);
and_8  g01772(n7294, n5198, new_n2149);
xor_4  g01773(new_n2149, new_n2148, new_n2150);
xor_4  g01774(new_n2150, new_n2147, new_n2151);
and_8  g01775(new_n2003, new_n2002, new_n2152);
or_8   g01776(new_n2003, new_n2002, new_n2153);
and_8  g01777(new_n2153, new_n2001, new_n2154);
or_8   g01778(new_n2154, new_n2152, new_n2155);
xor_4  g01779(new_n2155, new_n2151, new_n2156);
nand_5 g01780(n10174, n7354, new_n2157);
and_8  g01781(n4928, n2464, new_n2158);
and_8  g01782(n11311, n4141, new_n2159);
xor_4  g01783(new_n2159, new_n2158, new_n2160);
and_8  g01784(n4005, n3172, new_n2161);
and_8  g01785(n7236, n1906, new_n2162);
xnor_4 g01786(new_n2162, new_n2161, new_n2163);
xor_4  g01787(new_n2163, new_n2160, new_n2164);
xor_4  g01788(new_n2164, new_n2157, new_n2165);
xor_4  g01789(new_n2165, new_n2156, new_n2166);
xor_4  g01790(new_n2166, new_n2144, new_n2167);
nor_6  g01791(new_n2167, new_n2135, new_n2168);
and_8  g01792(new_n2167, new_n2135, new_n2169);
or_8   g01793(new_n2169, new_n2168, new_n2170);
or_8   g01794(new_n1964, new_n1947, new_n2171);
and_8  g01795(new_n1963, new_n2171, new_n2172);
and_8  g01796(n9080, n2509, new_n2173);
or_8   g01797(new_n1507, new_n1506, new_n2174);
or_8   g01798(new_n1508, new_n1505, new_n2175);
and_8  g01799(new_n2175, new_n2174, new_n2176);
not_8  g01800(n2508, new_n2177);
not_8  g01801(n5240, new_n2178);
or_8   g01802(new_n2178, new_n2177, new_n2179);
and_8  g01803(n11757, n2585, new_n2180);
and_8  g01804(n12706, n1333, new_n2181);
xor_4  g01805(new_n2181, new_n2180, new_n2182);
xor_4  g01806(new_n2182, new_n2179, new_n2183);
xor_4  g01807(new_n2183, new_n2176, new_n2184);
xor_4  g01808(new_n2184, new_n2173, new_n2185);
xor_4  g01809(new_n2185, new_n2172, new_n2186);
not_8  g01810(new_n2186, new_n2187);
or_8   g01811(new_n2187, new_n2170, new_n2188);
xor_4  g01812(new_n2167, new_n2135, new_n2189);
or_8   g01813(new_n2186, new_n2189, new_n2190);
and_8  g01814(new_n2190, new_n2188, new_n2191);
and_8  g01815(new_n1936, new_n1935, new_n2192);
and_8  g01816(new_n1938, new_n1933, new_n2193);
or_8   g01817(new_n2193, new_n2192, new_n2194);
nand_5 g01818(new_n1499, new_n1498, new_n2195);
and_8  g01819(new_n1522, new_n2195, new_n2196);
xor_4  g01820(new_n2196, new_n2194, new_n2197);
or_8   g01821(new_n1922, new_n1917, new_n2198);
not_8  g01822(new_n1923, new_n2199);
or_8   g01823(new_n1932, new_n2199, new_n2200);
and_8  g01824(new_n2200, new_n2198, new_n2201);
and_8  g01825(n12704, n6358, new_n2202);
and_8  g01826(n3146, n1512, new_n2203);
xor_4  g01827(new_n2203, new_n2202, new_n2204);
and_8  g01828(n5105, n4187, new_n2205);
and_8  g01829(n6294, n2802, new_n2206);
xor_4  g01830(new_n2206, new_n2205, new_n2207);
and_8  g01831(n9400, n8236, new_n2208);
and_8  g01832(n1980, n1471, new_n2209);
xor_4  g01833(new_n2209, new_n2208, new_n2210);
xor_4  g01834(new_n2210, new_n2207, new_n2211);
xor_4  g01835(new_n2211, new_n2204, new_n2212);
nand_5 g01836(n12720, n11821, new_n2213);
and_8  g01837(n4938, n1564, new_n2214);
and_8  g01838(n5694, n4805, new_n2215);
xor_4  g01839(new_n2215, new_n2214, new_n2216);
xor_4  g01840(new_n2216, new_n2213, new_n2217);
xor_4  g01841(new_n2217, new_n2212, new_n2218);
or_8   g01842(new_n1950, new_n1949, new_n2219);
or_8   g01843(new_n1951, new_n1948, new_n2220);
and_8  g01844(new_n2220, new_n2219, new_n2221);
nand_5 g01845(new_n1503, new_n1502, new_n2222);
or_8   g01846(new_n1509, new_n1504, new_n2223);
and_8  g01847(new_n2223, new_n2222, new_n2224);
xor_4  g01848(new_n2224, new_n2221, new_n2225);
xor_4  g01849(new_n2225, new_n2218, new_n2226_1);
nor_6  g01850(new_n2226_1, new_n2201, new_n2227);
and_8  g01851(new_n2226_1, new_n2201, new_n2228);
or_8   g01852(new_n2228, new_n2227, new_n2229);
not_8  g01853(new_n2021, new_n2230);
or_8   g01854(new_n2024_1, new_n2018, new_n2231);
and_8  g01855(new_n2231, new_n2230, new_n2232);
nor_6  g01856(new_n2017, new_n2008, new_n2233);
or_8   g01857(new_n2233, new_n2006, new_n2234);
and_8  g01858(new_n1955, new_n1954, new_n2235);
nor_6  g01859(new_n1961, new_n1956, new_n2236);
or_8   g01860(new_n2236, new_n2235, new_n2237);
and_8  g01861(n4203, n1209, new_n2238);
and_8  g01862(n6826, n6038, new_n2239);
and_8  g01863(n5283, n5069, new_n2240);
xor_4  g01864(new_n2240, new_n2239, new_n2241);
xor_4  g01865(new_n2241, new_n2238, new_n2242);
not_8  g01866(new_n2242, new_n2243);
or_8   g01867(new_n2243, new_n2237, new_n2244);
nor_6  g01868(new_n2236, new_n2235, new_n2245);
or_8   g01869(new_n2242, new_n2245, new_n2246);
and_8  g01870(new_n2246, new_n2244, new_n2247);
or_8   g01871(new_n2014, new_n2013, new_n2248);
or_8   g01872(new_n2015, new_n2012, new_n2249);
and_8  g01873(new_n2249, new_n2248, new_n2250);
nor_6  g01874(new_n1959, new_n1958, new_n2251);
and_8  g01875(new_n1960, new_n1957, new_n2252);
or_8   g01876(new_n2252, new_n2251, new_n2253_1);
and_8  g01877(new_n1920, new_n1919, new_n2254);
or_8   g01878(new_n1920, new_n1919, new_n2255);
and_8  g01879(new_n2255, new_n1918, new_n2256);
or_8   g01880(new_n2256, new_n2254, new_n2257);
xor_4  g01881(new_n2257, new_n2253_1, new_n2258);
and_8  g01882(new_n2258, new_n2250, new_n2259);
nor_6  g01883(new_n2258, new_n2250, new_n2260);
or_8   g01884(new_n2260, new_n2259, new_n2261);
xor_4  g01885(new_n2261, new_n2247, new_n2262);
and_8  g01886(new_n2262, new_n2234, new_n2263);
not_8  g01887(new_n2234, new_n2264);
xor_4  g01888(new_n2258, new_n2250, new_n2265);
xor_4  g01889(new_n2265, new_n2247, new_n2266);
and_8  g01890(new_n2266, new_n2264, new_n2267);
or_8   g01891(new_n2267, new_n2263, new_n2268);
or_8   g01892(new_n2268, new_n2232, new_n2269);
or_8   g01893(new_n2025, new_n2021, new_n2270);
nor_6  g01894(new_n2267, new_n2263, new_n2271);
or_8   g01895(new_n2271, new_n2270, new_n2272);
and_8  g01896(new_n2272, new_n2269, new_n2273);
xor_4  g01897(new_n2273, new_n2229, new_n2274);
and_8  g01898(new_n2274, new_n2197, new_n2275);
nor_6  g01899(new_n2193, new_n2192, new_n2276);
xor_4  g01900(new_n2196, new_n2276, new_n2277);
xor_4  g01901(new_n2226_1, new_n2201, new_n2278_1);
xor_4  g01902(new_n2273, new_n2278_1, new_n2279);
and_8  g01903(new_n2279, new_n2277, new_n2280);
or_8   g01904(new_n2280, new_n2275, new_n2281);
or_8   g01905(new_n2281, new_n2191, new_n2282);
xor_4  g01906(new_n2186, new_n2170, new_n2283);
or_8   g01907(new_n2279, new_n2277, new_n2284);
or_8   g01908(new_n2274, new_n2197, new_n2285);
and_8  g01909(new_n2285, new_n2284, new_n2286);
or_8   g01910(new_n2286, new_n2283, new_n2287);
and_8  g01911(new_n2287, new_n2282, new_n2288);
and_8  g01912(new_n2288, new_n2134, new_n2289);
nor_6  g01913(new_n2288, new_n2134, new_n2290);
or_8   g01914(new_n2290, new_n2289, new_n2291);
and_8  g01915(new_n2291, new_n2115, new_n2292);
or_8   g01916(new_n2040, new_n2030, new_n2293);
xor_4  g01917(new_n2288, new_n2134, new_n2294);
and_8  g01918(new_n2294, new_n2293, new_n2295);
or_8   g01919(new_n2295, new_n2292, new_n2296);
nand_5 g01920(new_n1925, new_n1924, new_n2297);
or_8   g01921(new_n1931, new_n1926, new_n2298);
and_8  g01922(new_n2298, new_n2297, new_n2299);
and_8  g01923(n6877, n783, new_n2300);
and_8  g01924(n8028, n4722, new_n2301_1);
xor_4  g01925(new_n2301_1, new_n2300, new_n2302);
xor_4  g01926(new_n2302, new_n2299, new_n2303);
not_8  g01927(new_n1621, new_n2304);
and_8  g01928(new_n1939, new_n2304, new_n2305);
xor_4  g01929(new_n1939, new_n2304, new_n2306);
not_8  g01930(new_n1593, new_n2307);
xor_4  g01931(new_n1625, new_n1594, new_n2308);
and_8  g01932(new_n2308, new_n2307, new_n2309);
or_8   g01933(new_n2309, new_n1626, new_n2310);
and_8  g01934(new_n2310, new_n2306, new_n2311);
or_8   g01935(new_n2311, new_n2305, new_n2312);
nand_5 g01936(n10848, n7646, new_n2313);
not_8  g01937(new_n2313, new_n2314);
or_8   g01938(new_n2314, new_n2312, new_n2315);
not_8  g01939(new_n2305, new_n2316_1);
or_8   g01940(new_n1943, new_n1940, new_n2317);
and_8  g01941(new_n2317, new_n2316_1, new_n2318);
or_8   g01942(new_n2313, new_n2318, new_n2319);
and_8  g01943(new_n2319, new_n2315, new_n2320);
and_8  g01944(new_n2320, new_n2303, new_n2321);
not_8  g01945(new_n2303, new_n2322);
and_8  g01946(new_n2313, new_n2318, new_n2323);
and_8  g01947(new_n2314, new_n2312, new_n2324);
or_8   g01948(new_n2324, new_n2323, new_n2325);
and_8  g01949(new_n2325, new_n2322, new_n2326);
or_8   g01950(new_n2326, new_n2321, new_n2327);
or_8   g01951(new_n2027, new_n1804, new_n2328);
not_8  g01952(new_n2028, new_n2329);
or_8   g01953(new_n2329, new_n1999, new_n2330);
and_8  g01954(new_n2330, new_n2328, new_n2331);
and_8  g01955(new_n1519, new_n1514, new_n2332);
and_8  g01956(new_n1520, new_n1510_1, new_n2333);
or_8   g01957(new_n2333, new_n2332, new_n2334);
or_8   g01958(new_n1929, new_n1928, new_n2335);
or_8   g01959(new_n1930, new_n1927, new_n2336);
and_8  g01960(new_n2336, new_n2335, new_n2337);
nand_5 g01961(n12753, n7500, new_n2338);
and_8  g01962(new_n1517, new_n1516, new_n2339);
or_8   g01963(new_n1517, new_n1516, new_n2340);
and_8  g01964(new_n2340, new_n1515, new_n2341);
or_8   g01965(new_n2341, new_n2339, new_n2342);
xor_4  g01966(new_n2342, new_n2338, new_n2343);
xor_4  g01967(new_n2343, new_n2337, new_n2344);
xor_4  g01968(new_n2344, new_n2334, new_n2345);
xor_4  g01969(new_n2345, new_n2331, new_n2346);
xor_4  g01970(new_n2346, new_n2327, new_n2347_1);
and_8  g01971(new_n2347_1, new_n2296, new_n2348);
nor_6  g01972(new_n2347_1, new_n2296, new_n2349);
or_8   g01973(new_n2349, new_n2348, new_n2350);
or_8   g01974(new_n2350, new_n2114, new_n2351);
and_8  g01975(new_n2057, new_n2043, new_n2352);
xor_4  g01976(new_n2347_1, new_n2296, new_n2353);
or_8   g01977(new_n2353, new_n2352, new_n2354);
and_8  g01978(new_n2354, new_n2351, new_n2355);
xor_4  g01979(new_n2355, new_n2113, n671);
and_8  g01980(n11917, n4312, new_n2357);
and_8  g01981(n12705, n4921, new_n2358);
and_8  g01982(n12025, n9956, new_n2359);
xor_4  g01983(new_n2359, new_n2358, new_n2360);
xor_4  g01984(new_n2360, new_n2357, new_n2361);
and_8  g01985(n12705, n9956, new_n2362);
and_8  g01986(n11917, n1097, new_n2363);
or_8   g01987(new_n2363, new_n2362, new_n2364);
and_8  g01988(new_n2363, new_n2362, new_n2365);
and_8  g01989(n4921, n4312, new_n2366);
or_8   g01990(new_n2366, new_n2365, new_n2367);
nand_5 g01991(new_n2367, new_n2364, new_n2368);
xnor_4 g01992(new_n2368, new_n2361, new_n2369);
and_8  g01993(n5964, n2577, new_n2370);
and_8  g01994(n3842, n1097, new_n2371);
xor_4  g01995(new_n2371, new_n2370, new_n2372);
xor_4  g01996(new_n2372, new_n2369, new_n2373);
and_8  g01997(n5964, n3842, new_n2374);
and_8  g01998(n9956, n4312, new_n2375);
and_8  g01999(n11917, n5964, new_n2376);
or_8   g02000(new_n2376, new_n2375, new_n2377);
and_8  g02001(new_n2376, new_n2375, new_n2378);
and_8  g02002(n4921, n1097, new_n2379);
or_8   g02003(new_n2379, new_n2378, new_n2380);
and_8  g02004(new_n2380, new_n2377, new_n2381);
and_8  g02005(new_n2381, new_n2374, new_n2382);
xor_4  g02006(new_n2381, new_n2374, new_n2383_1);
xor_4  g02007(new_n2363, new_n2362, new_n2384);
xor_4  g02008(new_n2384, new_n2366, new_n2385);
and_8  g02009(new_n2385, new_n2383_1, new_n2386);
or_8   g02010(new_n2386, new_n2382, new_n2387);
xor_4  g02011(new_n2387, new_n2373, new_n2388);
and_8  g02012(n5305, n2577, new_n2389);
not_8  g02013(new_n2389, new_n2390);
xnor_4 g02014(new_n2385, new_n2383_1, new_n2391);
nand_5 g02015(new_n2391, new_n2390, new_n2392);
xor_4  g02016(new_n2391, new_n2389, new_n2393_1);
and_8  g02017(n5305, n3842, new_n2394);
and_8  g02018(n9956, n1097, new_n2395);
and_8  g02019(n11917, n5305, new_n2396);
and_8  g02020(new_n2396, new_n2395, new_n2397);
or_8   g02021(new_n2396, new_n2395, new_n2398);
and_8  g02022(n5964, n4921, new_n2399);
and_8  g02023(new_n2399, new_n2398, new_n2400);
or_8   g02024(new_n2400, new_n2397, new_n2401);
and_8  g02025(new_n2401, new_n2394, new_n2402);
xor_4  g02026(new_n2401, new_n2394, new_n2403);
xor_4  g02027(new_n2376, new_n2375, new_n2404);
xor_4  g02028(new_n2404, new_n2379, new_n2405);
and_8  g02029(new_n2405, new_n2403, new_n2406);
or_8   g02030(new_n2406, new_n2402, new_n2407);
or_8   g02031(new_n2407, new_n2393_1, new_n2408);
and_8  g02032(new_n2408, new_n2392, new_n2409);
and_8  g02033(new_n2409, new_n2388, new_n2410);
nor_6  g02034(new_n2360, new_n2357, new_n2411);
and_8  g02035(new_n2368, new_n2361, new_n2412);
or_8   g02036(new_n2412, new_n2411, new_n2413);
and_8  g02037(n9637, n5964, new_n2414);
and_8  g02038(n2577, n1097, new_n2415);
and_8  g02039(n5305, n1835, new_n2416);
xnor_4 g02040(new_n2416, new_n2415, new_n2417);
xor_4  g02041(new_n2417, new_n2414, new_n2418);
xor_4  g02042(new_n2418, new_n2413, new_n2419);
and_8  g02043(new_n2359, new_n2358, new_n2420);
and_8  g02044(n4312, n3842, new_n2421);
xnor_4 g02045(new_n2421, new_n2420, new_n2422);
nand_5 g02046(n12025, n4921, new_n2423);
and_8  g02047(n12705, n11917, new_n2424);
and_8  g02048(n11257, n9956, new_n2425_1);
xnor_4 g02049(new_n2425_1, new_n2424, new_n2426);
xor_4  g02050(new_n2426, new_n2423, new_n2427);
xor_4  g02051(new_n2427, new_n2422, new_n2428);
xor_4  g02052(new_n2428, new_n2419, new_n2429);
nand_5 g02053(new_n2372, new_n2369, new_n2430);
nand_5 g02054(new_n2371, new_n2370, new_n2431_1);
and_8  g02055(new_n2387, new_n2373, new_n2432);
xor_4  g02056(new_n2432, new_n2431_1, new_n2433_1);
and_8  g02057(new_n2433_1, new_n2430, new_n2434_1);
xor_4  g02058(new_n2434_1, new_n2429, new_n2435);
xor_4  g02059(new_n2435, new_n2410, new_n2436);
and_8  g02060(n9637, n5305, new_n2437);
xor_4  g02061(new_n2409, new_n2388, new_n2438);
and_8  g02062(new_n2438, new_n2437, new_n2439);
xor_4  g02063(new_n2405, new_n2403, new_n2440);
not_8  g02064(new_n2440, new_n2441);
xor_4  g02065(new_n2396, new_n2395, new_n2442);
and_8  g02066(n9956, n5964, new_n2443);
and_8  g02067(n5305, n4921, new_n2444);
nand_5 g02068(new_n2444, new_n2443, new_n2445);
or_8   g02069(new_n2445, new_n2442, new_n2446);
or_8   g02070(new_n2446, new_n2441, new_n2447);
xor_4  g02071(new_n2407, new_n2393_1, new_n2448);
nor_6  g02072(new_n2448, new_n2447, new_n2449);
xor_4  g02073(new_n2438, new_n2437, new_n2450);
and_8  g02074(new_n2450, new_n2449, new_n2451);
or_8   g02075(new_n2451, new_n2439, new_n2452);
xor_4  g02076(new_n2452, new_n2436, new_n2453);
not_8  g02077(new_n2453, new_n2454);
and_8  g02078(n8759, n8065, new_n2455);
not_8  g02079(new_n2455, new_n2456);
and_8  g02080(n7436, n6126, new_n2457);
not_8  g02081(new_n2457, new_n2458);
and_8  g02082(n9241, n3719, new_n2459);
and_8  g02083(n8276, n3602, new_n2460);
xor_4  g02084(new_n2460, new_n2459, new_n2461);
xor_4  g02085(new_n2461, new_n2458, new_n2462);
and_8  g02086(n8276, n3719, new_n2463);
and_8  g02087(n12299, n6126, new_n2464_1);
or_8   g02088(new_n2464_1, new_n2463, new_n2465);
and_8  g02089(new_n2464_1, new_n2463, new_n2466);
and_8  g02090(n7436, n3602, new_n2467);
or_8   g02091(new_n2467, new_n2466, new_n2468);
and_8  g02092(new_n2468, new_n2465, new_n2469);
xor_4  g02093(new_n2469, new_n2462, new_n2470);
and_8  g02094(n10439, n6776, new_n2471);
and_8  g02095(n12299, n8595, new_n2472);
xor_4  g02096(new_n2472, new_n2471, new_n2473);
not_8  g02097(new_n2473, new_n2474);
or_8   g02098(new_n2474, new_n2470, new_n2475);
xor_4  g02099(new_n2461, new_n2457, new_n2476);
xor_4  g02100(new_n2469, new_n2476, new_n2477);
or_8   g02101(new_n2473, new_n2477, new_n2478);
and_8  g02102(new_n2478, new_n2475, new_n2479);
and_8  g02103(n8595, n6776, new_n2480);
and_8  g02104(n7436, n3719, new_n2481);
and_8  g02105(n6776, n6126, new_n2482);
or_8   g02106(new_n2482, new_n2481, new_n2483);
and_8  g02107(new_n2482, new_n2481, new_n2484);
and_8  g02108(n12299, n3602, new_n2485);
or_8   g02109(new_n2485, new_n2484, new_n2486);
and_8  g02110(new_n2486, new_n2483, new_n2487);
and_8  g02111(new_n2487, new_n2480, new_n2488);
xnor_4 g02112(new_n2487, new_n2480, new_n2489);
xnor_4 g02113(new_n2464_1, new_n2463, new_n2490);
xor_4  g02114(new_n2490, new_n2467, new_n2491);
nor_6  g02115(new_n2491, new_n2489, new_n2492);
or_8   g02116(new_n2492, new_n2488, new_n2493);
and_8  g02117(new_n2493, new_n2479, new_n2494);
nor_6  g02118(new_n2493, new_n2479, new_n2495);
or_8   g02119(new_n2495, new_n2494, new_n2496);
not_8  g02120(new_n2496, new_n2497);
and_8  g02121(n10439, n8759, new_n2498_1);
not_8  g02122(new_n2498_1, new_n2499);
and_8  g02123(new_n2491, new_n2489, new_n2500);
or_8   g02124(new_n2500, new_n2492, new_n2501);
and_8  g02125(new_n2501, new_n2499, new_n2502);
xor_4  g02126(new_n2491, new_n2489, new_n2503);
or_8   g02127(new_n2503, new_n2498_1, new_n2504);
or_8   g02128(new_n2501, new_n2499, new_n2505);
and_8  g02129(new_n2505, new_n2504, new_n2506);
and_8  g02130(n8759, n8595, new_n2507_1);
and_8  g02131(n12299, n3719, new_n2508_1);
and_8  g02132(n8759, n6126, new_n2509_1);
and_8  g02133(new_n2509_1, new_n2508_1, new_n2510);
or_8   g02134(new_n2509_1, new_n2508_1, new_n2511);
and_8  g02135(n6776, n3602, new_n2512_1);
and_8  g02136(new_n2512_1, new_n2511, new_n2513);
or_8   g02137(new_n2513, new_n2510, new_n2514);
and_8  g02138(new_n2514, new_n2507_1, new_n2515_1);
xor_4  g02139(new_n2514, new_n2507_1, new_n2516);
xor_4  g02140(new_n2482, new_n2481, new_n2517);
xor_4  g02141(new_n2517, new_n2485, new_n2518);
and_8  g02142(new_n2518, new_n2516, new_n2519);
or_8   g02143(new_n2519, new_n2515_1, new_n2520);
not_8  g02144(new_n2520, new_n2521);
and_8  g02145(new_n2521, new_n2506, new_n2522_1);
or_8   g02146(new_n2522_1, new_n2502, new_n2523);
xor_4  g02147(new_n2523, new_n2497, new_n2524);
or_8   g02148(new_n2524, new_n2456, new_n2525);
xnor_4 g02149(new_n2518, new_n2516, new_n2526);
xnor_4 g02150(new_n2509_1, new_n2508_1, new_n2527);
and_8  g02151(n6776, n3719, new_n2528);
and_8  g02152(n8759, n3602, new_n2529);
and_8  g02153(new_n2529, new_n2528, new_n2530_1);
and_8  g02154(new_n2530_1, new_n2527, new_n2531);
not_8  g02155(new_n2531, new_n2532);
or_8   g02156(new_n2532, new_n2526, new_n2533);
and_8  g02157(new_n2503, new_n2498_1, new_n2534);
or_8   g02158(new_n2534, new_n2502, new_n2535);
xor_4  g02159(new_n2520, new_n2535, new_n2536);
or_8   g02160(new_n2536, new_n2533, new_n2537);
or_8   g02161(new_n2523, new_n2496, new_n2538);
or_8   g02162(new_n2520, new_n2535, new_n2539);
and_8  g02163(new_n2539, new_n2504, new_n2540);
or_8   g02164(new_n2540, new_n2497, new_n2541);
and_8  g02165(new_n2541, new_n2538, new_n2542);
xor_4  g02166(new_n2542, new_n2456, new_n2543);
or_8   g02167(new_n2543, new_n2537, new_n2544);
and_8  g02168(new_n2544, new_n2525, new_n2545);
not_8  g02169(new_n2538, new_n2546);
and_8  g02170(new_n2461, new_n2457, new_n2547);
and_8  g02171(new_n2469, new_n2476, new_n2548);
nor_6  g02172(new_n2548, new_n2547, new_n2549);
and_8  g02173(n8065, n6776, new_n2550);
and_8  g02174(n12299, n10439, new_n2551_1);
and_8  g02175(n10391, n8759, new_n2552);
xnor_4 g02176(new_n2552, new_n2551_1, new_n2553);
xor_4  g02177(new_n2553, new_n2550, new_n2554);
and_8  g02178(new_n2554, new_n2549, new_n2555);
nor_6  g02179(new_n2554, new_n2549, new_n2556);
or_8   g02180(new_n2556, new_n2555, new_n2557);
and_8  g02181(new_n2460, new_n2459, new_n2558_1);
and_8  g02182(n8595, n7436, new_n2559);
xnor_4 g02183(new_n2559, new_n2558_1, new_n2560);
and_8  g02184(n9241, n3602, new_n2561);
and_8  g02185(n8276, n6126, new_n2562);
and_8  g02186(n10510, n3719, new_n2563);
xnor_4 g02187(new_n2563, new_n2562, new_n2564_1);
xor_4  g02188(new_n2564_1, new_n2561, new_n2565);
xor_4  g02189(new_n2565, new_n2560, new_n2566);
xor_4  g02190(new_n2566, new_n2557, new_n2567);
not_8  g02191(new_n2567, new_n2568);
not_8  g02192(new_n2475, new_n2569);
and_8  g02193(new_n2472, new_n2471, new_n2570);
xor_4  g02194(new_n2494, new_n2570, new_n2571);
or_8   g02195(new_n2571, new_n2569, new_n2572);
xor_4  g02196(new_n2572, new_n2568, new_n2573);
and_8  g02197(new_n2573, new_n2546, new_n2574);
xor_4  g02198(new_n2572, new_n2567, new_n2575);
and_8  g02199(new_n2575, new_n2538, new_n2576);
or_8   g02200(new_n2576, new_n2574, new_n2577_1);
xor_4  g02201(new_n2577_1, new_n2545, new_n2578);
not_8  g02202(new_n2578, new_n2579);
and_8  g02203(n12648, n4826, new_n2580);
and_8  g02204(n10545, n7733, new_n2581_1);
and_8  g02205(n12925, n7690, new_n2582);
xor_4  g02206(new_n2582, new_n2581_1, new_n2583);
and_8  g02207(new_n2583, new_n2580, new_n2584);
nor_6  g02208(new_n2583, new_n2580, new_n2585_1);
or_8   g02209(new_n2585_1, new_n2584, new_n2586);
and_8  g02210(n12925, n10545, new_n2587);
and_8  g02211(n4826, n2530, new_n2588);
nor_6  g02212(new_n2588, new_n2587, new_n2589);
and_8  g02213(n12648, n7733, new_n2590);
not_8  g02214(new_n2590, new_n2591);
xor_4  g02215(new_n2588, new_n2587, new_n2592);
and_8  g02216(new_n2592, new_n2591, new_n2593);
or_8   g02217(new_n2593, new_n2589, new_n2594);
xor_4  g02218(new_n2594, new_n2586, new_n2595);
and_8  g02219(n8476, n4970, new_n2596);
and_8  g02220(n7610, n2530, new_n2597);
xor_4  g02221(new_n2597, new_n2596, new_n2598);
xor_4  g02222(new_n2598, new_n2595, new_n2599);
nand_5 g02223(n8476, n7610, new_n2600);
not_8  g02224(new_n2600, new_n2601);
and_8  g02225(n12925, n12648, new_n2602);
and_8  g02226(n8476, n4826, new_n2603);
or_8   g02227(new_n2603, new_n2602, new_n2604);
and_8  g02228(n7733, n2530, new_n2605);
xnor_4 g02229(new_n2603, new_n2602, new_n2606);
or_8   g02230(new_n2606, new_n2605, new_n2607);
and_8  g02231(new_n2607, new_n2604, new_n2608);
and_8  g02232(new_n2608, new_n2601, new_n2609);
not_8  g02233(new_n2609, new_n2610);
xor_4  g02234(new_n2608, new_n2600, new_n2611);
xor_4  g02235(new_n2592, new_n2591, new_n2612);
or_8   g02236(new_n2612, new_n2611, new_n2613);
and_8  g02237(new_n2613, new_n2610, new_n2614);
xor_4  g02238(new_n2614, new_n2599, new_n2615);
and_8  g02239(n5331, n4970, new_n2616);
and_8  g02240(n7610, n5331, new_n2617);
and_8  g02241(n12925, n2530, new_n2618);
and_8  g02242(n5331, n4826, new_n2619);
or_8   g02243(new_n2619, new_n2618, new_n2620);
and_8  g02244(new_n2619, new_n2618, new_n2621);
and_8  g02245(n8476, n7733, new_n2622);
or_8   g02246(new_n2622, new_n2621, new_n2623);
and_8  g02247(new_n2623, new_n2620, new_n2624_1);
and_8  g02248(new_n2624_1, new_n2617, new_n2625);
xor_4  g02249(new_n2624_1, new_n2617, new_n2626);
nor_6  g02250(new_n2606, new_n2605, new_n2627);
and_8  g02251(new_n2606, new_n2605, new_n2628);
or_8   g02252(new_n2628, new_n2627, new_n2629);
and_8  g02253(new_n2629, new_n2626, new_n2630);
or_8   g02254(new_n2630, new_n2625, new_n2631);
nor_6  g02255(new_n2631, new_n2616, new_n2632);
xor_4  g02256(new_n2608, new_n2601, new_n2633);
xor_4  g02257(new_n2612, new_n2633, new_n2634);
xor_4  g02258(new_n2631, new_n2616, new_n2635);
and_8  g02259(new_n2635, new_n2634, new_n2636);
or_8   g02260(new_n2636, new_n2632, new_n2637);
or_8   g02261(new_n2637, new_n2615, new_n2638);
nand_5 g02262(new_n2598, new_n2595, new_n2639);
not_8  g02263(new_n2639, new_n2640);
nand_5 g02264(new_n2597, new_n2596, new_n2641);
not_8  g02265(new_n2641, new_n2642);
not_8  g02266(new_n2612, new_n2643);
and_8  g02267(new_n2643, new_n2633, new_n2644);
or_8   g02268(new_n2644, new_n2609, new_n2645);
and_8  g02269(new_n2645, new_n2599, new_n2646);
xor_4  g02270(new_n2646, new_n2642, new_n2647);
or_8   g02271(new_n2647, new_n2640, new_n2648);
and_8  g02272(new_n2582, new_n2581_1, new_n2649);
and_8  g02273(n12648, n7610, new_n2650);
xnor_4 g02274(new_n2650, new_n2649, new_n2651);
and_8  g02275(n7733, n7690, new_n2652);
and_8  g02276(n10545, n4826, new_n2653);
and_8  g02277(n12925, n3616, new_n2654);
xnor_4 g02278(new_n2654, new_n2653, new_n2655);
xor_4  g02279(new_n2655, new_n2652, new_n2656);
xor_4  g02280(new_n2656, new_n2651, new_n2657);
nand_5 g02281(new_n2583, new_n2580, new_n2658);
or_8   g02282(new_n2594, new_n2586, new_n2659);
and_8  g02283(new_n2659, new_n2658, new_n2660);
and_8  g02284(n8476, n503, new_n2661);
and_8  g02285(n4970, n2530, new_n2662);
and_8  g02286(n10965, n5331, new_n2663);
xnor_4 g02287(new_n2663, new_n2662, new_n2664);
xor_4  g02288(new_n2664, new_n2661, new_n2665);
xor_4  g02289(new_n2665, new_n2660, new_n2666);
xor_4  g02290(new_n2666, new_n2657, new_n2667);
and_8  g02291(new_n2667, new_n2648, new_n2668);
xor_4  g02292(new_n2646, new_n2641, new_n2669);
and_8  g02293(new_n2669, new_n2639, new_n2670);
not_8  g02294(new_n2667, new_n2671);
and_8  g02295(new_n2671, new_n2670, new_n2672);
or_8   g02296(new_n2672, new_n2668, new_n2673);
nor_6  g02297(new_n2673, new_n2638, new_n2674);
and_8  g02298(new_n2673, new_n2638, new_n2675);
nor_6  g02299(new_n2675, new_n2674, new_n2676);
and_8  g02300(n5331, n503, new_n2677);
xor_4  g02301(new_n2645, new_n2599, new_n2678);
not_8  g02302(new_n2632, new_n2679_1);
xor_4  g02303(new_n2612, new_n2611, new_n2680);
and_8  g02304(new_n2631, new_n2616, new_n2681);
or_8   g02305(new_n2681, new_n2632, new_n2682);
or_8   g02306(new_n2682, new_n2680, new_n2683);
and_8  g02307(new_n2683, new_n2679_1, new_n2684);
or_8   g02308(new_n2684, new_n2678, new_n2685);
and_8  g02309(new_n2685, new_n2638, new_n2686);
and_8  g02310(new_n2686, new_n2677, new_n2687);
xor_4  g02311(new_n2629, new_n2626, new_n2688);
not_8  g02312(n12925, new_n2689);
or_8   g02313(new_n2689, new_n695, new_n2690);
and_8  g02314(new_n2690, new_n2622, new_n2691);
nor_6  g02315(new_n2691, new_n2620, new_n2692);
or_8   g02316(new_n2692, new_n2621, new_n2693);
and_8  g02317(new_n2693, new_n2622, new_n2694);
and_8  g02318(new_n2694, new_n2688, new_n2695);
not_8  g02319(new_n2695, new_n2696);
xor_4  g02320(new_n2635, new_n2634, new_n2697);
nor_6  g02321(new_n2697, new_n2696, new_n2698);
xor_4  g02322(new_n2686, new_n2677, new_n2699);
and_8  g02323(new_n2699, new_n2698, new_n2700);
or_8   g02324(new_n2700, new_n2687, new_n2701);
and_8  g02325(new_n2701, new_n2676, new_n2702);
or_8   g02326(new_n2675, new_n2674, new_n2703);
not_8  g02327(new_n2687, new_n2704);
or_8   g02328(new_n2697, new_n2696, new_n2705);
not_8  g02329(new_n2677, new_n2706);
xor_4  g02330(new_n2686, new_n2706, new_n2707);
or_8   g02331(new_n2707, new_n2705, new_n2708_1);
and_8  g02332(new_n2708_1, new_n2704, new_n2709);
and_8  g02333(new_n2709, new_n2703, new_n2710);
or_8   g02334(new_n2710, new_n2702, new_n2711);
and_8  g02335(n4086, n2393, new_n2712);
and_8  g02336(n5860, n405, new_n2713);
and_8  g02337(n8433, n3986, new_n2714);
xor_4  g02338(new_n2714, new_n2713, new_n2715);
xor_4  g02339(new_n2715, new_n2712, new_n2716);
and_8  g02340(n8433, n5860, new_n2717);
and_8  g02341(n11892, n4086, new_n2718);
or_8   g02342(new_n2718, new_n2717, new_n2719);
and_8  g02343(n2393, n405, new_n2720);
xnor_4 g02344(new_n2718, new_n2717, new_n2721);
or_8   g02345(new_n2721, new_n2720, new_n2722);
and_8  g02346(new_n2722, new_n2719, new_n2723);
and_8  g02347(new_n2723, new_n2716, new_n2724);
nor_6  g02348(new_n2723, new_n2716, new_n2725);
or_8   g02349(new_n2725, new_n2724, new_n2726);
and_8  g02350(n7388, n6611, new_n2727);
and_8  g02351(n11892, n217, new_n2728);
xor_4  g02352(new_n2728, new_n2727, new_n2729);
not_8  g02353(new_n2729, new_n2730);
or_8   g02354(new_n2730, new_n2726, new_n2731);
xor_4  g02355(new_n2723, new_n2716, new_n2732);
or_8   g02356(new_n2729, new_n2732, new_n2733);
and_8  g02357(new_n2733, new_n2731, new_n2734);
and_8  g02358(n7388, n217, new_n2735);
and_8  g02359(n8433, n2393, new_n2736);
and_8  g02360(n7388, n4086, new_n2737);
or_8   g02361(new_n2737, new_n2736, new_n2738);
and_8  g02362(n11892, n405, new_n2739);
nor_6  g02363(new_n2737, new_n2736, new_n2740);
and_8  g02364(new_n2737, new_n2736, new_n2741);
or_8   g02365(new_n2741, new_n2740, new_n2742);
or_8   g02366(new_n2742, new_n2739, new_n2743);
and_8  g02367(new_n2743, new_n2738, new_n2744);
and_8  g02368(new_n2744, new_n2735, new_n2745);
xor_4  g02369(new_n2744, new_n2735, new_n2746);
not_8  g02370(n405, new_n2747);
not_8  g02371(n2393, new_n2748);
or_8   g02372(new_n2748, new_n2747, new_n2749_1);
xor_4  g02373(new_n2721, new_n2749_1, new_n2750);
and_8  g02374(new_n2750, new_n2746, new_n2751);
or_8   g02375(new_n2751, new_n2745, new_n2752);
and_8  g02376(new_n2752, new_n2734, new_n2753);
nor_6  g02377(new_n2752, new_n2734, new_n2754);
or_8   g02378(new_n2754, new_n2753, new_n2755);
and_8  g02379(n7965, n6611, new_n2756);
not_8  g02380(new_n2756, new_n2757);
nor_6  g02381(new_n2744, new_n2735, new_n2758);
or_8   g02382(new_n2758, new_n2745, new_n2759);
xor_4  g02383(new_n2721, new_n2720, new_n2760);
and_8  g02384(new_n2760, new_n2759, new_n2761);
or_8   g02385(new_n2761, new_n2751, new_n2762);
or_8   g02386(new_n2762, new_n2757, new_n2763);
xor_4  g02387(new_n2762, new_n2756, new_n2764);
and_8  g02388(n7965, n217, new_n2765);
and_8  g02389(n11892, n8433, new_n2766);
and_8  g02390(n7965, n4086, new_n2767);
and_8  g02391(new_n2767, new_n2766, new_n2768);
or_8   g02392(new_n2767, new_n2766, new_n2769);
and_8  g02393(n7388, n405, new_n2770);
and_8  g02394(new_n2770, new_n2769, new_n2771);
or_8   g02395(new_n2771, new_n2768, new_n2772);
and_8  g02396(new_n2772, new_n2765, new_n2773);
xor_4  g02397(new_n2772, new_n2765, new_n2774);
xnor_4 g02398(new_n2742, new_n2739, new_n2775);
and_8  g02399(new_n2775, new_n2774, new_n2776);
or_8   g02400(new_n2776, new_n2773, new_n2777);
not_8  g02401(new_n2777, new_n2778);
or_8   g02402(new_n2778, new_n2764, new_n2779);
and_8  g02403(new_n2779, new_n2763, new_n2780);
or_8   g02404(new_n2780, new_n2755, new_n2781);
and_8  g02405(new_n2728, new_n2727, new_n2782);
and_8  g02406(new_n2753, new_n2782, new_n2783);
nor_6  g02407(new_n2753, new_n2782, new_n2784);
or_8   g02408(new_n2784, new_n2783, new_n2785);
and_8  g02409(new_n2785, new_n2731, new_n2786);
not_8  g02410(new_n2786, new_n2787);
and_8  g02411(new_n2714, new_n2713, new_n2788);
and_8  g02412(n2393, n217, new_n2789);
xnor_4 g02413(new_n2789, new_n2788, new_n2790);
and_8  g02414(n3986, n405, new_n2791);
and_8  g02415(n5860, n4086, new_n2792);
and_8  g02416(n8433, n5857, new_n2793);
xnor_4 g02417(new_n2793, new_n2792, new_n2794);
xor_4  g02418(new_n2794, new_n2791, new_n2795);
xnor_4 g02419(new_n2795, new_n2790, new_n2796);
and_8  g02420(new_n2715, new_n2712, new_n2797);
nor_6  g02421(new_n2724, new_n2797, new_n2798);
and_8  g02422(n11296, n7965, new_n2799);
and_8  g02423(n11892, n6611, new_n2800);
and_8  g02424(n7388, n6359, new_n2801);
xnor_4 g02425(new_n2801, new_n2800, new_n2802_1);
xor_4  g02426(new_n2802_1, new_n2799, new_n2803);
xor_4  g02427(new_n2803, new_n2798, new_n2804);
nor_6  g02428(new_n2804, new_n2796, new_n2805);
and_8  g02429(new_n2804, new_n2796, new_n2806);
or_8   g02430(new_n2806, new_n2805, new_n2807);
and_8  g02431(new_n2807, new_n2787, new_n2808);
not_8  g02432(new_n2807, new_n2809);
and_8  g02433(new_n2809, new_n2786, new_n2810);
or_8   g02434(new_n2810, new_n2808, new_n2811);
or_8   g02435(new_n2811, new_n2781, new_n2812);
xor_4  g02436(new_n2752, new_n2734, new_n2813);
nor_6  g02437(new_n2762, new_n2757, new_n2814);
xor_4  g02438(new_n2762, new_n2757, new_n2815);
and_8  g02439(new_n2777, new_n2815, new_n2816);
or_8   g02440(new_n2816, new_n2814, new_n2817);
and_8  g02441(new_n2817, new_n2813, new_n2818_1);
or_8   g02442(new_n2809, new_n2786, new_n2819);
or_8   g02443(new_n2807, new_n2787, new_n2820);
and_8  g02444(new_n2820, new_n2819, new_n2821);
or_8   g02445(new_n2821, new_n2818_1, new_n2822);
and_8  g02446(new_n2822, new_n2812, new_n2823);
and_8  g02447(n7965, n6359, new_n2824);
not_8  g02448(new_n2824, new_n2825);
and_8  g02449(new_n2780, new_n2755, new_n2826);
or_8   g02450(new_n2826, new_n2818_1, new_n2827);
or_8   g02451(new_n2827, new_n2825, new_n2828);
nor_6  g02452(new_n2775, new_n2774, new_n2829);
or_8   g02453(new_n2829, new_n2776, new_n2830);
xnor_4 g02454(new_n2767, new_n2766, new_n2831);
and_8  g02455(n8433, n7388, new_n2832);
and_8  g02456(n7965, n405, new_n2833);
and_8  g02457(new_n2833, new_n2832, new_n2834);
nand_5 g02458(new_n2834, new_n2831, new_n2835);
or_8   g02459(new_n2835, new_n2830, new_n2836);
xor_4  g02460(new_n2778, new_n2815, new_n2837);
or_8   g02461(new_n2837, new_n2836, new_n2838);
or_8   g02462(new_n2817, new_n2813, new_n2839);
and_8  g02463(new_n2839, new_n2781, new_n2840);
and_8  g02464(new_n2840, new_n2824, new_n2841);
and_8  g02465(new_n2827, new_n2825, new_n2842);
or_8   g02466(new_n2842, new_n2841, new_n2843);
or_8   g02467(new_n2843, new_n2838, new_n2844);
and_8  g02468(new_n2844, new_n2828, new_n2845);
xor_4  g02469(new_n2845, new_n2823, new_n2846);
and_8  g02470(new_n2846, new_n2711, new_n2847);
or_8   g02471(new_n2709, new_n2703, new_n2848);
or_8   g02472(new_n2701, new_n2676, new_n2849);
and_8  g02473(new_n2849, new_n2848, new_n2850);
not_8  g02474(new_n2838, new_n2851);
or_8   g02475(new_n2840, new_n2824, new_n2852);
and_8  g02476(new_n2852, new_n2828, new_n2853);
and_8  g02477(new_n2853, new_n2851, new_n2854);
or_8   g02478(new_n2854, new_n2841, new_n2855);
xor_4  g02479(new_n2855, new_n2823, new_n2856);
and_8  g02480(new_n2856, new_n2850, new_n2857);
or_8   g02481(new_n2857, new_n2847, new_n2858);
or_8   g02482(new_n2699, new_n2698, new_n2859);
and_8  g02483(new_n2859, new_n2708_1, new_n2860);
xor_4  g02484(new_n2853, new_n2851, new_n2861);
or_8   g02485(new_n2861, new_n2860, new_n2862);
not_8  g02486(new_n2836, new_n2863);
xor_4  g02487(new_n2778, new_n2764, new_n2864);
or_8   g02488(new_n2864, new_n2863, new_n2865);
and_8  g02489(new_n2865, new_n2838, new_n2866);
nor_6  g02490(new_n2694, new_n2688, new_n2867);
or_8   g02491(new_n2867, new_n2695, new_n2868);
not_8  g02492(new_n2868, new_n2869);
xor_4  g02493(new_n2835, new_n2830, new_n2870);
or_8   g02494(new_n2870, new_n2869, new_n2871);
and_8  g02495(n12925, n5331, new_n2872);
and_8  g02496(n8433, n7965, new_n2873);
and_8  g02497(new_n2873, new_n2872, new_n2874);
xor_4  g02498(new_n2833, new_n2832, new_n2875);
or_8   g02499(new_n2875, new_n2874, new_n2876);
xnor_4 g02500(new_n2875, new_n2874, new_n2877);
and_8  g02501(n12925, n8476, new_n2878);
and_8  g02502(n7733, n5331, new_n2879_1);
xor_4  g02503(new_n2879_1, new_n2878, new_n2880);
or_8   g02504(new_n2880, new_n2877, new_n2881);
and_8  g02505(new_n2881, new_n2876, new_n2882);
and_8  g02506(new_n2691, new_n2620, new_n2883);
nor_6  g02507(new_n2883, new_n2693, new_n2884);
or_8   g02508(new_n2884, new_n2882, new_n2885);
or_8   g02509(new_n2883, new_n2693, new_n2886);
xor_4  g02510(new_n2886, new_n2882, new_n2887);
not_8  g02511(new_n2873, new_n2888);
nand_5 g02512(new_n2888, new_n2770, new_n2889);
nand_5 g02513(new_n2889, new_n2831, new_n2890);
not_8  g02514(new_n2889, new_n2891);
nand_5 g02515(new_n2891, new_n2769, new_n2892);
and_8  g02516(new_n2892, new_n2890, new_n2893);
or_8   g02517(new_n2893, new_n2887, new_n2894);
and_8  g02518(new_n2894, new_n2885, new_n2895);
not_8  g02519(new_n2870, new_n2896);
xor_4  g02520(new_n2896, new_n2869, new_n2897);
or_8   g02521(new_n2897, new_n2895, new_n2898);
and_8  g02522(new_n2898, new_n2871, new_n2899);
nor_6  g02523(new_n2899, new_n2866, new_n2900);
xor_4  g02524(new_n2697, new_n2695, new_n2901);
xor_4  g02525(new_n2899, new_n2866, new_n2902_1);
and_8  g02526(new_n2902_1, new_n2901, new_n2903);
nor_6  g02527(new_n2903, new_n2900, new_n2904);
and_8  g02528(new_n2707, new_n2705, new_n2905);
or_8   g02529(new_n2905, new_n2700, new_n2906);
xor_4  g02530(new_n2853, new_n2838, new_n2907);
and_8  g02531(new_n2907, new_n2906, new_n2908);
and_8  g02532(new_n2861, new_n2860, new_n2909);
or_8   g02533(new_n2909, new_n2908, new_n2910);
or_8   g02534(new_n2910, new_n2904, new_n2911);
and_8  g02535(new_n2911, new_n2862, new_n2912);
or_8   g02536(new_n2912, new_n2858, new_n2913);
or_8   g02537(new_n2856, new_n2850, new_n2914);
or_8   g02538(new_n2846, new_n2711, new_n2915);
and_8  g02539(new_n2915, new_n2914, new_n2916);
or_8   g02540(new_n2903, new_n2900, new_n2917);
or_8   g02541(new_n2907, new_n2906, new_n2918);
and_8  g02542(new_n2918, new_n2862, new_n2919);
and_8  g02543(new_n2919, new_n2917, new_n2920);
or_8   g02544(new_n2920, new_n2908, new_n2921);
or_8   g02545(new_n2921, new_n2916, new_n2922);
and_8  g02546(new_n2922, new_n2913, new_n2923);
xor_4  g02547(new_n2923, new_n2579, new_n2924);
not_8  g02548(new_n2537, new_n2925);
xor_4  g02549(new_n2542, new_n2455, new_n2926);
xor_4  g02550(new_n2926, new_n2925, new_n2927);
not_8  g02551(new_n2927, new_n2928);
or_8   g02552(new_n2919, new_n2917, new_n2929);
and_8  g02553(new_n2929, new_n2911, new_n2930);
and_8  g02554(new_n2930, new_n2928, new_n2931);
and_8  g02555(new_n2910, new_n2904, new_n2932);
or_8   g02556(new_n2932, new_n2920, new_n2933);
or_8   g02557(new_n2933, new_n2927, new_n2934);
or_8   g02558(new_n2930, new_n2928, new_n2935);
and_8  g02559(new_n2935, new_n2934, new_n2936);
xor_4  g02560(new_n2536, new_n2533, new_n2937);
not_8  g02561(new_n2937, new_n2938);
not_8  g02562(new_n2901, new_n2939);
and_8  g02563(new_n2899, new_n2866, new_n2940);
or_8   g02564(new_n2940, new_n2900, new_n2941);
or_8   g02565(new_n2941, new_n2939, new_n2942);
or_8   g02566(new_n2902_1, new_n2901, new_n2943);
and_8  g02567(new_n2943, new_n2942, new_n2944);
or_8   g02568(new_n2944, new_n2938, new_n2945);
xor_4  g02569(new_n2944, new_n2937, new_n2946);
xor_4  g02570(new_n2532, new_n2526, new_n2947);
xor_4  g02571(new_n2896, new_n2868, new_n2948);
xor_4  g02572(new_n2948, new_n2895, new_n2949);
and_8  g02573(new_n2949, new_n2947, new_n2950);
not_8  g02574(new_n2950, new_n2951);
nor_6  g02575(new_n2949, new_n2947, new_n2952);
or_8   g02576(new_n2952, new_n2950, new_n2953);
xor_4  g02577(new_n2893, new_n2887, new_n2954);
and_8  g02578(n8759, n3719, new_n2955);
not_8  g02579(new_n2955, new_n2956);
and_8  g02580(new_n2956, new_n2512_1, new_n2957);
not_8  g02581(new_n2957, new_n2958);
and_8  g02582(new_n2958, new_n2527, new_n2959);
and_8  g02583(new_n2957, new_n2511, new_n2960);
or_8   g02584(new_n2960, new_n2959, new_n2961);
nor_6  g02585(new_n2961, new_n2954, new_n2962);
not_8  g02586(new_n2962, new_n2963);
and_8  g02587(new_n2961, new_n2954, new_n2964);
or_8   g02588(new_n2964, new_n2962, new_n2965);
xnor_4 g02589(new_n2880, new_n2877, new_n2966);
xor_4  g02590(new_n2529, new_n2528, new_n2967);
and_8  g02591(new_n2967, new_n2966, new_n2968);
xor_4  g02592(new_n2873, new_n2872, new_n2969);
and_8  g02593(new_n2969, new_n2955, new_n2970);
xor_4  g02594(new_n2967, new_n2966, new_n2971);
and_8  g02595(new_n2971, new_n2970, new_n2972);
or_8   g02596(new_n2972, new_n2968, new_n2973);
not_8  g02597(new_n2973, new_n2974);
or_8   g02598(new_n2974, new_n2965, new_n2975);
and_8  g02599(new_n2975, new_n2963, new_n2976);
or_8   g02600(new_n2976, new_n2953, new_n2977);
and_8  g02601(new_n2977, new_n2951, new_n2978);
or_8   g02602(new_n2978, new_n2946, new_n2979);
and_8  g02603(new_n2979, new_n2945, new_n2980);
and_8  g02604(new_n2980, new_n2936, new_n2981);
nor_6  g02605(new_n2981, new_n2931, new_n2982);
and_8  g02606(new_n2982, new_n2924, new_n2983);
xor_4  g02607(new_n2923, new_n2578, new_n2984);
or_8   g02608(new_n2981, new_n2931, new_n2985);
and_8  g02609(new_n2985, new_n2984, new_n2986);
or_8   g02610(new_n2986, new_n2983, new_n2987);
or_8   g02611(new_n2987, new_n2454, new_n2988);
or_8   g02612(new_n2985, new_n2984, new_n2989);
or_8   g02613(new_n2982, new_n2924, new_n2990);
and_8  g02614(new_n2990, new_n2989, new_n2991);
and_8  g02615(new_n2991, new_n2453, new_n2992);
and_8  g02616(new_n2987, new_n2454, new_n2993);
or_8   g02617(new_n2993, new_n2992, new_n2994);
xor_4  g02618(new_n2450, new_n2449, new_n2995);
and_8  g02619(new_n2933, new_n2927, new_n2996);
or_8   g02620(new_n2996, new_n2931, new_n2997);
xor_4  g02621(new_n2980, new_n2997, new_n2998);
and_8  g02622(new_n2998, new_n2995, new_n2999);
not_8  g02623(new_n2999, new_n3000);
xor_4  g02624(new_n2448, new_n2447, new_n3001);
xor_4  g02625(new_n2944, new_n2938, new_n3002);
nor_6  g02626(new_n2976, new_n2953, new_n3003);
or_8   g02627(new_n3003, new_n2950, new_n3004);
or_8   g02628(new_n3004, new_n3002, new_n3005);
and_8  g02629(new_n3005, new_n2979, new_n3006);
nor_6  g02630(new_n3006, new_n3001, new_n3007);
xor_4  g02631(new_n3006, new_n3001, new_n3008);
xor_4  g02632(new_n2446, new_n2440, new_n3009);
and_8  g02633(new_n2976, new_n2953, new_n3010);
or_8   g02634(new_n3010, new_n3003, new_n3011);
and_8  g02635(new_n3011, new_n3009, new_n3012);
not_8  g02636(new_n2965, new_n3013);
xor_4  g02637(new_n2973, new_n3013, new_n3014);
and_8  g02638(n9956, n5305, new_n3015);
not_8  g02639(new_n3015, new_n3016);
nand_5 g02640(new_n3016, new_n2399, new_n3017);
not_8  g02641(new_n3017, new_n3018);
nor_6  g02642(new_n3018, new_n2442, new_n3019);
not_8  g02643(new_n3019, new_n3020);
nand_5 g02644(new_n3018, new_n2398, new_n3021);
nand_5 g02645(new_n3021, new_n3020, new_n3022_1);
not_8  g02646(new_n3022_1, new_n3023);
or_8   g02647(new_n3023, new_n3014, new_n3024);
nor_6  g02648(new_n3023, new_n3014, new_n3025);
and_8  g02649(new_n3023, new_n3014, new_n3026);
or_8   g02650(new_n3026, new_n3025, new_n3027);
xor_4  g02651(new_n2969, new_n2955, new_n3028);
and_8  g02652(new_n3028, new_n3015, new_n3029);
xor_4  g02653(new_n2444, new_n2443, new_n3030);
or_8   g02654(new_n3030, new_n3029, new_n3031);
xor_4  g02655(new_n2971, new_n2970, new_n3032);
xnor_4 g02656(new_n3030, new_n3029, new_n3033);
or_8   g02657(new_n3033, new_n3032, new_n3034);
and_8  g02658(new_n3034, new_n3031, new_n3035);
or_8   g02659(new_n3035, new_n3027, new_n3036);
and_8  g02660(new_n3036, new_n3024, new_n3037);
not_8  g02661(new_n3009, new_n3038);
xor_4  g02662(new_n2976, new_n2953, new_n3039);
and_8  g02663(new_n3039, new_n3038, new_n3040);
or_8   g02664(new_n3040, new_n3012, new_n3041);
nor_6  g02665(new_n3041, new_n3037, new_n3042);
or_8   g02666(new_n3042, new_n3012, new_n3043);
and_8  g02667(new_n3043, new_n3008, new_n3044);
or_8   g02668(new_n3044, new_n3007, new_n3045);
not_8  g02669(new_n2995, new_n3046);
xor_4  g02670(new_n2980, new_n2936, new_n3047);
and_8  g02671(new_n3047, new_n3046, new_n3048);
or_8   g02672(new_n3048, new_n2999, new_n3049);
or_8   g02673(new_n3049, new_n3045, new_n3050);
and_8  g02674(new_n3050, new_n3000, new_n3051);
or_8   g02675(new_n3051, new_n2994, new_n3052);
and_8  g02676(new_n3052, new_n2988, new_n3053);
nor_6  g02677(new_n2923, new_n2579, new_n3054);
or_8   g02678(new_n2983, new_n3054, new_n3055);
nand_5 g02679(new_n2650, new_n2649, new_n3056);
or_8   g02680(new_n2656, new_n2651, new_n3057);
and_8  g02681(new_n3057, new_n3056, new_n3058);
or_8   g02682(new_n2654, new_n2653, new_n3059);
or_8   g02683(new_n2655, new_n2652, new_n3060);
and_8  g02684(new_n3060, new_n3059, new_n3061);
not_8  g02685(n4970, new_n3062);
or_8   g02686(new_n702, new_n3062, new_n3063);
and_8  g02687(n11296, n7388, new_n3064);
and_8  g02688(n9241, n6126, new_n3065);
xor_4  g02689(new_n3065, new_n3064, new_n3066);
xor_4  g02690(new_n3066, new_n3063, new_n3067);
xor_4  g02691(new_n3067, new_n3061, new_n3068);
xor_4  g02692(new_n3068, new_n3058, new_n3069);
or_8   g02693(new_n2793, new_n2792, new_n3070);
or_8   g02694(new_n2794, new_n2791, new_n3071_1);
and_8  g02695(new_n3071_1, new_n3070, new_n3072);
or_8   g02696(new_n2801, new_n2800, new_n3073);
or_8   g02697(new_n2802_1, new_n2799, new_n3074);
and_8  g02698(new_n3074, new_n3073, new_n3075);
xor_4  g02699(new_n3075, new_n3072, new_n3076);
and_8  g02700(n11892, n6359, new_n3077);
and_8  g02701(n7546, n5331, new_n3078);
xor_4  g02702(new_n3078, new_n3077, new_n3079);
xor_4  g02703(new_n3079, new_n3076, new_n3080);
nand_5 g02704(new_n2559, new_n2558_1, new_n3081);
or_8   g02705(new_n2565, new_n2560, new_n3082);
and_8  g02706(new_n3082, new_n3081, new_n3083);
and_8  g02707(n8595, n8276, new_n3084);
and_8  g02708(n6611, n2393, new_n3085);
xor_4  g02709(new_n3085, new_n3084, new_n3086);
and_8  g02710(n12925, n4499, new_n3087);
and_8  g02711(n11536, n5305, new_n3088);
xor_4  g02712(new_n3088, new_n3087, new_n3089);
xnor_4 g02713(new_n3089, new_n3086, new_n3090);
xor_4  g02714(new_n3090, new_n3083, new_n3091);
xor_4  g02715(new_n3091, new_n3080, new_n3092);
nand_5 g02716(new_n2789, new_n2788, new_n3093);
or_8   g02717(new_n2795, new_n2790, new_n3094);
and_8  g02718(new_n3094, new_n3093, new_n3095);
or_8   g02719(new_n2663, new_n2662, new_n3096);
or_8   g02720(new_n2664, new_n2661, new_n3097);
and_8  g02721(new_n3097, new_n3096, new_n3098);
and_8  g02722(n4086, n3986, new_n3099);
and_8  g02723(n7733, n3616, new_n3100);
xor_4  g02724(new_n3100, new_n3099, new_n3101);
xor_4  g02725(new_n3101, new_n3098, new_n3102);
xor_4  g02726(new_n3102, new_n3095, new_n3103);
xor_4  g02727(new_n3103, new_n3092, new_n3104);
xor_4  g02728(new_n3104, new_n3069, new_n3105);
and_8  g02729(new_n2821, new_n2818_1, new_n3106);
and_8  g02730(new_n2855, new_n2823, new_n3107);
or_8   g02731(new_n3107, new_n3106, new_n3108);
nand_5 g02732(n5860, n217, new_n3109);
not_8  g02733(new_n3109, new_n3110);
xor_4  g02734(new_n3110, new_n3108, new_n3111);
and_8  g02735(new_n2542, new_n2455, new_n3112);
and_8  g02736(new_n2926, new_n2925, new_n3113);
or_8   g02737(new_n3113, new_n3112, new_n3114);
nor_6  g02738(new_n2576, new_n2574, new_n3115);
and_8  g02739(new_n3115, new_n3114, new_n3116);
or_8   g02740(new_n3116, new_n2574, new_n3117);
nor_6  g02741(new_n2665, new_n2660, new_n3118);
and_8  g02742(new_n2666, new_n2657, new_n3119);
or_8   g02743(new_n3119, new_n3118, new_n3120);
and_8  g02744(n12299, n8065, new_n3121);
and_8  g02745(n10510, n3602, new_n3122);
xor_4  g02746(new_n3122, new_n3121, new_n3123);
and_8  g02747(n10644, n3719, new_n3124_1);
and_8  g02748(n7965, n1357, new_n3125);
xor_4  g02749(new_n3125, new_n3124_1, new_n3126);
and_8  g02750(n10439, n7436, new_n3127);
and_8  g02751(n8759, n4190, new_n3128);
xor_4  g02752(new_n3128, new_n3127, new_n3129);
xnor_4 g02753(new_n3129, new_n3126, new_n3130);
xor_4  g02754(new_n3130, new_n3123, new_n3131);
or_8   g02755(new_n2416, new_n2415, new_n3132);
or_8   g02756(new_n2417, new_n2414, new_n3133);
and_8  g02757(new_n3133, new_n3132, new_n3134);
and_8  g02758(n9637, n1097, new_n3135);
xor_4  g02759(new_n3135, new_n3134, new_n3136);
xor_4  g02760(new_n3136, new_n3131, new_n3137);
xor_4  g02761(new_n3137, new_n3120, new_n3138);
not_8  g02762(new_n2555, new_n3139);
or_8   g02763(new_n2566, new_n2557, new_n3140);
and_8  g02764(new_n3140, new_n3139, new_n3141);
and_8  g02765(new_n2418, new_n2413, new_n3142);
and_8  g02766(new_n2428, new_n2419, new_n3143);
or_8   g02767(new_n3143, new_n3142, new_n3144);
xor_4  g02768(new_n3144, new_n3141, new_n3145);
xor_4  g02769(new_n3145, new_n3138, new_n3146_1);
and_8  g02770(new_n2494, new_n2570, new_n3147);
and_8  g02771(new_n2572, new_n2568, new_n3148);
or_8   g02772(new_n3148, new_n3147, new_n3149);
or_8   g02773(new_n2552, new_n2551_1, new_n3150);
or_8   g02774(new_n2553, new_n2550, new_n3151);
and_8  g02775(new_n3151, new_n3150, new_n3152);
and_8  g02776(n4312, n2577, new_n3153);
xor_4  g02777(new_n3153, new_n3152, new_n3154);
and_8  g02778(new_n2563, new_n2562, new_n3155);
or_8   g02779(new_n2563, new_n2562, new_n3156);
and_8  g02780(new_n3156, new_n2561, new_n3157);
or_8   g02781(new_n3157, new_n3155, new_n3158);
and_8  g02782(n11257, n4921, new_n3159);
and_8  g02783(n12705, n3842, new_n3160);
xnor_4 g02784(new_n3160, new_n3159, new_n3161);
xor_4  g02785(new_n3161, new_n3158, new_n3162);
xor_4  g02786(new_n3162, new_n3154, new_n3163);
not_8  g02787(new_n3163, new_n3164);
and_8  g02788(n8433, n45, new_n3165);
and_8  g02789(n12025, n11917, new_n3166);
xor_4  g02790(new_n3166, new_n3165, new_n3167);
or_8   g02791(new_n2425_1, new_n2424, new_n3168);
not_8  g02792(new_n2423, new_n3169);
or_8   g02793(new_n2426, new_n3169, new_n3170);
and_8  g02794(new_n3170, new_n3168, new_n3171);
and_8  g02795(n5964, n1835, new_n3172_1);
and_8  g02796(n5857, n405, new_n3173);
xor_4  g02797(new_n3173, new_n3172_1, new_n3174);
not_8  g02798(new_n3174, new_n3175);
xor_4  g02799(new_n3175, new_n3171, new_n3176);
xor_4  g02800(new_n3176, new_n3167, new_n3177);
or_8   g02801(new_n2421, new_n2420, new_n3178);
or_8   g02802(new_n2427, new_n2422, new_n3179);
and_8  g02803(new_n3179, new_n3178, new_n3180);
and_8  g02804(n10391, n6776, new_n3181);
xor_4  g02805(new_n3181, new_n3180, new_n3182);
and_8  g02806(new_n3182, new_n3177, new_n3183);
nor_6  g02807(new_n3182, new_n3177, new_n3184);
or_8   g02808(new_n3184, new_n3183, new_n3185);
xor_4  g02809(new_n3185, new_n3164, new_n3186);
or_8   g02810(new_n3186, new_n3149, new_n3187);
nor_6  g02811(new_n3148, new_n3147, new_n3188);
xor_4  g02812(new_n3185, new_n3163, new_n3189);
or_8   g02813(new_n3189, new_n3188, new_n3190);
and_8  g02814(new_n3190, new_n3187, new_n3191);
xor_4  g02815(new_n3191, new_n3146_1, new_n3192);
or_8   g02816(new_n3192, new_n3117, new_n3193);
not_8  g02817(new_n2574, new_n3194);
or_8   g02818(new_n2577_1, new_n2545, new_n3195);
and_8  g02819(new_n3195, new_n3194, new_n3196);
and_8  g02820(new_n3191, new_n3146_1, new_n3197);
nor_6  g02821(new_n3191, new_n3146_1, new_n3198);
or_8   g02822(new_n3198, new_n3197, new_n3199);
or_8   g02823(new_n3199, new_n3196, new_n3200);
and_8  g02824(new_n3200, new_n3193, new_n3201);
or_8   g02825(new_n3201, new_n3111, new_n3202);
xor_4  g02826(new_n3109, new_n3108, new_n3203);
and_8  g02827(new_n3199, new_n3196, new_n3204);
and_8  g02828(new_n3192, new_n3117, new_n3205);
or_8   g02829(new_n3205, new_n3204, new_n3206);
or_8   g02830(new_n3206, new_n3203, new_n3207);
and_8  g02831(new_n3207, new_n3202, new_n3208);
xor_4  g02832(new_n3208, new_n3105, new_n3209);
and_8  g02833(new_n2913, new_n2914, new_n3210);
or_8   g02834(new_n2808, new_n2783, new_n3211);
not_8  g02835(new_n2431_1, new_n3212);
nand_5 g02836(new_n2432, new_n3212, new_n3213);
or_8   g02837(new_n2434_1, new_n2429, new_n3214_1);
and_8  g02838(new_n3214_1, new_n3213, new_n3215);
xor_4  g02839(new_n3215, new_n3211, new_n3216);
xor_4  g02840(new_n3216, new_n3210, new_n3217);
and_8  g02841(new_n3217, new_n3209, new_n3218);
not_8  g02842(new_n3105, new_n3219);
xor_4  g02843(new_n3208, new_n3219, new_n3220);
not_8  g02844(new_n3216, new_n3221);
xor_4  g02845(new_n3221, new_n3210, new_n3222);
and_8  g02846(new_n3222, new_n3220, new_n3223);
or_8   g02847(new_n3223, new_n3218, new_n3224);
or_8   g02848(new_n3224, new_n3055, new_n3225);
or_8   g02849(new_n2923, new_n2579, new_n3226);
and_8  g02850(new_n2989, new_n3226, new_n3227);
or_8   g02851(new_n3222, new_n3220, new_n3228);
or_8   g02852(new_n3217, new_n3209, new_n3229);
and_8  g02853(new_n3229, new_n3228, new_n3230_1);
or_8   g02854(new_n3230_1, new_n3227, new_n3231);
and_8  g02855(new_n3231, new_n3225, new_n3232);
or_8   g02856(new_n2702, new_n2674, new_n3233);
and_8  g02857(new_n2435, new_n2410, new_n3234);
and_8  g02858(new_n2452, new_n2436, new_n3235);
or_8   g02859(new_n3235, new_n3234, new_n3236);
xor_4  g02860(new_n3236, new_n3233, new_n3237);
and_8  g02861(new_n2646, new_n2642, new_n3238);
nor_6  g02862(new_n2668, new_n3238, new_n3239);
and_8  g02863(new_n2803, new_n2798, new_n3240);
or_8   g02864(new_n2806, new_n3240, new_n3241);
and_8  g02865(n10547, n9956, new_n3242);
and_8  g02866(n10965, n8476, new_n3243);
and_8  g02867(n7690, n4826, new_n3244);
xor_4  g02868(new_n3244, new_n3243, new_n3245);
and_8  g02869(n10545, n7610, new_n3246);
and_8  g02870(n2530, n503, new_n3247);
xnor_4 g02871(new_n3247, new_n3246, new_n3248);
xor_4  g02872(new_n3248, new_n3245, new_n3249);
xor_4  g02873(new_n3249, new_n3242, new_n3250);
xor_4  g02874(new_n3250, new_n3241, new_n3251);
xor_4  g02875(new_n3251, new_n3239, new_n3252);
xor_4  g02876(new_n3252, new_n3237, new_n3253);
xor_4  g02877(new_n3253, new_n3232, new_n3254);
and_8  g02878(new_n3254, new_n3053, new_n3255);
nor_6  g02879(new_n3051, new_n2994, new_n3256);
or_8   g02880(new_n3256, new_n2992, new_n3257);
nor_6  g02881(new_n3253, new_n3232, new_n3258);
and_8  g02882(new_n3253, new_n3232, new_n3259);
or_8   g02883(new_n3259, new_n3258, new_n3260);
and_8  g02884(new_n3260, new_n3257, new_n3261);
or_8   g02885(new_n3261, new_n3255, n837);
and_8  g02886(n11917, n11757, new_n3263);
and_8  g02887(n9956, n5240, new_n3264);
and_8  g02888(n11757, n4921, new_n3265);
and_8  g02889(n11917, n3172, new_n3266);
xnor_4 g02890(new_n3266, new_n3264, new_n3267);
or_8   g02891(new_n3267, new_n3265, new_n3268);
and_8  g02892(new_n3268, new_n3264, new_n3269);
nor_6  g02893(new_n3269, new_n3263, new_n3270);
and_8  g02894(n4921, n3172, new_n3271);
or_8   g02895(new_n3271, new_n3269, new_n3272_1);
and_8  g02896(new_n3272_1, new_n3263, new_n3273);
or_8   g02897(new_n3273, new_n3270, new_n3274);
and_8  g02898(n5240, n4921, new_n3275);
and_8  g02899(n11821, n9956, new_n3276);
xnor_4 g02900(new_n3276, new_n3275, new_n3277);
xor_4  g02901(new_n3277, new_n3274, new_n3278);
and_8  g02902(n2577, n1333, new_n3279);
and_8  g02903(n3842, n3172, new_n3280);
xor_4  g02904(new_n3280, new_n3279, new_n3281);
xor_4  g02905(new_n3281, new_n3278, new_n3282);
and_8  g02906(n3842, n1333, new_n3283);
and_8  g02907(n11757, n9956, new_n3284);
and_8  g02908(n11917, n1333, new_n3285);
or_8   g02909(new_n3285, new_n3284, new_n3286);
and_8  g02910(new_n3285, new_n3284, new_n3287_1);
or_8   g02911(new_n3287_1, new_n3271, new_n3288);
and_8  g02912(new_n3288, new_n3286, new_n3289);
and_8  g02913(new_n3289, new_n3283, new_n3290);
xnor_4 g02914(new_n3267, new_n3265, new_n3291);
xor_4  g02915(new_n3289, new_n3283, new_n3292);
and_8  g02916(new_n3292, new_n3291, new_n3293);
or_8   g02917(new_n3293, new_n3290, new_n3294);
xor_4  g02918(new_n3294, new_n3282, new_n3295);
and_8  g02919(n7862, n2577, new_n3296);
not_8  g02920(new_n3296, new_n3297);
nor_6  g02921(new_n3292, new_n3291, new_n3298);
or_8   g02922(new_n3298, new_n3293, new_n3299);
nor_6  g02923(new_n3299, new_n3297, new_n3300);
and_8  g02924(n7862, n3842, new_n3301);
and_8  g02925(n9956, n3172, new_n3302);
and_8  g02926(n11917, n7862, new_n3303);
and_8  g02927(new_n3303, new_n3302, new_n3304);
or_8   g02928(new_n3303, new_n3302, new_n3305);
and_8  g02929(n4921, n1333, new_n3306);
and_8  g02930(new_n3306, new_n3305, new_n3307);
or_8   g02931(new_n3307, new_n3304, new_n3308);
and_8  g02932(new_n3308, new_n3301, new_n3309);
xor_4  g02933(new_n3308, new_n3301, new_n3310);
xor_4  g02934(new_n3285, new_n3284, new_n3311);
xor_4  g02935(new_n3311, new_n3271, new_n3312);
and_8  g02936(new_n3312, new_n3310, new_n3313);
or_8   g02937(new_n3313, new_n3309, new_n3314);
xor_4  g02938(new_n3299, new_n3297, new_n3315);
and_8  g02939(new_n3315, new_n3314, new_n3316);
or_8   g02940(new_n3316, new_n3300, new_n3317);
and_8  g02941(new_n3317, new_n3295, new_n3318);
not_8  g02942(new_n3318, new_n3319);
not_8  g02943(new_n3273, new_n3320);
or_8   g02944(new_n3277, new_n3274, new_n3321);
and_8  g02945(new_n3321, new_n3320, new_n3322);
and_8  g02946(n9637, n1333, new_n3323);
and_8  g02947(n3172, n2577, new_n3324);
and_8  g02948(n7862, n1835, new_n3325);
xnor_4 g02949(new_n3325, new_n3324, new_n3326);
xor_4  g02950(new_n3326, new_n3323, new_n3327);
xor_4  g02951(new_n3327, new_n3322, new_n3328);
and_8  g02952(new_n3276, new_n3275, new_n3329);
and_8  g02953(n11757, n3842, new_n3330);
xnor_4 g02954(new_n3330, new_n3329, new_n3331);
and_8  g02955(n11821, n4921, new_n3332);
and_8  g02956(n9956, n9080, new_n3333);
and_8  g02957(n11917, n5240, new_n3334);
xnor_4 g02958(new_n3334, new_n3333, new_n3335);
xor_4  g02959(new_n3335, new_n3332, new_n3336);
xnor_4 g02960(new_n3336, new_n3331, new_n3337);
xor_4  g02961(new_n3337, new_n3328, new_n3338);
not_8  g02962(new_n3338, new_n3339_1);
nand_5 g02963(new_n3281, new_n3278, new_n3340);
nand_5 g02964(new_n3280, new_n3279, new_n3341);
and_8  g02965(new_n3294, new_n3282, new_n3342_1);
xor_4  g02966(new_n3342_1, new_n3341, new_n3343);
and_8  g02967(new_n3343, new_n3340, new_n3344);
xor_4  g02968(new_n3344, new_n3339_1, new_n3345);
and_8  g02969(new_n3345, new_n3319, new_n3346);
xor_4  g02970(new_n3344, new_n3338, new_n3347);
and_8  g02971(new_n3347, new_n3318, new_n3348);
or_8   g02972(new_n3348, new_n3346, new_n3349);
and_8  g02973(n9637, n7862, new_n3350);
not_8  g02974(new_n3350, new_n3351);
nor_6  g02975(new_n3317, new_n3295, new_n3352);
or_8   g02976(new_n3352, new_n3318, new_n3353);
or_8   g02977(new_n3353, new_n3351, new_n3354);
xor_4  g02978(new_n3312, new_n3310, new_n3355);
xor_4  g02979(new_n3303, new_n3302, new_n3356);
not_8  g02980(new_n3356, new_n3357);
and_8  g02981(n9956, n1333, new_n3358);
and_8  g02982(n7862, n4921, new_n3359);
and_8  g02983(new_n3359, new_n3358, new_n3360);
nand_5 g02984(new_n3360, new_n3357, new_n3361);
not_8  g02985(new_n3361, new_n3362);
and_8  g02986(new_n3362, new_n3355, new_n3363);
xor_4  g02987(new_n3315, new_n3314, new_n3364);
and_8  g02988(new_n3364, new_n3363, new_n3365);
not_8  g02989(new_n3365, new_n3366);
xor_4  g02990(new_n3317, new_n3295, new_n3367);
and_8  g02991(new_n3367, new_n3350, new_n3368);
and_8  g02992(new_n3353, new_n3351, new_n3369);
or_8   g02993(new_n3369, new_n3368, new_n3370);
or_8   g02994(new_n3370, new_n3366, new_n3371);
and_8  g02995(new_n3371, new_n3354, new_n3372);
xor_4  g02996(new_n3372, new_n3349, new_n3373);
or_8   g02997(new_n3367, new_n3350, new_n3374);
and_8  g02998(new_n3374, new_n3354, new_n3375);
xor_4  g02999(new_n3375, new_n3365, new_n3376);
and_8  g03000(n8595, n6877, new_n3377);
and_8  g03001(n6877, n6126, new_n3378);
and_8  g03002(n3719, n2464, new_n3379);
nor_6  g03003(new_n3379, new_n3378, new_n3380);
not_8  g03004(new_n3380, new_n3381);
and_8  g03005(n6877, n3719, new_n3382);
and_8  g03006(n6126, n2464, new_n3383);
and_8  g03007(new_n3383, new_n3382, new_n3384);
and_8  g03008(n9400, n3602, new_n3385);
or_8   g03009(new_n3385, new_n3384, new_n3386);
and_8  g03010(new_n3386, new_n3381, new_n3387);
xor_4  g03011(new_n3387, new_n3377, new_n3388);
and_8  g03012(n3602, n2464, new_n3389);
and_8  g03013(n9400, n6126, new_n3390);
and_8  g03014(n11311, n3719, new_n3391);
xor_4  g03015(new_n3391, new_n3390, new_n3392);
xor_4  g03016(new_n3392, new_n3389, new_n3393);
xnor_4 g03017(new_n3393, new_n3388, new_n3394);
not_8  g03018(new_n3385, new_n3395);
or_8   g03019(new_n3395, new_n3382, new_n3396);
or_8   g03020(new_n3384, new_n3380, new_n3397);
and_8  g03021(new_n3397, new_n3396, new_n3398);
not_8  g03022(new_n3398, new_n3399);
or_8   g03023(new_n3399, new_n3395, new_n3400);
nor_6  g03024(new_n3400, new_n3394, new_n3401);
nand_5 g03025(n10439, n6877, new_n3402);
and_8  g03026(n9400, n8595, new_n3403);
or_8   g03027(new_n3391, new_n3390, new_n3404);
and_8  g03028(new_n3391, new_n3390, new_n3405);
or_8   g03029(new_n3405, new_n3389, new_n3406);
and_8  g03030(new_n3406, new_n3404, new_n3407);
xnor_4 g03031(new_n3407, new_n3403, new_n3408);
and_8  g03032(n11311, n3602, new_n3409);
and_8  g03033(n4187, n3719, new_n3410);
xnor_4 g03034(new_n3410, new_n3383, new_n3411);
and_8  g03035(new_n3411, new_n3409, new_n3412);
nor_6  g03036(new_n3411, new_n3409, new_n3413);
or_8   g03037(new_n3413, new_n3412, new_n3414);
xor_4  g03038(new_n3414, new_n3408, new_n3415);
nor_6  g03039(new_n3415, new_n3402, new_n3416);
and_8  g03040(new_n3415, new_n3402, new_n3417);
or_8   g03041(new_n3417, new_n3416, new_n3418);
and_8  g03042(new_n3387, new_n3377, new_n3419);
and_8  g03043(new_n3393, new_n3388, new_n3420);
or_8   g03044(new_n3420, new_n3419, new_n3421);
not_8  g03045(new_n3421, new_n3422);
xor_4  g03046(new_n3422, new_n3418, new_n3423);
nand_5 g03047(new_n3423, new_n3401, new_n3424);
nand_5 g03048(n8065, n6877, new_n3425);
not_8  g03049(new_n3425, new_n3426);
and_8  g03050(n11311, n6126, new_n3427);
and_8  g03051(n4203, n3719, new_n3428);
and_8  g03052(n4187, n3602, new_n3429);
xor_4  g03053(new_n3429, new_n3428, new_n3430);
xor_4  g03054(new_n3430, new_n3427, new_n3431);
or_8   g03055(new_n3410, new_n3383, new_n3432);
or_8   g03056(new_n3411, new_n3409, new_n3433);
and_8  g03057(new_n3433, new_n3432, new_n3434);
xor_4  g03058(new_n3434, new_n3431, new_n3435);
and_8  g03059(n10439, n9400, new_n3436);
and_8  g03060(n8595, n2464, new_n3437);
xor_4  g03061(new_n3437, new_n3436, new_n3438);
xor_4  g03062(new_n3438, new_n3435, new_n3439);
and_8  g03063(new_n3407, new_n3403, new_n3440);
not_8  g03064(new_n3408, new_n3441);
and_8  g03065(new_n3414, new_n3441, new_n3442);
or_8   g03066(new_n3442, new_n3440, new_n3443);
and_8  g03067(new_n3443, new_n3439, new_n3444);
nor_6  g03068(new_n3443, new_n3439, new_n3445);
or_8   g03069(new_n3445, new_n3444, new_n3446);
nor_6  g03070(new_n3422, new_n3418, new_n3447);
nor_6  g03071(new_n3447, new_n3416, new_n3448);
or_8   g03072(new_n3448, new_n3446, new_n3449);
xor_4  g03073(new_n3443, new_n3439, new_n3450);
or_8   g03074(new_n3447, new_n3416, new_n3451);
or_8   g03075(new_n3451, new_n3450, new_n3452);
and_8  g03076(new_n3452, new_n3449, new_n3453);
xor_4  g03077(new_n3453, new_n3426, new_n3454);
nor_6  g03078(new_n3454, new_n3424, new_n3455);
and_8  g03079(new_n3454, new_n3424, new_n3456_1);
or_8   g03080(new_n3456_1, new_n3455, new_n3457);
xor_4  g03081(new_n3423, new_n3401, new_n3458);
xor_4  g03082(new_n3400, new_n3394, new_n3459);
or_8   g03083(new_n3396, new_n3380, new_n3460);
nand_5 g03084(new_n3460, new_n3399, new_n3461);
and_8  g03085(n8433, n7236, new_n3462);
and_8  g03086(n12925, n4805, new_n3463);
and_8  g03087(new_n3463, new_n3462, new_n3464);
and_8  g03088(n7733, n4805, new_n3465);
and_8  g03089(n12925, n11478, new_n3466);
xor_4  g03090(new_n3466, new_n3465, new_n3467);
nor_6  g03091(new_n3467, new_n3464, new_n3468);
xor_4  g03092(new_n3467, new_n3464, new_n3469);
and_8  g03093(n7236, n405, new_n3470);
and_8  g03094(n8433, n3992, new_n3471);
xnor_4 g03095(new_n3471, new_n3470, new_n3472);
and_8  g03096(new_n3472, new_n3469, new_n3473);
or_8   g03097(new_n3473, new_n3468, new_n3474);
and_8  g03098(n3992, n405, new_n3475);
not_8  g03099(new_n3475, new_n3476);
or_8   g03100(new_n3476, new_n3462, new_n3477);
and_8  g03101(n8433, n8384, new_n3478);
and_8  g03102(n7236, n4086, new_n3479);
or_8   g03103(new_n3479, new_n3478, new_n3480);
not_8  g03104(new_n3480, new_n3481);
and_8  g03105(new_n3481, new_n3477, new_n3482);
and_8  g03106(new_n3479, new_n3478, new_n3483);
or_8   g03107(new_n3483, new_n3482, new_n3484);
nor_6  g03108(new_n3481, new_n3477, new_n3485);
or_8   g03109(new_n3485, new_n3484, new_n3486);
xor_4  g03110(new_n3486, new_n3474, new_n3487);
and_8  g03111(n11478, n7733, new_n3488);
not_8  g03112(new_n3488, new_n3489);
or_8   g03113(new_n3489, new_n3463, new_n3490);
and_8  g03114(n12925, n5283, new_n3491);
and_8  g03115(n4826, n4805, new_n3492);
or_8   g03116(new_n3492, new_n3491, new_n3493);
or_8   g03117(new_n3493, new_n3490, new_n3494);
not_8  g03118(new_n3490, new_n3495);
xnor_4 g03119(new_n3492, new_n3491, new_n3496);
or_8   g03120(new_n3496, new_n3495, new_n3497);
and_8  g03121(new_n3497, new_n3494, new_n3498);
xor_4  g03122(new_n3498, new_n3487, new_n3499);
or_8   g03123(new_n3499, new_n3461, new_n3500);
not_8  g03124(new_n3500, new_n3501);
xor_4  g03125(new_n3499, new_n3461, new_n3502);
xnor_4 g03126(new_n3472, new_n3469, new_n3503);
and_8  g03127(n9400, n3719, new_n3504);
and_8  g03128(n6877, n3602, new_n3505);
xor_4  g03129(new_n3505, new_n3504, new_n3506);
and_8  g03130(new_n3506, new_n3503, new_n3507);
xor_4  g03131(new_n3463, new_n3462, new_n3508);
and_8  g03132(new_n3508, new_n3382, new_n3509);
xor_4  g03133(new_n3506, new_n3503, new_n3510);
and_8  g03134(new_n3510, new_n3509, new_n3511);
or_8   g03135(new_n3511, new_n3507, new_n3512);
and_8  g03136(new_n3512, new_n3502, new_n3513);
or_8   g03137(new_n3513, new_n3501, new_n3514);
or_8   g03138(new_n3514, new_n3459, new_n3515);
and_8  g03139(n7610, n4805, new_n3516);
and_8  g03140(new_n3492, new_n3491, new_n3517);
and_8  g03141(new_n3493, new_n3488, new_n3518);
or_8   g03142(new_n3518, new_n3517, new_n3519);
xnor_4 g03143(new_n3519, new_n3516, new_n3520);
and_8  g03144(n7733, n5283, new_n3521);
and_8  g03145(n12925, n137, new_n3522);
and_8  g03146(n11478, n4826, new_n3523);
xnor_4 g03147(new_n3523, new_n3522, new_n3524);
and_8  g03148(new_n3524, new_n3521, new_n3525);
or_8   g03149(new_n3524, new_n3521, new_n3526);
not_8  g03150(new_n3526, new_n3527);
or_8   g03151(new_n3527, new_n3525, new_n3528);
xor_4  g03152(new_n3528, new_n3520, new_n3529);
and_8  g03153(new_n3466, new_n3465, new_n3530);
nand_5 g03154(new_n3496, new_n3530, new_n3531);
xor_4  g03155(new_n3531, new_n3529, new_n3532);
and_8  g03156(n7236, n217, new_n3533);
or_8   g03157(new_n3483, new_n3475, new_n3534);
and_8  g03158(new_n3534, new_n3480, new_n3535);
xnor_4 g03159(new_n3535, new_n3533, new_n3536);
and_8  g03160(n8384, n405, new_n3537);
and_8  g03161(n8433, n6358, new_n3538);
and_8  g03162(n4086, n3992, new_n3539);
xnor_4 g03163(new_n3539, new_n3538, new_n3540);
and_8  g03164(new_n3540, new_n3537, new_n3541);
or_8   g03165(new_n3540, new_n3537, new_n3542);
not_8  g03166(new_n3542, new_n3543);
or_8   g03167(new_n3543, new_n3541, new_n3544);
xor_4  g03168(new_n3544, new_n3536, new_n3545);
nand_5 g03169(new_n3484, new_n3475, new_n3546);
xor_4  g03170(new_n3546, new_n3545, new_n3547);
and_8  g03171(new_n3547, new_n3532, new_n3548);
nor_6  g03172(new_n3531, new_n3529, new_n3549);
and_8  g03173(new_n3531, new_n3529, new_n3550);
or_8   g03174(new_n3550, new_n3549, new_n3551);
nor_6  g03175(new_n3546, new_n3545, new_n3552);
and_8  g03176(new_n3546, new_n3545, new_n3553);
or_8   g03177(new_n3553, new_n3552, new_n3554);
and_8  g03178(new_n3554, new_n3551, new_n3555);
or_8   g03179(new_n3555, new_n3548, new_n3556);
and_8  g03180(new_n3486, new_n3474, new_n3557);
and_8  g03181(new_n3498, new_n3487, new_n3558);
nor_6  g03182(new_n3558, new_n3557, new_n3559);
xnor_4 g03183(new_n3559, new_n3556, new_n3560);
xnor_4 g03184(new_n3400, new_n3394, new_n3561);
nor_6  g03185(new_n3498, new_n3487, new_n3562);
or_8   g03186(new_n3562, new_n3558, new_n3563);
xor_4  g03187(new_n3563, new_n3461, new_n3564);
nor_6  g03188(new_n3511, new_n3507, new_n3565);
or_8   g03189(new_n3565, new_n3564, new_n3566);
and_8  g03190(new_n3566, new_n3500, new_n3567);
and_8  g03191(new_n3567, new_n3561, new_n3568);
and_8  g03192(new_n3514, new_n3459, new_n3569);
or_8   g03193(new_n3569, new_n3568, new_n3570);
or_8   g03194(new_n3570, new_n3560, new_n3571);
and_8  g03195(new_n3571, new_n3515, new_n3572);
or_8   g03196(new_n3572, new_n3458, new_n3573);
and_8  g03197(new_n3572, new_n3458, new_n3574);
not_8  g03198(n6611, new_n3575);
not_8  g03199(n7236, new_n3576);
or_8   g03200(new_n3576, new_n3575, new_n3577);
and_8  g03201(n3992, n217, new_n3578);
or_8   g03202(new_n3539, new_n3538, new_n3579);
and_8  g03203(new_n3542, new_n3579, new_n3580);
and_8  g03204(new_n3580, new_n3578, new_n3581);
nor_6  g03205(new_n3580, new_n3578, new_n3582);
or_8   g03206(new_n3582, new_n3581, new_n3583);
and_8  g03207(n6358, n405, new_n3584);
and_8  g03208(n8384, n4086, new_n3585);
and_8  g03209(n8433, n5198, new_n3586);
xnor_4 g03210(new_n3586, new_n3585, new_n3587);
xor_4  g03211(new_n3587, new_n3584, new_n3588);
nor_6  g03212(new_n3588, new_n3583, new_n3589);
and_8  g03213(new_n3588, new_n3583, new_n3590);
or_8   g03214(new_n3590, new_n3589, new_n3591);
nor_6  g03215(new_n3591, new_n3577, new_n3592);
and_8  g03216(new_n3591, new_n3577, new_n3593);
or_8   g03217(new_n3593, new_n3592, new_n3594);
and_8  g03218(new_n3535, new_n3533, new_n3595);
not_8  g03219(new_n3536, new_n3596);
and_8  g03220(new_n3544, new_n3596, new_n3597);
nor_6  g03221(new_n3597, new_n3595, new_n3598);
xor_4  g03222(new_n3598, new_n3594, new_n3599);
xor_4  g03223(new_n3599, new_n3552, new_n3600);
not_8  g03224(n4805, new_n3601);
or_8   g03225(new_n3062, new_n3601, new_n3602_1);
and_8  g03226(n11478, n7610, new_n3603);
or_8   g03227(new_n3523, new_n3522, new_n3604);
and_8  g03228(new_n3526, new_n3604, new_n3605);
and_8  g03229(new_n3605, new_n3603, new_n3606);
nor_6  g03230(new_n3605, new_n3603, new_n3607);
or_8   g03231(new_n3607, new_n3606, new_n3608);
and_8  g03232(n7733, n137, new_n3609);
and_8  g03233(n5283, n4826, new_n3610);
and_8  g03234(n12925, n6294, new_n3611);
xnor_4 g03235(new_n3611, new_n3610, new_n3612);
xor_4  g03236(new_n3612, new_n3609, new_n3613);
nor_6  g03237(new_n3613, new_n3608, new_n3614);
and_8  g03238(new_n3613, new_n3608, new_n3615);
or_8   g03239(new_n3615, new_n3614, new_n3616_1);
nor_6  g03240(new_n3616_1, new_n3602_1, new_n3617);
and_8  g03241(new_n3616_1, new_n3602_1, new_n3618);
or_8   g03242(new_n3618, new_n3617, new_n3619);
and_8  g03243(new_n3519, new_n3516, new_n3620);
not_8  g03244(new_n3520, new_n3621);
and_8  g03245(new_n3528, new_n3621, new_n3622);
nor_6  g03246(new_n3622, new_n3620, new_n3623);
or_8   g03247(new_n3623, new_n3619, new_n3624);
xor_4  g03248(new_n3616_1, new_n3602_1, new_n3625);
or_8   g03249(new_n3622, new_n3620, new_n3626);
or_8   g03250(new_n3626, new_n3625, new_n3627_1);
and_8  g03251(new_n3627_1, new_n3624, new_n3628);
and_8  g03252(new_n3628, new_n3549, new_n3629);
not_8  g03253(new_n3549, new_n3630);
and_8  g03254(new_n3626, new_n3625, new_n3631);
and_8  g03255(new_n3623, new_n3619, new_n3632);
or_8   g03256(new_n3632, new_n3631, new_n3633);
and_8  g03257(new_n3633, new_n3630, new_n3634);
or_8   g03258(new_n3634, new_n3629, new_n3635);
nor_6  g03259(new_n3559, new_n3556, new_n3636);
or_8   g03260(new_n3636, new_n3555, new_n3637);
or_8   g03261(new_n3637, new_n3635, new_n3638);
or_8   g03262(new_n3633, new_n3630, new_n3639);
or_8   g03263(new_n3628, new_n3549, new_n3640);
and_8  g03264(new_n3640, new_n3639, new_n3641);
not_8  g03265(new_n3555, new_n3642);
or_8   g03266(new_n3559, new_n3556, new_n3643);
and_8  g03267(new_n3643, new_n3642, new_n3644);
or_8   g03268(new_n3644, new_n3641, new_n3645);
and_8  g03269(new_n3645, new_n3638, new_n3646);
xor_4  g03270(new_n3646, new_n3600, new_n3647);
or_8   g03271(new_n3647, new_n3574, new_n3648);
and_8  g03272(new_n3648, new_n3573, new_n3649);
nor_6  g03273(new_n3649, new_n3457, new_n3650);
and_8  g03274(new_n3649, new_n3457, new_n3651);
or_8   g03275(new_n3651, new_n3650, new_n3652);
and_8  g03276(new_n3599, new_n3552, new_n3653);
and_8  g03277(n7236, n6359, new_n3654_1);
and_8  g03278(n6358, n4086, new_n3655);
or_8   g03279(new_n3586, new_n3585, new_n3656);
or_8   g03280(new_n3587, new_n3584, new_n3657);
and_8  g03281(new_n3657, new_n3656, new_n3658);
xor_4  g03282(new_n3658, new_n3655, new_n3659);
and_8  g03283(n5198, n405, new_n3660);
and_8  g03284(n8433, n1471, new_n3661_1);
xor_4  g03285(new_n3661_1, new_n3660, new_n3662);
or_8   g03286(new_n3662, new_n3659, new_n3663);
and_8  g03287(new_n3658, new_n3655, new_n3664);
nor_6  g03288(new_n3658, new_n3655, new_n3665);
or_8   g03289(new_n3665, new_n3664, new_n3666);
not_8  g03290(new_n3662, new_n3667);
or_8   g03291(new_n3667, new_n3666, new_n3668);
and_8  g03292(new_n3668, new_n3663, new_n3669);
and_8  g03293(n8384, n217, new_n3670);
and_8  g03294(n6611, n3992, new_n3671);
xor_4  g03295(new_n3671, new_n3670, new_n3672);
xor_4  g03296(new_n3672, new_n3669, new_n3673);
or_8   g03297(new_n3589, new_n3581, new_n3674);
and_8  g03298(new_n3674, new_n3673, new_n3675);
and_8  g03299(new_n3672, new_n3669, new_n3676);
nor_6  g03300(new_n3672, new_n3669, new_n3677_1);
or_8   g03301(new_n3677_1, new_n3676, new_n3678);
not_8  g03302(new_n3674, new_n3679);
and_8  g03303(new_n3679, new_n3678, new_n3680);
or_8   g03304(new_n3680, new_n3675, new_n3681);
not_8  g03305(new_n3592, new_n3682);
or_8   g03306(new_n3598, new_n3594, new_n3683);
and_8  g03307(new_n3683, new_n3682, new_n3684);
or_8   g03308(new_n3684, new_n3681, new_n3685);
or_8   g03309(new_n3679, new_n3678, new_n3686);
or_8   g03310(new_n3674, new_n3673, new_n3687);
and_8  g03311(new_n3687, new_n3686, new_n3688);
xor_4  g03312(new_n3591, new_n3577, new_n3689);
or_8   g03313(new_n3597, new_n3595, new_n3690);
and_8  g03314(new_n3690, new_n3689, new_n3691);
or_8   g03315(new_n3691, new_n3592, new_n3692);
or_8   g03316(new_n3692, new_n3688, new_n3693);
and_8  g03317(new_n3693, new_n3685, new_n3694);
and_8  g03318(new_n3694, new_n3654_1, new_n3695);
not_8  g03319(new_n3654_1, new_n3696);
and_8  g03320(new_n3692, new_n3688, new_n3697);
and_8  g03321(new_n3684, new_n3681, new_n3698);
or_8   g03322(new_n3698, new_n3697, new_n3699);
and_8  g03323(new_n3699, new_n3696, new_n3700);
or_8   g03324(new_n3700, new_n3695, new_n3701);
and_8  g03325(new_n3701, new_n3653, new_n3702);
nor_6  g03326(new_n3701, new_n3653, new_n3703);
or_8   g03327(new_n3703, new_n3702, new_n3704);
and_8  g03328(n4805, n503, new_n3705);
and_8  g03329(n4826, n137, new_n3706);
and_8  g03330(n7733, n6294, new_n3707);
and_8  g03331(n12925, n6797, new_n3708);
xor_4  g03332(new_n3708, new_n3707, new_n3709);
xor_4  g03333(new_n3709, new_n3706, new_n3710);
or_8   g03334(new_n3611, new_n3610, new_n3711);
or_8   g03335(new_n3612, new_n3609, new_n3712);
and_8  g03336(new_n3712, new_n3711, new_n3713);
xor_4  g03337(new_n3713, new_n3710, new_n3714);
and_8  g03338(n11478, n4970, new_n3715);
and_8  g03339(n7610, n5283, new_n3716);
xor_4  g03340(new_n3716, new_n3715, new_n3717);
xor_4  g03341(new_n3717, new_n3714, new_n3718);
or_8   g03342(new_n3614, new_n3606, new_n3719_1);
and_8  g03343(new_n3719_1, new_n3718, new_n3720);
nor_6  g03344(new_n3719_1, new_n3718, new_n3721);
or_8   g03345(new_n3721, new_n3720, new_n3722);
not_8  g03346(new_n3617, new_n3723);
and_8  g03347(new_n3624, new_n3723, new_n3724);
or_8   g03348(new_n3724, new_n3722, new_n3725);
xor_4  g03349(new_n3719_1, new_n3718, new_n3726);
or_8   g03350(new_n3631, new_n3617, new_n3727);
or_8   g03351(new_n3727, new_n3726, new_n3728);
and_8  g03352(new_n3728, new_n3725, new_n3729);
and_8  g03353(new_n3729, new_n3705, new_n3730);
not_8  g03354(new_n3705, new_n3731);
and_8  g03355(new_n3727, new_n3726, new_n3732);
and_8  g03356(new_n3724, new_n3722, new_n3733);
or_8   g03357(new_n3733, new_n3732, new_n3734);
and_8  g03358(new_n3734, new_n3731, new_n3735);
or_8   g03359(new_n3735, new_n3730, new_n3736);
xor_4  g03360(new_n3736, new_n3639, new_n3737);
and_8  g03361(new_n3737, new_n3704, new_n3738);
xor_4  g03362(new_n3701, new_n3653, new_n3739);
xor_4  g03363(new_n3736, new_n3629, new_n3740);
and_8  g03364(new_n3740, new_n3739, new_n3741);
or_8   g03365(new_n3741, new_n3738, new_n3742);
xor_4  g03366(new_n3644, new_n3635, new_n3743);
or_8   g03367(new_n3743, new_n3600, new_n3744);
and_8  g03368(new_n3744, new_n3645, new_n3745);
xor_4  g03369(new_n3745, new_n3742, new_n3746);
or_8   g03370(new_n3746, new_n3652, new_n3747);
xor_4  g03371(new_n3649, new_n3457, new_n3748);
and_8  g03372(new_n3745, new_n3742, new_n3749);
nor_6  g03373(new_n3745, new_n3742, new_n3750);
or_8   g03374(new_n3750, new_n3749, new_n3751);
or_8   g03375(new_n3751, new_n3748, new_n3752);
and_8  g03376(new_n3752, new_n3747, new_n3753);
or_8   g03377(new_n3753, new_n3376, new_n3754_1);
and_8  g03378(new_n3753, new_n3376, new_n3755);
xor_4  g03379(new_n3364, new_n3363, new_n3756);
not_8  g03380(new_n3756, new_n3757);
xor_4  g03381(new_n3743, new_n3600, new_n3758);
not_8  g03382(new_n3458, new_n3759);
xor_4  g03383(new_n3559, new_n3556, new_n3760);
or_8   g03384(new_n3567, new_n3561, new_n3761);
and_8  g03385(new_n3761, new_n3515, new_n3762);
and_8  g03386(new_n3762, new_n3760, new_n3763);
or_8   g03387(new_n3763, new_n3568, new_n3764);
or_8   g03388(new_n3764, new_n3759, new_n3765);
and_8  g03389(new_n3765, new_n3573, new_n3766);
xor_4  g03390(new_n3766, new_n3758, new_n3767);
or_8   g03391(new_n3767, new_n3757, new_n3768);
not_8  g03392(new_n3768, new_n3769);
xor_4  g03393(new_n3361, new_n3355, new_n3770);
xor_4  g03394(new_n3762, new_n3760, new_n3771);
nor_6  g03395(new_n3771, new_n3770, new_n3772);
xor_4  g03396(new_n3512, new_n3564, new_n3773);
and_8  g03397(n9956, n7862, new_n3774);
not_8  g03398(new_n3774, new_n3775);
and_8  g03399(new_n3775, new_n3306, new_n3776);
or_8   g03400(new_n3776, new_n3356, new_n3777);
nand_5 g03401(new_n3776, new_n3305, new_n3778);
nand_5 g03402(new_n3778, new_n3777, new_n3779);
nand_5 g03403(new_n3779, new_n3773, new_n3780);
not_8  g03404(new_n3779, new_n3781);
xor_4  g03405(new_n3781, new_n3773, new_n3782);
xor_4  g03406(new_n3508, new_n3382, new_n3783);
and_8  g03407(new_n3783, new_n3774, new_n3784);
xor_4  g03408(new_n3359, new_n3358, new_n3785);
or_8   g03409(new_n3785, new_n3784, new_n3786);
xor_4  g03410(new_n3510, new_n3509, new_n3787);
xnor_4 g03411(new_n3785, new_n3784, new_n3788);
or_8   g03412(new_n3788, new_n3787, new_n3789);
and_8  g03413(new_n3789, new_n3786, new_n3790);
or_8   g03414(new_n3790, new_n3782, new_n3791);
and_8  g03415(new_n3791, new_n3780, new_n3792);
xor_4  g03416(new_n3771, new_n3770, new_n3793);
and_8  g03417(new_n3793, new_n3792, new_n3794);
or_8   g03418(new_n3794, new_n3772, new_n3795);
xor_4  g03419(new_n3766, new_n3647, new_n3796);
or_8   g03420(new_n3796, new_n3756, new_n3797);
and_8  g03421(new_n3797, new_n3768, new_n3798);
and_8  g03422(new_n3798, new_n3795, new_n3799);
or_8   g03423(new_n3799, new_n3769, new_n3800);
or_8   g03424(new_n3800, new_n3755, new_n3801);
and_8  g03425(new_n3801, new_n3754_1, new_n3802);
nor_6  g03426(new_n3802, new_n3373, new_n3803);
and_8  g03427(new_n3802, new_n3373, new_n3804);
or_8   g03428(new_n3804, new_n3803, new_n3805);
and_8  g03429(n9400, n8065, new_n3806);
and_8  g03430(n10439, n2464, new_n3807);
and_8  g03431(n10391, n6877, new_n3808);
xnor_4 g03432(new_n3808, new_n3807, new_n3809);
xor_4  g03433(new_n3809, new_n3806, new_n3810);
and_8  g03434(new_n3430, new_n3427, new_n3811);
and_8  g03435(new_n3434, new_n3431, new_n3812);
nor_6  g03436(new_n3812, new_n3811, new_n3813);
xor_4  g03437(new_n3813, new_n3810, new_n3814);
and_8  g03438(new_n3429, new_n3428, new_n3815);
and_8  g03439(n11311, n8595, new_n3816);
xnor_4 g03440(new_n3816, new_n3815, new_n3817);
and_8  g03441(n4203, n3602, new_n3818);
and_8  g03442(n6126, n4187, new_n3819);
and_8  g03443(n12753, n3719, new_n3820);
xnor_4 g03444(new_n3820, new_n3819, new_n3821);
xor_4  g03445(new_n3821, new_n3818, new_n3822);
xor_4  g03446(new_n3822, new_n3817, new_n3823);
not_8  g03447(new_n3823, new_n3824);
xor_4  g03448(new_n3824, new_n3814, new_n3825);
and_8  g03449(new_n3438, new_n3435, new_n3826);
and_8  g03450(new_n3437, new_n3436, new_n3827);
xor_4  g03451(new_n3444, new_n3827, new_n3828);
or_8   g03452(new_n3828, new_n3826, new_n3829);
xor_4  g03453(new_n3829, new_n3825, new_n3830);
and_8  g03454(new_n3830, new_n3449, new_n3831);
not_8  g03455(new_n3449, new_n3832);
not_8  g03456(new_n3825, new_n3833);
xor_4  g03457(new_n3829, new_n3833, new_n3834);
and_8  g03458(new_n3834, new_n3832, new_n3835);
or_8   g03459(new_n3835, new_n3831, new_n3836);
nor_6  g03460(new_n3453, new_n3426, new_n3837);
or_8   g03461(new_n3456_1, new_n3837, new_n3838);
xor_4  g03462(new_n3838, new_n3836, new_n3839);
not_8  g03463(new_n3839, new_n3840);
and_8  g03464(n10965, n4805, new_n3841);
and_8  g03465(n5283, n4970, new_n3842_1);
and_8  g03466(n11478, n503, new_n3843);
xnor_4 g03467(new_n3843, new_n3842_1, new_n3844);
xor_4  g03468(new_n3844, new_n3841, new_n3845);
and_8  g03469(new_n3709, new_n3706, new_n3846);
and_8  g03470(new_n3713, new_n3710, new_n3847);
or_8   g03471(new_n3847, new_n3846, new_n3848);
xor_4  g03472(new_n3848, new_n3845, new_n3849_1);
and_8  g03473(new_n3708, new_n3707, new_n3850);
and_8  g03474(n7610, n137, new_n3851);
xnor_4 g03475(new_n3851, new_n3850, new_n3852);
and_8  g03476(n7733, n6797, new_n3853);
and_8  g03477(n6294, n4826, new_n3854);
and_8  g03478(n12925, n3146, new_n3855);
xnor_4 g03479(new_n3855, new_n3854, new_n3856);
xor_4  g03480(new_n3856, new_n3853, new_n3857);
xor_4  g03481(new_n3857, new_n3852, new_n3858);
xor_4  g03482(new_n3858, new_n3849_1, new_n3859);
and_8  g03483(new_n3717, new_n3714, new_n3860);
and_8  g03484(new_n3716, new_n3715, new_n3861);
xor_4  g03485(new_n3720, new_n3861, new_n3862);
nor_6  g03486(new_n3862, new_n3860, new_n3863);
or_8   g03487(new_n3863, new_n3859, new_n3864);
not_8  g03488(new_n3859, new_n3865_1);
or_8   g03489(new_n3862, new_n3860, new_n3866);
or_8   g03490(new_n3866, new_n3865_1, new_n3867);
and_8  g03491(new_n3867, new_n3864, new_n3868);
or_8   g03492(new_n3868, new_n3732, new_n3869);
and_8  g03493(new_n3866, new_n3865_1, new_n3870);
and_8  g03494(new_n3863, new_n3859, new_n3871);
or_8   g03495(new_n3871, new_n3870, new_n3872);
or_8   g03496(new_n3872, new_n3725, new_n3873);
and_8  g03497(new_n3873, new_n3869, new_n3874);
or_8   g03498(new_n3729, new_n3705, new_n3875);
or_8   g03499(new_n3736, new_n3629, new_n3876);
and_8  g03500(new_n3876, new_n3875, new_n3877);
nor_6  g03501(new_n3877, new_n3874, new_n3878);
and_8  g03502(new_n3877, new_n3874, new_n3879);
or_8   g03503(new_n3879, new_n3878, new_n3880);
and_8  g03504(n11296, n7236, new_n3881);
and_8  g03505(n8384, n6611, new_n3882);
and_8  g03506(n6359, n3992, new_n3883);
xnor_4 g03507(new_n3883, new_n3882, new_n3884);
xor_4  g03508(new_n3884, new_n3881, new_n3885);
and_8  g03509(new_n3662, new_n3659, new_n3886);
or_8   g03510(new_n3886, new_n3664, new_n3887);
xor_4  g03511(new_n3887, new_n3885, new_n3888);
and_8  g03512(new_n3661_1, new_n3660, new_n3889);
and_8  g03513(n6358, n217, new_n3890);
xnor_4 g03514(new_n3890, new_n3889, new_n3891);
and_8  g03515(n1471, n405, new_n3892);
and_8  g03516(n5198, n4086, new_n3893);
and_8  g03517(n8433, n7646, new_n3894);
xnor_4 g03518(new_n3894, new_n3893, new_n3895);
xor_4  g03519(new_n3895, new_n3892, new_n3896);
xor_4  g03520(new_n3896, new_n3891, new_n3897);
nor_6  g03521(new_n3897, new_n3888, new_n3898);
and_8  g03522(new_n3897, new_n3888, new_n3899);
or_8   g03523(new_n3899, new_n3898, new_n3900);
not_8  g03524(new_n3900, new_n3901);
not_8  g03525(new_n3676, new_n3902);
nand_5 g03526(new_n3671, new_n3670, new_n3903);
not_8  g03527(new_n3903, new_n3904);
and_8  g03528(new_n3675, new_n3904, new_n3905);
and_8  g03529(new_n3686, new_n3903, new_n3906);
or_8   g03530(new_n3906, new_n3905, new_n3907);
and_8  g03531(new_n3907, new_n3902, new_n3908);
or_8   g03532(new_n3908, new_n3901, new_n3909);
or_8   g03533(new_n3686, new_n3903, new_n3910);
or_8   g03534(new_n3675, new_n3904, new_n3911);
and_8  g03535(new_n3911, new_n3910, new_n3912);
or_8   g03536(new_n3912, new_n3676, new_n3913);
or_8   g03537(new_n3913, new_n3900, new_n3914);
and_8  g03538(new_n3914, new_n3909, new_n3915);
xor_4  g03539(new_n3915, new_n3685, new_n3916);
or_8   g03540(new_n3703, new_n3700, new_n3917);
and_8  g03541(new_n3917, new_n3916, new_n3918);
xor_4  g03542(new_n3915, new_n3697, new_n3919);
nor_6  g03543(new_n3703, new_n3700, new_n3920);
and_8  g03544(new_n3920, new_n3919, new_n3921);
or_8   g03545(new_n3921, new_n3918, new_n3922);
or_8   g03546(new_n3922, new_n3880, new_n3923);
xor_4  g03547(new_n3877, new_n3874, new_n3924);
or_8   g03548(new_n3920, new_n3919, new_n3925);
or_8   g03549(new_n3917, new_n3916, new_n3926);
and_8  g03550(new_n3926, new_n3925, new_n3927);
or_8   g03551(new_n3927, new_n3924, new_n3928);
and_8  g03552(new_n3928, new_n3923, new_n3929);
or_8   g03553(new_n3737, new_n3704, new_n3930);
or_8   g03554(new_n3745, new_n3742, new_n3931);
and_8  g03555(new_n3931, new_n3930, new_n3932_1);
and_8  g03556(new_n3932_1, new_n3929, new_n3933);
nor_6  g03557(new_n3932_1, new_n3929, new_n3934);
or_8   g03558(new_n3934, new_n3933, new_n3935);
or_8   g03559(new_n3935, new_n3840, new_n3936);
xor_4  g03560(new_n3932_1, new_n3929, new_n3937);
or_8   g03561(new_n3937, new_n3839, new_n3938);
and_8  g03562(new_n3938, new_n3936, new_n3939);
and_8  g03563(new_n3751, new_n3748, new_n3940);
nor_6  g03564(new_n3940, new_n3651, new_n3941);
and_8  g03565(new_n3941, new_n3939, new_n3942);
and_8  g03566(new_n3937, new_n3839, new_n3943);
and_8  g03567(new_n3935, new_n3840, new_n3944);
or_8   g03568(new_n3944, new_n3943, new_n3945);
or_8   g03569(new_n3940, new_n3651, new_n3946);
and_8  g03570(new_n3946, new_n3945, new_n3947);
nor_6  g03571(new_n3947, new_n3942, new_n3948);
xor_4  g03572(new_n3948, new_n3805, n844);
and_8  g03573(n7456, n6687, new_n3950);
and_8  g03574(n12591, n6687, new_n3951);
and_8  g03575(n4189, n1798, new_n3952);
or_8   g03576(new_n3952, new_n3951, new_n3953);
and_8  g03577(n6687, n1798, new_n3954);
and_8  g03578(n12591, n4189, new_n3955);
and_8  g03579(new_n3955, new_n3954, new_n3956);
and_8  g03580(n3932, n2564, new_n3957);
or_8   g03581(new_n3957, new_n3956, new_n3958);
and_8  g03582(new_n3958, new_n3953, new_n3959);
xor_4  g03583(new_n3959, new_n3950, new_n3960);
and_8  g03584(n4189, n3932, new_n3961);
and_8  g03585(n12591, n2564, new_n3962);
and_8  g03586(n6770, n1798, new_n3963);
xor_4  g03587(new_n3963, new_n3962, new_n3964);
xor_4  g03588(new_n3964, new_n3961, new_n3965);
xor_4  g03589(new_n3965, new_n3960, new_n3966);
not_8  g03590(new_n3954, new_n3967);
nand_5 g03591(new_n3957, new_n3967, new_n3968);
not_8  g03592(new_n3956, new_n3969);
nand_5 g03593(new_n3969, new_n3953, new_n3970);
and_8  g03594(new_n3970, new_n3968, new_n3971);
and_8  g03595(new_n3971, new_n3957, new_n3972);
xor_4  g03596(new_n3972, new_n3966, new_n3973);
not_8  g03597(new_n3973, new_n3974);
not_8  g03598(new_n3968, new_n3975);
and_8  g03599(new_n3975, new_n3953, new_n3976);
or_8   g03600(new_n3976, new_n3971, new_n3977);
and_8  g03601(n8336, n6703, new_n3978);
and_8  g03602(n11876, n11222, new_n3979);
and_8  g03603(n12069, n5645, new_n3980);
xor_4  g03604(new_n3980, new_n3979, new_n3981);
and_8  g03605(new_n3981, new_n3978, new_n3982);
and_8  g03606(n9640, n8336, new_n3983);
and_8  g03607(n10928, n6703, new_n3984);
xor_4  g03608(new_n3984, new_n3983, new_n3985);
nand_5 g03609(new_n3985, new_n3982, new_n3986_1);
and_8  g03610(new_n3980, new_n3979, new_n3987);
and_8  g03611(n12391, n5645, new_n3988);
and_8  g03612(n12069, n1067, new_n3989);
xor_4  g03613(new_n3989, new_n3988, new_n3990);
xor_4  g03614(new_n3990, new_n3987, new_n3991);
and_8  g03615(n11222, n10898, new_n3992_1);
and_8  g03616(n11876, n11153, new_n3993);
xnor_4 g03617(new_n3993, new_n3992_1, new_n3994);
xor_4  g03618(new_n3994, new_n3991, new_n3995);
xor_4  g03619(new_n3985, new_n3982, new_n3996);
not_8  g03620(new_n3996, new_n3997);
or_8   g03621(new_n3997, new_n3995, new_n3998);
and_8  g03622(new_n3998, new_n3986_1, new_n3999);
not_8  g03623(n9640, new_n4000);
not_8  g03624(n10928, new_n4001);
or_8   g03625(new_n4001, new_n4000, new_n4002);
or_8   g03626(new_n4002, new_n3978, new_n4003);
and_8  g03627(n6986, n6703, new_n4004);
and_8  g03628(n8336, n3022, new_n4005_1);
or_8   g03629(new_n4005_1, new_n4004, new_n4006);
not_8  g03630(new_n4006, new_n4007);
and_8  g03631(n6986, n3022, new_n4008);
and_8  g03632(new_n4008, new_n3978, new_n4009);
or_8   g03633(new_n4009, new_n4007, new_n4010);
nand_5 g03634(new_n4010, new_n4003, new_n4011);
or_8   g03635(new_n4007, new_n4003, new_n4012);
and_8  g03636(new_n4012, new_n4011, new_n4013);
xor_4  g03637(new_n4013, new_n3999, new_n4014);
nand_5 g03638(new_n3989, new_n3988, new_n4015);
and_8  g03639(n12069, n8665, new_n4016);
and_8  g03640(n12391, n1067, new_n4017);
and_8  g03641(n7891, n5645, new_n4018);
nor_6  g03642(new_n4018, new_n4017, new_n4019);
and_8  g03643(new_n4018, new_n4017, new_n4020);
or_8   g03644(new_n4020, new_n4019, new_n4021);
xor_4  g03645(new_n4021, new_n4016, new_n4022);
xnor_4 g03646(new_n4022, new_n4015, new_n4023);
nor_6  g03647(new_n3990, new_n3987, new_n4024);
and_8  g03648(new_n3994, new_n3991, new_n4025);
nor_6  g03649(new_n4025, new_n4024, new_n4026);
not_8  g03650(n10898, new_n4027);
not_8  g03651(n11153, new_n4028);
or_8   g03652(new_n4028, new_n4027, new_n4029);
nor_6  g03653(new_n4029, new_n3979, new_n4030);
and_8  g03654(n11876, n5314, new_n4031);
and_8  g03655(n11222, n3754, new_n4032);
or_8   g03656(new_n4032, new_n4031, new_n4033);
nor_6  g03657(new_n4033, new_n4030, new_n4034);
and_8  g03658(n5314, n3754, new_n4035);
and_8  g03659(new_n4035, new_n3979, new_n4036);
or_8   g03660(new_n4036, new_n4034, new_n4037);
and_8  g03661(new_n4033, new_n4030, new_n4038);
nor_6  g03662(new_n4038, new_n4037, new_n4039);
xor_4  g03663(new_n4039, new_n4026, new_n4040);
xnor_4 g03664(new_n4040, new_n4023, new_n4041);
xor_4  g03665(new_n4041, new_n4014, new_n4042);
or_8   g03666(new_n4042, new_n3977, new_n4043);
xor_4  g03667(new_n3981, new_n3978, new_n4044);
and_8  g03668(new_n4044, new_n3954, new_n4045);
and_8  g03669(n2564, n1798, new_n4046);
and_8  g03670(n6687, n3932, new_n4047);
xor_4  g03671(new_n4047, new_n4046, new_n4048);
or_8   g03672(new_n4048, new_n4045, new_n4049);
not_8  g03673(new_n4049, new_n4050);
xor_4  g03674(new_n3996, new_n3995, new_n4051);
xor_4  g03675(new_n4048, new_n4045, new_n4052);
and_8  g03676(new_n4052, new_n4051, new_n4053);
or_8   g03677(new_n4053, new_n4050, new_n4054);
not_8  g03678(new_n4043, new_n4055);
and_8  g03679(new_n4042, new_n3977, new_n4056);
or_8   g03680(new_n4056, new_n4055, new_n4057);
or_8   g03681(new_n4057, new_n4054, new_n4058);
and_8  g03682(new_n4058, new_n4043, new_n4059);
xor_4  g03683(new_n4059, new_n3974, new_n4060);
or_8   g03684(new_n4022, new_n4015, new_n4061);
and_8  g03685(n12069, n11922, new_n4062);
or_8   g03686(new_n4018, new_n4017, new_n4063);
or_8   g03687(new_n4021, new_n4016, new_n4064);
and_8  g03688(new_n4064, new_n4063, new_n4065);
and_8  g03689(new_n4065, new_n4062, new_n4066);
nor_6  g03690(new_n4065, new_n4062, new_n4067);
or_8   g03691(new_n4067, new_n4066, new_n4068);
and_8  g03692(n7160, n5645, new_n4069);
and_8  g03693(n7891, n1067, new_n4070);
and_8  g03694(n12391, n8665, new_n4071);
nor_6  g03695(new_n4071, new_n4070, new_n4072);
and_8  g03696(new_n4071, new_n4070, new_n4073);
or_8   g03697(new_n4073, new_n4072, new_n4074);
xor_4  g03698(new_n4074, new_n4069, new_n4075);
nor_6  g03699(new_n4075, new_n4068, new_n4076);
and_8  g03700(new_n4075, new_n4068, new_n4077);
or_8   g03701(new_n4077, new_n4076, new_n4078);
and_8  g03702(new_n4078, new_n4061, new_n4079);
nor_6  g03703(new_n4078, new_n4061, new_n4080);
or_8   g03704(new_n4080, new_n4079, new_n4081);
and_8  g03705(n11222, n2749, new_n4082);
and_8  g03706(n11153, n10898, new_n4083);
or_8   g03707(new_n4036, new_n4083, new_n4084);
and_8  g03708(new_n4084, new_n4033, new_n4085);
xor_4  g03709(new_n4085, new_n4082, new_n4086_1);
and_8  g03710(n10898, n5314, new_n4087);
and_8  g03711(n11153, n3754, new_n4088_1);
and_8  g03712(n11876, n996, new_n4089);
nor_6  g03713(new_n4089, new_n4088_1, new_n4090);
and_8  g03714(new_n4089, new_n4088_1, new_n4091);
or_8   g03715(new_n4091, new_n4090, new_n4092);
and_8  g03716(new_n4092, new_n4087, new_n4093);
nor_6  g03717(new_n4092, new_n4087, new_n4094_1);
or_8   g03718(new_n4094_1, new_n4093, new_n4095);
and_8  g03719(new_n4095, new_n4086_1, new_n4096);
nor_6  g03720(new_n4095, new_n4086_1, new_n4097);
or_8   g03721(new_n4097, new_n4096, new_n4098);
nor_6  g03722(new_n4036, new_n4034, new_n4099);
or_8   g03723(new_n4099, new_n4029, new_n4100);
nor_6  g03724(new_n4100, new_n4098, new_n4101);
and_8  g03725(new_n4100, new_n4098, new_n4102);
or_8   g03726(new_n4102, new_n4101, new_n4103);
xor_4  g03727(new_n4103, new_n4081, new_n4104);
nor_6  g03728(new_n4039, new_n4026, new_n4105);
and_8  g03729(new_n4040, new_n4023, new_n4106);
or_8   g03730(new_n4106, new_n4105, new_n4107);
xor_4  g03731(new_n4107, new_n4104, new_n4108);
not_8  g03732(new_n4108, new_n4109);
and_8  g03733(n11023, n8336, new_n4110);
and_8  g03734(n10928, n9640, new_n4111);
or_8   g03735(new_n4009, new_n4111, new_n4112);
and_8  g03736(new_n4112, new_n4006, new_n4113);
xor_4  g03737(new_n4113, new_n4110, new_n4114);
and_8  g03738(n9640, n6986, new_n4115);
and_8  g03739(n10928, n3022, new_n4116);
and_8  g03740(n6703, n2226, new_n4117);
xor_4  g03741(new_n4117, new_n4116, new_n4118);
xor_4  g03742(new_n4118, new_n4115, new_n4119);
xor_4  g03743(new_n4119, new_n4114, new_n4120);
nor_6  g03744(new_n4011, new_n4002, new_n4121);
xor_4  g03745(new_n4121, new_n4120, new_n4122);
not_8  g03746(new_n3999, new_n4123);
or_8   g03747(new_n4013, new_n4123, new_n4124);
or_8   g03748(new_n4041, new_n4014, new_n4125);
and_8  g03749(new_n4125, new_n4124, new_n4126);
xor_4  g03750(new_n4126, new_n4122, new_n4127);
xor_4  g03751(new_n4127, new_n4109, new_n4128);
xor_4  g03752(new_n4128, new_n4060, n911);
and_8  g03753(n6687, n3842, new_n4130);
and_8  g03754(n11917, n6687, new_n4131);
and_8  g03755(n9956, n4189, new_n4132);
or_8   g03756(new_n4132, new_n4131, new_n4133);
and_8  g03757(n9956, n6687, new_n4134);
and_8  g03758(n11917, n4189, new_n4135);
and_8  g03759(new_n4135, new_n4134, new_n4136);
and_8  g03760(n4921, n2564, new_n4137);
or_8   g03761(new_n4137, new_n4136, new_n4138);
and_8  g03762(new_n4138, new_n4133, new_n4139);
xor_4  g03763(new_n4139, new_n4130, new_n4140);
and_8  g03764(n4921, n4189, new_n4141_1);
and_8  g03765(n11917, n2564, new_n4142);
and_8  g03766(n9956, n6770, new_n4143);
xor_4  g03767(new_n4143, new_n4142, new_n4144);
xor_4  g03768(new_n4144, new_n4141_1, new_n4145);
xor_4  g03769(new_n4145, new_n4140, new_n4146);
not_8  g03770(new_n4136, new_n4147);
nand_5 g03771(new_n4147, new_n4133, new_n4148);
and_8  g03772(n9956, n2564, new_n4149);
and_8  g03773(n6687, n4921, new_n4150);
and_8  g03774(new_n4150, new_n4149, new_n4151);
and_8  g03775(new_n4151, new_n4148, new_n4152);
and_8  g03776(new_n4152, new_n4146, new_n4153);
and_8  g03777(n6687, n2577, new_n4154);
and_8  g03778(new_n4139, new_n4130, new_n4155_1);
and_8  g03779(new_n4145, new_n4140, new_n4156);
or_8   g03780(new_n4156, new_n4155_1, new_n4157);
xnor_4 g03781(new_n4157, new_n4154, new_n4158);
and_8  g03782(n3842, n2564, new_n4159_1);
or_8   g03783(new_n4143, new_n4142, new_n4160);
and_8  g03784(new_n4143, new_n4142, new_n4161);
or_8   g03785(new_n4161, new_n4141_1, new_n4162);
and_8  g03786(new_n4162, new_n4160, new_n4163);
xor_4  g03787(new_n4163, new_n4159_1, new_n4164);
and_8  g03788(n6770, n4921, new_n4165);
and_8  g03789(n9956, n9920, new_n4166);
xnor_4 g03790(new_n4166, new_n4135, new_n4167);
xnor_4 g03791(new_n4167, new_n4165, new_n4168);
and_8  g03792(new_n4168, new_n4164, new_n4169);
nor_6  g03793(new_n4168, new_n4164, new_n4170);
or_8   g03794(new_n4170, new_n4169, new_n4171);
xor_4  g03795(new_n4171, new_n4158, new_n4172);
xnor_4 g03796(new_n4172, new_n4153, new_n4173);
xor_4  g03797(new_n4152, new_n4146, new_n4174);
and_8  g03798(n8595, n8336, new_n4175);
and_8  g03799(n8336, n6126, new_n4176);
and_8  g03800(n6986, n3719, new_n4177);
or_8   g03801(new_n4177, new_n4176, new_n4178);
and_8  g03802(n8336, n3719, new_n4179);
and_8  g03803(n6986, n6126, new_n4180);
and_8  g03804(new_n4180, new_n4179, new_n4181);
and_8  g03805(n10928, n3602, new_n4182);
or_8   g03806(new_n4182, new_n4181, new_n4183);
and_8  g03807(new_n4183, new_n4178, new_n4184);
xor_4  g03808(new_n4184, new_n4175, new_n4185);
and_8  g03809(n6986, n3602, new_n4186);
and_8  g03810(n10928, n6126, new_n4187_1);
and_8  g03811(n3719, n2226, new_n4188);
xor_4  g03812(new_n4188, new_n4187_1, new_n4189_1);
xor_4  g03813(new_n4189_1, new_n4186, new_n4190_1);
xnor_4 g03814(new_n4190_1, new_n4185, new_n4191);
not_8  g03815(new_n4182, new_n4192);
or_8   g03816(new_n4192, new_n4179, new_n4193);
not_8  g03817(new_n4178, new_n4194);
or_8   g03818(new_n4181, new_n4194, new_n4195);
and_8  g03819(new_n4195, new_n4193, new_n4196);
not_8  g03820(new_n4196, new_n4197);
or_8   g03821(new_n4197, new_n4192, new_n4198);
xor_4  g03822(new_n4198, new_n4191, new_n4199);
and_8  g03823(n12069, n7610, new_n4200);
and_8  g03824(n12069, n4826, new_n4201);
and_8  g03825(n12925, n7891, new_n4202);
or_8   g03826(new_n4202, new_n4201, new_n4203_1);
and_8  g03827(n12925, n12069, new_n4204);
and_8  g03828(n7891, n4826, new_n4205);
and_8  g03829(new_n4205, new_n4204, new_n4206);
and_8  g03830(n12391, n7733, new_n4207);
or_8   g03831(new_n4207, new_n4206, new_n4208);
and_8  g03832(new_n4208, new_n4203_1, new_n4209);
xor_4  g03833(new_n4209, new_n4200, new_n4210);
and_8  g03834(n7891, n7733, new_n4211);
and_8  g03835(n12925, n7160, new_n4212);
and_8  g03836(n12391, n4826, new_n4213);
nor_6  g03837(new_n4213, new_n4212, new_n4214);
and_8  g03838(new_n4213, new_n4212, new_n4215);
or_8   g03839(new_n4215, new_n4214, new_n4216);
and_8  g03840(new_n4216, new_n4211, new_n4217);
nor_6  g03841(new_n4216, new_n4211, new_n4218);
or_8   g03842(new_n4218, new_n4217, new_n4219);
xor_4  g03843(new_n4219, new_n4210, new_n4220);
nor_6  g03844(new_n4202, new_n4201, new_n4221);
or_8   g03845(new_n4206, new_n4221, new_n4222);
and_8  g03846(n12925, n12391, new_n4223);
and_8  g03847(n12069, n7733, new_n4224);
and_8  g03848(new_n4224, new_n4223, new_n4225);
nand_5 g03849(new_n4225, new_n4222, new_n4226_1);
xor_4  g03850(new_n4226_1, new_n4220, new_n4227);
and_8  g03851(n11222, n217, new_n4228);
and_8  g03852(n8433, n5314, new_n4229);
and_8  g03853(n11222, n4086, new_n4230_1);
or_8   g03854(new_n4230_1, new_n4229, new_n4231);
and_8  g03855(new_n4230_1, new_n4229, new_n4232);
and_8  g03856(n11153, n405, new_n4233);
or_8   g03857(new_n4233, new_n4232, new_n4234);
and_8  g03858(new_n4234, new_n4231, new_n4235);
xor_4  g03859(new_n4235, new_n4228, new_n4236);
and_8  g03860(n5314, n405, new_n4237);
and_8  g03861(n8433, n996, new_n4238);
and_8  g03862(n11153, n4086, new_n4239);
xor_4  g03863(new_n4239, new_n4238, new_n4240);
xor_4  g03864(new_n4240, new_n4237, new_n4241);
xor_4  g03865(new_n4241, new_n4236, new_n4242);
not_8  g03866(n8433, new_n4243);
not_8  g03867(n11222, new_n4244);
or_8   g03868(new_n4244, new_n4243, new_n4245);
and_8  g03869(new_n4245, new_n4233, new_n4246);
nor_6  g03870(new_n4246, new_n4231, new_n4247);
or_8   g03871(new_n4247, new_n4232, new_n4248);
and_8  g03872(new_n4248, new_n4233, new_n4249);
and_8  g03873(new_n4249, new_n4242, new_n4250);
nor_6  g03874(new_n4249, new_n4242, new_n4251);
or_8   g03875(new_n4251, new_n4250, new_n4252);
nor_6  g03876(new_n4252, new_n4227, new_n4253);
and_8  g03877(new_n4252, new_n4227, new_n4254);
or_8   g03878(new_n4254, new_n4253, new_n4255);
and_8  g03879(n11222, n8433, new_n4256);
and_8  g03880(new_n4256, new_n4204, new_n4257);
and_8  g03881(n11153, n8433, new_n4258);
and_8  g03882(n11222, n405, new_n4259);
xor_4  g03883(new_n4259, new_n4258, new_n4260);
or_8   g03884(new_n4260, new_n4257, new_n4261);
xor_4  g03885(new_n4260, new_n4257, new_n4262);
not_8  g03886(new_n4262, new_n4263);
xor_4  g03887(new_n4224, new_n4223, new_n4264);
or_8   g03888(new_n4264, new_n4263, new_n4265);
and_8  g03889(new_n4265, new_n4261, new_n4266);
and_8  g03890(new_n4246, new_n4231, new_n4267);
nor_6  g03891(new_n4267, new_n4248, new_n4268);
nor_6  g03892(new_n4268, new_n4266, new_n4269);
xor_4  g03893(new_n4268, new_n4266, new_n4270);
not_8  g03894(new_n4204, new_n4271);
nand_5 g03895(new_n4207, new_n4271, new_n4272);
and_8  g03896(new_n4272, new_n4222, new_n4273);
nor_6  g03897(new_n4272, new_n4221, new_n4274);
or_8   g03898(new_n4274, new_n4273, new_n4275);
and_8  g03899(new_n4275, new_n4270, new_n4276);
nor_6  g03900(new_n4276, new_n4269, new_n4277);
and_8  g03901(new_n4277, new_n4255, new_n4278);
nor_6  g03902(new_n4277, new_n4255, new_n4279);
or_8   g03903(new_n4279, new_n4278, new_n4280);
and_8  g03904(new_n4280, new_n4199, new_n4281);
nor_6  g03905(new_n4280, new_n4199, new_n4282);
or_8   g03906(new_n4282, new_n4281, new_n4283);
or_8   g03907(new_n4193, new_n4194, new_n4284);
nand_5 g03908(new_n4284, new_n4197, new_n4285);
xor_4  g03909(new_n4275, new_n4270, new_n4286);
or_8   g03910(new_n4286, new_n4285, new_n4287);
not_8  g03911(new_n4287, new_n4288);
and_8  g03912(new_n4286, new_n4285, new_n4289);
or_8   g03913(new_n4289, new_n4288, new_n4290);
xor_4  g03914(new_n4264, new_n4262, new_n4291);
and_8  g03915(n10928, n3719, new_n4292);
and_8  g03916(n8336, n3602, new_n4293);
xor_4  g03917(new_n4293, new_n4292, new_n4294);
and_8  g03918(new_n4294, new_n4291, new_n4295);
xor_4  g03919(new_n4256, new_n4204, new_n4296);
and_8  g03920(new_n4296, new_n4179, new_n4297);
xor_4  g03921(new_n4294, new_n4291, new_n4298);
and_8  g03922(new_n4298, new_n4297, new_n4299);
or_8   g03923(new_n4299, new_n4295, new_n4300_1);
not_8  g03924(new_n4300_1, new_n4301);
or_8   g03925(new_n4301, new_n4290, new_n4302);
and_8  g03926(new_n4302, new_n4287, new_n4303);
or_8   g03927(new_n4303, new_n4283, new_n4304);
xor_4  g03928(new_n4280, new_n4199, new_n4305);
xor_4  g03929(new_n4286, new_n4285, new_n4306);
and_8  g03930(new_n4300_1, new_n4306, new_n4307);
or_8   g03931(new_n4307, new_n4288, new_n4308);
or_8   g03932(new_n4308, new_n4305, new_n4309);
and_8  g03933(new_n4309, new_n4304, new_n4310);
or_8   g03934(new_n4310, new_n4174, new_n4311);
and_8  g03935(new_n4301, new_n4290, new_n4312_1);
nor_6  g03936(new_n4312_1, new_n4307, new_n4313);
not_8  g03937(new_n4148, new_n4314);
not_8  g03938(new_n4134, new_n4315);
and_8  g03939(new_n4137, new_n4315, new_n4316);
or_8   g03940(new_n4316, new_n4314, new_n4317);
nand_5 g03941(new_n4316, new_n4133, new_n4318);
nand_5 g03942(new_n4318, new_n4317, new_n4319);
not_8  g03943(new_n4319, new_n4320);
or_8   g03944(new_n4320, new_n4313, new_n4321);
or_8   g03945(new_n4312_1, new_n4307, new_n4322);
and_8  g03946(new_n4319, new_n4322, new_n4323);
and_8  g03947(new_n4320, new_n4313, new_n4324);
or_8   g03948(new_n4324, new_n4323, new_n4325);
xor_4  g03949(new_n4296, new_n4179, new_n4326_1);
and_8  g03950(new_n4326_1, new_n4134, new_n4327);
xor_4  g03951(new_n4150, new_n4149, new_n4328);
or_8   g03952(new_n4328, new_n4327, new_n4329);
xor_4  g03953(new_n4298, new_n4297, new_n4330);
xnor_4 g03954(new_n4328, new_n4327, new_n4331);
or_8   g03955(new_n4331, new_n4330, new_n4332);
and_8  g03956(new_n4332, new_n4329, new_n4333_1);
or_8   g03957(new_n4333_1, new_n4325, new_n4334);
and_8  g03958(new_n4334, new_n4321, new_n4335);
not_8  g03959(new_n4174, new_n4336);
and_8  g03960(new_n4308, new_n4305, new_n4337);
and_8  g03961(new_n4303, new_n4283, new_n4338);
or_8   g03962(new_n4338, new_n4337, new_n4339);
and_8  g03963(new_n4339, new_n4336, new_n4340);
and_8  g03964(new_n4310, new_n4174, new_n4341);
or_8   g03965(new_n4341, new_n4340, new_n4342);
or_8   g03966(new_n4342, new_n4335, new_n4343);
and_8  g03967(new_n4343, new_n4311, new_n4344);
xor_4  g03968(new_n4344, new_n4173, new_n4345);
nor_6  g03969(new_n4198, new_n4191, new_n4346);
and_8  g03970(n10439, n8336, new_n4347);
and_8  g03971(new_n4184, new_n4175, new_n4348);
and_8  g03972(new_n4190_1, new_n4185, new_n4349);
or_8   g03973(new_n4349, new_n4348, new_n4350);
xnor_4 g03974(new_n4350, new_n4347, new_n4351);
and_8  g03975(n10928, n8595, new_n4352);
or_8   g03976(new_n4188, new_n4187_1, new_n4353);
and_8  g03977(new_n4188, new_n4187_1, new_n4354);
or_8   g03978(new_n4354, new_n4186, new_n4355);
and_8  g03979(new_n4355, new_n4353, new_n4356);
xor_4  g03980(new_n4356, new_n4352, new_n4357);
and_8  g03981(n3602, n2226, new_n4358);
and_8  g03982(n3719, n1094, new_n4359);
xnor_4 g03983(new_n4359, new_n4180, new_n4360);
xnor_4 g03984(new_n4360, new_n4358, new_n4361);
and_8  g03985(new_n4361, new_n4357, new_n4362);
nor_6  g03986(new_n4361, new_n4357, new_n4363);
or_8   g03987(new_n4363, new_n4362, new_n4364);
xor_4  g03988(new_n4364, new_n4351, new_n4365);
xor_4  g03989(new_n4365, new_n4346, new_n4366);
and_8  g03990(n11222, n6611, new_n4367);
nand_5 g03991(n11153, n217, new_n4368);
not_8  g03992(new_n4368, new_n4369);
and_8  g03993(n996, n405, new_n4370_1);
and_8  g03994(n5314, n4086, new_n4371);
and_8  g03995(n8433, n5767, new_n4372);
xor_4  g03996(new_n4372, new_n4371, new_n4373);
xor_4  g03997(new_n4373, new_n4370_1, new_n4374);
and_8  g03998(new_n4374, new_n4369, new_n4375);
not_8  g03999(n996, new_n4376);
or_8   g04000(new_n4376, new_n2747, new_n4377);
xor_4  g04001(new_n4373, new_n4377, new_n4378_1);
and_8  g04002(new_n4378_1, new_n4368, new_n4379);
or_8   g04003(new_n4379, new_n4375, new_n4380);
or_8   g04004(new_n4239, new_n4238, new_n4381);
and_8  g04005(new_n4239, new_n4238, new_n4382);
or_8   g04006(new_n4382, new_n4237, new_n4383);
nand_5 g04007(new_n4383, new_n4381, new_n4384);
or_8   g04008(new_n4384, new_n4380, new_n4385);
nor_6  g04009(new_n4379, new_n4375, new_n4386);
not_8  g04010(new_n4384, new_n4387);
or_8   g04011(new_n4387, new_n4386, new_n4388);
and_8  g04012(new_n4388, new_n4385, new_n4389);
xor_4  g04013(new_n4389, new_n4367, new_n4390);
and_8  g04014(new_n4235, new_n4228, new_n4391);
and_8  g04015(new_n4241, new_n4236, new_n4392);
or_8   g04016(new_n4392, new_n4391, new_n4393);
xor_4  g04017(new_n4393, new_n4390, new_n4394);
xor_4  g04018(new_n4394, new_n4250, new_n4395);
not_8  g04019(new_n4226_1, new_n4396);
nand_5 g04020(new_n4396, new_n4220, new_n4397_1);
not_8  g04021(n12069, new_n4398);
or_8   g04022(new_n4398, new_n3062, new_n4399);
and_8  g04023(n12391, n7610, new_n4400);
or_8   g04024(new_n4213, new_n4212, new_n4401);
or_8   g04025(new_n4216, new_n4211, new_n4402);
and_8  g04026(new_n4402, new_n4401, new_n4403);
xor_4  g04027(new_n4403, new_n4400, new_n4404);
and_8  g04028(n7733, n7160, new_n4405);
and_8  g04029(n12925, n4828, new_n4406);
xnor_4 g04030(new_n4406, new_n4205, new_n4407);
and_8  g04031(new_n4407, new_n4405, new_n4408);
nor_6  g04032(new_n4407, new_n4405, new_n4409);
or_8   g04033(new_n4409, new_n4408, new_n4410);
and_8  g04034(new_n4410, new_n4404, new_n4411);
and_8  g04035(new_n4403, new_n4400, new_n4412);
nor_6  g04036(new_n4403, new_n4400, new_n4413);
or_8   g04037(new_n4413, new_n4412, new_n4414);
xor_4  g04038(new_n4407, new_n4405, new_n4415);
and_8  g04039(new_n4415, new_n4414, new_n4416);
or_8   g04040(new_n4416, new_n4411, new_n4417);
nor_6  g04041(new_n4417, new_n4399, new_n4418);
and_8  g04042(new_n4417, new_n4399, new_n4419);
or_8   g04043(new_n4419, new_n4418, new_n4420);
and_8  g04044(new_n4209, new_n4200, new_n4421);
and_8  g04045(new_n4219, new_n4210, new_n4422);
or_8   g04046(new_n4422, new_n4421, new_n4423);
xor_4  g04047(new_n4423, new_n4420, new_n4424);
nor_6  g04048(new_n4424, new_n4397_1, new_n4425);
and_8  g04049(new_n4424, new_n4397_1, new_n4426);
or_8   g04050(new_n4426, new_n4425, new_n4427);
or_8   g04051(new_n4279, new_n4254, new_n4428);
nor_6  g04052(new_n4428, new_n4427, new_n4429);
and_8  g04053(new_n4428, new_n4427, new_n4430);
or_8   g04054(new_n4430, new_n4429, new_n4431);
xor_4  g04055(new_n4431, new_n4395, new_n4432);
xor_4  g04056(new_n4432, new_n4366, new_n4433);
or_8   g04057(new_n4337, new_n4281, new_n4434);
not_8  g04058(new_n4434, new_n4435);
and_8  g04059(new_n4435, new_n4433, new_n4436_1);
not_8  g04060(new_n4366, new_n4437);
xor_4  g04061(new_n4432, new_n4437, new_n4438);
and_8  g04062(new_n4434, new_n4438, new_n4439);
or_8   g04063(new_n4439, new_n4436_1, new_n4440);
xor_4  g04064(new_n4440, new_n4345, n992);
and_8  g04065(n7265, n6687, new_n4442);
and_8  g04066(n8336, n7946, new_n4443);
and_8  g04067(n11222, n9763, new_n4444);
and_8  g04068(n12069, n2558, new_n4445);
xor_4  g04069(new_n4445, new_n4444, new_n4446);
xor_4  g04070(new_n4446, new_n4443, new_n4447);
xor_4  g04071(new_n4447, new_n4442, n1020);
xor_4  g04072(new_n2109, new_n2104, n1136);
xnor_4 g04073(new_n4342, new_n4335, n1138);
and_8  g04074(n12591, n11757, new_n4451);
and_8  g04075(n5240, n3932, new_n4452);
and_8  g04076(n11821, n1798, new_n4453);
xor_4  g04077(new_n4453, new_n4452, new_n4454);
xor_4  g04078(new_n4454, new_n4451, new_n4455);
and_8  g04079(n5240, n1798, new_n4456);
and_8  g04080(n12591, n3172, new_n4457);
or_8   g04081(new_n4457, new_n4456, new_n4458);
and_8  g04082(new_n4457, new_n4456, new_n4459);
and_8  g04083(n11757, n3932, new_n4460);
or_8   g04084(new_n4460, new_n4459, new_n4461);
and_8  g04085(new_n4461, new_n4458, new_n4462);
xor_4  g04086(new_n4462, new_n4455, new_n4463);
and_8  g04087(n7456, n1333, new_n4464);
and_8  g04088(n11757, n1798, new_n4465);
and_8  g04089(n12591, n1333, new_n4466);
or_8   g04090(new_n4466, new_n4465, new_n4467);
and_8  g04091(new_n4466, new_n4465, new_n4468);
and_8  g04092(n3932, n3172, new_n4469);
or_8   g04093(new_n4469, new_n4468, new_n4470);
and_8  g04094(new_n4470, new_n4467, new_n4471);
and_8  g04095(new_n4471, new_n4464, new_n4472);
xnor_4 g04096(new_n4471, new_n4464, new_n4473);
xnor_4 g04097(new_n4457, new_n4456, new_n4474);
xor_4  g04098(new_n4474, new_n4460, new_n4475);
nor_6  g04099(new_n4475, new_n4473, new_n4476);
or_8   g04100(new_n4476, new_n4472, new_n4477);
and_8  g04101(n11662, n1333, new_n4478);
and_8  g04102(n7456, n3172, new_n4479);
xor_4  g04103(new_n4479, new_n4478, new_n4480);
xor_4  g04104(new_n4480, new_n4477, new_n4481);
and_8  g04105(new_n4481, new_n4463, new_n4482);
not_8  g04106(new_n4463, new_n4483);
not_8  g04107(new_n4480, new_n4484);
xor_4  g04108(new_n4484, new_n4477, new_n4485);
and_8  g04109(new_n4485, new_n4483, new_n4486);
or_8   g04110(new_n4486, new_n4482, new_n4487);
and_8  g04111(n11662, n7862, new_n4488);
not_8  g04112(new_n4488, new_n4489);
and_8  g04113(new_n4475, new_n4473, new_n4490);
or_8   g04114(new_n4490, new_n4476, new_n4491);
and_8  g04115(new_n4491, new_n4489, new_n4492);
xor_4  g04116(new_n4491, new_n4489, new_n4493);
and_8  g04117(n7862, n7456, new_n4494);
and_8  g04118(n3172, n1798, new_n4495);
and_8  g04119(n12591, n7862, new_n4496);
and_8  g04120(new_n4496, new_n4495, new_n4497);
or_8   g04121(new_n4496, new_n4495, new_n4498);
and_8  g04122(n3932, n1333, new_n4499_1);
and_8  g04123(new_n4499_1, new_n4498, new_n4500);
or_8   g04124(new_n4500, new_n4497, new_n4501);
and_8  g04125(new_n4501, new_n4494, new_n4502);
xor_4  g04126(new_n4501, new_n4494, new_n4503);
xor_4  g04127(new_n4466, new_n4465, new_n4504);
xor_4  g04128(new_n4504, new_n4469, new_n4505);
and_8  g04129(new_n4505, new_n4503, new_n4506);
or_8   g04130(new_n4506, new_n4502, new_n4507);
not_8  g04131(new_n4507, new_n4508);
and_8  g04132(new_n4508, new_n4493, new_n4509);
or_8   g04133(new_n4509, new_n4492, new_n4510);
or_8   g04134(new_n4510, new_n4487, new_n4511);
not_8  g04135(new_n4511, new_n4512);
and_8  g04136(new_n4454, new_n4451, new_n4513);
and_8  g04137(new_n4462, new_n4455, new_n4514);
or_8   g04138(new_n4514, new_n4513, new_n4515);
and_8  g04139(n10327, n1333, new_n4516_1);
and_8  g04140(n11662, n3172, new_n4517);
and_8  g04141(n9583, n7862, new_n4518);
xnor_4 g04142(new_n4518, new_n4517, new_n4519);
xor_4  g04143(new_n4519, new_n4516_1, new_n4520);
xor_4  g04144(new_n4520, new_n4515, new_n4521);
and_8  g04145(new_n4453, new_n4452, new_n4522);
and_8  g04146(n11757, n7456, new_n4523);
xnor_4 g04147(new_n4523, new_n4522, new_n4524);
and_8  g04148(n11821, n3932, new_n4525);
and_8  g04149(n12591, n5240, new_n4526);
and_8  g04150(n9080, n1798, new_n4527);
xnor_4 g04151(new_n4527, new_n4526, new_n4528);
xor_4  g04152(new_n4528, new_n4525, new_n4529);
xor_4  g04153(new_n4529, new_n4524, new_n4530);
xor_4  g04154(new_n4530, new_n4521, new_n4531);
nand_5 g04155(new_n4480, new_n4477, new_n4532);
and_8  g04156(new_n4479, new_n4478, new_n4533);
and_8  g04157(new_n4482, new_n4533, new_n4534);
not_8  g04158(new_n4533, new_n4535);
or_8   g04159(new_n4485, new_n4483, new_n4536);
and_8  g04160(new_n4536, new_n4535, new_n4537);
or_8   g04161(new_n4537, new_n4534, new_n4538);
and_8  g04162(new_n4538, new_n4532, new_n4539);
xor_4  g04163(new_n4539, new_n4531, new_n4540);
and_8  g04164(new_n4540, new_n4512, new_n4541);
not_8  g04165(new_n4531, new_n4542);
xor_4  g04166(new_n4539, new_n4542, new_n4543);
and_8  g04167(new_n4543, new_n4511, new_n4544);
or_8   g04168(new_n4544, new_n4541, new_n4545);
and_8  g04169(n10327, n7862, new_n4546);
or_8   g04170(new_n4481, new_n4463, new_n4547);
and_8  g04171(new_n4547, new_n4536, new_n4548);
not_8  g04172(new_n4492, new_n4549);
xor_4  g04173(new_n4491, new_n4488, new_n4550);
or_8   g04174(new_n4507, new_n4550, new_n4551);
and_8  g04175(new_n4551, new_n4549, new_n4552);
or_8   g04176(new_n4552, new_n4548, new_n4553_1);
and_8  g04177(new_n4553_1, new_n4511, new_n4554);
and_8  g04178(new_n4554, new_n4546, new_n4555);
not_8  g04179(new_n4555, new_n4556);
xnor_4 g04180(new_n4505, new_n4503, new_n4557);
xnor_4 g04181(new_n4496, new_n4495, new_n4558);
and_8  g04182(n1798, n1333, new_n4559);
and_8  g04183(n7862, n3932, new_n4560);
and_8  g04184(new_n4560, new_n4559, new_n4561);
and_8  g04185(new_n4561, new_n4558, new_n4562);
not_8  g04186(new_n4562, new_n4563);
or_8   g04187(new_n4563, new_n4557, new_n4564);
xor_4  g04188(new_n4507, new_n4550, new_n4565);
or_8   g04189(new_n4565, new_n4564, new_n4566);
nor_6  g04190(new_n4554, new_n4546, new_n4567);
or_8   g04191(new_n4567, new_n4555, new_n4568);
or_8   g04192(new_n4568, new_n4566, new_n4569);
and_8  g04193(new_n4569, new_n4556, new_n4570);
xor_4  g04194(new_n4570, new_n4545, new_n4571);
and_8  g04195(n11311, n3022, new_n4572);
and_8  g04196(n9640, n4187, new_n4573);
and_8  g04197(n6703, n4203, new_n4574);
xor_4  g04198(new_n4574, new_n4573, new_n4575);
xor_4  g04199(new_n4575, new_n4572, new_n4576);
and_8  g04200(n6703, n4187, new_n4577);
and_8  g04201(n3022, n2464, new_n4578);
or_8   g04202(new_n4578, new_n4577, new_n4579);
and_8  g04203(new_n4578, new_n4577, new_n4580);
and_8  g04204(n11311, n9640, new_n4581);
or_8   g04205(new_n4581, new_n4580, new_n4582);
and_8  g04206(new_n4582, new_n4579, new_n4583);
xor_4  g04207(new_n4583, new_n4576, new_n4584);
and_8  g04208(n10451, n9400, new_n4585);
and_8  g04209(n11023, n2464, new_n4586);
xor_4  g04210(new_n4586, new_n4585, new_n4587);
xor_4  g04211(new_n4587, new_n4584, new_n4588);
and_8  g04212(n11023, n9400, new_n4589);
and_8  g04213(n11311, n6703, new_n4590);
and_8  g04214(n9400, n3022, new_n4591);
or_8   g04215(new_n4591, new_n4590, new_n4592);
and_8  g04216(new_n4591, new_n4590, new_n4593);
and_8  g04217(n9640, n2464, new_n4594);
or_8   g04218(new_n4594, new_n4593, new_n4595);
and_8  g04219(new_n4595, new_n4592, new_n4596);
and_8  g04220(new_n4596, new_n4589, new_n4597);
xnor_4 g04221(new_n4596, new_n4589, new_n4598);
xnor_4 g04222(new_n4578, new_n4577, new_n4599);
xor_4  g04223(new_n4599, new_n4581, new_n4600);
nor_6  g04224(new_n4600, new_n4598, new_n4601);
or_8   g04225(new_n4601, new_n4597, new_n4602);
and_8  g04226(new_n4602, new_n4588, new_n4603);
nor_6  g04227(new_n4602, new_n4588, new_n4604);
or_8   g04228(new_n4604, new_n4603, new_n4605);
and_8  g04229(n10451, n6877, new_n4606);
not_8  g04230(new_n4606, new_n4607);
and_8  g04231(new_n4600, new_n4598, new_n4608);
or_8   g04232(new_n4608, new_n4601, new_n4609);
or_8   g04233(new_n4609, new_n4607, new_n4610);
and_8  g04234(n11023, n6877, new_n4611);
and_8  g04235(n6703, n2464, new_n4612);
and_8  g04236(n6877, n3022, new_n4613);
or_8   g04237(new_n4613, new_n4612, new_n4614);
and_8  g04238(new_n4613, new_n4612, new_n4615);
and_8  g04239(n9640, n9400, new_n4616);
or_8   g04240(new_n4616, new_n4615, new_n4617);
and_8  g04241(new_n4617, new_n4614, new_n4618);
and_8  g04242(new_n4618, new_n4611, new_n4619);
xor_4  g04243(new_n4618, new_n4611, new_n4620);
xor_4  g04244(new_n4591, new_n4590, new_n4621);
xor_4  g04245(new_n4621, new_n4594, new_n4622);
and_8  g04246(new_n4622, new_n4620, new_n4623);
or_8   g04247(new_n4623, new_n4619, new_n4624);
not_8  g04248(new_n4624, new_n4625);
xor_4  g04249(new_n4609, new_n4606, new_n4626);
or_8   g04250(new_n4626, new_n4625, new_n4627);
and_8  g04251(new_n4627, new_n4610, new_n4628);
or_8   g04252(new_n4628, new_n4605, new_n4629);
not_8  g04253(new_n4629, new_n4630);
and_8  g04254(new_n4575, new_n4572, new_n4631);
and_8  g04255(new_n4583, new_n4576, new_n4632);
or_8   g04256(new_n4632, new_n4631, new_n4633);
and_8  g04257(n10278, n9400, new_n4634_1);
and_8  g04258(n10451, n2464, new_n4635);
and_8  g04259(n11423, n6877, new_n4636);
xnor_4 g04260(new_n4636, new_n4635, new_n4637);
xor_4  g04261(new_n4637, new_n4634_1, new_n4638);
xor_4  g04262(new_n4638, new_n4633, new_n4639);
and_8  g04263(new_n4574, new_n4573, new_n4640);
and_8  g04264(n11311, n11023, new_n4641);
xnor_4 g04265(new_n4641, new_n4640, new_n4642);
and_8  g04266(n9640, n4203, new_n4643);
and_8  g04267(n4187, n3022, new_n4644);
and_8  g04268(n12753, n6703, new_n4645);
xnor_4 g04269(new_n4645, new_n4644, new_n4646);
xor_4  g04270(new_n4646, new_n4643, new_n4647);
xor_4  g04271(new_n4647, new_n4642, new_n4648);
xor_4  g04272(new_n4648, new_n4639, new_n4649);
not_8  g04273(new_n4649, new_n4650);
and_8  g04274(new_n4587, new_n4584, new_n4651);
and_8  g04275(new_n4586, new_n4585, new_n4652);
xor_4  g04276(new_n4603, new_n4652, new_n4653);
or_8   g04277(new_n4653, new_n4651, new_n4654);
xor_4  g04278(new_n4654, new_n4650, new_n4655);
and_8  g04279(new_n4655, new_n4630, new_n4656);
xor_4  g04280(new_n4654, new_n4649, new_n4657);
and_8  g04281(new_n4657, new_n4629, new_n4658);
or_8   g04282(new_n4658, new_n4656, new_n4659);
and_8  g04283(n10278, n6877, new_n4660);
xor_4  g04284(new_n4602, new_n4588, new_n4661);
not_8  g04285(new_n4610, new_n4662);
xor_4  g04286(new_n4609, new_n4607, new_n4663);
and_8  g04287(new_n4663, new_n4624, new_n4664);
or_8   g04288(new_n4664, new_n4662, new_n4665);
or_8   g04289(new_n4665, new_n4661, new_n4666);
and_8  g04290(new_n4666, new_n4629, new_n4667);
and_8  g04291(new_n4667, new_n4660, new_n4668);
not_8  g04292(new_n4668, new_n4669);
xor_4  g04293(new_n4622, new_n4620, new_n4670);
and_8  g04294(n6877, n6703, new_n4671);
not_8  g04295(new_n4671, new_n4672);
nand_5 g04296(new_n4672, new_n4616, new_n4673);
xnor_4 g04297(new_n4613, new_n4612, new_n4674);
and_8  g04298(new_n4674, new_n4673, new_n4675);
and_8  g04299(new_n4675, new_n4616, new_n4676);
nand_5 g04300(new_n4676, new_n4670, new_n4677);
not_8  g04301(new_n4677, new_n4678);
xor_4  g04302(new_n4663, new_n4624, new_n4679);
and_8  g04303(new_n4679, new_n4678, new_n4680);
not_8  g04304(new_n4680, new_n4681);
nor_6  g04305(new_n4667, new_n4660, new_n4682);
or_8   g04306(new_n4682, new_n4668, new_n4683);
or_8   g04307(new_n4683, new_n4681, new_n4684);
and_8  g04308(new_n4684, new_n4669, new_n4685);
xor_4  g04309(new_n4685, new_n4659, new_n4686_1);
and_8  g04310(n12826, n4805, new_n4687);
and_8  g04311(n8665, n137, new_n4688);
and_8  g04312(n6294, n1067, new_n4689_1);
and_8  g04313(n6797, n5645, new_n4690);
xor_4  g04314(new_n4690, new_n4689_1, new_n4691);
xor_4  g04315(new_n4691, new_n4688, new_n4692);
and_8  g04316(n6294, n5645, new_n4693);
and_8  g04317(n8665, n5283, new_n4694);
or_8   g04318(new_n4694, new_n4693, new_n4695);
and_8  g04319(n1067, n137, new_n4696);
xor_4  g04320(new_n4694, new_n4693, new_n4697);
not_8  g04321(new_n4697, new_n4698);
or_8   g04322(new_n4698, new_n4696, new_n4699);
and_8  g04323(new_n4699, new_n4695, new_n4700);
xor_4  g04324(new_n4700, new_n4692, new_n4701);
and_8  g04325(n11922, n11478, new_n4702);
and_8  g04326(n5283, n1067, new_n4703);
and_8  g04327(n11478, n8665, new_n4704);
or_8   g04328(new_n4704, new_n4703, new_n4705);
and_8  g04329(n5645, n137, new_n4706);
nor_6  g04330(new_n4704, new_n4703, new_n4707);
and_8  g04331(new_n4704, new_n4703, new_n4708);
or_8   g04332(new_n4708, new_n4707, new_n4709);
or_8   g04333(new_n4709, new_n4706, new_n4710);
and_8  g04334(new_n4710, new_n4705, new_n4711);
and_8  g04335(new_n4711, new_n4702, new_n4712);
xor_4  g04336(new_n4697, new_n4696, new_n4713);
not_8  g04337(new_n4702, new_n4714);
nor_6  g04338(new_n4709, new_n4706, new_n4715);
or_8   g04339(new_n4715, new_n4707, new_n4716);
or_8   g04340(new_n4716, new_n4714, new_n4717);
or_8   g04341(new_n4711, new_n4702, new_n4718);
and_8  g04342(new_n4718, new_n4717, new_n4719);
and_8  g04343(new_n4719, new_n4713, new_n4720);
or_8   g04344(new_n4720, new_n4712, new_n4721);
and_8  g04345(n11478, n2551, new_n4722_1);
and_8  g04346(n11922, n5283, new_n4723);
xor_4  g04347(new_n4723, new_n4722_1, new_n4724);
xor_4  g04348(new_n4724, new_n4721, new_n4725);
and_8  g04349(new_n4725, new_n4701, new_n4726);
and_8  g04350(new_n4700, new_n4692, new_n4727);
nor_6  g04351(new_n4700, new_n4692, new_n4728);
or_8   g04352(new_n4728, new_n4727, new_n4729);
not_8  g04353(new_n4696, new_n4730);
xor_4  g04354(new_n4697, new_n4730, new_n4731);
and_8  g04355(new_n4716, new_n4714, new_n4732);
or_8   g04356(new_n4732, new_n4712, new_n4733_1);
or_8   g04357(new_n4733_1, new_n4731, new_n4734);
and_8  g04358(new_n4734, new_n4717, new_n4735);
xor_4  g04359(new_n4724, new_n4735, new_n4736);
and_8  g04360(new_n4736, new_n4729, new_n4737);
or_8   g04361(new_n4737, new_n4726, new_n4738);
and_8  g04362(n4805, n2551, new_n4739);
and_8  g04363(n11922, n4805, new_n4740);
and_8  g04364(n5645, n5283, new_n4741);
and_8  g04365(n8665, n4805, new_n4742);
and_8  g04366(new_n4742, new_n4741, new_n4743);
or_8   g04367(new_n4742, new_n4741, new_n4744);
and_8  g04368(n11478, n1067, new_n4745);
and_8  g04369(new_n4745, new_n4744, new_n4746);
or_8   g04370(new_n4746, new_n4743, new_n4747);
and_8  g04371(new_n4747, new_n4740, new_n4748);
nor_6  g04372(new_n4747, new_n4740, new_n4749);
or_8   g04373(new_n4749, new_n4748, new_n4750);
xor_4  g04374(new_n4709, new_n4706, new_n4751);
nor_6  g04375(new_n4751, new_n4750, new_n4752);
or_8   g04376(new_n4752, new_n4748, new_n4753);
nor_6  g04377(new_n4753, new_n4739, new_n4754);
xor_4  g04378(new_n4719, new_n4731, new_n4755);
xor_4  g04379(new_n4753, new_n4739, new_n4756);
and_8  g04380(new_n4756, new_n4755, new_n4757_1);
or_8   g04381(new_n4757_1, new_n4754, new_n4758);
or_8   g04382(new_n4758, new_n4738, new_n4759);
or_8   g04383(new_n4736, new_n4729, new_n4760);
or_8   g04384(new_n4725, new_n4701, new_n4761);
and_8  g04385(new_n4761, new_n4760, new_n4762);
or_8   g04386(new_n4753, new_n4739, new_n4763);
xor_4  g04387(new_n4719, new_n4713, new_n4764);
and_8  g04388(new_n4753, new_n4739, new_n4765);
or_8   g04389(new_n4765, new_n4754, new_n4766);
or_8   g04390(new_n4766, new_n4764, new_n4767);
and_8  g04391(new_n4767, new_n4763, new_n4768);
or_8   g04392(new_n4768, new_n4762, new_n4769);
and_8  g04393(new_n4769, new_n4759, new_n4770);
and_8  g04394(new_n4770, new_n4687, new_n4771);
xor_4  g04395(new_n4751, new_n4750, new_n4772);
xnor_4 g04396(new_n4742, new_n4741, new_n4773);
and_8  g04397(n4805, n1067, new_n4774);
and_8  g04398(n11478, n5645, new_n4775);
and_8  g04399(new_n4775, new_n4774, new_n4776);
and_8  g04400(new_n4776, new_n4773, new_n4777);
and_8  g04401(new_n4777, new_n4772, new_n4778);
not_8  g04402(new_n4778, new_n4779);
xor_4  g04403(new_n4766, new_n4764, new_n4780);
or_8   g04404(new_n4780, new_n4779, new_n4781);
not_8  g04405(new_n4781, new_n4782);
not_8  g04406(new_n4687, new_n4783);
and_8  g04407(new_n4768, new_n4762, new_n4784);
and_8  g04408(new_n4758, new_n4738, new_n4785);
or_8   g04409(new_n4785, new_n4784, new_n4786);
or_8   g04410(new_n4786, new_n4783, new_n4787);
or_8   g04411(new_n4770, new_n4687, new_n4788);
and_8  g04412(new_n4788, new_n4787, new_n4789);
and_8  g04413(new_n4789, new_n4782, new_n4790);
nor_6  g04414(new_n4790, new_n4771, new_n4791);
and_8  g04415(n12826, n11478, new_n4792);
and_8  g04416(n5283, n2551, new_n4793);
and_8  g04417(n4805, n4094, new_n4794);
xnor_4 g04418(new_n4794, new_n4793, new_n4795);
xor_4  g04419(new_n4795, new_n4792, new_n4796);
and_8  g04420(new_n4691, new_n4688, new_n4797);
or_8   g04421(new_n4727, new_n4797, new_n4798);
xor_4  g04422(new_n4798, new_n4796, new_n4799);
and_8  g04423(new_n4690, new_n4689_1, new_n4800);
and_8  g04424(n11922, n137, new_n4801);
xnor_4 g04425(new_n4801, new_n4800, new_n4802);
and_8  g04426(n6797, n1067, new_n4803);
and_8  g04427(n8665, n6294, new_n4804);
and_8  g04428(n5645, n3146, new_n4805_1);
xnor_4 g04429(new_n4805_1, new_n4804, new_n4806);
xor_4  g04430(new_n4806, new_n4803, new_n4807);
xor_4  g04431(new_n4807, new_n4802, new_n4808);
xor_4  g04432(new_n4808, new_n4799, new_n4809);
nand_5 g04433(new_n4724, new_n4721, new_n4810);
nand_5 g04434(new_n4723, new_n4722_1, new_n4811);
not_8  g04435(new_n4811, new_n4812);
and_8  g04436(new_n4726, new_n4812, new_n4813);
and_8  g04437(new_n4760, new_n4811, new_n4814);
or_8   g04438(new_n4814, new_n4813, new_n4815);
and_8  g04439(new_n4815, new_n4810, new_n4816);
or_8   g04440(new_n4816, new_n4809, new_n4817_1);
nor_6  g04441(new_n4808, new_n4799, new_n4818);
and_8  g04442(new_n4808, new_n4799, new_n4819);
or_8   g04443(new_n4819, new_n4818, new_n4820);
not_8  g04444(new_n4810, new_n4821);
or_8   g04445(new_n4760, new_n4811, new_n4822);
or_8   g04446(new_n4726, new_n4812, new_n4823);
and_8  g04447(new_n4823, new_n4822, new_n4824);
or_8   g04448(new_n4824, new_n4821, new_n4825);
or_8   g04449(new_n4825, new_n4820, new_n4826_1);
and_8  g04450(new_n4826_1, new_n4817_1, new_n4827);
xor_4  g04451(new_n4827, new_n4759, new_n4828_1);
or_8   g04452(new_n4828_1, new_n4791, new_n4829);
or_8   g04453(new_n4790, new_n4771, new_n4830);
xor_4  g04454(new_n4827, new_n4784, new_n4831);
or_8   g04455(new_n4831, new_n4830, new_n4832);
and_8  g04456(new_n4832, new_n4829, new_n4833);
and_8  g04457(n3992, n2749, new_n4834);
and_8  g04458(n11876, n6358, new_n4835);
and_8  g04459(n3992, n3754, new_n4836);
or_8   g04460(new_n4836, new_n4835, new_n4837);
and_8  g04461(n10898, n8384, new_n4838);
nor_6  g04462(new_n4836, new_n4835, new_n4839);
and_8  g04463(new_n4836, new_n4835, new_n4840);
or_8   g04464(new_n4840, new_n4839, new_n4841);
or_8   g04465(new_n4841, new_n4838, new_n4842);
and_8  g04466(new_n4842, new_n4837, new_n4843);
and_8  g04467(new_n4843, new_n4834, new_n4844);
not_8  g04468(new_n4834, new_n4845);
nor_6  g04469(new_n4841, new_n4838, new_n4846);
or_8   g04470(new_n4846, new_n4839, new_n4847);
or_8   g04471(new_n4847, new_n4845, new_n4848);
or_8   g04472(new_n4843, new_n4834, new_n4849);
and_8  g04473(new_n4849, new_n4848, new_n4850);
and_8  g04474(n10898, n6358, new_n4851);
and_8  g04475(n11876, n5198, new_n4852);
and_8  g04476(n8384, n3754, new_n4853);
xor_4  g04477(new_n4853, new_n4852, new_n4854);
xor_4  g04478(new_n4854, new_n4851, new_n4855);
and_8  g04479(new_n4855, new_n4850, new_n4856);
or_8   g04480(new_n4856, new_n4844, new_n4857);
and_8  g04481(n8384, n2749, new_n4858);
and_8  g04482(n3992, n159, new_n4859);
xor_4  g04483(new_n4859, new_n4858, new_n4860);
xor_4  g04484(new_n4860, new_n4857, new_n4861);
nand_5 g04485(n6358, n3754, new_n4862);
and_8  g04486(n10898, n5198, new_n4863);
and_8  g04487(n11876, n1471, new_n4864);
xor_4  g04488(new_n4864, new_n4863, new_n4865);
xor_4  g04489(new_n4865, new_n4862, new_n4866);
or_8   g04490(new_n4853, new_n4852, new_n4867);
xnor_4 g04491(new_n4853, new_n4852, new_n4868);
or_8   g04492(new_n4868, new_n4851, new_n4869);
and_8  g04493(new_n4869, new_n4867, new_n4870);
not_8  g04494(new_n4870, new_n4871);
xor_4  g04495(new_n4871, new_n4866, new_n4872);
and_8  g04496(new_n4872, new_n4861, new_n4873);
and_8  g04497(new_n4847, new_n4845, new_n4874);
or_8   g04498(new_n4874, new_n4844, new_n4875);
not_8  g04499(new_n4851, new_n4876);
xor_4  g04500(new_n4854, new_n4876, new_n4877);
or_8   g04501(new_n4877, new_n4875, new_n4878);
and_8  g04502(new_n4878, new_n4848, new_n4879);
xor_4  g04503(new_n4860, new_n4879, new_n4880);
xor_4  g04504(new_n4870, new_n4866, new_n4881);
and_8  g04505(new_n4881, new_n4880, new_n4882);
or_8   g04506(new_n4882, new_n4873, new_n4883);
and_8  g04507(n7236, n159, new_n4884);
and_8  g04508(n7236, n2749, new_n4885);
and_8  g04509(n11876, n8384, new_n4886);
and_8  g04510(n7236, n3754, new_n4887);
or_8   g04511(new_n4887, new_n4886, new_n4888);
and_8  g04512(n11876, n7236, new_n4889);
and_8  g04513(new_n4889, new_n4853, new_n4890);
and_8  g04514(n10898, n3992, new_n4891);
or_8   g04515(new_n4891, new_n4890, new_n4892);
and_8  g04516(new_n4892, new_n4888, new_n4893);
and_8  g04517(new_n4893, new_n4885, new_n4894);
xor_4  g04518(new_n4893, new_n4885, new_n4895);
and_8  g04519(new_n4841, new_n4838, new_n4896);
or_8   g04520(new_n4896, new_n4846, new_n4897);
and_8  g04521(new_n4897, new_n4895, new_n4898);
or_8   g04522(new_n4898, new_n4894, new_n4899);
nor_6  g04523(new_n4899, new_n4884, new_n4900);
xor_4  g04524(new_n4877, new_n4850, new_n4901);
xor_4  g04525(new_n4899, new_n4884, new_n4902);
and_8  g04526(new_n4902, new_n4901, new_n4903_1);
or_8   g04527(new_n4903_1, new_n4900, new_n4904);
or_8   g04528(new_n4904, new_n4883, new_n4905);
and_8  g04529(new_n4864, new_n4863, new_n4906);
and_8  g04530(n6358, n2749, new_n4907);
xnor_4 g04531(new_n4907, new_n4906, new_n4908);
and_8  g04532(n10898, n1471, new_n4909);
and_8  g04533(n5198, n3754, new_n4910);
and_8  g04534(n11876, n7646, new_n4911);
xnor_4 g04535(new_n4911, new_n4910, new_n4912);
xor_4  g04536(new_n4912, new_n4909, new_n4913);
nor_6  g04537(new_n4913, new_n4908, new_n4914);
and_8  g04538(new_n4913, new_n4908, new_n4915);
or_8   g04539(new_n4915, new_n4914, new_n4916);
and_8  g04540(n6358, n3754, new_n4917);
or_8   g04541(new_n4865, new_n4917, new_n4918);
or_8   g04542(new_n4870, new_n4866, new_n4919);
and_8  g04543(new_n4919, new_n4918, new_n4920);
and_8  g04544(n3992, n1510, new_n4921_1);
not_8  g04545(new_n4921_1, new_n4922);
and_8  g04546(n8384, n159, new_n4923);
and_8  g04547(n12247, n7236, new_n4924);
xnor_4 g04548(new_n4924, new_n4923, new_n4925);
xor_4  g04549(new_n4925, new_n4922, new_n4926);
xor_4  g04550(new_n4926, new_n4920, new_n4927);
xor_4  g04551(new_n4927, new_n4916, new_n4928_1);
nand_5 g04552(new_n4860, new_n4857, new_n4929);
nand_5 g04553(new_n4859, new_n4858, new_n4930);
not_8  g04554(new_n4930, new_n4931);
and_8  g04555(new_n4873, new_n4931, new_n4932);
or_8   g04556(new_n4881, new_n4880, new_n4933);
and_8  g04557(new_n4933, new_n4930, new_n4934);
or_8   g04558(new_n4934, new_n4932, new_n4935);
and_8  g04559(new_n4935, new_n4929, new_n4936);
or_8   g04560(new_n4936, new_n4928_1, new_n4937);
nor_6  g04561(new_n4927, new_n4916, new_n4938_1);
and_8  g04562(new_n4927, new_n4916, new_n4939);
or_8   g04563(new_n4939, new_n4938_1, new_n4940);
not_8  g04564(new_n4929, new_n4941);
or_8   g04565(new_n4933, new_n4930, new_n4942);
or_8   g04566(new_n4873, new_n4931, new_n4943);
and_8  g04567(new_n4943, new_n4942, new_n4944);
or_8   g04568(new_n4944, new_n4941, new_n4945);
or_8   g04569(new_n4945, new_n4940, new_n4946);
and_8  g04570(new_n4946, new_n4937, new_n4947);
xor_4  g04571(new_n4947, new_n4905, new_n4948);
and_8  g04572(n7236, n1510, new_n4949);
or_8   g04573(new_n4872, new_n4861, new_n4950);
and_8  g04574(new_n4950, new_n4933, new_n4951);
nor_6  g04575(new_n4903_1, new_n4900, new_n4952);
or_8   g04576(new_n4952, new_n4951, new_n4953);
and_8  g04577(new_n4953, new_n4905, new_n4954);
and_8  g04578(new_n4954, new_n4949, new_n4955);
nor_6  g04579(new_n4897, new_n4895, new_n4956);
or_8   g04580(new_n4956, new_n4898, new_n4957);
nor_6  g04581(new_n4887, new_n4886, new_n4958);
or_8   g04582(new_n4890, new_n4958, new_n4959);
and_8  g04583(n11876, n3992, new_n4960);
and_8  g04584(n10898, n7236, new_n4961);
and_8  g04585(new_n4961, new_n4960, new_n4962);
nand_5 g04586(new_n4962, new_n4959, new_n4963);
or_8   g04587(new_n4963, new_n4957, new_n4964);
xor_4  g04588(new_n4902, new_n4901, new_n4965);
or_8   g04589(new_n4965, new_n4964, new_n4966);
not_8  g04590(new_n4966, new_n4967);
not_8  g04591(new_n4949, new_n4968);
and_8  g04592(new_n4952, new_n4951, new_n4969);
and_8  g04593(new_n4904, new_n4883, new_n4970_1);
or_8   g04594(new_n4970_1, new_n4969, new_n4971_1);
or_8   g04595(new_n4971_1, new_n4968, new_n4972);
or_8   g04596(new_n4954, new_n4949, new_n4973);
and_8  g04597(new_n4973, new_n4972, new_n4974);
and_8  g04598(new_n4974, new_n4967, new_n4975);
nor_6  g04599(new_n4975, new_n4955, new_n4976);
or_8   g04600(new_n4976, new_n4948, new_n4977);
xor_4  g04601(new_n4947, new_n4969, new_n4978);
or_8   g04602(new_n4975, new_n4955, new_n4979);
or_8   g04603(new_n4979, new_n4978, new_n4980);
and_8  g04604(new_n4980, new_n4977, new_n4981);
or_8   g04605(new_n4981, new_n4833, new_n4982);
and_8  g04606(new_n4831, new_n4830, new_n4983);
and_8  g04607(new_n4828_1, new_n4791, new_n4984);
or_8   g04608(new_n4984, new_n4983, new_n4985);
and_8  g04609(new_n4979, new_n4978, new_n4986);
and_8  g04610(new_n4976, new_n4948, new_n4987);
or_8   g04611(new_n4987, new_n4986, new_n4988);
or_8   g04612(new_n4988, new_n4985, new_n4989);
and_8  g04613(new_n4989, new_n4982, new_n4990);
xor_4  g04614(new_n4789, new_n4782, new_n4991);
xor_4  g04615(new_n4974, new_n4967, new_n4992);
or_8   g04616(new_n4992, new_n4991, new_n4993);
xor_4  g04617(new_n4789, new_n4781, new_n4994);
xor_4  g04618(new_n4974, new_n4966, new_n4995);
and_8  g04619(new_n4995, new_n4994, new_n4996);
and_8  g04620(new_n4992, new_n4991, new_n4997);
or_8   g04621(new_n4997, new_n4996, new_n4998);
xor_4  g04622(new_n4965, new_n4964, new_n4999);
xor_4  g04623(new_n4777, new_n4772, new_n5000);
xor_4  g04624(new_n4963, new_n4957, new_n5001);
or_8   g04625(new_n5001, new_n5000, new_n5002);
xor_4  g04626(new_n4961, new_n4960, new_n5003);
xor_4  g04627(new_n4775, new_n4774, new_n5004);
nor_6  g04628(new_n5004, new_n5003, new_n5005);
not_8  g04629(new_n4889, new_n5006);
not_8  g04630(n5645, new_n5007);
or_8   g04631(new_n5007, new_n3601, new_n5008);
or_8   g04632(new_n5008, new_n5006, new_n5009);
xor_4  g04633(new_n5004, new_n5003, new_n5010);
and_8  g04634(new_n5010, new_n5009, new_n5011);
or_8   g04635(new_n5011, new_n5005, new_n5012);
and_8  g04636(new_n5008, new_n4745, new_n5013);
not_8  g04637(new_n5013, new_n5014);
or_8   g04638(new_n5014, new_n4744, new_n5015);
or_8   g04639(new_n5013, new_n4773, new_n5016);
and_8  g04640(new_n5016, new_n5015, new_n5017);
and_8  g04641(new_n5017, new_n5012, new_n5018);
xor_4  g04642(new_n5017, new_n5012, new_n5019);
nand_5 g04643(new_n4891, new_n5006, new_n5020);
and_8  g04644(new_n5020, new_n4959, new_n5021);
nor_6  g04645(new_n5020, new_n4958, new_n5022);
or_8   g04646(new_n5022, new_n5021, new_n5023);
and_8  g04647(new_n5023, new_n5019, new_n5024);
or_8   g04648(new_n5024, new_n5018, new_n5025);
not_8  g04649(new_n5025, new_n5026);
nor_6  g04650(new_n5001, new_n5000, new_n5027);
and_8  g04651(new_n5001, new_n5000, new_n5028);
or_8   g04652(new_n5028, new_n5027, new_n5029);
or_8   g04653(new_n5029, new_n5026, new_n5030_1);
and_8  g04654(new_n5030_1, new_n5002, new_n5031);
or_8   g04655(new_n5031, new_n4999, new_n5032);
xor_4  g04656(new_n4780, new_n4779, new_n5033);
and_8  g04657(new_n4965, new_n4964, new_n5034_1);
or_8   g04658(new_n5034_1, new_n4967, new_n5035);
xor_4  g04659(new_n5031, new_n5035, new_n5036);
or_8   g04660(new_n5036, new_n5033, new_n5037);
and_8  g04661(new_n5037, new_n5032, new_n5038);
or_8   g04662(new_n5038, new_n4998, new_n5039);
and_8  g04663(new_n5039, new_n4993, new_n5040);
xor_4  g04664(new_n5040, new_n4990, new_n5041);
or_8   g04665(new_n5041, new_n4686_1, new_n5042);
or_8   g04666(new_n4657, new_n4629, new_n5043);
or_8   g04667(new_n4655, new_n4630, new_n5044);
and_8  g04668(new_n5044, new_n5043, new_n5045);
xor_4  g04669(new_n4685, new_n5045, new_n5046);
and_8  g04670(new_n4988, new_n4985, new_n5047);
and_8  g04671(new_n4981, new_n4833, new_n5048);
or_8   g04672(new_n5048, new_n5047, new_n5049);
xor_4  g04673(new_n5040, new_n5049, new_n5050);
or_8   g04674(new_n5050, new_n5046, new_n5051);
and_8  g04675(new_n5051, new_n5042, new_n5052);
xor_4  g04676(new_n4683, new_n4680, new_n5053);
or_8   g04677(new_n4995, new_n4994, new_n5054);
and_8  g04678(new_n5054, new_n4993, new_n5055);
nor_6  g04679(new_n5031, new_n4999, new_n5056);
not_8  g04680(new_n5033, new_n5057);
xor_4  g04681(new_n5031, new_n4999, new_n5058);
and_8  g04682(new_n5058, new_n5057, new_n5059);
or_8   g04683(new_n5059, new_n5056, new_n5060);
or_8   g04684(new_n5060, new_n5055, new_n5061);
and_8  g04685(new_n5061, new_n5039, new_n5062);
and_8  g04686(new_n5062, new_n5053, new_n5063);
xor_4  g04687(new_n4679, new_n4678, new_n5064);
not_8  g04688(new_n5064, new_n5065);
xor_4  g04689(new_n4676, new_n4670, new_n5066);
not_8  g04690(new_n5066, new_n5067);
xor_4  g04691(new_n5001, new_n5000, new_n5068);
or_8   g04692(new_n5068, new_n5025, new_n5069_1);
and_8  g04693(new_n5069_1, new_n5030_1, new_n5070);
or_8   g04694(new_n5070, new_n5067, new_n5071);
xor_4  g04695(new_n5070, new_n5066, new_n5072);
nor_6  g04696(new_n5023, new_n5019, new_n5073);
or_8   g04697(new_n5073, new_n5024, new_n5074);
not_8  g04698(new_n4673, new_n5075);
and_8  g04699(new_n5075, new_n4614, new_n5076);
nor_6  g04700(new_n5076, new_n4675, new_n5077);
and_8  g04701(new_n5077, new_n5074, new_n5078);
xor_4  g04702(new_n5023, new_n5019, new_n5079);
or_8   g04703(new_n5076, new_n4675, new_n5080);
or_8   g04704(new_n5080, new_n5079, new_n5081);
or_8   g04705(new_n5077, new_n5074, new_n5082);
and_8  g04706(new_n5082, new_n5081, new_n5083);
xnor_4 g04707(new_n5010, new_n5009, new_n5084);
and_8  g04708(n9400, n6703, new_n5085);
and_8  g04709(n9640, n6877, new_n5086);
xor_4  g04710(new_n5086, new_n5085, new_n5087);
and_8  g04711(new_n5087, new_n5084, new_n5088);
xor_4  g04712(new_n5008, new_n5006, new_n5089);
and_8  g04713(new_n5089, new_n4671, new_n5090);
xor_4  g04714(new_n5087, new_n5084, new_n5091);
and_8  g04715(new_n5091, new_n5090, new_n5092);
or_8   g04716(new_n5092, new_n5088, new_n5093);
and_8  g04717(new_n5093, new_n5083, new_n5094_1);
nor_6  g04718(new_n5094_1, new_n5078, new_n5095);
or_8   g04719(new_n5095, new_n5072, new_n5096);
and_8  g04720(new_n5096, new_n5071, new_n5097);
and_8  g04721(new_n5097, new_n5065, new_n5098);
xor_4  g04722(new_n5036, new_n5033, new_n5099);
and_8  g04723(new_n5068, new_n5025, new_n5100);
and_8  g04724(new_n5029, new_n5026, new_n5101);
or_8   g04725(new_n5101, new_n5100, new_n5102);
and_8  g04726(new_n5102, new_n5066, new_n5103);
xor_4  g04727(new_n5102, new_n5066, new_n5104);
or_8   g04728(new_n5094_1, new_n5078, new_n5105_1);
and_8  g04729(new_n5105_1, new_n5104, new_n5106);
or_8   g04730(new_n5106, new_n5103, new_n5107);
or_8   g04731(new_n5107, new_n5064, new_n5108);
or_8   g04732(new_n5097, new_n5065, new_n5109);
and_8  g04733(new_n5109, new_n5108, new_n5110);
and_8  g04734(new_n5110, new_n5099, new_n5111);
or_8   g04735(new_n5111, new_n5098, new_n5112);
xor_4  g04736(new_n4683, new_n4681, new_n5113);
and_8  g04737(new_n5060, new_n5055, new_n5114);
and_8  g04738(new_n5038, new_n4998, new_n5115);
or_8   g04739(new_n5115, new_n5114, new_n5116);
or_8   g04740(new_n5116, new_n5113, new_n5117);
or_8   g04741(new_n5062, new_n5053, new_n5118);
and_8  g04742(new_n5118, new_n5117, new_n5119);
and_8  g04743(new_n5119, new_n5112, new_n5120);
or_8   g04744(new_n5120, new_n5063, new_n5121);
and_8  g04745(new_n5121, new_n5052, new_n5122);
and_8  g04746(new_n5050, new_n5046, new_n5123);
and_8  g04747(new_n5041, new_n4686_1, new_n5124);
or_8   g04748(new_n5124, new_n5123, new_n5125);
nor_6  g04749(new_n5120, new_n5063, new_n5126);
and_8  g04750(new_n5126, new_n5125, new_n5127);
or_8   g04751(new_n5127, new_n5122, new_n5128);
and_8  g04752(new_n5128, new_n4571, new_n5129);
not_8  g04753(new_n4571, new_n5130);
or_8   g04754(new_n5126, new_n5125, new_n5131);
or_8   g04755(new_n5121, new_n5052, new_n5132_1);
and_8  g04756(new_n5132_1, new_n5131, new_n5133);
or_8   g04757(new_n5133, new_n5130, new_n5134);
or_8   g04758(new_n5128, new_n4571, new_n5135);
and_8  g04759(new_n5135, new_n5134, new_n5136);
xor_4  g04760(new_n4568, new_n4566, new_n5137);
nor_6  g04761(new_n5119, new_n5112, new_n5138);
or_8   g04762(new_n5138, new_n5120, new_n5139);
and_8  g04763(new_n5139, new_n5137, new_n5140);
xor_4  g04764(new_n4565, new_n4564, new_n5141);
not_8  g04765(new_n5099, new_n5142);
xor_4  g04766(new_n5110, new_n5142, new_n5143);
or_8   g04767(new_n5143, new_n5141, new_n5144);
and_8  g04768(new_n5107, new_n5064, new_n5145);
or_8   g04769(new_n5145, new_n5098, new_n5146);
or_8   g04770(new_n5146, new_n5142, new_n5147);
or_8   g04771(new_n5110, new_n5099, new_n5148);
and_8  g04772(new_n5148, new_n5147, new_n5149);
xor_4  g04773(new_n5149, new_n5141, new_n5150);
xor_4  g04774(new_n4563, new_n4557, new_n5151);
xor_4  g04775(new_n5095, new_n5072, new_n5152);
nor_6  g04776(new_n5152, new_n5151, new_n5153_1);
not_8  g04777(new_n5153_1, new_n5154);
xor_4  g04778(new_n5093, new_n5083, new_n5155);
not_8  g04779(new_n4558, new_n5156);
and_8  g04780(n7862, n1798, new_n5157);
not_8  g04781(new_n5157, new_n5158);
and_8  g04782(new_n5158, new_n4499_1, new_n5159);
or_8   g04783(new_n5159, new_n5156, new_n5160);
nand_5 g04784(new_n5159, new_n4498, new_n5161);
and_8  g04785(new_n5161, new_n5160, new_n5162);
or_8   g04786(new_n5162, new_n5155, new_n5163);
xor_4  g04787(new_n5162, new_n5155, new_n5164);
not_8  g04788(new_n5164, new_n5165);
xor_4  g04789(new_n5089, new_n4671, new_n5166);
and_8  g04790(new_n5166, new_n5157, new_n5167);
xor_4  g04791(new_n4560, new_n4559, new_n5168);
or_8   g04792(new_n5168, new_n5167, new_n5169);
xor_4  g04793(new_n5091, new_n5090, new_n5170);
xor_4  g04794(new_n5168, new_n5167, new_n5171);
not_8  g04795(new_n5171, new_n5172);
or_8   g04796(new_n5172, new_n5170, new_n5173);
and_8  g04797(new_n5173, new_n5169, new_n5174);
or_8   g04798(new_n5174, new_n5165, new_n5175);
and_8  g04799(new_n5175, new_n5163, new_n5176);
and_8  g04800(new_n5152, new_n5151, new_n5177);
or_8   g04801(new_n5177, new_n5153_1, new_n5178);
or_8   g04802(new_n5178, new_n5176, new_n5179);
and_8  g04803(new_n5179, new_n5154, new_n5180);
or_8   g04804(new_n5180, new_n5150, new_n5181);
and_8  g04805(new_n5181, new_n5144, new_n5182);
not_8  g04806(new_n5137, new_n5183);
xor_4  g04807(new_n5119, new_n5112, new_n5184);
or_8   g04808(new_n5184, new_n5183, new_n5185);
or_8   g04809(new_n5139, new_n5137, new_n5186);
and_8  g04810(new_n5186, new_n5185, new_n5187);
and_8  g04811(new_n5187, new_n5182, new_n5188);
or_8   g04812(new_n5188, new_n5140, new_n5189);
and_8  g04813(new_n5189, new_n5136, new_n5190);
or_8   g04814(new_n5190, new_n5129, new_n5191_1);
xor_4  g04815(new_n4667, new_n4660, new_n5192);
and_8  g04816(new_n5192, new_n4680, new_n5193);
or_8   g04817(new_n5193, new_n4668, new_n5194);
and_8  g04818(new_n5194, new_n5045, new_n5195);
or_8   g04819(new_n5195, new_n4656, new_n5196);
nand_5 g04820(n7862, n753, new_n5197);
not_8  g04821(new_n4798, new_n5198_1);
and_8  g04822(new_n5198_1, new_n4796, new_n5199);
or_8   g04823(new_n4818, new_n5199, new_n5200);
xor_4  g04824(new_n5200, new_n5197, new_n5201);
nand_5 g04825(new_n4801, new_n4800, new_n5202);
or_8   g04826(new_n4807, new_n4802, new_n5203);
and_8  g04827(new_n5203, new_n5202, new_n5204);
and_8  g04828(n3146, n1067, new_n5205);
and_8  g04829(n2551, n137, new_n5206);
xor_4  g04830(new_n5206, new_n5205, new_n5207);
and_8  g04831(n12826, n5283, new_n5208);
and_8  g04832(n8665, n6797, new_n5209);
xor_4  g04833(new_n5209, new_n5208, new_n5210);
xnor_4 g04834(new_n5210, new_n5207, new_n5211);
xor_4  g04835(new_n5211, new_n5204, new_n5212_1);
and_8  g04836(new_n4907, new_n4906, new_n5213);
or_8   g04837(new_n4914, new_n5213, new_n5214);
or_8   g04838(new_n4924, new_n4923, new_n5215);
or_8   g04839(new_n4925, new_n4921_1, new_n5216);
and_8  g04840(new_n5216, new_n5215, new_n5217);
and_8  g04841(n8384, n1510, new_n5218);
and_8  g04842(n5198, n2749, new_n5219);
xor_4  g04843(new_n5219, new_n5218, new_n5220);
xnor_4 g04844(new_n5220, new_n5217, new_n5221);
xor_4  g04845(new_n5221, new_n5214, new_n5222);
xor_4  g04846(new_n5222, new_n5212_1, new_n5223);
xor_4  g04847(new_n5223, new_n5201, new_n5224);
not_8  g04848(new_n5224, new_n5225);
or_8   g04849(new_n5225, new_n5196, new_n5226);
or_8   g04850(new_n4685, new_n4659, new_n5227);
and_8  g04851(new_n5227, new_n5043, new_n5228);
or_8   g04852(new_n5224, new_n5228, new_n5229);
and_8  g04853(new_n5229, new_n5226, new_n5230);
not_8  g04854(new_n4534, new_n5231);
or_8   g04855(new_n4539, new_n4531, new_n5232);
and_8  g04856(new_n5232, new_n5231, new_n5233);
and_8  g04857(new_n4817_1, new_n4822, new_n5234);
xor_4  g04858(new_n5234, new_n5233, new_n5235);
and_8  g04859(n12511, n7236, new_n5236);
and_8  g04860(n6826, n1798, new_n5237);
xor_4  g04861(new_n5237, new_n5236, new_n5238);
or_8   g04862(new_n4805_1, new_n4804, new_n5239);
or_8   g04863(new_n4806, new_n4803, new_n5240_1);
and_8  g04864(new_n5240_1, new_n5239, new_n5241);
or_8   g04865(new_n4911, new_n4910, new_n5242);
or_8   g04866(new_n4912, new_n4909, new_n5243);
and_8  g04867(new_n5243, new_n5242, new_n5244);
xor_4  g04868(new_n5244, new_n5241, new_n5245);
xor_4  g04869(new_n5245, new_n5238, new_n5246);
and_8  g04870(n6358, n159, new_n5247);
or_8   g04871(new_n4795, new_n4792, new_n5248);
and_8  g04872(new_n5248, new_n4793, new_n5249);
and_8  g04873(n11478, n4094, new_n5250);
nand_5 g04874(new_n5250, new_n5249, new_n5251);
and_8  g04875(new_n5250, new_n4783, new_n5252);
or_8   g04876(new_n5252, new_n5249, new_n5253);
and_8  g04877(new_n5253, new_n5251, new_n5254);
xor_4  g04878(new_n5254, new_n5247, new_n5255);
xor_4  g04879(new_n5255, new_n5246, new_n5256);
not_8  g04880(new_n5256, new_n5257_1);
xor_4  g04881(new_n5257_1, new_n5235, new_n5258);
and_8  g04882(new_n5258, new_n5230, new_n5259);
and_8  g04883(new_n5224, new_n5228, new_n5260);
and_8  g04884(new_n5225, new_n5196, new_n5261);
or_8   g04885(new_n5261, new_n5260, new_n5262);
xor_4  g04886(new_n5256, new_n5235, new_n5263);
and_8  g04887(new_n5263, new_n5262, new_n5264);
or_8   g04888(new_n5264, new_n5259, new_n5265);
and_8  g04889(new_n4937, new_n4942, new_n5266);
and_8  g04890(n5645, n4938, new_n5267);
and_8  g04891(n10898, n7646, new_n5268);
xor_4  g04892(new_n5268, new_n5267, new_n5269);
xnor_4 g04893(new_n5269, new_n5266, new_n5270);
xor_4  g04894(new_n5270, new_n5265, new_n5271);
nor_6  g04895(new_n5040, new_n5049, new_n5272);
or_8   g04896(new_n5272, new_n5047, new_n5273);
and_8  g04897(n11922, n6294, new_n5274);
nand_5 g04898(new_n4827, new_n4784, new_n5275);
and_8  g04899(new_n4829, new_n5275, new_n5276);
xor_4  g04900(new_n5276, new_n5274, new_n5277);
or_8   g04901(new_n4543, new_n4511, new_n5278);
or_8   g04902(new_n4570, new_n4545, new_n5279);
and_8  g04903(new_n5279, new_n5278, new_n5280);
and_8  g04904(new_n4603, new_n4652, new_n5281);
and_8  g04905(new_n4654, new_n4650, new_n5282);
or_8   g04906(new_n5282, new_n5281, new_n5283_1);
xnor_4 g04907(new_n4637, new_n4634_1, new_n5284);
or_8   g04908(new_n5284, new_n4633, new_n5285);
or_8   g04909(new_n4648, new_n4639, new_n5286);
and_8  g04910(new_n5286, new_n5285, new_n5287);
nand_5 g04911(new_n4645, new_n4644, new_n5288);
or_8   g04912(new_n4645, new_n4644, new_n5289);
nand_5 g04913(new_n5289, new_n4643, new_n5290);
and_8  g04914(new_n5290, new_n5288, new_n5291);
and_8  g04915(n4203, n3022, new_n5292);
and_8  g04916(n11023, n4187, new_n5293);
xor_4  g04917(new_n5293, new_n5292, new_n5294);
xor_4  g04918(new_n5294, new_n5291, new_n5295);
and_8  g04919(n7456, n5240, new_n5296);
and_8  g04920(n12753, n9640, new_n5297);
xor_4  g04921(new_n5297, new_n5296, new_n5298);
and_8  g04922(n9583, n1333, new_n5299);
and_8  g04923(n12591, n11821, new_n5300);
xor_4  g04924(new_n5300, new_n5299, new_n5301);
xnor_4 g04925(new_n5301, new_n5298, new_n5302);
xor_4  g04926(new_n5302, new_n5295, new_n5303);
xor_4  g04927(new_n5303, new_n5287, new_n5304);
xnor_4 g04928(new_n4519, new_n4516_1, new_n5305_1);
or_8   g04929(new_n5305_1, new_n4515, new_n5306);
or_8   g04930(new_n4530, new_n4521, new_n5307);
and_8  g04931(new_n5307, new_n5306, new_n5308);
nand_5 g04932(n9080, n3932, new_n5309);
and_8  g04933(n10174, n6703, new_n5310);
and_8  g04934(n6877, n2278, new_n5311);
xor_4  g04935(new_n5311, new_n5310, new_n5312);
xor_4  g04936(new_n5312, new_n5309, new_n5313);
xor_4  g04937(new_n5313, new_n5308, new_n5314_1);
xor_4  g04938(new_n5314_1, new_n5304, new_n5315);
xor_4  g04939(new_n5315, new_n5283_1, new_n5316);
not_8  g04940(new_n5316, new_n5317);
or_8   g04941(new_n5317, new_n5280, new_n5318);
or_8   g04942(new_n4540, new_n4512, new_n5319_1);
and_8  g04943(new_n5319_1, new_n5278, new_n5320_1);
not_8  g04944(new_n4566, new_n5321);
xor_4  g04945(new_n4554, new_n4546, new_n5322);
and_8  g04946(new_n5322, new_n5321, new_n5323);
or_8   g04947(new_n5323, new_n4555, new_n5324);
and_8  g04948(new_n5324, new_n5320_1, new_n5325);
or_8   g04949(new_n5325, new_n4541, new_n5326);
or_8   g04950(new_n5316, new_n5326, new_n5327);
and_8  g04951(new_n5327, new_n5318, new_n5328);
nor_6  g04952(new_n5328, new_n5277, new_n5329);
and_8  g04953(new_n5328, new_n5277, new_n5330);
or_8   g04954(new_n5330, new_n5329, new_n5331_1);
or_8   g04955(new_n5331_1, new_n5273, new_n5332);
nor_6  g04956(new_n5272, new_n5047, new_n5333);
xor_4  g04957(new_n5328, new_n5277, new_n5334);
or_8   g04958(new_n5334, new_n5333, new_n5335);
and_8  g04959(new_n5335, new_n5332, new_n5336);
xor_4  g04960(new_n5336, new_n5271, new_n5337);
xor_4  g04961(new_n5337, new_n5191_1, new_n5338);
nor_6  g04962(new_n4926, new_n4920, new_n5339);
or_8   g04963(new_n4939, new_n5339, new_n5340);
nand_5 g04964(new_n4523, new_n4522, new_n5341);
or_8   g04965(new_n4529, new_n4524, new_n5342);
and_8  g04966(new_n5342, new_n5341, new_n5343);
and_8  g04967(new_n4636, new_n4635, new_n5344);
or_8   g04968(new_n4636, new_n4635, new_n5345);
and_8  g04969(new_n5345, new_n4634_1, new_n5346);
or_8   g04970(new_n5346, new_n5344, new_n5347);
xor_4  g04971(new_n5347, new_n5343, new_n5348);
or_8   g04972(new_n4518, new_n4517, new_n5349);
or_8   g04973(new_n4519, new_n4516_1, new_n5350);
and_8  g04974(new_n5350, new_n5349, new_n5351);
and_8  g04975(new_n4527, new_n4526, new_n5352);
or_8   g04976(new_n4527, new_n4526, new_n5353);
and_8  g04977(new_n5353, new_n4525, new_n5354);
or_8   g04978(new_n5354, new_n5352, new_n5355);
and_8  g04979(n10278, n2464, new_n5356);
and_8  g04980(n11757, n11662, new_n5357);
xor_4  g04981(new_n5357, new_n5356, new_n5358);
and_8  g04982(n10327, n3172, new_n5359);
and_8  g04983(n11423, n9400, new_n5360);
xor_4  g04984(new_n5360, new_n5359, new_n5361);
xor_4  g04985(new_n5361, new_n5358, new_n5362);
xor_4  g04986(new_n5362, new_n5355, new_n5363);
xor_4  g04987(new_n5363, new_n5351, new_n5364);
xor_4  g04988(new_n5364, new_n5348, new_n5365);
xor_4  g04989(new_n5365, new_n5340, new_n5366);
and_8  g04990(n3754, n1471, new_n5367);
and_8  g04991(n11311, n10451, new_n5368);
xor_4  g04992(new_n5368, new_n5367, new_n5369);
nand_5 g04993(new_n4641, new_n4640, new_n5370);
or_8   g04994(new_n4647, new_n4642, new_n5371);
and_8  g04995(new_n5371, new_n5370, new_n5372);
nand_5 g04996(n11876, n4722, new_n5373);
and_8  g04997(n10685, n4805, new_n5374);
and_8  g04998(n12247, n3992, new_n5375);
xor_4  g04999(new_n5375, new_n5374, new_n5376);
xor_4  g05000(new_n5376, new_n5373, new_n5377);
xor_4  g05001(new_n5377, new_n5372, new_n5378);
xor_4  g05002(new_n5378, new_n5369, new_n5379);
xor_4  g05003(new_n5379, new_n5366, new_n5380);
nand_5 g05004(new_n4947, new_n4969, new_n5381);
and_8  g05005(new_n4977, new_n5381, new_n5382);
and_8  g05006(new_n5131, new_n5042, new_n5383);
xor_4  g05007(new_n5383, new_n5382, new_n5384);
xor_4  g05008(new_n5384, new_n5380, new_n5385);
and_8  g05009(new_n5385, new_n5338, new_n5386);
and_8  g05010(new_n5133, new_n5130, new_n5387);
or_8   g05011(new_n5387, new_n5129, new_n5388);
not_8  g05012(new_n5144, new_n5389);
not_8  g05013(new_n5141, new_n5390);
xor_4  g05014(new_n5149, new_n5390, new_n5391);
nor_6  g05015(new_n5178, new_n5176, new_n5392);
or_8   g05016(new_n5392, new_n5153_1, new_n5393);
and_8  g05017(new_n5393, new_n5391, new_n5394);
or_8   g05018(new_n5394, new_n5389, new_n5395);
and_8  g05019(new_n5184, new_n5183, new_n5396);
or_8   g05020(new_n5396, new_n5140, new_n5397);
or_8   g05021(new_n5397, new_n5395, new_n5398);
and_8  g05022(new_n5398, new_n5185, new_n5399);
or_8   g05023(new_n5399, new_n5388, new_n5400);
and_8  g05024(new_n5400, new_n5134, new_n5401);
xor_4  g05025(new_n5337, new_n5401, new_n5402);
not_8  g05026(new_n5380, new_n5403);
xor_4  g05027(new_n5384, new_n5403, new_n5404);
and_8  g05028(new_n5404, new_n5402, new_n5405);
or_8   g05029(new_n5405, new_n5386, n1269);
and_8  g05030(n10223, n4312, new_n5407);
and_8  g05031(n12705, n7265, new_n5408);
and_8  g05032(n4312, n2879, new_n5409);
xnor_4 g05033(new_n5408, new_n1060, new_n5410);
or_8   g05034(new_n5410, new_n5409, new_n5411_1);
and_8  g05035(new_n5411_1, new_n5408, new_n5412);
nor_6  g05036(new_n5412, new_n5407, new_n5413);
or_8   g05037(new_n5412, new_n1066, new_n5414);
and_8  g05038(new_n5414, new_n5407, new_n5415);
or_8   g05039(new_n5415, new_n5413, new_n5416);
and_8  g05040(n12025, n7265, new_n5417);
and_8  g05041(n12705, n2879, new_n5418);
xnor_4 g05042(new_n5418, new_n5417, new_n5419);
xor_4  g05043(new_n5419, new_n5416, new_n5420);
and_8  g05044(n9195, n5964, new_n5421);
and_8  g05045(n4634, n1097, new_n5422);
xor_4  g05046(new_n5422, new_n5421, new_n5423);
xor_4  g05047(new_n5423, new_n5420, new_n5424);
and_8  g05048(n5964, n4634, new_n5425);
or_8   g05049(new_n1068, new_n1067_1, new_n5426);
and_8  g05050(new_n1068, new_n1067_1, new_n5427);
or_8   g05051(new_n5427, new_n1066, new_n5428);
and_8  g05052(new_n5428, new_n5426, new_n5429);
and_8  g05053(new_n5429, new_n5425, new_n5430);
xnor_4 g05054(new_n5410, new_n5409, new_n5431);
xor_4  g05055(new_n5429, new_n5425, new_n5432);
and_8  g05056(new_n5432, new_n5431, new_n5433);
or_8   g05057(new_n5433, new_n5430, new_n5434);
xor_4  g05058(new_n5434, new_n5424, new_n5435_1);
and_8  g05059(n9195, n5305, new_n5436);
and_8  g05060(new_n1064, new_n1055, new_n5437);
and_8  g05061(new_n1070, new_n1065, new_n5438);
or_8   g05062(new_n5438, new_n5437, new_n5439);
or_8   g05063(new_n5439, new_n5436, new_n5440);
nor_6  g05064(new_n5432, new_n5431, new_n5441);
or_8   g05065(new_n5441, new_n5433, new_n5442);
xor_4  g05066(new_n5439, new_n5436, new_n5443);
nand_5 g05067(new_n5443, new_n5442, new_n5444);
and_8  g05068(new_n5444, new_n5440, new_n5445);
and_8  g05069(new_n5445, new_n5435_1, new_n5446);
not_8  g05070(new_n5446, new_n5447);
not_8  g05071(new_n5415, new_n5448);
or_8   g05072(new_n5419, new_n5416, new_n5449);
and_8  g05073(new_n5449, new_n5448, new_n5450);
and_8  g05074(n5964, n2253, new_n5451);
and_8  g05075(n9195, n1097, new_n5452);
and_8  g05076(n5305, n3865, new_n5453);
xnor_4 g05077(new_n5453, new_n5452, new_n5454);
xor_4  g05078(new_n5454, new_n5451, new_n5455);
xor_4  g05079(new_n5455, new_n5450, new_n5456);
and_8  g05080(new_n5418, new_n5417, new_n5457);
and_8  g05081(n4634, n4312, new_n5458);
xnor_4 g05082(new_n5458, new_n5457, new_n5459);
and_8  g05083(n12025, n2879, new_n5460);
and_8  g05084(n11257, n7265, new_n5461);
and_8  g05085(n12705, n10223, new_n5462);
xnor_4 g05086(new_n5462, new_n5461, new_n5463);
xor_4  g05087(new_n5463, new_n5460, new_n5464);
xnor_4 g05088(new_n5464, new_n5459, new_n5465);
xnor_4 g05089(new_n5465, new_n5456, new_n5466);
nand_5 g05090(new_n5423, new_n5420, new_n5467);
not_8  g05091(new_n5467, new_n5468);
nand_5 g05092(new_n5422, new_n5421, new_n5469);
not_8  g05093(new_n5469, new_n5470);
and_8  g05094(new_n5434, new_n5424, new_n5471);
xor_4  g05095(new_n5471, new_n5470, new_n5472);
or_8   g05096(new_n5472, new_n5468, new_n5473);
and_8  g05097(new_n5473, new_n5466, new_n5474);
nor_6  g05098(new_n5473, new_n5466, new_n5475);
or_8   g05099(new_n5475, new_n5474, new_n5476);
and_8  g05100(new_n5476, new_n5447, new_n5477);
xor_4  g05101(new_n5473, new_n5466, new_n5478);
and_8  g05102(new_n5478, new_n5446, new_n5479);
or_8   g05103(new_n5479, new_n5477, new_n5480);
and_8  g05104(n5305, n2253, new_n5481);
not_8  g05105(new_n5481, new_n5482);
nor_6  g05106(new_n5445, new_n5435_1, new_n5483);
or_8   g05107(new_n5483, new_n5446, new_n5484);
or_8   g05108(new_n5484, new_n5482, new_n5485);
nand_5 g05109(new_n1078, new_n1071, new_n5486);
xor_4  g05110(new_n5443, new_n5442, new_n5487);
or_8   g05111(new_n5487, new_n5486, new_n5488);
xor_4  g05112(new_n5445, new_n5435_1, new_n5489);
and_8  g05113(new_n5489, new_n5481, new_n5490);
and_8  g05114(new_n5484, new_n5482, new_n5491);
or_8   g05115(new_n5491, new_n5490, new_n5492);
or_8   g05116(new_n5492, new_n5488, new_n5493);
and_8  g05117(new_n5493, new_n5485, new_n5494);
xor_4  g05118(new_n5494, new_n5480, new_n5495);
not_8  g05119(new_n5495, new_n5496);
not_8  g05120(new_n5488, new_n5497);
or_8   g05121(new_n5489, new_n5481, new_n5498);
and_8  g05122(new_n5498, new_n5485, new_n5499);
xor_4  g05123(new_n5499, new_n5497, new_n5500);
not_8  g05124(new_n5500, new_n5501);
nor_6  g05125(new_n1181, new_n1179, new_n5502);
and_8  g05126(n12145, n8759, new_n5503);
and_8  g05127(new_n1172, new_n1169, new_n5504);
and_8  g05128(new_n1178, new_n1173, new_n5505);
or_8   g05129(new_n5505, new_n5504, new_n5506);
xnor_4 g05130(new_n5506, new_n5503, new_n5507);
and_8  g05131(n6776, n2522, new_n5508);
or_8   g05132(new_n1176, new_n1175, new_n5509);
and_8  g05133(new_n1176, new_n1175, new_n5510);
or_8   g05134(new_n5510, new_n1174, new_n5511);
and_8  g05135(new_n5511, new_n5509, new_n5512);
xor_4  g05136(new_n5512, new_n5508, new_n5513);
and_8  g05137(n7436, n2024, new_n5514);
and_8  g05138(n12299, n9189, new_n5515);
and_8  g05139(n8276, n7946, new_n5516);
xnor_4 g05140(new_n5516, new_n5515, new_n5517);
xnor_4 g05141(new_n5517, new_n5514, new_n5518);
and_8  g05142(new_n5518, new_n5513, new_n5519);
nor_6  g05143(new_n5518, new_n5513, new_n5520);
or_8   g05144(new_n5520, new_n5519, new_n5521);
xor_4  g05145(new_n5521, new_n5507, new_n5522);
and_8  g05146(new_n5522, new_n5502, new_n5523);
not_8  g05147(new_n5523, new_n5524);
and_8  g05148(n12221, n8759, new_n5525);
not_8  g05149(new_n5525, new_n5526);
and_8  g05150(new_n5512, new_n5508, new_n5527);
or_8   g05151(new_n5519, new_n5527, new_n5528);
and_8  g05152(n12145, n6776, new_n5529);
and_8  g05153(n12299, n2522, new_n5530);
xor_4  g05154(new_n5530, new_n5529, new_n5531);
xor_4  g05155(new_n5531, new_n5528, new_n5532);
and_8  g05156(n9189, n7436, new_n5533);
or_8   g05157(new_n5517, new_n5514, new_n5534);
and_8  g05158(new_n5534, new_n5516, new_n5535);
nor_6  g05159(new_n5535, new_n5533, new_n5536);
or_8   g05160(new_n5535, new_n1174, new_n5537);
and_8  g05161(new_n5537, new_n5533, new_n5538);
or_8   g05162(new_n5538, new_n5536, new_n5539);
and_8  g05163(n8276, n2024, new_n5540);
and_8  g05164(n9241, n7946, new_n5541);
xnor_4 g05165(new_n5541, new_n5540, new_n5542);
xor_4  g05166(new_n5542, new_n5539, new_n5543);
and_8  g05167(new_n5543, new_n5532, new_n5544);
not_8  g05168(new_n5531, new_n5545);
xor_4  g05169(new_n5545, new_n5528, new_n5546);
not_8  g05170(new_n5543, new_n5547);
and_8  g05171(new_n5547, new_n5546, new_n5548);
or_8   g05172(new_n5548, new_n5544, new_n5549);
and_8  g05173(new_n5506, new_n5503, new_n5550);
nor_6  g05174(new_n5521, new_n5507, new_n5551);
or_8   g05175(new_n5551, new_n5550, new_n5552);
not_8  g05176(new_n5552, new_n5553);
or_8   g05177(new_n5553, new_n5549, new_n5554);
or_8   g05178(new_n5547, new_n5546, new_n5555);
or_8   g05179(new_n5543, new_n5532, new_n5556);
and_8  g05180(new_n5556, new_n5555, new_n5557);
or_8   g05181(new_n5552, new_n5557, new_n5558);
and_8  g05182(new_n5558, new_n5554, new_n5559);
xor_4  g05183(new_n5559, new_n5526, new_n5560);
or_8   g05184(new_n5560, new_n5524, new_n5561);
xor_4  g05185(new_n5559, new_n5525, new_n5562);
or_8   g05186(new_n5562, new_n5523, new_n5563);
and_8  g05187(new_n5563, new_n5561, new_n5564);
nor_6  g05188(new_n5522, new_n5502, new_n5565);
or_8   g05189(new_n5565, new_n5523, new_n5566);
not_8  g05190(new_n5566, new_n5567);
and_8  g05191(new_n1206, new_n1204, new_n5568);
not_8  g05192(new_n5568, new_n5569);
and_8  g05193(n6016, n5331, new_n5570);
and_8  g05194(n8476, n521, new_n5571);
or_8   g05195(new_n1197, new_n1196, new_n5572);
or_8   g05196(new_n1200, new_n1195, new_n5573);
and_8  g05197(new_n5573, new_n5572, new_n5574);
and_8  g05198(new_n5574, new_n5571, new_n5575);
not_8  g05199(new_n5571, new_n5576);
or_8   g05200(new_n1202, new_n1198_1, new_n5577);
and_8  g05201(new_n5577, new_n5576, new_n5578);
or_8   g05202(new_n5578, new_n5575, new_n5579_1);
and_8  g05203(n12648, n2498, new_n5580);
not_8  g05204(new_n5580, new_n5581);
and_8  g05205(n10545, n2558, new_n5582);
xor_4  g05206(new_n5582, new_n1142, new_n5583);
xor_4  g05207(new_n5583, new_n5581, new_n5584);
or_8   g05208(new_n5584, new_n5579_1, new_n5585);
or_8   g05209(new_n5577, new_n5576, new_n5586);
or_8   g05210(new_n5574, new_n5571, new_n5587);
and_8  g05211(new_n5587, new_n5586, new_n5588);
xor_4  g05212(new_n5583, new_n5580, new_n5589);
or_8   g05213(new_n5589, new_n5588, new_n5590);
and_8  g05214(new_n5590, new_n5585, new_n5591);
xor_4  g05215(new_n5591, new_n5570, new_n5592);
and_8  g05216(new_n1193, new_n1190, new_n5593);
and_8  g05217(new_n1203, new_n1194, new_n5594);
or_8   g05218(new_n5594, new_n5593, new_n5595);
and_8  g05219(new_n5595, new_n5592, new_n5596);
not_8  g05220(new_n5570, new_n5597);
xor_4  g05221(new_n5591, new_n5597, new_n5598);
not_8  g05222(new_n5595, new_n5599);
and_8  g05223(new_n5599, new_n5598, new_n5600);
or_8   g05224(new_n5600, new_n5596, new_n5601);
or_8   g05225(new_n5601, new_n5569, new_n5602);
or_8   g05226(new_n5599, new_n5598, new_n5603);
or_8   g05227(new_n5595, new_n5592, new_n5604);
and_8  g05228(new_n5604, new_n5603, new_n5605);
or_8   g05229(new_n5605, new_n5568, new_n5606);
and_8  g05230(new_n5606, new_n5602, new_n5607);
not_8  g05231(new_n1227, new_n5608);
and_8  g05232(n7965, n7270, new_n5609);
and_8  g05233(n7388, n806, new_n5610);
or_8   g05234(new_n1216, new_n1215, new_n5611);
or_8   g05235(new_n1219, new_n1214, new_n5612);
and_8  g05236(new_n5612, new_n5611, new_n5613);
and_8  g05237(new_n5613, new_n5610, new_n5614);
not_8  g05238(new_n5610, new_n5615);
or_8   g05239(new_n1221, new_n1217, new_n5616);
and_8  g05240(new_n5616, new_n5615, new_n5617);
or_8   g05241(new_n5617, new_n5614, new_n5618);
and_8  g05242(n9111, n2393, new_n5619);
not_8  g05243(new_n5619, new_n5620);
and_8  g05244(n9763, n5860, new_n5621);
xor_4  g05245(new_n5621, new_n1122, new_n5622);
xor_4  g05246(new_n5622, new_n5620, new_n5623);
or_8   g05247(new_n5623, new_n5618, new_n5624);
or_8   g05248(new_n5616, new_n5615, new_n5625);
or_8   g05249(new_n5613, new_n5610, new_n5626);
and_8  g05250(new_n5626, new_n5625, new_n5627);
xor_4  g05251(new_n5622, new_n5619, new_n5628);
or_8   g05252(new_n5628, new_n5627, new_n5629);
and_8  g05253(new_n5629, new_n5624, new_n5630);
xor_4  g05254(new_n5630, new_n5609, new_n5631);
and_8  g05255(new_n1212, new_n1208, new_n5632);
or_8   g05256(new_n1223, new_n5632, new_n5633);
and_8  g05257(new_n5633, new_n5631, new_n5634);
not_8  g05258(new_n5609, new_n5635);
xor_4  g05259(new_n5630, new_n5635, new_n5636);
not_8  g05260(new_n5633, new_n5637);
and_8  g05261(new_n5637, new_n5636, new_n5638);
or_8   g05262(new_n5638, new_n5634, new_n5639);
or_8   g05263(new_n5639, new_n5608, new_n5640);
or_8   g05264(new_n5637, new_n5636, new_n5641_1);
or_8   g05265(new_n5633, new_n5631, new_n5642);
and_8  g05266(new_n5642, new_n5641_1, new_n5643);
or_8   g05267(new_n5643, new_n1227, new_n5644);
and_8  g05268(new_n5644, new_n5640, new_n5645_1);
and_8  g05269(new_n5645_1, new_n5607, new_n5646);
and_8  g05270(new_n5605, new_n5568, new_n5647);
and_8  g05271(new_n5601, new_n5569, new_n5648);
or_8   g05272(new_n5648, new_n5647, new_n5649);
and_8  g05273(new_n5643, new_n1227, new_n5650);
and_8  g05274(new_n5639, new_n5608, new_n5651);
or_8   g05275(new_n5651, new_n5650, new_n5652);
and_8  g05276(new_n5652, new_n5649, new_n5653);
or_8   g05277(new_n5653, new_n5646, new_n5654);
not_8  g05278(new_n1229, new_n5655);
or_8   g05279(new_n5655, new_n1207, new_n5656);
or_8   g05280(new_n1234, new_n1230, new_n5657);
and_8  g05281(new_n5657, new_n5656, new_n5658);
and_8  g05282(new_n5658, new_n5654, new_n5659);
nor_6  g05283(new_n5658, new_n5654, new_n5660);
or_8   g05284(new_n5660, new_n5659, new_n5661);
and_8  g05285(new_n5661, new_n5567, new_n5662);
xor_4  g05286(new_n1186, new_n1182, new_n5663);
not_8  g05287(new_n1235, new_n5664);
and_8  g05288(new_n5664, new_n5663, new_n5665);
or_8   g05289(new_n5665, new_n1187, new_n5666);
xor_4  g05290(new_n5658, new_n5654, new_n5667);
or_8   g05291(new_n5667, new_n5566, new_n5668);
or_8   g05292(new_n5661, new_n5567, new_n5669);
and_8  g05293(new_n5669, new_n5668, new_n5670_1);
and_8  g05294(new_n5670_1, new_n5666, new_n5671);
or_8   g05295(new_n5671, new_n5662, new_n5672);
or_8   g05296(new_n5672, new_n5564, new_n5673);
and_8  g05297(new_n5562, new_n5523, new_n5674);
and_8  g05298(new_n5560, new_n5524, new_n5675);
or_8   g05299(new_n5675, new_n5674, new_n5676);
not_8  g05300(new_n1187, new_n5677);
or_8   g05301(new_n1235, new_n1189, new_n5678);
and_8  g05302(new_n5678, new_n5677, new_n5679);
and_8  g05303(new_n5667, new_n5566, new_n5680);
or_8   g05304(new_n5680, new_n5662, new_n5681);
or_8   g05305(new_n5681, new_n5679, new_n5682);
and_8  g05306(new_n5682, new_n5668, new_n5683);
or_8   g05307(new_n5683, new_n5676, new_n5684);
and_8  g05308(new_n5684, new_n5673, new_n5685);
and_8  g05309(n5798, n5331, new_n5686);
and_8  g05310(n12648, n5579, new_n5687);
and_8  g05311(n10545, n2498, new_n5688);
and_8  g05312(n7690, n2558, new_n5689);
xor_4  g05313(new_n5689, new_n5688, new_n5690);
xor_4  g05314(new_n5690, new_n5687, new_n5691);
or_8   g05315(new_n5582, new_n1142, new_n5692);
and_8  g05316(new_n5582, new_n1142, new_n5693_1);
or_8   g05317(new_n5693_1, new_n5580, new_n5694_1);
and_8  g05318(new_n5694_1, new_n5692, new_n5695);
and_8  g05319(new_n5695, new_n5691, new_n5696);
nor_6  g05320(new_n5695, new_n5691, new_n5697);
or_8   g05321(new_n5697, new_n5696, new_n5698);
and_8  g05322(n8476, n6016, new_n5699);
and_8  g05323(n2530, n521, new_n5700);
xor_4  g05324(new_n5700, new_n5699, new_n5701);
not_8  g05325(new_n5701, new_n5702);
or_8   g05326(new_n5702, new_n5698, new_n5703);
xor_4  g05327(new_n5695, new_n5691, new_n5704);
or_8   g05328(new_n5701, new_n5704, new_n5705);
and_8  g05329(new_n5705, new_n5703, new_n5706);
and_8  g05330(new_n5589, new_n5588, new_n5707);
or_8   g05331(new_n5707, new_n5575, new_n5708);
and_8  g05332(new_n5708, new_n5706, new_n5709);
nor_6  g05333(new_n5708, new_n5706, new_n5710);
or_8   g05334(new_n5710, new_n5709, new_n5711);
and_8  g05335(new_n5591, new_n5570, new_n5712);
nor_6  g05336(new_n5596, new_n5712, new_n5713);
xor_4  g05337(new_n5713, new_n5711, new_n5714);
and_8  g05338(new_n5714, new_n5686, new_n5715);
not_8  g05339(new_n5686, new_n5716);
or_8   g05340(new_n5596, new_n5712, new_n5717);
xor_4  g05341(new_n5717, new_n5711, new_n5718);
and_8  g05342(new_n5718, new_n5716, new_n5719);
or_8   g05343(new_n5719, new_n5715, new_n5720);
xor_4  g05344(new_n5720, new_n5647, new_n5721);
and_8  g05345(n7965, n5153, new_n5722);
and_8  g05346(n3342, n2393, new_n5723);
and_8  g05347(n9763, n3986, new_n5724);
and_8  g05348(n9111, n5860, new_n5725);
xor_4  g05349(new_n5725, new_n5724, new_n5726);
and_8  g05350(new_n5726, new_n5723, new_n5727);
nor_6  g05351(new_n5726, new_n5723, new_n5728);
or_8   g05352(new_n5728, new_n5727, new_n5729);
or_8   g05353(new_n5621, new_n1122, new_n5730);
and_8  g05354(new_n5621, new_n1122, new_n5731);
or_8   g05355(new_n5731, new_n5619, new_n5732);
and_8  g05356(new_n5732, new_n5730, new_n5733);
xor_4  g05357(new_n5733, new_n5729, new_n5734);
and_8  g05358(n7388, n7270, new_n5735);
and_8  g05359(n11892, n806, new_n5736);
xor_4  g05360(new_n5736, new_n5735, new_n5737);
not_8  g05361(new_n5737, new_n5738);
or_8   g05362(new_n5738, new_n5734, new_n5739);
xor_4  g05363(new_n5726, new_n5723, new_n5740);
xor_4  g05364(new_n5733, new_n5740, new_n5741);
or_8   g05365(new_n5737, new_n5741, new_n5742);
and_8  g05366(new_n5742, new_n5739, new_n5743);
and_8  g05367(new_n5628, new_n5627, new_n5744);
or_8   g05368(new_n5744, new_n5614, new_n5745);
and_8  g05369(new_n5745, new_n5743, new_n5746);
nor_6  g05370(new_n5745, new_n5743, new_n5747);
or_8   g05371(new_n5747, new_n5746, new_n5748);
and_8  g05372(new_n5630, new_n5609, new_n5749);
nor_6  g05373(new_n5634, new_n5749, new_n5750);
xor_4  g05374(new_n5750, new_n5748, new_n5751);
and_8  g05375(new_n5751, new_n5722, new_n5752);
not_8  g05376(new_n5722, new_n5753);
nor_6  g05377(new_n5750, new_n5748, new_n5754);
and_8  g05378(new_n5750, new_n5748, new_n5755);
or_8   g05379(new_n5755, new_n5754, new_n5756);
and_8  g05380(new_n5756, new_n5753, new_n5757);
or_8   g05381(new_n5757, new_n5752, new_n5758);
xor_4  g05382(new_n5758, new_n5650, new_n5759);
or_8   g05383(new_n5759, new_n5721, new_n5760_1);
xor_4  g05384(new_n5720, new_n5602, new_n5761);
xor_4  g05385(new_n5758, new_n5640, new_n5762);
or_8   g05386(new_n5762, new_n5761, new_n5763);
and_8  g05387(new_n5763, new_n5760_1, new_n5764);
or_8   g05388(new_n5660, new_n5653, new_n5765);
or_8   g05389(new_n5765, new_n5764, new_n5766);
and_8  g05390(new_n5762, new_n5761, new_n5767_1);
and_8  g05391(new_n5759, new_n5721, new_n5768);
or_8   g05392(new_n5768, new_n5767_1, new_n5769);
not_8  g05393(new_n5765, new_n5770);
or_8   g05394(new_n5770, new_n5769, new_n5771);
and_8  g05395(new_n5771, new_n5766, new_n5772);
xor_4  g05396(new_n5772, new_n5685, new_n5773);
and_8  g05397(new_n5773, new_n5501, new_n5774);
and_8  g05398(new_n5683, new_n5676, new_n5775);
and_8  g05399(new_n5672, new_n5564, new_n5776);
or_8   g05400(new_n5776, new_n5775, new_n5777);
xor_4  g05401(new_n5772, new_n5777, new_n5778);
or_8   g05402(new_n5778, new_n5500, new_n5779);
or_8   g05403(new_n5773, new_n5501, new_n5780);
and_8  g05404(new_n5780, new_n5779, new_n5781);
xor_4  g05405(new_n5487, new_n5486, new_n5782);
xor_4  g05406(new_n5670_1, new_n5666, new_n5783);
nor_6  g05407(new_n5783, new_n5782, new_n5784);
nor_6  g05408(new_n1237, new_n1168, new_n5785);
or_8   g05409(new_n5785, new_n1166, new_n5786);
and_8  g05410(new_n5783, new_n5782, new_n5787);
or_8   g05411(new_n5787, new_n5784, new_n5788);
nor_6  g05412(new_n5788, new_n5786, new_n5789);
or_8   g05413(new_n5789, new_n5784, new_n5790);
and_8  g05414(new_n5790, new_n5781, new_n5791);
or_8   g05415(new_n5791, new_n5774, new_n5792);
or_8   g05416(new_n5792, new_n5496, new_n5793);
and_8  g05417(new_n5778, new_n5500, new_n5794);
or_8   g05418(new_n5794, new_n5774, new_n5795);
not_8  g05419(new_n5784, new_n5796);
or_8   g05420(new_n5788, new_n5786, new_n5797);
and_8  g05421(new_n5797, new_n5796, new_n5798_1);
or_8   g05422(new_n5798_1, new_n5795, new_n5799);
and_8  g05423(new_n5799, new_n5779, new_n5800);
or_8   g05424(new_n5800, new_n5495, new_n5801);
and_8  g05425(new_n5801, new_n5793, new_n5802);
xor_4  g05426(new_n5553, new_n5557, new_n5803);
or_8   g05427(new_n5803, new_n5526, new_n5804);
and_8  g05428(new_n5561, new_n5804, new_n5805);
not_8  g05429(new_n5554, new_n5806);
not_8  g05430(new_n5538, new_n5807);
or_8   g05431(new_n5542, new_n5539, new_n5808);
and_8  g05432(new_n5808, new_n5807, new_n5809);
and_8  g05433(n12221, n6776, new_n5810);
and_8  g05434(n12299, n12145, new_n5811);
and_8  g05435(n10217, n8759, new_n5812);
xnor_4 g05436(new_n5812, new_n5811, new_n5813);
xor_4  g05437(new_n5813, new_n5810, new_n5814_1);
xnor_4 g05438(new_n5814_1, new_n5809, new_n5815);
and_8  g05439(new_n5541, new_n5540, new_n5816);
and_8  g05440(n7436, n2522, new_n5817);
xnor_4 g05441(new_n5817, new_n5816, new_n5818);
and_8  g05442(n9241, n2024, new_n5819);
and_8  g05443(n10510, n7946, new_n5820);
and_8  g05444(n9189, n8276, new_n5821);
xnor_4 g05445(new_n5821, new_n5820, new_n5822);
xor_4  g05446(new_n5822, new_n5819, new_n5823);
xor_4  g05447(new_n5823, new_n5818, new_n5824);
nor_6  g05448(new_n5824, new_n5815, new_n5825);
and_8  g05449(new_n5824, new_n5815, new_n5826);
or_8   g05450(new_n5826, new_n5825, new_n5827);
not_8  g05451(new_n5827, new_n5828);
nand_5 g05452(new_n5531, new_n5528, new_n5829);
nand_5 g05453(new_n5530, new_n5529, new_n5830);
nor_6  g05454(new_n5555, new_n5830, new_n5831);
and_8  g05455(new_n5555, new_n5830, new_n5832);
or_8   g05456(new_n5832, new_n5831, new_n5833);
and_8  g05457(new_n5833, new_n5829, new_n5834);
xor_4  g05458(new_n5834, new_n5828, new_n5835);
or_8   g05459(new_n5835, new_n5806, new_n5836);
xor_4  g05460(new_n5834, new_n5827, new_n5837);
or_8   g05461(new_n5837, new_n5554, new_n5838);
and_8  g05462(new_n5838, new_n5836, new_n5839);
xor_4  g05463(new_n5839, new_n5805, new_n5840);
or_8   g05464(new_n5772, new_n5777, new_n5841);
and_8  g05465(new_n5841, new_n5684, new_n5842);
and_8  g05466(new_n5842, new_n5840, new_n5843);
nor_6  g05467(new_n5842, new_n5840, new_n5844);
or_8   g05468(new_n5844, new_n5843, new_n5845);
or_8   g05469(new_n5713, new_n5711, new_n5846);
and_8  g05470(n8476, n5798, new_n5847);
and_8  g05471(n6016, n2530, new_n5848);
and_8  g05472(n5331, n2347, new_n5849);
xnor_4 g05473(new_n5849, new_n5848, new_n5850);
xor_4  g05474(new_n5850, new_n5847, new_n5851);
and_8  g05475(new_n5690, new_n5687, new_n5852);
or_8   g05476(new_n5696, new_n5852, new_n5853);
xor_4  g05477(new_n5853, new_n5851, new_n5854);
and_8  g05478(new_n5689, new_n5688, new_n5855);
and_8  g05479(n12648, n521, new_n5856);
xnor_4 g05480(new_n5856, new_n5855, new_n5857_1);
and_8  g05481(n7690, n2498, new_n5858);
and_8  g05482(n10545, n5579, new_n5859);
and_8  g05483(n3616, n2558, new_n5860_1);
xnor_4 g05484(new_n5860_1, new_n5859, new_n5861);
xor_4  g05485(new_n5861, new_n5858, new_n5862);
xor_4  g05486(new_n5862, new_n5857_1, new_n5863);
or_8   g05487(new_n5863, new_n5854, new_n5864);
not_8  g05488(new_n5864, new_n5865);
and_8  g05489(new_n5863, new_n5854, new_n5866);
or_8   g05490(new_n5866, new_n5865, new_n5867);
not_8  g05491(new_n5703, new_n5868);
and_8  g05492(new_n5700, new_n5699, new_n5869);
xor_4  g05493(new_n5709, new_n5869, new_n5870);
or_8   g05494(new_n5870, new_n5868, new_n5871);
xor_4  g05495(new_n5871, new_n5867, new_n5872);
xor_4  g05496(new_n5872, new_n5846, new_n5873);
not_8  g05497(new_n5715, new_n5874);
or_8   g05498(new_n5720, new_n5602, new_n5875);
and_8  g05499(new_n5875, new_n5874, new_n5876);
xor_4  g05500(new_n5876, new_n5873, new_n5877);
and_8  g05501(new_n5733, new_n5740, new_n5878);
nor_6  g05502(new_n5878, new_n5727, new_n5879);
and_8  g05503(n7388, n5153, new_n5880);
and_8  g05504(n11892, n7270, new_n5881);
and_8  g05505(n7965, n2507, new_n5882);
xnor_4 g05506(new_n5882, new_n5881, new_n5883);
xor_4  g05507(new_n5883, new_n5880, new_n5884);
xor_4  g05508(new_n5884, new_n5879, new_n5885);
and_8  g05509(new_n5725, new_n5724, new_n5886);
and_8  g05510(n2393, n806, new_n5887);
xnor_4 g05511(new_n5887, new_n5886, new_n5888);
and_8  g05512(n9111, n3986, new_n5889);
and_8  g05513(n5860, n3342, new_n5890);
and_8  g05514(n9763, n5857, new_n5891);
xnor_4 g05515(new_n5891, new_n5890, new_n5892);
xor_4  g05516(new_n5892, new_n5889, new_n5893);
xor_4  g05517(new_n5893, new_n5888, new_n5894);
xor_4  g05518(new_n5894, new_n5885, new_n5895);
not_8  g05519(new_n5739, new_n5896);
and_8  g05520(new_n5736, new_n5735, new_n5897);
xor_4  g05521(new_n5746, new_n5897, new_n5898);
or_8   g05522(new_n5898, new_n5896, new_n5899);
xor_4  g05523(new_n5899, new_n5895, new_n5900);
xor_4  g05524(new_n5900, new_n5754, new_n5901);
not_8  g05525(new_n5757, new_n5902);
or_8   g05526(new_n5758, new_n5650, new_n5903);
and_8  g05527(new_n5903, new_n5902, new_n5904);
xor_4  g05528(new_n5904, new_n5901, new_n5905);
and_8  g05529(new_n5905, new_n5877, new_n5906);
and_8  g05530(new_n5876, new_n5873, new_n5907);
nor_6  g05531(new_n5876, new_n5873, new_n5908);
or_8   g05532(new_n5908, new_n5907, new_n5909);
nor_6  g05533(new_n5904, new_n5901, new_n5910);
and_8  g05534(new_n5904, new_n5901, new_n5911);
or_8   g05535(new_n5911, new_n5910, new_n5912);
and_8  g05536(new_n5912, new_n5909, new_n5913);
or_8   g05537(new_n5913, new_n5906, new_n5914);
and_8  g05538(new_n5771, new_n5763, new_n5915);
nor_6  g05539(new_n5915, new_n5914, new_n5916);
and_8  g05540(new_n5915, new_n5914, new_n5917);
or_8   g05541(new_n5917, new_n5916, new_n5918);
xor_4  g05542(new_n5918, new_n5845, new_n5919);
and_8  g05543(new_n5919, new_n5802, new_n5920);
nor_6  g05544(new_n5919, new_n5802, new_n5921);
or_8   g05545(new_n5921, new_n5920, n1523);
and_8  g05546(n6687, n4634, new_n5923);
and_8  g05547(n10223, n4189, new_n5924);
and_8  g05548(new_n5924, new_n4442, new_n5925);
and_8  g05549(n10223, n6687, new_n5926);
and_8  g05550(n7265, n4189, new_n5927);
or_8   g05551(new_n5927, new_n5926, new_n5928);
and_8  g05552(n2879, n2564, new_n5929);
and_8  g05553(new_n5929, new_n5928, new_n5930);
or_8   g05554(new_n5930, new_n5925, new_n5931);
xor_4  g05555(new_n5931, new_n5923, new_n5932);
and_8  g05556(n4189, n2879, new_n5933);
and_8  g05557(n10223, n2564, new_n5934_1);
and_8  g05558(n7265, n6770, new_n5935);
xnor_4 g05559(new_n5935, new_n5934_1, new_n5936);
xnor_4 g05560(new_n5936, new_n5933, new_n5937);
xnor_4 g05561(new_n5937, new_n5932, new_n5938);
not_8  g05562(new_n5928, new_n5939);
or_8   g05563(new_n5939, new_n5925, new_n5940);
and_8  g05564(n7265, n2564, new_n5941);
and_8  g05565(n6687, n2879, new_n5942);
and_8  g05566(new_n5942, new_n5941, new_n5943);
nand_5 g05567(new_n5943, new_n5940, new_n5944);
nor_6  g05568(new_n5944, new_n5938, new_n5945);
and_8  g05569(n9195, n6687, new_n5946);
and_8  g05570(n4634, n2564, new_n5947);
and_8  g05571(n6770, n2879, new_n5948);
and_8  g05572(n9920, n7265, new_n5949);
xor_4  g05573(new_n5949, new_n5924, new_n5950);
xor_4  g05574(new_n5950, new_n5948, new_n5951);
xor_4  g05575(new_n5951, new_n5947, new_n5952);
or_8   g05576(new_n5935, new_n5934_1, new_n5953);
or_8   g05577(new_n5936, new_n5933, new_n5954);
and_8  g05578(new_n5954, new_n5953, new_n5955);
xor_4  g05579(new_n5955, new_n5952, new_n5956);
xor_4  g05580(new_n5956, new_n5946, new_n5957);
and_8  g05581(new_n5931, new_n5923, new_n5958);
and_8  g05582(new_n5937, new_n5932, new_n5959);
or_8   g05583(new_n5959, new_n5958, new_n5960);
xor_4  g05584(new_n5960, new_n5957, new_n5961);
xor_4  g05585(new_n5961, new_n5945, new_n5962);
not_8  g05586(new_n5962, new_n5963);
and_8  g05587(n8336, n2522, new_n5964_1);
and_8  g05588(n9189, n8336, new_n5965);
and_8  g05589(n7946, n6986, new_n5966);
or_8   g05590(new_n5966, new_n5965, new_n5967);
and_8  g05591(n9189, n6986, new_n5968);
and_8  g05592(new_n5968, new_n4443, new_n5969);
and_8  g05593(n10928, n2024, new_n5970);
or_8   g05594(new_n5970, new_n5969, new_n5971);
and_8  g05595(new_n5971, new_n5967, new_n5972);
xor_4  g05596(new_n5972, new_n5964_1, new_n5973);
and_8  g05597(n6986, n2024, new_n5974);
and_8  g05598(n10928, n9189, new_n5975);
and_8  g05599(n7946, n2226, new_n5976);
xor_4  g05600(new_n5976, new_n5975, new_n5977);
xor_4  g05601(new_n5977, new_n5974, new_n5978);
xnor_4 g05602(new_n5978, new_n5973, new_n5979);
not_8  g05603(new_n5970, new_n5980);
or_8   g05604(new_n5980, new_n4443, new_n5981);
not_8  g05605(new_n5967, new_n5982);
or_8   g05606(new_n5969, new_n5982, new_n5983);
and_8  g05607(new_n5983, new_n5981, new_n5984);
not_8  g05608(new_n5984, new_n5985);
or_8   g05609(new_n5985, new_n5980, new_n5986);
nor_6  g05610(new_n5986, new_n5979, new_n5987);
nand_5 g05611(n12145, n8336, new_n5988);
and_8  g05612(n10928, n2522, new_n5989);
or_8   g05613(new_n5976, new_n5975, new_n5990);
and_8  g05614(new_n5976, new_n5975, new_n5991);
or_8   g05615(new_n5991, new_n5974, new_n5992);
and_8  g05616(new_n5992, new_n5990, new_n5993);
xor_4  g05617(new_n5993, new_n5989, new_n5994);
and_8  g05618(n2226, n2024, new_n5995);
and_8  g05619(n7946, n1094, new_n5996);
xor_4  g05620(new_n5996, new_n5968, new_n5997);
xor_4  g05621(new_n5997, new_n5995, new_n5998);
and_8  g05622(new_n5998, new_n5994, new_n5999);
nor_6  g05623(new_n5998, new_n5994, new_n6000);
or_8   g05624(new_n6000, new_n5999, new_n6001);
xor_4  g05625(new_n6001, new_n5988, new_n6002);
and_8  g05626(new_n5972, new_n5964_1, new_n6003);
and_8  g05627(new_n5978, new_n5973, new_n6004);
or_8   g05628(new_n6004, new_n6003, new_n6005);
xor_4  g05629(new_n6005, new_n6002, new_n6006);
xor_4  g05630(new_n6006, new_n5987, new_n6007);
xor_4  g05631(new_n5986, new_n5979, new_n6008);
and_8  g05632(n12069, n521, new_n6009);
and_8  g05633(n7891, n5579, new_n6010);
and_8  g05634(new_n6010, new_n4445, new_n6011);
and_8  g05635(n12069, n5579, new_n6012);
and_8  g05636(n7891, n2558, new_n6013);
or_8   g05637(new_n6013, new_n6012, new_n6014);
and_8  g05638(n12391, n2498, new_n6015);
and_8  g05639(new_n6015, new_n6014, new_n6016_1);
or_8   g05640(new_n6016_1, new_n6011, new_n6017);
xor_4  g05641(new_n6017, new_n6009, new_n6018);
and_8  g05642(n7891, n2498, new_n6019);
and_8  g05643(n12391, n5579, new_n6020);
and_8  g05644(n7160, n2558, new_n6021);
xor_4  g05645(new_n6021, new_n6020, new_n6022);
xor_4  g05646(new_n6022, new_n6019, new_n6023);
and_8  g05647(new_n6023, new_n6018, new_n6024);
nor_6  g05648(new_n6023, new_n6018, new_n6025);
or_8   g05649(new_n6025, new_n6024, new_n6026);
nor_6  g05650(new_n6013, new_n6012, new_n6027);
or_8   g05651(new_n6027, new_n6011, new_n6028);
and_8  g05652(n12391, n2558, new_n6029);
and_8  g05653(n12069, n2498, new_n6030);
and_8  g05654(new_n6030, new_n6029, new_n6031);
nand_5 g05655(new_n6031, new_n6028, new_n6032);
and_8  g05656(new_n6032, new_n6026, new_n6033);
nor_6  g05657(new_n6032, new_n6026, new_n6034);
or_8   g05658(new_n6034, new_n6033, new_n6035);
and_8  g05659(n11222, n806, new_n6036);
and_8  g05660(n11222, n3342, new_n6037);
and_8  g05661(n9763, n5314, new_n6038_1);
or_8   g05662(new_n6038_1, new_n6037, new_n6039);
and_8  g05663(n5314, n3342, new_n6040);
and_8  g05664(new_n6040, new_n4444, new_n6041);
and_8  g05665(n11153, n9111, new_n6042);
or_8   g05666(new_n6042, new_n6041, new_n6043);
and_8  g05667(new_n6043, new_n6039, new_n6044);
xor_4  g05668(new_n6044, new_n6036, new_n6045);
and_8  g05669(n9111, n5314, new_n6046);
and_8  g05670(n11153, n3342, new_n6047);
and_8  g05671(n9763, n996, new_n6048);
xor_4  g05672(new_n6048, new_n6047, new_n6049);
xor_4  g05673(new_n6049, new_n6046, new_n6050);
and_8  g05674(new_n6050, new_n6045, new_n6051);
nor_6  g05675(new_n6050, new_n6045, new_n6052);
or_8   g05676(new_n6052, new_n6051, new_n6053);
not_8  g05677(new_n6042, new_n6054);
not_8  g05678(new_n4444, new_n6055);
and_8  g05679(new_n6042, new_n6055, new_n6056);
nor_6  g05680(new_n6056, new_n6039, new_n6057);
nor_6  g05681(new_n6057, new_n6041, new_n6058);
or_8   g05682(new_n6058, new_n6054, new_n6059);
xor_4  g05683(new_n6059, new_n6053, new_n6060);
xor_4  g05684(new_n6060, new_n6035, new_n6061);
nand_5 g05685(new_n6056, new_n6039, new_n6062);
and_8  g05686(new_n6062, new_n6058, new_n6063);
and_8  g05687(new_n4445, new_n4444, new_n6064);
xor_4  g05688(new_n6030, new_n6029, new_n6065);
or_8   g05689(new_n6065, new_n6064, new_n6066);
xor_4  g05690(new_n6065, new_n6064, new_n6067);
not_8  g05691(new_n6067, new_n6068);
and_8  g05692(n11153, n9763, new_n6069);
and_8  g05693(n11222, n9111, new_n6070);
xor_4  g05694(new_n6070, new_n6069, new_n6071);
or_8   g05695(new_n6071, new_n6068, new_n6072);
and_8  g05696(new_n6072, new_n6066, new_n6073);
nor_6  g05697(new_n6073, new_n6063, new_n6074);
not_8  g05698(new_n6074, new_n6075);
and_8  g05699(new_n6073, new_n6063, new_n6076);
or_8   g05700(new_n6076, new_n6074, new_n6077);
not_8  g05701(new_n4445, new_n6078);
nand_5 g05702(new_n6015, new_n6078, new_n6079);
and_8  g05703(new_n6079, new_n6028, new_n6080);
nor_6  g05704(new_n6079, new_n6027, new_n6081);
or_8   g05705(new_n6081, new_n6080, new_n6082);
not_8  g05706(new_n6082, new_n6083);
or_8   g05707(new_n6083, new_n6077, new_n6084);
and_8  g05708(new_n6084, new_n6075, new_n6085);
and_8  g05709(new_n6085, new_n6061, new_n6086);
nor_6  g05710(new_n6059, new_n6053, new_n6087);
and_8  g05711(new_n6059, new_n6053, new_n6088);
or_8   g05712(new_n6088, new_n6087, new_n6089_1);
xor_4  g05713(new_n6089_1, new_n6035, new_n6090);
xor_4  g05714(new_n6073, new_n6063, new_n6091);
and_8  g05715(new_n6082, new_n6091, new_n6092);
or_8   g05716(new_n6092, new_n6074, new_n6093);
and_8  g05717(new_n6093, new_n6090, new_n6094);
or_8   g05718(new_n6094, new_n6086, new_n6095);
and_8  g05719(new_n6095, new_n6008, new_n6096);
xor_4  g05720(new_n6095, new_n6008, new_n6097);
or_8   g05721(new_n5981, new_n5982, new_n6098);
nand_5 g05722(new_n6098, new_n5985, new_n6099);
or_8   g05723(new_n6082, new_n6091, new_n6100);
and_8  g05724(new_n6100, new_n6084, new_n6101);
nor_6  g05725(new_n6101, new_n6099, new_n6102);
xor_4  g05726(new_n6101, new_n6099, new_n6103);
xor_4  g05727(new_n6071, new_n6067, new_n6104);
and_8  g05728(n10928, n7946, new_n6105);
and_8  g05729(n8336, n2024, new_n6106);
xor_4  g05730(new_n6106, new_n6105, new_n6107);
and_8  g05731(new_n6107, new_n6104, new_n6108);
and_8  g05732(new_n4446, new_n4443, new_n6109);
xor_4  g05733(new_n6107, new_n6104, new_n6110);
and_8  g05734(new_n6110, new_n6109, new_n6111);
or_8   g05735(new_n6111, new_n6108, new_n6112);
and_8  g05736(new_n6112, new_n6103, new_n6113);
or_8   g05737(new_n6113, new_n6102, new_n6114);
and_8  g05738(new_n6114, new_n6097, new_n6115);
or_8   g05739(new_n6115, new_n6096, new_n6116);
and_8  g05740(new_n6116, new_n6007, new_n6117);
not_8  g05741(new_n6007, new_n6118);
not_8  g05742(new_n6096, new_n6119);
nor_6  g05743(new_n6095, new_n6008, new_n6120);
or_8   g05744(new_n6120, new_n6096, new_n6121);
not_8  g05745(new_n6102, new_n6122);
and_8  g05746(new_n6101, new_n6099, new_n6123);
or_8   g05747(new_n6123, new_n6102, new_n6124);
not_8  g05748(new_n6112, new_n6125);
or_8   g05749(new_n6125, new_n6124, new_n6126_1);
and_8  g05750(new_n6126_1, new_n6122, new_n6127);
or_8   g05751(new_n6127, new_n6121, new_n6128);
and_8  g05752(new_n6128, new_n6119, new_n6129);
and_8  g05753(new_n6129, new_n6118, new_n6130);
or_8   g05754(new_n6130, new_n6117, new_n6131);
not_8  g05755(n6016, new_n6132);
or_8   g05756(new_n4398, new_n6132, new_n6133);
and_8  g05757(n12391, n521, new_n6134);
or_8   g05758(new_n6021, new_n6020, new_n6135);
and_8  g05759(new_n6021, new_n6020, new_n6136);
or_8   g05760(new_n6136, new_n6019, new_n6137);
and_8  g05761(new_n6137, new_n6135, new_n6138);
and_8  g05762(new_n6138, new_n6134, new_n6139);
nor_6  g05763(new_n6138, new_n6134, new_n6140);
or_8   g05764(new_n6140, new_n6139, new_n6141);
and_8  g05765(n7160, n2498, new_n6142);
and_8  g05766(n4828, n2558, new_n6143);
nor_6  g05767(new_n6143, new_n6010, new_n6144);
and_8  g05768(new_n6143, new_n6010, new_n6145);
or_8   g05769(new_n6145, new_n6144, new_n6146);
and_8  g05770(new_n6146, new_n6142, new_n6147);
nor_6  g05771(new_n6146, new_n6142, new_n6148);
or_8   g05772(new_n6148, new_n6147, new_n6149);
xor_4  g05773(new_n6149, new_n6141, new_n6150);
xor_4  g05774(new_n6150, new_n6133, new_n6151);
and_8  g05775(new_n6017, new_n6009, new_n6152);
or_8   g05776(new_n6024, new_n6152, new_n6153);
xor_4  g05777(new_n6153, new_n6151, new_n6154);
xor_4  g05778(new_n6154, new_n6034, new_n6155);
nand_5 g05779(n11222, n7270, new_n6156);
and_8  g05780(n11153, n806, new_n6157);
or_8   g05781(new_n6048, new_n6047, new_n6158);
and_8  g05782(new_n6048, new_n6047, new_n6159);
or_8   g05783(new_n6159, new_n6046, new_n6160);
and_8  g05784(new_n6160, new_n6158, new_n6161);
and_8  g05785(new_n6161, new_n6157, new_n6162);
nor_6  g05786(new_n6161, new_n6157, new_n6163);
or_8   g05787(new_n6163, new_n6162, new_n6164);
and_8  g05788(n9111, n996, new_n6165);
and_8  g05789(n9763, n5767, new_n6166);
xor_4  g05790(new_n6166, new_n6040, new_n6167);
xor_4  g05791(new_n6167, new_n6165, new_n6168);
xor_4  g05792(new_n6168, new_n6164, new_n6169);
nor_6  g05793(new_n6169, new_n6156, new_n6170);
and_8  g05794(new_n6169, new_n6156, new_n6171);
or_8   g05795(new_n6171, new_n6170, new_n6172);
and_8  g05796(new_n6044, new_n6036, new_n6173);
or_8   g05797(new_n6051, new_n6173, new_n6174);
not_8  g05798(new_n6174, new_n6175);
xor_4  g05799(new_n6175, new_n6172, new_n6176);
xor_4  g05800(new_n6176, new_n6087, new_n6177);
and_8  g05801(new_n6177, new_n6155, new_n6178);
nor_6  g05802(new_n6177, new_n6155, new_n6179);
or_8   g05803(new_n6179, new_n6178, new_n6180);
nand_5 g05804(new_n6089_1, new_n6035, new_n6181);
or_8   g05805(new_n6085, new_n6061, new_n6182);
and_8  g05806(new_n6182, new_n6181, new_n6183);
xor_4  g05807(new_n6183, new_n6180, new_n6184);
and_8  g05808(new_n6184, new_n6131, new_n6185);
or_8   g05809(new_n6129, new_n6118, new_n6186);
or_8   g05810(new_n6116, new_n6007, new_n6187);
and_8  g05811(new_n6187, new_n6186, new_n6188);
nor_6  g05812(new_n6183, new_n6180, new_n6189);
and_8  g05813(new_n6183, new_n6180, new_n6190);
or_8   g05814(new_n6190, new_n6189, new_n6191);
and_8  g05815(new_n6191, new_n6188, new_n6192_1);
or_8   g05816(new_n6192_1, new_n6185, new_n6193);
and_8  g05817(new_n6193, new_n5963, new_n6194);
or_8   g05818(new_n6191, new_n6188, new_n6195);
or_8   g05819(new_n6184, new_n6131, new_n6196);
and_8  g05820(new_n6196, new_n6195, new_n6197);
and_8  g05821(new_n6197, new_n5962, new_n6198);
or_8   g05822(new_n6198, new_n6194, new_n6199);
xor_4  g05823(new_n5944, new_n5938, new_n6200);
xor_4  g05824(new_n6127, new_n6121, new_n6201);
nor_6  g05825(new_n6201, new_n6200, new_n6202);
not_8  g05826(new_n6202, new_n6203);
xor_4  g05827(new_n6125, new_n6124, new_n6204);
not_8  g05828(new_n4442, new_n6205);
and_8  g05829(new_n5929, new_n6205, new_n6206);
not_8  g05830(new_n6206, new_n6207);
nand_5 g05831(new_n6207, new_n5940, new_n6208);
or_8   g05832(new_n6207, new_n5939, new_n6209);
nand_5 g05833(new_n6209, new_n6208, new_n6210);
not_8  g05834(new_n6210, new_n6211);
or_8   g05835(new_n6211, new_n6204, new_n6212);
xor_4  g05836(new_n6210, new_n6204, new_n6213);
and_8  g05837(new_n4447, new_n4442, new_n6214);
xor_4  g05838(new_n5942, new_n5941, new_n6215);
or_8   g05839(new_n6215, new_n6214, new_n6216);
xor_4  g05840(new_n6110, new_n6109, new_n6217);
xnor_4 g05841(new_n6215, new_n6214, new_n6218);
or_8   g05842(new_n6218, new_n6217, new_n6219);
and_8  g05843(new_n6219, new_n6216, new_n6220);
or_8   g05844(new_n6220, new_n6213, new_n6221);
and_8  g05845(new_n6221, new_n6212, new_n6222);
and_8  g05846(new_n6201, new_n6200, new_n6223);
or_8   g05847(new_n6223, new_n6202, new_n6224);
or_8   g05848(new_n6224, new_n6222, new_n6225);
and_8  g05849(new_n6225, new_n6203, new_n6226);
xnor_4 g05850(new_n6226, new_n6199, n1658);
and_8  g05851(n7862, n4634, new_n6228);
and_8  g05852(n10223, n7862, new_n6229);
and_8  g05853(n7265, n3172, new_n6230);
or_8   g05854(new_n6230, new_n6229, new_n6231);
nand_5 g05855(n7862, n7265, new_n6232);
not_8  g05856(new_n6232, new_n6233);
and_8  g05857(n10223, n3172, new_n6234);
and_8  g05858(new_n6234, new_n6233, new_n6235);
and_8  g05859(n2879, n1333, new_n6236);
or_8   g05860(new_n6236, new_n6235, new_n6237);
and_8  g05861(new_n6237, new_n6231, new_n6238);
xor_4  g05862(new_n6238, new_n6228, new_n6239);
and_8  g05863(n3172, n2879, new_n6240);
and_8  g05864(n10223, n1333, new_n6241);
and_8  g05865(n11757, n7265, new_n6242);
xor_4  g05866(new_n6242, new_n6241, new_n6243);
xor_4  g05867(new_n6243, new_n6240, new_n6244);
xor_4  g05868(new_n6244, new_n6239, new_n6245);
and_8  g05869(new_n6236, new_n6232, new_n6246);
nor_6  g05870(new_n6246, new_n6231, new_n6247);
or_8   g05871(new_n6247, new_n6235, new_n6248);
and_8  g05872(new_n6248, new_n6236, new_n6249);
xor_4  g05873(new_n6249, new_n6245, new_n6250);
nand_5 g05874(n6877, n2522, new_n6251);
not_8  g05875(new_n6251, new_n6252);
nand_5 g05876(n2464, n2024, new_n6253);
and_8  g05877(n9400, n9189, new_n6254_1);
and_8  g05878(n11311, n7946, new_n6255);
xnor_4 g05879(new_n6255, new_n6254_1, new_n6256);
xor_4  g05880(new_n6256, new_n6253, new_n6257);
and_8  g05881(new_n6257, new_n6252, new_n6258);
not_8  g05882(new_n6253, new_n6259);
xor_4  g05883(new_n6256, new_n6259, new_n6260);
and_8  g05884(new_n6260, new_n6251, new_n6261);
or_8   g05885(new_n6261, new_n6258, new_n6262);
and_8  g05886(n9189, n6877, new_n6263);
and_8  g05887(n7946, n2464, new_n6264);
or_8   g05888(new_n6264, new_n6263, new_n6265);
and_8  g05889(n7946, n6877, new_n6266);
and_8  g05890(n9189, n2464, new_n6267);
and_8  g05891(new_n6267, new_n6266, new_n6268);
and_8  g05892(n9400, n2024, new_n6269);
or_8   g05893(new_n6269, new_n6268, new_n6270);
nand_5 g05894(new_n6270, new_n6265, new_n6271);
or_8   g05895(new_n6271, new_n6262, new_n6272);
or_8   g05896(new_n6260, new_n6251, new_n6273_1);
or_8   g05897(new_n6257, new_n6252, new_n6274);
and_8  g05898(new_n6274, new_n6273_1, new_n6275);
not_8  g05899(new_n6271, new_n6276);
or_8   g05900(new_n6276, new_n6275, new_n6277);
and_8  g05901(new_n6277, new_n6272, new_n6278);
not_8  g05902(new_n6269, new_n6279);
or_8   g05903(new_n6279, new_n6266, new_n6280);
not_8  g05904(new_n6265, new_n6281);
or_8   g05905(new_n6268, new_n6281, new_n6282);
and_8  g05906(new_n6282, new_n6280, new_n6283);
and_8  g05907(new_n6283, new_n6269, new_n6284);
nor_6  g05908(new_n6284, new_n6278, new_n6285);
and_8  g05909(new_n6284, new_n6278, new_n6286);
or_8   g05910(new_n6286, new_n6285, new_n6287);
nor_6  g05911(new_n6280, new_n6281, new_n6288);
or_8   g05912(new_n6288, new_n6283, new_n6289);
not_8  g05913(new_n6289, new_n6290);
and_8  g05914(n4805, n2558, new_n6291);
and_8  g05915(n9763, n7236, new_n6292);
xor_4  g05916(new_n6292, new_n6291, new_n6293);
and_8  g05917(new_n6293, new_n6266, new_n6294_1);
and_8  g05918(n9400, n7946, new_n6295);
and_8  g05919(n6877, n2024, new_n6296);
xor_4  g05920(new_n6296, new_n6295, new_n6297);
and_8  g05921(new_n6297, new_n6294_1, new_n6298);
and_8  g05922(new_n6292, new_n6291, new_n6299);
and_8  g05923(n9111, n7236, new_n6300);
and_8  g05924(n9763, n3992, new_n6301);
xor_4  g05925(new_n6301, new_n6300, new_n6302);
and_8  g05926(new_n6302, new_n6299, new_n6303);
nor_6  g05927(new_n6302, new_n6299, new_n6304);
or_8   g05928(new_n6304, new_n6303, new_n6305);
and_8  g05929(n4805, n2498, new_n6306);
and_8  g05930(n11478, n2558, new_n6307);
xor_4  g05931(new_n6307, new_n6306, new_n6308);
not_8  g05932(new_n6308, new_n6309);
xor_4  g05933(new_n6309, new_n6305, new_n6310);
xor_4  g05934(new_n6297, new_n6294_1, new_n6311);
and_8  g05935(new_n6311, new_n6310, new_n6312);
or_8   g05936(new_n6312, new_n6298, new_n6313);
or_8   g05937(new_n6313, new_n6290, new_n6314);
not_8  g05938(new_n6304, new_n6315);
or_8   g05939(new_n6308, new_n6305, new_n6316);
and_8  g05940(new_n6316, new_n6315, new_n6317);
and_8  g05941(n11478, n2498, new_n6318);
not_8  g05942(new_n6318, new_n6319);
or_8   g05943(new_n6319, new_n6291, new_n6320);
and_8  g05944(n5283, n2558, new_n6321);
and_8  g05945(n5579, n4805, new_n6322);
or_8   g05946(new_n6322, new_n6321, new_n6323);
not_8  g05947(new_n6323, new_n6324);
and_8  g05948(new_n6322, new_n6321, new_n6325);
or_8   g05949(new_n6325, new_n6324, new_n6326);
and_8  g05950(new_n6326, new_n6320, new_n6327);
nor_6  g05951(new_n6324, new_n6320, new_n6328);
nor_6  g05952(new_n6328, new_n6327, new_n6329);
and_8  g05953(new_n6329, new_n6317, new_n6330);
nor_6  g05954(new_n6329, new_n6317, new_n6331);
or_8   g05955(new_n6331, new_n6330, new_n6332);
not_8  g05956(new_n6292, new_n6333);
and_8  g05957(n9111, n3992, new_n6334);
and_8  g05958(new_n6334, new_n6333, new_n6335);
and_8  g05959(n9763, n8384, new_n6336);
and_8  g05960(n7236, n3342, new_n6337);
nor_6  g05961(new_n6337, new_n6336, new_n6338);
nand_5 g05962(new_n6338, new_n6335, new_n6339);
and_8  g05963(new_n6337, new_n6336, new_n6340);
or_8   g05964(new_n6340, new_n6338, new_n6341);
or_8   g05965(new_n6341, new_n6335, new_n6342);
and_8  g05966(new_n6342, new_n6339, new_n6343);
xor_4  g05967(new_n6343, new_n6332, new_n6344);
xor_4  g05968(new_n6313, new_n6289, new_n6345);
or_8   g05969(new_n6345, new_n6344, new_n6346);
and_8  g05970(new_n6346, new_n6314, new_n6347);
xor_4  g05971(new_n6347, new_n6287, new_n6348);
and_8  g05972(n4805, n521, new_n6349);
or_8   g05973(new_n6325, new_n6318, new_n6350);
and_8  g05974(new_n6350, new_n6323, new_n6351);
xor_4  g05975(new_n6351, new_n6349, new_n6352);
and_8  g05976(n5283, n2498, new_n6353);
and_8  g05977(n2558, n137, new_n6354);
and_8  g05978(n11478, n5579, new_n6355);
xor_4  g05979(new_n6355, new_n6354, new_n6356);
xor_4  g05980(new_n6356, new_n6353, new_n6357);
xor_4  g05981(new_n6357, new_n6352, new_n6358_1);
and_8  g05982(new_n6327, new_n6318, new_n6359_1);
and_8  g05983(new_n6359_1, new_n6358_1, new_n6360);
nor_6  g05984(new_n6359_1, new_n6358_1, new_n6361);
or_8   g05985(new_n6361, new_n6360, new_n6362);
and_8  g05986(n7236, n806, new_n6363);
or_8   g05987(new_n6337, new_n6336, new_n6364);
and_8  g05988(new_n6364, new_n6334, new_n6365);
or_8   g05989(new_n6365, new_n6340, new_n6366);
xor_4  g05990(new_n6366, new_n6363, new_n6367);
and_8  g05991(n9111, n8384, new_n6368);
and_8  g05992(n9763, n6358, new_n6369);
and_8  g05993(n3992, n3342, new_n6370);
xor_4  g05994(new_n6370, new_n6369, new_n6371);
xor_4  g05995(new_n6371, new_n6368, new_n6372);
and_8  g05996(new_n6372, new_n6367, new_n6373);
nor_6  g05997(new_n6372, new_n6367, new_n6374);
or_8   g05998(new_n6374, new_n6373, new_n6375);
and_8  g05999(new_n6301, new_n6300, new_n6376);
nand_5 g06000(new_n6341, new_n6376, new_n6377);
xor_4  g06001(new_n6377, new_n6375, new_n6378);
xor_4  g06002(new_n6378, new_n6362, new_n6379);
not_8  g06003(new_n6332, new_n6380);
and_8  g06004(new_n6343, new_n6380, new_n6381);
nor_6  g06005(new_n6381, new_n6331, new_n6382);
xor_4  g06006(new_n6382, new_n6379, new_n6383);
xor_4  g06007(new_n6383, new_n6348, new_n6384);
and_8  g06008(new_n6384, new_n6250, new_n6385);
nor_6  g06009(new_n6384, new_n6250, new_n6386);
or_8   g06010(new_n6386, new_n6385, new_n6387);
and_8  g06011(new_n6246, new_n6231, new_n6388);
nor_6  g06012(new_n6388, new_n6248, new_n6389);
xnor_4 g06013(new_n6345, new_n6344, new_n6390);
and_8  g06014(new_n6390, new_n6389, new_n6391);
xor_4  g06015(new_n6293, new_n6266, new_n6392);
and_8  g06016(new_n6392, new_n6233, new_n6393);
and_8  g06017(n7265, n1333, new_n6394);
and_8  g06018(n7862, n2879, new_n6395);
xor_4  g06019(new_n6395, new_n6394, new_n6396);
or_8   g06020(new_n6396, new_n6393, new_n6397);
xor_4  g06021(new_n6311, new_n6310, new_n6398);
xnor_4 g06022(new_n6396, new_n6393, new_n6399);
or_8   g06023(new_n6399, new_n6398, new_n6400);
and_8  g06024(new_n6400, new_n6397, new_n6401);
xor_4  g06025(new_n6390, new_n6389, new_n6402);
and_8  g06026(new_n6402, new_n6401, new_n6403);
or_8   g06027(new_n6403, new_n6391, new_n6404);
xnor_4 g06028(new_n6404, new_n6387, n1847);
and_8  g06029(n5305, n1798, new_n6406);
and_8  g06030(n8759, n6703, new_n6407);
and_8  g06031(n5645, n5331, new_n6408);
and_8  g06032(n11876, n7965, new_n6409);
xor_4  g06033(new_n6409, new_n6408, new_n6410);
xor_4  g06034(new_n6410, new_n6407, new_n6411);
and_8  g06035(new_n6411, new_n6406, new_n6412);
and_8  g06036(n5305, n3932, new_n6413);
and_8  g06037(n5964, n1798, new_n6414);
xor_4  g06038(new_n6414, new_n6413, new_n6415);
xor_4  g06039(new_n6415, new_n6412, new_n6416);
and_8  g06040(new_n6410, new_n6407, new_n6417);
and_8  g06041(n9640, n8759, new_n6418);
and_8  g06042(n6776, n6703, new_n6419);
xor_4  g06043(new_n6419, new_n6418, new_n6420);
xor_4  g06044(new_n6420, new_n6417, new_n6421);
and_8  g06045(new_n6409, new_n6408, new_n6422);
and_8  g06046(n10898, n7965, new_n6423);
and_8  g06047(n11876, n7388, new_n6424);
xor_4  g06048(new_n6424, new_n6423, new_n6425);
xor_4  g06049(new_n6425, new_n6422, new_n6426);
and_8  g06050(n5331, n1067, new_n6427);
and_8  g06051(n8476, n5645, new_n6428);
xor_4  g06052(new_n6428, new_n6427, new_n6429_1);
xor_4  g06053(new_n6429_1, new_n6426, new_n6430);
xor_4  g06054(new_n6430, new_n6421, new_n6431_1);
xor_4  g06055(new_n6431_1, new_n6416, n2096);
xor_4  g06056(new_n3798, new_n3795, n2131);
and_8  g06057(n7456, n2564, new_n6434);
or_8   g06058(new_n3963, new_n3962, new_n6435);
and_8  g06059(new_n3963, new_n3962, new_n6436);
or_8   g06060(new_n6436, new_n3961, new_n6437);
and_8  g06061(new_n6437, new_n6435, new_n6438);
and_8  g06062(new_n6438, new_n6434, new_n6439);
xor_4  g06063(new_n6438, new_n6434, new_n6440);
and_8  g06064(n6770, n3932, new_n6441_1);
and_8  g06065(n9920, n1798, new_n6442);
xor_4  g06066(new_n6442, new_n3955, new_n6443);
xor_4  g06067(new_n6443, new_n6441_1, new_n6444);
and_8  g06068(new_n6444, new_n6440, new_n6445_1);
or_8   g06069(new_n6445_1, new_n6439, new_n6446);
and_8  g06070(n11662, n2564, new_n6447);
and_8  g06071(n7456, n4189, new_n6448);
xor_4  g06072(new_n6448, new_n6447, new_n6449);
not_8  g06073(new_n6449, new_n6450);
xor_4  g06074(new_n6450, new_n6446, new_n6451);
and_8  g06075(n12591, n6770, new_n6452);
and_8  g06076(n3627, n1798, new_n6453);
and_8  g06077(n9920, n3932, new_n6454);
xor_4  g06078(new_n6454, new_n6453, new_n6455);
xor_4  g06079(new_n6455, new_n6452, new_n6456);
or_8   g06080(new_n6442, new_n3955, new_n6457);
and_8  g06081(new_n6442, new_n3955, new_n6458);
or_8   g06082(new_n6458, new_n6441_1, new_n6459);
and_8  g06083(new_n6459, new_n6457, new_n6460);
xor_4  g06084(new_n6460, new_n6456, new_n6461);
xor_4  g06085(new_n6461, new_n6451, new_n6462);
and_8  g06086(n11662, n6687, new_n6463);
and_8  g06087(new_n3959, new_n3950, new_n6464);
and_8  g06088(new_n3965, new_n3960, new_n6465);
or_8   g06089(new_n6465, new_n6464, new_n6466);
nor_6  g06090(new_n6466, new_n6463, new_n6467);
xnor_4 g06091(new_n6444, new_n6440, new_n6468);
xor_4  g06092(new_n6466, new_n6463, new_n6469);
and_8  g06093(new_n6469, new_n6468, new_n6470);
or_8   g06094(new_n6470, new_n6467, new_n6471);
or_8   g06095(new_n6471, new_n6462, new_n6472);
and_8  g06096(new_n6455, new_n6452, new_n6473);
and_8  g06097(new_n6460, new_n6456, new_n6474);
or_8   g06098(new_n6474, new_n6473, new_n6475);
and_8  g06099(n10327, n2564, new_n6476);
and_8  g06100(n11662, n4189, new_n6477);
and_8  g06101(n9583, n6687, new_n6478);
xnor_4 g06102(new_n6478, new_n6477, new_n6479);
xor_4  g06103(new_n6479, new_n6476, new_n6480);
xor_4  g06104(new_n6480, new_n6475, new_n6481);
and_8  g06105(new_n6454, new_n6453, new_n6482);
and_8  g06106(n7456, n6770, new_n6483);
xnor_4 g06107(new_n6483, new_n6482, new_n6484);
and_8  g06108(n3932, n3627, new_n6485);
and_8  g06109(n12591, n9920, new_n6486);
and_8  g06110(n4516, n1798, new_n6487);
xnor_4 g06111(new_n6487, new_n6486, new_n6488);
xor_4  g06112(new_n6488, new_n6485, new_n6489);
xor_4  g06113(new_n6489, new_n6484, new_n6490);
xor_4  g06114(new_n6490, new_n6481, new_n6491);
not_8  g06115(new_n6491, new_n6492);
nand_5 g06116(new_n6449, new_n6446, new_n6493);
and_8  g06117(new_n6448, new_n6447, new_n6494);
not_8  g06118(new_n6461, new_n6495);
or_8   g06119(new_n6495, new_n6451, new_n6496);
xor_4  g06120(new_n6496, new_n6494, new_n6497);
and_8  g06121(new_n6497, new_n6493, new_n6498);
xor_4  g06122(new_n6498, new_n6492, new_n6499);
and_8  g06123(new_n6499, new_n6472, new_n6500);
not_8  g06124(new_n6472, new_n6501);
xor_4  g06125(new_n6498, new_n6491, new_n6502);
and_8  g06126(new_n6502, new_n6501, new_n6503);
or_8   g06127(new_n6503, new_n6500, new_n6504);
and_8  g06128(n10327, n6687, new_n6505);
xor_4  g06129(new_n6495, new_n6451, new_n6506);
not_8  g06130(new_n6471, new_n6507);
or_8   g06131(new_n6507, new_n6506, new_n6508);
and_8  g06132(new_n6508, new_n6472, new_n6509);
and_8  g06133(new_n6509, new_n6505, new_n6510);
nand_5 g06134(new_n3972, new_n3966, new_n6511);
xor_4  g06135(new_n6469, new_n6468, new_n6512);
nor_6  g06136(new_n6512, new_n6511, new_n6513);
xor_4  g06137(new_n6509, new_n6505, new_n6514);
and_8  g06138(new_n6514, new_n6513, new_n6515);
nor_6  g06139(new_n6515, new_n6510, new_n6516);
xor_4  g06140(new_n6516, new_n6504, new_n6517);
not_8  g06141(new_n6517, new_n6518);
and_8  g06142(n3022, n2226, new_n6519);
and_8  g06143(n9640, n1094, new_n6520);
and_8  g06144(n10678, n6703, new_n6521);
xor_4  g06145(new_n6521, new_n6520, new_n6522);
xor_4  g06146(new_n6522, new_n6519, new_n6523);
and_8  g06147(n6703, n1094, new_n6524);
or_8   g06148(new_n6524, new_n4008, new_n6525);
and_8  g06149(new_n6524, new_n4008, new_n6526);
and_8  g06150(n9640, n2226, new_n6527);
or_8   g06151(new_n6527, new_n6526, new_n6528);
and_8  g06152(new_n6528, new_n6525, new_n6529);
and_8  g06153(new_n6529, new_n6523, new_n6530);
nor_6  g06154(new_n6529, new_n6523, new_n6531);
or_8   g06155(new_n6531, new_n6530, new_n6532);
and_8  g06156(n10928, n10451, new_n6533);
and_8  g06157(n11023, n6986, new_n6534);
xor_4  g06158(new_n6534, new_n6533, new_n6535);
not_8  g06159(new_n6535, new_n6536);
or_8   g06160(new_n6536, new_n6532, new_n6537);
not_8  g06161(new_n6530, new_n6538);
or_8   g06162(new_n6529, new_n6523, new_n6539);
and_8  g06163(new_n6539, new_n6538, new_n6540);
or_8   g06164(new_n6535, new_n6540, new_n6541);
and_8  g06165(new_n6541, new_n6537, new_n6542);
and_8  g06166(n11023, n10928, new_n6543);
or_8   g06167(new_n4117, new_n4116, new_n6544);
and_8  g06168(new_n4117, new_n4116, new_n6545);
or_8   g06169(new_n6545, new_n4115, new_n6546);
and_8  g06170(new_n6546, new_n6544, new_n6547);
and_8  g06171(new_n6547, new_n6543, new_n6548);
xor_4  g06172(new_n6547, new_n6543, new_n6549);
xor_4  g06173(new_n6524, new_n4008, new_n6550);
xor_4  g06174(new_n6550, new_n6527, new_n6551);
and_8  g06175(new_n6551, new_n6549, new_n6552);
or_8   g06176(new_n6552, new_n6548, new_n6553);
and_8  g06177(new_n6553, new_n6542, new_n6554);
nor_6  g06178(new_n6553, new_n6542, new_n6555);
or_8   g06179(new_n6555, new_n6554, new_n6556);
and_8  g06180(n10451, n8336, new_n6557);
not_8  g06181(new_n6557, new_n6558);
nor_6  g06182(new_n6551, new_n6549, new_n6559);
or_8   g06183(new_n6559, new_n6552, new_n6560);
or_8   g06184(new_n6560, new_n6558, new_n6561);
not_8  g06185(new_n6561, new_n6562);
and_8  g06186(new_n4113, new_n4110, new_n6563);
and_8  g06187(new_n4119, new_n4114, new_n6564);
or_8   g06188(new_n6564, new_n6563, new_n6565);
xor_4  g06189(new_n6560, new_n6558, new_n6566);
and_8  g06190(new_n6566, new_n6565, new_n6567);
nor_6  g06191(new_n6567, new_n6562, new_n6568);
or_8   g06192(new_n6568, new_n6556, new_n6569);
not_8  g06193(new_n6569, new_n6570);
and_8  g06194(new_n6522, new_n6519, new_n6571);
or_8   g06195(new_n6530, new_n6571, new_n6572);
and_8  g06196(n10928, n10278, new_n6573);
and_8  g06197(n10451, n6986, new_n6574);
and_8  g06198(n11423, n8336, new_n6575);
xnor_4 g06199(new_n6575, new_n6574, new_n6576);
xor_4  g06200(new_n6576, new_n6573, new_n6577);
xor_4  g06201(new_n6577, new_n6572, new_n6578_1);
and_8  g06202(new_n6521, new_n6520, new_n6579);
and_8  g06203(n11023, n2226, new_n6580);
xnor_4 g06204(new_n6580, new_n6579, new_n6581);
not_8  g06205(n10678, new_n6582);
or_8   g06206(new_n6582, new_n4000, new_n6583);
and_8  g06207(n3022, n1094, new_n6584);
and_8  g06208(n7320, n6703, new_n6585);
xor_4  g06209(new_n6585, new_n6584, new_n6586);
xor_4  g06210(new_n6586, new_n6583, new_n6587);
xor_4  g06211(new_n6587, new_n6581, new_n6588);
nor_6  g06212(new_n6588, new_n6578_1, new_n6589);
and_8  g06213(new_n6588, new_n6578_1, new_n6590);
or_8   g06214(new_n6590, new_n6589, new_n6591);
not_8  g06215(new_n6537, new_n6592);
and_8  g06216(new_n6534, new_n6533, new_n6593);
xor_4  g06217(new_n6554, new_n6593, new_n6594);
or_8   g06218(new_n6594, new_n6592, new_n6595);
xor_4  g06219(new_n6595, new_n6591, new_n6596);
or_8   g06220(new_n6596, new_n6570, new_n6597);
and_8  g06221(new_n6595, new_n6591, new_n6598);
nor_6  g06222(new_n6595, new_n6591, new_n6599);
or_8   g06223(new_n6599, new_n6598, new_n6600);
or_8   g06224(new_n6600, new_n6569, new_n6601);
and_8  g06225(new_n6601, new_n6597, new_n6602);
and_8  g06226(n10278, n8336, new_n6603);
xor_4  g06227(new_n6553, new_n6542, new_n6604_1);
or_8   g06228(new_n6567, new_n6562, new_n6605);
or_8   g06229(new_n6605, new_n6604_1, new_n6606);
and_8  g06230(new_n6606, new_n6569, new_n6607);
or_8   g06231(new_n6607, new_n6603, new_n6608);
nand_5 g06232(new_n4121, new_n4120, new_n6609);
not_8  g06233(new_n6609, new_n6610);
xor_4  g06234(new_n6566, new_n6565, new_n6611_1);
and_8  g06235(new_n6611_1, new_n6610, new_n6612);
nor_6  g06236(new_n6607, new_n6603, new_n6613);
and_8  g06237(new_n6607, new_n6603, new_n6614);
or_8   g06238(new_n6614, new_n6613, new_n6615);
or_8   g06239(new_n6615, new_n6612, new_n6616);
and_8  g06240(new_n6616, new_n6608, new_n6617);
xnor_4 g06241(new_n6617, new_n6602, new_n6618);
and_8  g06242(n8665, n7160, new_n6619);
and_8  g06243(n4828, n1067, new_n6620);
and_8  g06244(n5645, n2515, new_n6621);
xor_4  g06245(new_n6621, new_n6620, new_n6622);
xor_4  g06246(new_n6622, new_n6619, new_n6623);
and_8  g06247(n5645, n4828, new_n6624);
and_8  g06248(n8665, n7891, new_n6625);
nor_6  g06249(new_n6625, new_n6624, new_n6626);
not_8  g06250(n1067, new_n6627);
not_8  g06251(n7160, new_n6628);
or_8   g06252(new_n6628, new_n6627, new_n6629);
xor_4  g06253(new_n6625, new_n6624, new_n6630);
and_8  g06254(new_n6630, new_n6629, new_n6631);
nor_6  g06255(new_n6631, new_n6626, new_n6632);
and_8  g06256(new_n6632, new_n6623, new_n6633);
and_8  g06257(new_n6622, new_n6619, new_n6634);
nor_6  g06258(new_n6622, new_n6619, new_n6635);
or_8   g06259(new_n6635, new_n6634, new_n6636);
or_8   g06260(new_n6631, new_n6626, new_n6637);
and_8  g06261(new_n6637, new_n6636, new_n6638);
or_8   g06262(new_n6638, new_n6633, new_n6639);
and_8  g06263(n12391, n2551, new_n6640);
and_8  g06264(n11922, n7891, new_n6641);
xor_4  g06265(new_n6641, new_n6640, new_n6642);
not_8  g06266(new_n6642, new_n6643);
or_8   g06267(new_n6643, new_n6639, new_n6644);
or_8   g06268(new_n6637, new_n6636, new_n6645_1);
or_8   g06269(new_n6632, new_n6623, new_n6646);
and_8  g06270(new_n6646, new_n6645_1, new_n6647);
or_8   g06271(new_n6642, new_n6647, new_n6648);
and_8  g06272(new_n6648, new_n6644, new_n6649);
and_8  g06273(n12391, n11922, new_n6650);
or_8   g06274(new_n4071, new_n4070, new_n6651);
or_8   g06275(new_n4074, new_n4069, new_n6652);
and_8  g06276(new_n6652, new_n6651, new_n6653);
and_8  g06277(new_n6653, new_n6650, new_n6654);
nor_6  g06278(new_n6630, new_n6629, new_n6655);
or_8   g06279(new_n6655, new_n6631, new_n6656);
xor_4  g06280(new_n6653, new_n6650, new_n6657);
and_8  g06281(new_n6657, new_n6656, new_n6658);
or_8   g06282(new_n6658, new_n6654, new_n6659);
and_8  g06283(new_n6659, new_n6649, new_n6660);
nor_6  g06284(new_n6659, new_n6649, new_n6661);
or_8   g06285(new_n6661, new_n6660, new_n6662);
not_8  g06286(n2551, new_n6663);
or_8   g06287(new_n4398, new_n6663, new_n6664);
nor_6  g06288(new_n6657, new_n6656, new_n6665);
or_8   g06289(new_n6665, new_n6658, new_n6666);
or_8   g06290(new_n6666, new_n6664, new_n6667);
and_8  g06291(new_n6666, new_n6664, new_n6668);
nor_6  g06292(new_n4076, new_n4066, new_n6669);
or_8   g06293(new_n6669, new_n6668, new_n6670);
and_8  g06294(new_n6670, new_n6667, new_n6671);
nor_6  g06295(new_n6671, new_n6662, new_n6672);
not_8  g06296(new_n6672, new_n6673);
or_8   g06297(new_n6633, new_n6634, new_n6674);
and_8  g06298(n12826, n12391, new_n6675);
and_8  g06299(n7891, n2551, new_n6676);
and_8  g06300(n12069, n4094, new_n6677);
xnor_4 g06301(new_n6677, new_n6676, new_n6678);
xor_4  g06302(new_n6678, new_n6675, new_n6679);
xor_4  g06303(new_n6679, new_n6674, new_n6680);
and_8  g06304(new_n6621, new_n6620, new_n6681);
and_8  g06305(n11922, n7160, new_n6682);
xor_4  g06306(new_n6682, new_n6681, new_n6683);
and_8  g06307(n2515, n1067, new_n6684);
and_8  g06308(n8665, n4828, new_n6685);
and_8  g06309(n5645, n1199, new_n6686);
or_8   g06310(new_n6686, new_n6685, new_n6687_1);
nand_5 g06311(new_n6686, new_n6685, new_n6688);
and_8  g06312(new_n6688, new_n6687_1, new_n6689_1);
xor_4  g06313(new_n6689_1, new_n6684, new_n6690);
xor_4  g06314(new_n6690, new_n6683, new_n6691);
xor_4  g06315(new_n6691, new_n6680, new_n6692);
not_8  g06316(new_n6644, new_n6693);
and_8  g06317(new_n6641, new_n6640, new_n6694);
xor_4  g06318(new_n6660, new_n6694, new_n6695);
nor_6  g06319(new_n6695, new_n6693, new_n6696);
nor_6  g06320(new_n6696, new_n6692, new_n6697);
and_8  g06321(new_n6696, new_n6692, new_n6698);
or_8   g06322(new_n6698, new_n6697, new_n6699);
and_8  g06323(new_n6699, new_n6673, new_n6700);
not_8  g06324(new_n6700, new_n6701);
or_8   g06325(new_n6699, new_n6673, new_n6702);
and_8  g06326(new_n6702, new_n6701, new_n6703_1);
and_8  g06327(n12826, n12069, new_n6704);
not_8  g06328(new_n6704, new_n6705);
and_8  g06329(new_n6671, new_n6662, new_n6706);
or_8   g06330(new_n6706, new_n6672, new_n6707);
and_8  g06331(new_n6707, new_n6705, new_n6708);
not_8  g06332(new_n4080, new_n6709);
or_8   g06333(new_n4076, new_n4066, new_n6710);
nor_6  g06334(new_n6666, new_n6664, new_n6711);
or_8   g06335(new_n6668, new_n6711, new_n6712);
xor_4  g06336(new_n6712, new_n6710, new_n6713);
or_8   g06337(new_n6713, new_n6709, new_n6714);
xor_4  g06338(new_n6707, new_n6705, new_n6715);
and_8  g06339(new_n6715, new_n6714, new_n6716);
nor_6  g06340(new_n6716, new_n6708, new_n6717);
xor_4  g06341(new_n6717, new_n6703_1, new_n6718);
not_8  g06342(new_n6718, new_n6719);
and_8  g06343(n3754, n996, new_n6720);
and_8  g06344(n10898, n5767, new_n6721);
and_8  g06345(n11876, n5319, new_n6722);
xor_4  g06346(new_n6722, new_n6721, new_n6723);
xor_4  g06347(new_n6723, new_n6720, new_n6724);
and_8  g06348(n10898, n996, new_n6725);
nor_6  g06349(new_n6725, new_n4035, new_n6726);
nand_5 g06350(n11876, n5767, new_n6727);
xor_4  g06351(new_n6725, new_n4035, new_n6728);
and_8  g06352(new_n6728, new_n6727, new_n6729);
nor_6  g06353(new_n6729, new_n6726, new_n6730);
and_8  g06354(new_n6730, new_n6724, new_n6731);
and_8  g06355(new_n6723, new_n6720, new_n6732);
nor_6  g06356(new_n6723, new_n6720, new_n6733);
or_8   g06357(new_n6733, new_n6732, new_n6734);
or_8   g06358(new_n6729, new_n6726, new_n6735);
and_8  g06359(new_n6735, new_n6734, new_n6736);
or_8   g06360(new_n6736, new_n6731, new_n6737);
and_8  g06361(n11153, n159, new_n6738);
and_8  g06362(n5314, n2749, new_n6739);
xor_4  g06363(new_n6739, new_n6738, new_n6740);
not_8  g06364(new_n6740, new_n6741);
or_8   g06365(new_n6741, new_n6737, new_n6742_1);
or_8   g06366(new_n6735, new_n6734, new_n6743);
or_8   g06367(new_n6730, new_n6724, new_n6744);
and_8  g06368(new_n6744, new_n6743, new_n6745);
or_8   g06369(new_n6740, new_n6745, new_n6746);
and_8  g06370(new_n6746, new_n6742_1, new_n6747);
and_8  g06371(n11153, n2749, new_n6748);
or_8   g06372(new_n4089, new_n4088_1, new_n6749);
or_8   g06373(new_n4092, new_n4087, new_n6750);
and_8  g06374(new_n6750, new_n6749, new_n6751);
and_8  g06375(new_n6751, new_n6748, new_n6752);
nor_6  g06376(new_n6751, new_n6748, new_n6753);
or_8   g06377(new_n6753, new_n6752, new_n6754);
xor_4  g06378(new_n6728, new_n6727, new_n6755);
nor_6  g06379(new_n6755, new_n6754, new_n6756);
or_8   g06380(new_n6756, new_n6752, new_n6757);
and_8  g06381(new_n6757, new_n6747, new_n6758);
nor_6  g06382(new_n6757, new_n6747, new_n6759);
or_8   g06383(new_n6759, new_n6758, new_n6760);
not_8  g06384(n159, new_n6761);
or_8   g06385(new_n4244, new_n6761, new_n6762);
and_8  g06386(new_n6755, new_n6754, new_n6763);
or_8   g06387(new_n6763, new_n6756, new_n6764);
or_8   g06388(new_n6764, new_n6762, new_n6765);
and_8  g06389(new_n6764, new_n6762, new_n6766);
and_8  g06390(new_n4085, new_n4082, new_n6767);
or_8   g06391(new_n4096, new_n6767, new_n6768);
not_8  g06392(new_n6768, new_n6769);
or_8   g06393(new_n6769, new_n6766, new_n6770_1);
and_8  g06394(new_n6770_1, new_n6765, new_n6771);
nor_6  g06395(new_n6771, new_n6760, new_n6772);
not_8  g06396(new_n6742_1, new_n6773);
and_8  g06397(new_n6739, new_n6738, new_n6774);
xor_4  g06398(new_n6758, new_n6774, new_n6775);
or_8   g06399(new_n6775, new_n6773, new_n6776_1);
or_8   g06400(new_n6731, new_n6732, new_n6777);
nand_5 g06401(n11153, n1510, new_n6778);
and_8  g06402(n5314, n159, new_n6779);
and_8  g06403(n12247, n11222, new_n6780);
xnor_4 g06404(new_n6780, new_n6779, new_n6781);
xor_4  g06405(new_n6781, new_n6778, new_n6782);
xor_4  g06406(new_n6782, new_n6777, new_n6783);
and_8  g06407(new_n6722, new_n6721, new_n6784);
and_8  g06408(n2749, n996, new_n6785);
xnor_4 g06409(new_n6785, new_n6784, new_n6786);
and_8  g06410(n10898, n5319, new_n6787);
and_8  g06411(n11876, n9457, new_n6788);
and_8  g06412(n5767, n3754, new_n6789);
xnor_4 g06413(new_n6789, new_n6788, new_n6790);
xor_4  g06414(new_n6790, new_n6787, new_n6791);
xor_4  g06415(new_n6791, new_n6786, new_n6792);
and_8  g06416(new_n6792, new_n6783, new_n6793);
nor_6  g06417(new_n6792, new_n6783, new_n6794);
or_8   g06418(new_n6794, new_n6793, new_n6795);
not_8  g06419(new_n6795, new_n6796);
xor_4  g06420(new_n6796, new_n6776_1, new_n6797_1);
or_8   g06421(new_n6797_1, new_n6772, new_n6798);
not_8  g06422(new_n6772, new_n6799);
xor_4  g06423(new_n6795, new_n6776_1, new_n6800);
or_8   g06424(new_n6800, new_n6799, new_n6801);
and_8  g06425(new_n6801, new_n6798, new_n6802);
and_8  g06426(n11222, n1510, new_n6803);
xor_4  g06427(new_n6771, new_n6760, new_n6804);
or_8   g06428(new_n6804, new_n6803, new_n6805);
xor_4  g06429(new_n6764, new_n6762, new_n6806_1);
xor_4  g06430(new_n6806_1, new_n6768, new_n6807);
and_8  g06431(new_n6807, new_n4101, new_n6808);
and_8  g06432(new_n6771, new_n6760, new_n6809_1);
or_8   g06433(new_n6809_1, new_n6772, new_n6810);
xor_4  g06434(new_n6810, new_n6803, new_n6811);
or_8   g06435(new_n6811, new_n6808, new_n6812);
and_8  g06436(new_n6812, new_n6805, new_n6813);
and_8  g06437(new_n6813, new_n6802, new_n6814);
and_8  g06438(new_n6800, new_n6799, new_n6815);
and_8  g06439(new_n6797_1, new_n6772, new_n6816);
or_8   g06440(new_n6816, new_n6815, new_n6817);
not_8  g06441(new_n6805, new_n6818);
not_8  g06442(new_n6808, new_n6819);
not_8  g06443(new_n6803, new_n6820);
xor_4  g06444(new_n6810, new_n6820, new_n6821);
and_8  g06445(new_n6821, new_n6819, new_n6822_1);
or_8   g06446(new_n6822_1, new_n6818, new_n6823);
and_8  g06447(new_n6823, new_n6817, new_n6824);
or_8   g06448(new_n6824, new_n6814, new_n6825);
or_8   g06449(new_n6821, new_n6819, new_n6826_1);
and_8  g06450(new_n6826_1, new_n6812, new_n6827);
xor_4  g06451(new_n6712, new_n6669, new_n6828);
and_8  g06452(new_n6828, new_n4080, new_n6829);
xor_4  g06453(new_n6707, new_n6704, new_n6830);
or_8   g06454(new_n6830, new_n6829, new_n6831);
or_8   g06455(new_n6715, new_n6714, new_n6832);
and_8  g06456(new_n6832, new_n6831, new_n6833);
or_8   g06457(new_n6833, new_n6827, new_n6834);
and_8  g06458(new_n6833, new_n6827, new_n6835);
and_8  g06459(new_n6713, new_n6709, new_n6836);
or_8   g06460(new_n6836, new_n6829, new_n6837);
and_8  g06461(new_n4103, new_n4081, new_n6838);
and_8  g06462(new_n4107, new_n4104, new_n6839);
or_8   g06463(new_n6839, new_n6838, new_n6840);
and_8  g06464(new_n6840, new_n6837, new_n6841);
nor_6  g06465(new_n6807, new_n4101, new_n6842);
or_8   g06466(new_n6842, new_n6808, new_n6843);
or_8   g06467(new_n6828, new_n4080, new_n6844);
and_8  g06468(new_n6844, new_n6714, new_n6845);
not_8  g06469(new_n4081, new_n6846);
xor_4  g06470(new_n4100, new_n4098, new_n6847);
or_8   g06471(new_n6847, new_n6846, new_n6848);
xor_4  g06472(new_n6847, new_n4081, new_n6849);
not_8  g06473(new_n4107, new_n6850);
or_8   g06474(new_n6850, new_n6849, new_n6851);
and_8  g06475(new_n6851, new_n6848, new_n6852);
or_8   g06476(new_n6852, new_n6845, new_n6853);
or_8   g06477(new_n6840, new_n6837, new_n6854);
and_8  g06478(new_n6854, new_n6853, new_n6855);
and_8  g06479(new_n6855, new_n6843, new_n6856);
or_8   g06480(new_n6856, new_n6841, new_n6857);
or_8   g06481(new_n6857, new_n6835, new_n6858);
and_8  g06482(new_n6858, new_n6834, new_n6859);
xor_4  g06483(new_n6859, new_n6825, new_n6860_1);
or_8   g06484(new_n6860_1, new_n6719, new_n6861);
nor_6  g06485(new_n6824, new_n6814, new_n6862);
xor_4  g06486(new_n6859, new_n6862, new_n6863);
or_8   g06487(new_n6863, new_n6718, new_n6864);
and_8  g06488(new_n6864, new_n6861, new_n6865);
nor_6  g06489(new_n6865, new_n6618, new_n6866);
and_8  g06490(new_n6865, new_n6618, new_n6867);
or_8   g06491(new_n6867, new_n6866, new_n6868);
xor_4  g06492(new_n6615, new_n6612, new_n6869);
not_8  g06493(new_n6869, new_n6870);
xor_4  g06494(new_n6611_1, new_n6609, new_n6871);
not_8  g06495(new_n6871, new_n6872);
xor_4  g06496(new_n6807, new_n4101, new_n6873);
xor_4  g06497(new_n6855, new_n6873, new_n6874);
and_8  g06498(new_n6874, new_n6872, new_n6875);
and_8  g06499(new_n4126, new_n4122, new_n6876);
and_8  g06500(new_n4127, new_n4109, new_n6877_1);
or_8   g06501(new_n6877_1, new_n6876, new_n6878);
xor_4  g06502(new_n6855, new_n6843, new_n6879);
or_8   g06503(new_n6879, new_n6871, new_n6880);
or_8   g06504(new_n6874, new_n6872, new_n6881);
and_8  g06505(new_n6881, new_n6880, new_n6882);
and_8  g06506(new_n6882, new_n6878, new_n6883);
or_8   g06507(new_n6883, new_n6875, new_n6884);
and_8  g06508(new_n6884, new_n6870, new_n6885);
not_8  g06509(new_n6876, new_n6886);
not_8  g06510(new_n4122, new_n6887);
xor_4  g06511(new_n4126, new_n6887, new_n6888);
or_8   g06512(new_n6888, new_n4108, new_n6889);
and_8  g06513(new_n6889, new_n6886, new_n6890);
and_8  g06514(new_n6879, new_n6871, new_n6891);
or_8   g06515(new_n6891, new_n6875, new_n6892);
or_8   g06516(new_n6892, new_n6890, new_n6893);
and_8  g06517(new_n6893, new_n6880, new_n6894);
or_8   g06518(new_n6894, new_n6869, new_n6895);
or_8   g06519(new_n6884, new_n6870, new_n6896);
and_8  g06520(new_n6896, new_n6895, new_n6897);
nor_6  g06521(new_n6833, new_n6827, new_n6898);
or_8   g06522(new_n6835, new_n6898, new_n6899);
xor_4  g06523(new_n6899, new_n6857, new_n6900);
and_8  g06524(new_n6900, new_n6897, new_n6901);
or_8   g06525(new_n6901, new_n6885, new_n6902);
xor_4  g06526(new_n6902, new_n6868, new_n6903);
or_8   g06527(new_n6903, new_n6518, new_n6904);
nor_6  g06528(new_n6901, new_n6885, new_n6905);
xor_4  g06529(new_n6905, new_n6868, new_n6906);
or_8   g06530(new_n6906, new_n6517, new_n6907);
and_8  g06531(new_n6907, new_n6904, new_n6908);
xor_4  g06532(new_n6514, new_n6513, new_n6909);
xor_4  g06533(new_n6900, new_n6897, new_n6910);
and_8  g06534(new_n6910, new_n6909, new_n6911);
or_8   g06535(new_n6910, new_n6909, new_n6912);
xor_4  g06536(new_n6512, new_n6511, new_n6913);
xor_4  g06537(new_n6882, new_n6878, new_n6914);
or_8   g06538(new_n6914, new_n6913, new_n6915);
nor_6  g06539(new_n4059, new_n3974, new_n6916);
and_8  g06540(new_n4128, new_n4060, new_n6917);
or_8   g06541(new_n6917, new_n6916, new_n6918);
not_8  g06542(new_n6913, new_n6919);
xor_4  g06543(new_n6914, new_n6919, new_n6920);
or_8   g06544(new_n6920, new_n6918, new_n6921);
and_8  g06545(new_n6921, new_n6915, new_n6922);
and_8  g06546(new_n6922, new_n6912, new_n6923);
or_8   g06547(new_n6923, new_n6911, new_n6924);
xor_4  g06548(new_n6924, new_n6908, n2301);
xor_4  g06549(new_n4057, new_n4054, n2316);
and_8  g06550(n4634, n1333, new_n6927);
or_8   g06551(new_n6242, new_n6241, new_n6928);
and_8  g06552(new_n6242, new_n6241, new_n6929);
or_8   g06553(new_n6929, new_n6240, new_n6930);
and_8  g06554(new_n6930, new_n6928, new_n6931);
and_8  g06555(new_n6931, new_n6927, new_n6932);
xor_4  g06556(new_n6931, new_n6927, new_n6933);
and_8  g06557(n11757, n2879, new_n6934);
and_8  g06558(n7265, n5240, new_n6935);
xor_4  g06559(new_n6935, new_n6234, new_n6936);
xor_4  g06560(new_n6936, new_n6934, new_n6937);
and_8  g06561(new_n6937, new_n6933, new_n6938);
or_8   g06562(new_n6938, new_n6932, new_n6939);
and_8  g06563(n4634, n3172, new_n6940);
and_8  g06564(n9195, n1333, new_n6941);
xor_4  g06565(new_n6941, new_n6940, new_n6942);
xnor_4 g06566(new_n6942, new_n6939, new_n6943);
and_8  g06567(n11757, n10223, new_n6944);
and_8  g06568(n5240, n2879, new_n6945);
and_8  g06569(n11821, n7265, new_n6946);
xor_4  g06570(new_n6946, new_n6945, new_n6947);
xnor_4 g06571(new_n6947, new_n6944, new_n6948);
or_8   g06572(new_n6935, new_n6234, new_n6949);
and_8  g06573(new_n6935, new_n6234, new_n6950);
or_8   g06574(new_n6950, new_n6934, new_n6951);
and_8  g06575(new_n6951, new_n6949, new_n6952);
xor_4  g06576(new_n6952, new_n6948, new_n6953);
xor_4  g06577(new_n6953, new_n6943, new_n6954);
nand_5 g06578(n9195, n7862, new_n6955);
xnor_4 g06579(new_n6937, new_n6933, new_n6956);
nor_6  g06580(new_n6956, new_n6955, new_n6957);
and_8  g06581(new_n6238, new_n6228, new_n6958);
and_8  g06582(new_n6244, new_n6239, new_n6959);
or_8   g06583(new_n6959, new_n6958, new_n6960);
xor_4  g06584(new_n6956, new_n6955, new_n6961);
and_8  g06585(new_n6961, new_n6960, new_n6962);
or_8   g06586(new_n6962, new_n6957, new_n6963);
nand_5 g06587(new_n6963, new_n6954, new_n6964);
nor_6  g06588(new_n6947, new_n6944, new_n6965);
nor_6  g06589(new_n6952, new_n6948, new_n6966);
or_8   g06590(new_n6966, new_n6965, new_n6967);
and_8  g06591(n2253, n1333, new_n6968);
and_8  g06592(n9195, n3172, new_n6969);
and_8  g06593(n7862, n3865, new_n6970);
xnor_4 g06594(new_n6970, new_n6969, new_n6971);
xor_4  g06595(new_n6971, new_n6968, new_n6972);
xor_4  g06596(new_n6972, new_n6967, new_n6973);
and_8  g06597(new_n6946, new_n6945, new_n6974);
and_8  g06598(n11757, n4634, new_n6975);
xor_4  g06599(new_n6975, new_n6974, new_n6976);
and_8  g06600(n11821, n2879, new_n6977);
and_8  g06601(n10223, n5240, new_n6978);
and_8  g06602(n9080, n7265, new_n6979);
xnor_4 g06603(new_n6979, new_n6978, new_n6980);
xor_4  g06604(new_n6980, new_n6977, new_n6981);
xor_4  g06605(new_n6981, new_n6976, new_n6982);
xnor_4 g06606(new_n6982, new_n6973, new_n6983);
nand_5 g06607(new_n6942, new_n6939, new_n6984);
nand_5 g06608(new_n6941, new_n6940, new_n6985);
nor_6  g06609(new_n6953, new_n6943, new_n6986_1);
xor_4  g06610(new_n6986_1, new_n6985, new_n6987);
and_8  g06611(new_n6987, new_n6984, new_n6988);
xor_4  g06612(new_n6988, new_n6983, new_n6989);
xor_4  g06613(new_n6989, new_n6964, new_n6990);
and_8  g06614(n7862, n2253, new_n6991);
xor_4  g06615(new_n6963, new_n6954, new_n6992);
and_8  g06616(new_n6992, new_n6991, new_n6993);
and_8  g06617(new_n6249, new_n6245, new_n6994);
xor_4  g06618(new_n6961, new_n6960, new_n6995);
and_8  g06619(new_n6995, new_n6994, new_n6996);
xor_4  g06620(new_n6992, new_n6991, new_n6997);
and_8  g06621(new_n6997, new_n6996, new_n6998);
or_8   g06622(new_n6998, new_n6993, new_n6999);
xor_4  g06623(new_n6999, new_n6990, new_n7000);
xor_4  g06624(new_n6997, new_n6996, new_n7001);
xor_4  g06625(new_n6995, new_n6994, new_n7002);
not_8  g06626(new_n6286, new_n7003);
and_8  g06627(n12145, n6877, new_n7004);
and_8  g06628(n9400, n2522, new_n7005);
and_8  g06629(n11311, n2024, new_n7006);
and_8  g06630(n7946, n4187, new_n7007);
xor_4  g06631(new_n7007, new_n6267, new_n7008);
xor_4  g06632(new_n7008, new_n7006, new_n7009);
xor_4  g06633(new_n7009, new_n7005, new_n7010);
not_8  g06634(new_n7010, new_n7011);
or_8   g06635(new_n6255, new_n6254_1, new_n7012);
or_8   g06636(new_n6256, new_n6259, new_n7013);
and_8  g06637(new_n7013, new_n7012, new_n7014);
xnor_4 g06638(new_n7014, new_n7011, new_n7015);
xor_4  g06639(new_n7015, new_n7004, new_n7016);
and_8  g06640(new_n6272, new_n6273_1, new_n7017);
not_8  g06641(new_n7017, new_n7018);
and_8  g06642(new_n7018, new_n7016, new_n7019);
and_8  g06643(new_n7015, new_n7004, new_n7020);
nor_6  g06644(new_n7015, new_n7004, new_n7021);
or_8   g06645(new_n7021, new_n7020, new_n7022);
and_8  g06646(new_n7017, new_n7022, new_n7023);
or_8   g06647(new_n7023, new_n7019, new_n7024);
nor_6  g06648(new_n7024, new_n7003, new_n7025);
and_8  g06649(new_n7024, new_n7003, new_n7026);
or_8   g06650(new_n7026, new_n7025, new_n7027);
xor_4  g06651(new_n6284, new_n6278, new_n7028);
and_8  g06652(new_n6347, new_n7028, new_n7029);
not_8  g06653(new_n7029, new_n7030);
or_8   g06654(new_n6383, new_n6348, new_n7031);
and_8  g06655(new_n7031, new_n7030, new_n7032);
and_8  g06656(new_n7032, new_n7027, new_n7033);
nor_6  g06657(new_n7026, new_n7025, new_n7034);
xor_4  g06658(new_n6347, new_n7028, new_n7035);
and_8  g06659(new_n6382, new_n6379, new_n7036);
nor_6  g06660(new_n6382, new_n6379, new_n7037);
or_8   g06661(new_n7037, new_n7036, new_n7038);
and_8  g06662(new_n7038, new_n7035, new_n7039);
or_8   g06663(new_n7039, new_n7029, new_n7040);
and_8  g06664(new_n7040, new_n7034, new_n7041);
or_8   g06665(new_n7041, new_n7033, new_n7042);
and_8  g06666(n11478, n521, new_n7043);
or_8   g06667(new_n6355, new_n6354, new_n7044);
and_8  g06668(new_n6355, new_n6354, new_n7045);
or_8   g06669(new_n7045, new_n6353, new_n7046);
and_8  g06670(new_n7046, new_n7044, new_n7047);
xnor_4 g06671(new_n7047, new_n7043, new_n7048);
and_8  g06672(n2498, n137, new_n7049);
and_8  g06673(n5579, n5283, new_n7050);
and_8  g06674(n6294, n2558, new_n7051);
xor_4  g06675(new_n7051, new_n7050, new_n7052);
xor_4  g06676(new_n7052, new_n7049, new_n7053);
xor_4  g06677(new_n7053, new_n7048, new_n7054);
and_8  g06678(n6016, n4805, new_n7055);
and_8  g06679(new_n6351, new_n6349, new_n7056);
and_8  g06680(new_n6357, new_n6352, new_n7057);
or_8   g06681(new_n7057, new_n7056, new_n7058);
nor_6  g06682(new_n7058, new_n7055, new_n7059);
and_8  g06683(new_n7058, new_n7055, new_n7060);
or_8   g06684(new_n7060, new_n7059, new_n7061);
xor_4  g06685(new_n7061, new_n7054, new_n7062);
xor_4  g06686(new_n7062, new_n6360, new_n7063);
or_8   g06687(new_n6377, new_n6375, new_n7064);
not_8  g06688(new_n7064, new_n7065);
and_8  g06689(n7270, n7236, new_n7066);
and_8  g06690(new_n6366, new_n6363, new_n7067);
or_8   g06691(new_n6373, new_n7067, new_n7068);
xor_4  g06692(new_n7068, new_n7066, new_n7069);
and_8  g06693(n3992, n806, new_n7070);
or_8   g06694(new_n6370, new_n6369, new_n7071);
and_8  g06695(new_n6370, new_n6369, new_n7072);
or_8   g06696(new_n7072, new_n6368, new_n7073);
and_8  g06697(new_n7073, new_n7071, new_n7074);
xnor_4 g06698(new_n7074, new_n7070, new_n7075);
and_8  g06699(n9111, n6358, new_n7076);
and_8  g06700(n8384, n3342, new_n7077);
and_8  g06701(n9763, n5198, new_n7078);
xnor_4 g06702(new_n7078, new_n7077, new_n7079);
xor_4  g06703(new_n7079, new_n7076, new_n7080);
nor_6  g06704(new_n7080, new_n7075, new_n7081);
and_8  g06705(new_n7080, new_n7075, new_n7082);
or_8   g06706(new_n7082, new_n7081, new_n7083);
xor_4  g06707(new_n7083, new_n7069, new_n7084);
not_8  g06708(new_n7084, new_n7085);
xor_4  g06709(new_n7085, new_n7065, new_n7086);
nor_6  g06710(new_n7086, new_n7063, new_n7087);
and_8  g06711(new_n7086, new_n7063, new_n7088);
or_8   g06712(new_n7088, new_n7087, new_n7089);
not_8  g06713(new_n6378, new_n7090);
and_8  g06714(new_n7090, new_n6362, new_n7091);
or_8   g06715(new_n7037, new_n7091, new_n7092);
not_8  g06716(new_n7092, new_n7093);
or_8   g06717(new_n7093, new_n7089, new_n7094);
xor_4  g06718(new_n7086, new_n7063, new_n7095);
or_8   g06719(new_n7092, new_n7095, new_n7096);
and_8  g06720(new_n7096, new_n7094, new_n7097);
xor_4  g06721(new_n7097, new_n7042, new_n7098);
or_8   g06722(new_n7098, new_n7002, new_n7099);
and_8  g06723(new_n7092, new_n7095, new_n7100);
and_8  g06724(new_n7093, new_n7089, new_n7101);
or_8   g06725(new_n7101, new_n7100, new_n7102);
or_8   g06726(new_n7102, new_n7042, new_n7103);
or_8   g06727(new_n7040, new_n7034, new_n7104);
or_8   g06728(new_n7032, new_n7027, new_n7105);
and_8  g06729(new_n7105, new_n7104, new_n7106);
or_8   g06730(new_n7097, new_n7106, new_n7107);
and_8  g06731(new_n7107, new_n7103, new_n7108);
xor_4  g06732(new_n7108, new_n7002, new_n7109);
nor_6  g06733(new_n6404, new_n6385, new_n7110);
nor_6  g06734(new_n7110, new_n6386, new_n7111);
or_8   g06735(new_n7111, new_n7109, new_n7112);
and_8  g06736(new_n7112, new_n7099, new_n7113);
or_8   g06737(new_n7113, new_n7001, new_n7114);
and_8  g06738(new_n7097, new_n7106, new_n7115);
or_8   g06739(new_n7115, new_n7033, new_n7116);
and_8  g06740(n12221, n6877, new_n7117);
not_8  g06741(new_n7117, new_n7118);
or_8   g06742(new_n7019, new_n7020, new_n7119);
or_8   g06743(new_n7009, new_n7005, new_n7120);
or_8   g06744(new_n7014, new_n7011, new_n7121);
and_8  g06745(new_n7121, new_n7120, new_n7122);
and_8  g06746(n11311, n9189, new_n7123);
and_8  g06747(n7946, n4203, new_n7124);
and_8  g06748(n4187, n2024, new_n7125);
xor_4  g06749(new_n7125, new_n7124, new_n7126);
xor_4  g06750(new_n7126, new_n7123, new_n7127);
or_8   g06751(new_n7007, new_n6267, new_n7128);
and_8  g06752(new_n7007, new_n6267, new_n7129);
or_8   g06753(new_n7129, new_n7006, new_n7130);
nand_5 g06754(new_n7130, new_n7128, new_n7131);
and_8  g06755(new_n7131, new_n7127, new_n7132);
nor_6  g06756(new_n7131, new_n7127, new_n7133);
or_8   g06757(new_n7133, new_n7132, new_n7134);
and_8  g06758(n12145, n9400, new_n7135);
and_8  g06759(n2522, n2464, new_n7136);
xor_4  g06760(new_n7136, new_n7135, new_n7137);
xor_4  g06761(new_n7137, new_n7134, new_n7138);
xor_4  g06762(new_n7138, new_n7122, new_n7139);
and_8  g06763(new_n7139, new_n7119, new_n7140);
nor_6  g06764(new_n7139, new_n7119, new_n7141);
or_8   g06765(new_n7141, new_n7140, new_n7142);
or_8   g06766(new_n7142, new_n7118, new_n7143);
xor_4  g06767(new_n7139, new_n7119, new_n7144);
or_8   g06768(new_n7144, new_n7117, new_n7145);
and_8  g06769(new_n7145, new_n7143, new_n7146);
xor_4  g06770(new_n7146, new_n7025, new_n7147);
xor_4  g06771(new_n7147, new_n7116, new_n7148);
or_8   g06772(new_n7084, new_n7064, new_n7149);
not_8  g06773(new_n7149, new_n7150);
and_8  g06774(n7236, n5153, new_n7151);
not_8  g06775(new_n7151, new_n7152);
and_8  g06776(n6358, n3342, new_n7153);
and_8  g06777(n9111, n5198, new_n7154);
and_8  g06778(n9763, n1471, new_n7155);
xor_4  g06779(new_n7155, new_n7154, new_n7156);
xor_4  g06780(new_n7156, new_n7153, new_n7157);
or_8   g06781(new_n7078, new_n7077, new_n7158);
or_8   g06782(new_n7079, new_n7076, new_n7159_1);
and_8  g06783(new_n7159_1, new_n7158, new_n7160_1);
xor_4  g06784(new_n7160_1, new_n7157, new_n7161);
and_8  g06785(n7270, n3992, new_n7162);
and_8  g06786(n8384, n806, new_n7163);
xor_4  g06787(new_n7163, new_n7162, new_n7164);
xor_4  g06788(new_n7164, new_n7161, new_n7165);
and_8  g06789(new_n7074, new_n7070, new_n7166);
or_8   g06790(new_n7081, new_n7166, new_n7167);
not_8  g06791(new_n7167, new_n7168);
xor_4  g06792(new_n7168, new_n7165, new_n7169);
nor_6  g06793(new_n7068, new_n7066, new_n7170);
and_8  g06794(new_n7083, new_n7069, new_n7171);
or_8   g06795(new_n7171, new_n7170, new_n7172);
or_8   g06796(new_n7172, new_n7169, new_n7173);
xor_4  g06797(new_n7167, new_n7165, new_n7174);
not_8  g06798(new_n7172, new_n7175);
or_8   g06799(new_n7175, new_n7174, new_n7176);
and_8  g06800(new_n7176, new_n7173, new_n7177);
xor_4  g06801(new_n7177, new_n7152, new_n7178);
and_8  g06802(new_n7178, new_n7150, new_n7179);
xor_4  g06803(new_n7177, new_n7151, new_n7180);
and_8  g06804(new_n7180, new_n7149, new_n7181);
or_8   g06805(new_n7181, new_n7179, new_n7182);
and_8  g06806(new_n7062, new_n6360, new_n7183);
not_8  g06807(new_n7183, new_n7184);
and_8  g06808(n5798, n4805, new_n7185);
and_8  g06809(n5579, n137, new_n7186);
and_8  g06810(n6797, n2558, new_n7187);
and_8  g06811(n6294, n2498, new_n7188);
xor_4  g06812(new_n7188, new_n7187, new_n7189);
xor_4  g06813(new_n7189, new_n7186, new_n7190);
or_8   g06814(new_n7051, new_n7050, new_n7191);
and_8  g06815(new_n7051, new_n7050, new_n7192);
or_8   g06816(new_n7192, new_n7049, new_n7193_1);
and_8  g06817(new_n7193_1, new_n7191, new_n7194);
xor_4  g06818(new_n7194, new_n7190, new_n7195);
and_8  g06819(n11478, n6016, new_n7196);
and_8  g06820(n5283, n521, new_n7197);
xor_4  g06821(new_n7197, new_n7196, new_n7198);
xor_4  g06822(new_n7198, new_n7195, new_n7199);
and_8  g06823(new_n7047, new_n7043, new_n7200);
not_8  g06824(new_n7048, new_n7201);
and_8  g06825(new_n7053, new_n7201, new_n7202);
or_8   g06826(new_n7202, new_n7200, new_n7203);
and_8  g06827(new_n7203, new_n7199, new_n7204);
nor_6  g06828(new_n7203, new_n7199, new_n7205);
or_8   g06829(new_n7205, new_n7204, new_n7206);
not_8  g06830(new_n7054, new_n7207);
nor_6  g06831(new_n7061, new_n7207, new_n7208);
or_8   g06832(new_n7208, new_n7059, new_n7209);
or_8   g06833(new_n7209, new_n7206, new_n7210);
xor_4  g06834(new_n7203, new_n7199, new_n7211);
nor_6  g06835(new_n7208, new_n7059, new_n7212);
or_8   g06836(new_n7212, new_n7211, new_n7213);
and_8  g06837(new_n7213, new_n7210, new_n7214);
xor_4  g06838(new_n7214, new_n7185, new_n7215);
and_8  g06839(new_n7215, new_n7184, new_n7216);
not_8  g06840(new_n7185, new_n7217);
xor_4  g06841(new_n7214, new_n7217, new_n7218);
and_8  g06842(new_n7218, new_n7183, new_n7219);
or_8   g06843(new_n7219, new_n7216, new_n7220);
or_8   g06844(new_n7220, new_n7182, new_n7221);
or_8   g06845(new_n7180, new_n7149, new_n7222);
or_8   g06846(new_n7178, new_n7150, new_n7223);
and_8  g06847(new_n7223, new_n7222, new_n7224);
or_8   g06848(new_n7218, new_n7183, new_n7225);
or_8   g06849(new_n7215, new_n7184, new_n7226);
and_8  g06850(new_n7226, new_n7225, new_n7227);
or_8   g06851(new_n7227, new_n7224, new_n7228);
and_8  g06852(new_n7228, new_n7221, new_n7229);
or_8   g06853(new_n7100, new_n7087, new_n7230);
and_8  g06854(new_n7230, new_n7229, new_n7231);
and_8  g06855(new_n7227, new_n7224, new_n7232);
and_8  g06856(new_n7220, new_n7182, new_n7233);
or_8   g06857(new_n7233, new_n7232, new_n7234);
not_8  g06858(new_n7230, new_n7235);
and_8  g06859(new_n7235, new_n7234, new_n7236_1);
nor_6  g06860(new_n7236_1, new_n7231, new_n7237);
or_8   g06861(new_n7237, new_n7148, new_n7238);
and_8  g06862(new_n7103, new_n7104, new_n7239);
xor_4  g06863(new_n7147, new_n7239, new_n7240);
or_8   g06864(new_n7236_1, new_n7231, new_n7241);
or_8   g06865(new_n7241, new_n7240, new_n7242);
and_8  g06866(new_n7242, new_n7238, new_n7243);
not_8  g06867(new_n7001, new_n7244);
not_8  g06868(new_n7002, new_n7245);
and_8  g06869(new_n7108, new_n7245, new_n7246);
xor_4  g06870(new_n7108, new_n7245, new_n7247);
or_8   g06871(new_n7110, new_n6386, new_n7248);
and_8  g06872(new_n7248, new_n7247, new_n7249);
or_8   g06873(new_n7249, new_n7246, new_n7250);
and_8  g06874(new_n7250, new_n7244, new_n7251);
and_8  g06875(new_n7113, new_n7001, new_n7252);
or_8   g06876(new_n7252, new_n7251, new_n7253);
or_8   g06877(new_n7253, new_n7243, new_n7254);
and_8  g06878(new_n7254, new_n7114, new_n7255);
or_8   g06879(new_n7255, new_n7000, new_n7256);
not_8  g06880(new_n7000, new_n7257);
xor_4  g06881(new_n7255, new_n7257, new_n7258);
not_8  g06882(new_n7140, new_n7259);
nor_6  g06883(new_n7126, new_n7123, new_n7260);
or_8   g06884(new_n7132, new_n7260, new_n7261);
and_8  g06885(n12221, n9400, new_n7262);
and_8  g06886(n12145, n2464, new_n7263);
and_8  g06887(n10217, n6877, new_n7264);
xnor_4 g06888(new_n7264, new_n7263, new_n7265_1);
xor_4  g06889(new_n7265_1, new_n7262, new_n7266);
xor_4  g06890(new_n7266, new_n7261, new_n7267);
and_8  g06891(new_n7125, new_n7124, new_n7268);
and_8  g06892(n11311, n2522, new_n7269);
xnor_4 g06893(new_n7269, new_n7268, new_n7270_1);
and_8  g06894(n4203, n2024, new_n7271);
and_8  g06895(n9189, n4187, new_n7272);
and_8  g06896(n12753, n7946, new_n7273);
xnor_4 g06897(new_n7273, new_n7272, new_n7274);
xor_4  g06898(new_n7274, new_n7271, new_n7275);
xor_4  g06899(new_n7275, new_n7270_1, new_n7276);
not_8  g06900(new_n7276, new_n7277);
xor_4  g06901(new_n7277, new_n7267, new_n7278);
nand_5 g06902(new_n7137, new_n7134, new_n7279);
nand_5 g06903(new_n7136, new_n7135, new_n7280);
or_8   g06904(new_n7137, new_n7134, new_n7281);
and_8  g06905(new_n7281, new_n7122, new_n7282);
xor_4  g06906(new_n7282, new_n7280, new_n7283);
and_8  g06907(new_n7283, new_n7279, new_n7284);
xnor_4 g06908(new_n7284, new_n7278, new_n7285);
xor_4  g06909(new_n7285, new_n7259, new_n7286);
not_8  g06910(new_n7143, new_n7287);
and_8  g06911(new_n7146, new_n7025, new_n7288);
or_8   g06912(new_n7288, new_n7287, new_n7289);
xor_4  g06913(new_n7289, new_n7286, new_n7290);
not_8  g06914(new_n7290, new_n7291);
and_8  g06915(n4805, n2347, new_n7292);
and_8  g06916(n6016, n5283, new_n7293);
and_8  g06917(n11478, n5798, new_n7294_1);
xnor_4 g06918(new_n7294_1, new_n7293, new_n7295);
xor_4  g06919(new_n7295, new_n7292, new_n7296);
nand_5 g06920(new_n7189, new_n7186, new_n7297);
nand_5 g06921(new_n7194, new_n7190, new_n7298);
and_8  g06922(new_n7298, new_n7297, new_n7299);
xor_4  g06923(new_n7299, new_n7296, new_n7300);
and_8  g06924(new_n7188, new_n7187, new_n7301);
and_8  g06925(n521, n137, new_n7302);
xnor_4 g06926(new_n7302, new_n7301, new_n7303);
and_8  g06927(n6797, n2498, new_n7304);
and_8  g06928(n6294, n5579, new_n7305);
and_8  g06929(n3146, n2558, new_n7306);
xnor_4 g06930(new_n7306, new_n7305, new_n7307);
xor_4  g06931(new_n7307, new_n7304, new_n7308);
xor_4  g06932(new_n7308, new_n7303, new_n7309);
xor_4  g06933(new_n7309, new_n7300, new_n7310);
nand_5 g06934(new_n7198, new_n7195, new_n7311);
not_8  g06935(new_n7311, new_n7312);
and_8  g06936(new_n7197, new_n7196, new_n7313);
xor_4  g06937(new_n7204, new_n7313, new_n7314);
or_8   g06938(new_n7314, new_n7312, new_n7315);
and_8  g06939(new_n7315, new_n7310, new_n7316);
not_8  g06940(new_n7296, new_n7317);
xor_4  g06941(new_n7299, new_n7317, new_n7318);
xor_4  g06942(new_n7309, new_n7318, new_n7319);
not_8  g06943(new_n7313, new_n7320_1);
xor_4  g06944(new_n7204, new_n7320_1, new_n7321);
and_8  g06945(new_n7321, new_n7311, new_n7322);
and_8  g06946(new_n7322, new_n7319, new_n7323);
or_8   g06947(new_n7323, new_n7316, new_n7324);
or_8   g06948(new_n7324, new_n7210, new_n7325);
not_8  g06949(new_n7210, new_n7326);
or_8   g06950(new_n7322, new_n7319, new_n7327);
or_8   g06951(new_n7315, new_n7310, new_n7328);
and_8  g06952(new_n7328, new_n7327, new_n7329);
or_8   g06953(new_n7329, new_n7326, new_n7330);
and_8  g06954(new_n7330, new_n7325, new_n7331);
and_8  g06955(new_n7214, new_n7185, new_n7332);
not_8  g06956(new_n7332, new_n7333);
xor_4  g06957(new_n7212, new_n7206, new_n7334);
and_8  g06958(new_n7334, new_n7217, new_n7335);
or_8   g06959(new_n7335, new_n7184, new_n7336);
and_8  g06960(new_n7336, new_n7333, new_n7337);
xor_4  g06961(new_n7337, new_n7331, new_n7338);
not_8  g06962(new_n7173, new_n7339);
nand_5 g06963(new_n7164, new_n7161, new_n7340);
and_8  g06964(new_n7163, new_n7162, new_n7341);
and_8  g06965(new_n7167, new_n7165, new_n7342);
and_8  g06966(new_n7342, new_n7341, new_n7343);
nor_6  g06967(new_n7342, new_n7341, new_n7344);
or_8   g06968(new_n7344, new_n7343, new_n7345);
and_8  g06969(new_n7345, new_n7340, new_n7346);
and_8  g06970(new_n7155, new_n7154, new_n7347);
and_8  g06971(n6358, n806, new_n7348);
xnor_4 g06972(new_n7348, new_n7347, new_n7349);
and_8  g06973(n9111, n1471, new_n7350);
and_8  g06974(n5198, n3342, new_n7351);
and_8  g06975(n9763, n7646, new_n7352);
xnor_4 g06976(new_n7352, new_n7351, new_n7353);
xor_4  g06977(new_n7353, new_n7350, new_n7354_1);
xnor_4 g06978(new_n7354_1, new_n7349, new_n7355);
and_8  g06979(new_n7156, new_n7153, new_n7356);
and_8  g06980(new_n7160_1, new_n7157, new_n7357);
nor_6  g06981(new_n7357, new_n7356, new_n7358);
and_8  g06982(n5153, n3992, new_n7359);
and_8  g06983(n8384, n7270, new_n7360);
and_8  g06984(n7236, n2507, new_n7361);
xnor_4 g06985(new_n7361, new_n7360, new_n7362);
xor_4  g06986(new_n7362, new_n7359, new_n7363);
xor_4  g06987(new_n7363, new_n7358, new_n7364);
xor_4  g06988(new_n7364, new_n7355, new_n7365);
or_8   g06989(new_n7365, new_n7346, new_n7366);
not_8  g06990(new_n7340, new_n7367);
xor_4  g06991(new_n7342, new_n7341, new_n7368);
or_8   g06992(new_n7368, new_n7367, new_n7369);
not_8  g06993(new_n7365, new_n7370);
or_8   g06994(new_n7370, new_n7369, new_n7371);
and_8  g06995(new_n7371, new_n7366, new_n7372);
and_8  g06996(new_n7372, new_n7339, new_n7373);
and_8  g06997(new_n7370, new_n7369, new_n7374);
and_8  g06998(new_n7365, new_n7346, new_n7375);
or_8   g06999(new_n7375, new_n7374, new_n7376);
and_8  g07000(new_n7376, new_n7173, new_n7377);
or_8   g07001(new_n7377, new_n7373, new_n7378);
or_8   g07002(new_n7177, new_n7151, new_n7379);
and_8  g07003(new_n7177, new_n7151, new_n7380);
or_8   g07004(new_n7380, new_n7150, new_n7381);
and_8  g07005(new_n7381, new_n7379, new_n7382);
xor_4  g07006(new_n7382, new_n7378, new_n7383);
and_8  g07007(new_n7383, new_n7338, new_n7384);
not_8  g07008(new_n7336, new_n7385);
or_8   g07009(new_n7385, new_n7332, new_n7386);
xor_4  g07010(new_n7386, new_n7331, new_n7387);
or_8   g07011(new_n7376, new_n7173, new_n7388_1);
or_8   g07012(new_n7372, new_n7339, new_n7389);
and_8  g07013(new_n7389, new_n7388_1, new_n7390);
xor_4  g07014(new_n7382, new_n7390, new_n7391);
and_8  g07015(new_n7391, new_n7387, new_n7392);
or_8   g07016(new_n7392, new_n7384, new_n7393);
or_8   g07017(new_n7235, new_n7234, new_n7394);
and_8  g07018(new_n7394, new_n7221, new_n7395);
or_8   g07019(new_n7395, new_n7393, new_n7396);
or_8   g07020(new_n7391, new_n7387, new_n7397);
or_8   g07021(new_n7383, new_n7338, new_n7398);
and_8  g07022(new_n7398, new_n7397, new_n7399);
or_8   g07023(new_n7231, new_n7232, new_n7400);
or_8   g07024(new_n7400, new_n7399, new_n7401);
and_8  g07025(new_n7401, new_n7396, new_n7402);
xor_4  g07026(new_n7402, new_n7291, new_n7403);
and_8  g07027(new_n7147, new_n7239, new_n7404);
and_8  g07028(new_n7241, new_n7240, new_n7405);
or_8   g07029(new_n7405, new_n7404, new_n7406);
and_8  g07030(new_n7406, new_n7403, new_n7407);
xor_4  g07031(new_n7402, new_n7290, new_n7408);
not_8  g07032(new_n7404, new_n7409);
and_8  g07033(new_n7238, new_n7409, new_n7410);
and_8  g07034(new_n7410, new_n7408, new_n7411);
nor_6  g07035(new_n7411, new_n7407, new_n7412);
or_8   g07036(new_n7412, new_n7258, new_n7413);
and_8  g07037(new_n7413, new_n7256, new_n7414);
nor_6  g07038(new_n7402, new_n7291, new_n7415);
or_8   g07039(new_n7407, new_n7415, new_n7416);
nand_5 g07040(n4805, n1576, new_n7417);
nand_5 g07041(new_n7204, new_n7313, new_n7418);
and_8  g07042(new_n7327, new_n7418, new_n7419);
xor_4  g07043(new_n7419, new_n7417, new_n7420);
not_8  g07044(new_n7420, new_n7421);
or_8   g07045(new_n7421, new_n7416, new_n7422);
or_8   g07046(new_n7402, new_n7291, new_n7423);
or_8   g07047(new_n7410, new_n7408, new_n7424);
and_8  g07048(new_n7424, new_n7423, new_n7425);
or_8   g07049(new_n7420, new_n7425, new_n7426);
and_8  g07050(new_n7426, new_n7422, new_n7427);
or_8   g07051(new_n7285, new_n7259, new_n7428);
not_8  g07052(new_n7428, new_n7429);
and_8  g07053(new_n7289, new_n7286, new_n7430);
nor_6  g07054(new_n7430, new_n7429, new_n7431);
and_8  g07055(new_n7382, new_n7390, new_n7432);
or_8   g07056(new_n7432, new_n7373, new_n7433);
and_8  g07057(new_n7266, new_n7261, new_n7434);
and_8  g07058(new_n7277, new_n7267, new_n7435);
or_8   g07059(new_n7435, new_n7434, new_n7436_1);
and_8  g07060(n9189, n4203, new_n7437);
and_8  g07061(n4187, n2522, new_n7438);
xor_4  g07062(new_n7438, new_n7437, new_n7439);
and_8  g07063(n9763, n4722, new_n7440);
and_8  g07064(n10217, n9400, new_n7441);
xor_4  g07065(new_n7441, new_n7440, new_n7442);
xor_4  g07066(new_n7442, new_n7439, new_n7443);
and_8  g07067(n9111, n7646, new_n7444);
and_8  g07068(n12221, n2464, new_n7445);
and_8  g07069(n12145, n11311, new_n7446);
xor_4  g07070(new_n7446, new_n7445, new_n7447);
xor_4  g07071(new_n7447, new_n7444, new_n7448);
xor_4  g07072(new_n7448, new_n7443, new_n7449);
xor_4  g07073(new_n7449, new_n7436_1, new_n7450);
xor_4  g07074(new_n7450, new_n7433, new_n7451);
xor_4  g07075(new_n7451, new_n7431, new_n7452);
not_8  g07076(new_n7280, new_n7453);
nand_5 g07077(new_n7282, new_n7453, new_n7454);
or_8   g07078(new_n7284, new_n7278, new_n7455);
nand_5 g07079(new_n7455, new_n7454, new_n7456_1);
or_8   g07080(new_n7374, new_n7343, new_n7457);
xor_4  g07081(new_n7457, new_n7456_1, new_n7458);
and_8  g07082(n11821, n10223, new_n7459);
and_8  g07083(n9080, n2879, new_n7460);
xor_4  g07084(new_n7460, new_n7459, new_n7461);
and_8  g07085(n11757, n9195, new_n7462);
and_8  g07086(n7862, n2512, new_n7463);
xor_4  g07087(new_n7463, new_n7462, new_n7464);
xor_4  g07088(new_n7464, new_n7461, new_n7465);
and_8  g07089(new_n6970, new_n6969, new_n7466);
or_8   g07090(new_n6970, new_n6969, new_n7467);
and_8  g07091(new_n7467, new_n6968, new_n7468);
or_8   g07092(new_n7468, new_n7466, new_n7469);
xor_4  g07093(new_n7469, new_n7465, new_n7470);
nand_5 g07094(n12753, n2024, new_n7471);
and_8  g07095(n3865, n1333, new_n7472);
and_8  g07096(n5240, n4634, new_n7473);
xor_4  g07097(new_n7473, new_n7472, new_n7474);
xor_4  g07098(new_n7474, new_n7471, new_n7475);
xor_4  g07099(new_n7475, new_n7470, new_n7476);
xor_4  g07100(new_n7476, new_n7458, new_n7477);
not_8  g07101(new_n7477, new_n7478);
not_8  g07102(new_n6985, new_n7479);
and_8  g07103(new_n6986_1, new_n7479, new_n7480);
not_8  g07104(new_n6988, new_n7481);
and_8  g07105(new_n7481, new_n6983, new_n7482);
or_8   g07106(new_n7482, new_n7480, new_n7483);
not_8  g07107(new_n7483, new_n7484);
and_8  g07108(new_n6972, new_n6967, new_n7485);
and_8  g07109(new_n6982, new_n6973, new_n7486);
or_8   g07110(new_n7486, new_n7485, new_n7487);
and_8  g07111(new_n7269, new_n7268, new_n7488);
nor_6  g07112(new_n7275, new_n7270_1, new_n7489);
or_8   g07113(new_n7489, new_n7488, new_n7490);
and_8  g07114(n8384, n5153, new_n7491);
and_8  g07115(n7270, n6358, new_n7492);
xor_4  g07116(new_n7492, new_n7491, new_n7493);
nand_5 g07117(new_n7273, new_n7272, new_n7494);
or_8   g07118(new_n7273, new_n7272, new_n7495);
nand_5 g07119(new_n7495, new_n7271, new_n7496);
and_8  g07120(new_n7496, new_n7494, new_n7497);
xnor_4 g07121(new_n7497, new_n7493, new_n7498);
xor_4  g07122(new_n7498, new_n7490, new_n7499);
xor_4  g07123(new_n7499, new_n7487, new_n7500_1);
and_8  g07124(n5198, n806, new_n7501);
and_8  g07125(n3992, n2507, new_n7502);
xor_4  g07126(new_n7502, new_n7501, new_n7503);
and_8  g07127(n7823, n6877, new_n7504);
and_8  g07128(n3342, n1471, new_n7505);
xor_4  g07129(new_n7505, new_n7504, new_n7506);
xor_4  g07130(new_n7506, new_n7503, new_n7507);
and_8  g07131(new_n7352, new_n7351, new_n7508);
or_8   g07132(new_n7352, new_n7351, new_n7509);
and_8  g07133(new_n7509, new_n7350, new_n7510);
or_8   g07134(new_n7510, new_n7508, new_n7511);
xor_4  g07135(new_n7511, new_n7507, new_n7512);
xor_4  g07136(new_n7512, new_n7500_1, new_n7513);
and_8  g07137(new_n7363, new_n7358, new_n7514);
and_8  g07138(new_n7364, new_n7355, new_n7515);
or_8   g07139(new_n7515, new_n7514, new_n7516);
or_8   g07140(new_n7264, new_n7263, new_n7517);
or_8   g07141(new_n7265_1, new_n7262, new_n7518);
and_8  g07142(new_n7518, new_n7517, new_n7519);
and_8  g07143(n7236, n6431, new_n7520);
and_8  g07144(n10174, n7946, new_n7521);
xor_4  g07145(new_n7521, new_n7520, new_n7522);
xor_4  g07146(new_n7522, new_n7519, new_n7523_1);
xor_4  g07147(new_n7523_1, new_n7516, new_n7524);
xor_4  g07148(new_n7524, new_n7513, new_n7525);
xor_4  g07149(new_n7525, new_n7484, new_n7526);
or_8   g07150(new_n7526, new_n7478, new_n7527);
xor_4  g07151(new_n7525, new_n7483, new_n7528);
or_8   g07152(new_n7528, new_n7477, new_n7529);
and_8  g07153(new_n7529, new_n7527, new_n7530);
xor_4  g07154(new_n7530, new_n7452, new_n7531);
and_8  g07155(new_n7400, new_n7399, new_n7532);
or_8   g07156(new_n7532, new_n7384, new_n7533);
nor_6  g07157(new_n6989, new_n6964, new_n7534);
and_8  g07158(new_n6999, new_n6990, new_n7535);
or_8   g07159(new_n7535, new_n7534, new_n7536);
not_8  g07160(new_n7325, new_n7537);
and_8  g07161(new_n7386, new_n7331, new_n7538);
nor_6  g07162(new_n7538, new_n7537, new_n7539);
nand_5 g07163(new_n7348, new_n7347, new_n7540);
or_8   g07164(new_n7354_1, new_n7349, new_n7541);
nand_5 g07165(new_n7541, new_n7540, new_n7542);
nand_5 g07166(new_n7302, new_n7301, new_n7543);
or_8   g07167(new_n7308, new_n7303, new_n7544);
and_8  g07168(new_n7544, new_n7543, new_n7545);
xor_4  g07169(new_n7545, new_n7542, new_n7546_1);
or_8   g07170(new_n6975, new_n6974, new_n7547);
nand_5 g07171(new_n6981, new_n6976, new_n7548);
and_8  g07172(new_n7548, new_n7547, new_n7549);
nand_5 g07173(n3172, n2253, new_n7550);
and_8  g07174(n6797, n5579, new_n7551);
and_8  g07175(n5798, n5283, new_n7552);
xor_4  g07176(new_n7552, new_n7551, new_n7553);
xor_4  g07177(new_n7553, new_n7550, new_n7554);
xor_4  g07178(new_n7554, new_n7549, new_n7555);
or_8   g07179(new_n7294_1, new_n7293, new_n7556);
or_8   g07180(new_n7295, new_n7292, new_n7557);
and_8  g07181(new_n7557, new_n7556, new_n7558);
or_8   g07182(new_n7306, new_n7305, new_n7559);
or_8   g07183(new_n7307, new_n7304, new_n7560);
and_8  g07184(new_n7560, new_n7559, new_n7561);
xor_4  g07185(new_n7561, new_n7558, new_n7562);
and_8  g07186(n11478, n2347, new_n7563);
and_8  g07187(n3146, n2498, new_n7564);
xor_4  g07188(new_n7564, new_n7563, new_n7565);
xor_4  g07189(new_n7565, new_n7562, new_n7566);
xor_4  g07190(new_n7566, new_n7555, new_n7567);
xor_4  g07191(new_n7567, new_n7546_1, new_n7568_1);
nand_5 g07192(new_n7299, new_n7296, new_n7569);
or_8   g07193(new_n7309, new_n7318, new_n7570);
and_8  g07194(new_n7570, new_n7569, new_n7571);
or_8   g07195(new_n6979, new_n6978, new_n7572);
or_8   g07196(new_n6980, new_n6977, new_n7573);
and_8  g07197(new_n7573, new_n7572, new_n7574);
nand_5 g07198(n6016, n137, new_n7575);
and_8  g07199(n7265, n6826, new_n7576);
and_8  g07200(n6294, n521, new_n7577);
xor_4  g07201(new_n7577, new_n7576, new_n7578);
xor_4  g07202(new_n7578, new_n7575, new_n7579);
xor_4  g07203(new_n7579, new_n7574, new_n7580);
not_8  g07204(n4938, new_n7581);
or_8   g07205(new_n7581, new_n1134, new_n7582);
or_8   g07206(new_n7361, new_n7360, new_n7583);
or_8   g07207(new_n7362, new_n7359, new_n7584);
and_8  g07208(new_n7584, new_n7583, new_n7585);
xor_4  g07209(new_n7585, new_n7582, new_n7586);
xor_4  g07210(new_n7586, new_n7580, new_n7587);
xor_4  g07211(new_n7587, new_n7571, new_n7588);
not_8  g07212(new_n7588, new_n7589);
or_8   g07213(new_n7589, new_n7568_1, new_n7590);
not_8  g07214(new_n7546_1, new_n7591);
xor_4  g07215(new_n7567, new_n7591, new_n7592);
or_8   g07216(new_n7588, new_n7592, new_n7593);
and_8  g07217(new_n7593, new_n7590, new_n7594);
xor_4  g07218(new_n7594, new_n7539, new_n7595);
or_8   g07219(new_n7595, new_n7536, new_n7596);
not_8  g07220(new_n7536, new_n7597);
or_8   g07221(new_n7538, new_n7537, new_n7598);
xor_4  g07222(new_n7594, new_n7598, new_n7599);
or_8   g07223(new_n7599, new_n7597, new_n7600);
and_8  g07224(new_n7600, new_n7596, new_n7601);
xor_4  g07225(new_n7601, new_n7533, new_n7602);
or_8   g07226(new_n7602, new_n7531, new_n7603);
or_8   g07227(new_n7430, new_n7429, new_n7604);
xor_4  g07228(new_n7451, new_n7604, new_n7605);
xor_4  g07229(new_n7530, new_n7605, new_n7606);
and_8  g07230(new_n7396, new_n7397, new_n7607);
xor_4  g07231(new_n7601, new_n7607, new_n7608);
or_8   g07232(new_n7608, new_n7606, new_n7609);
and_8  g07233(new_n7609, new_n7603, new_n7610_1);
and_8  g07234(new_n7610_1, new_n7427, new_n7611);
and_8  g07235(new_n7420, new_n7425, new_n7612);
and_8  g07236(new_n7421, new_n7416, new_n7613);
or_8   g07237(new_n7613, new_n7612, new_n7614);
and_8  g07238(new_n7608, new_n7606, new_n7615);
and_8  g07239(new_n7602, new_n7531, new_n7616);
or_8   g07240(new_n7616, new_n7615, new_n7617);
and_8  g07241(new_n7617, new_n7614, new_n7618);
or_8   g07242(new_n7618, new_n7611, new_n7619);
or_8   g07243(new_n7619, new_n7414, new_n7620);
nor_6  g07244(new_n7255, new_n7000, new_n7621);
xor_4  g07245(new_n7255, new_n7000, new_n7622);
or_8   g07246(new_n7411, new_n7407, new_n7623);
and_8  g07247(new_n7623, new_n7622, new_n7624);
or_8   g07248(new_n7624, new_n7621, new_n7625);
or_8   g07249(new_n7617, new_n7614, new_n7626);
or_8   g07250(new_n7610_1, new_n7427, new_n7627);
and_8  g07251(new_n7627, new_n7626, new_n7628);
or_8   g07252(new_n7628, new_n7625, new_n7629);
and_8  g07253(new_n7629, new_n7620, n2383);
xnor_4 g07254(new_n6220, new_n6213, n2425);
xor_4  g07255(new_n3051, new_n2994, n2431);
xnor_4 g07256(new_n2100, new_n2098, n2434);
xor_4  g07257(new_n5171, new_n5170, n2581);
xor_4  g07258(new_n6910, new_n6909, new_n7635);
xor_4  g07259(new_n7635, new_n6922, n2624);
and_8  g07260(n11917, n6770, new_n7637);
and_8  g07261(n9920, n4921, new_n7638);
and_8  g07262(n9956, n3627, new_n7639);
xor_4  g07263(new_n7639, new_n7638, new_n7640);
xor_4  g07264(new_n7640, new_n7637, new_n7641);
or_8   g07265(new_n4166, new_n4135, new_n7642);
or_8   g07266(new_n4167, new_n4165, new_n7643);
and_8  g07267(new_n7643, new_n7642, new_n7644);
xor_4  g07268(new_n7644, new_n7641, new_n7645);
and_8  g07269(n2577, n2564, new_n7646_1);
and_8  g07270(n4189, n3842, new_n7647);
xor_4  g07271(new_n7647, new_n7646_1, new_n7648);
xor_4  g07272(new_n7648, new_n7645, new_n7649);
and_8  g07273(new_n4163, new_n4159_1, new_n7650);
or_8   g07274(new_n4169, new_n7650, new_n7651);
and_8  g07275(new_n7651, new_n7649, new_n7652);
nor_6  g07276(new_n7651, new_n7649, new_n7653);
or_8   g07277(new_n7653, new_n7652, new_n7654);
and_8  g07278(new_n4157, new_n4154, new_n7655);
nor_6  g07279(new_n4171, new_n4158, new_n7656);
or_8   g07280(new_n7656, new_n7655, new_n7657);
not_8  g07281(new_n7657, new_n7658);
or_8   g07282(new_n7658, new_n7654, new_n7659);
and_8  g07283(new_n7639, new_n7638, new_n7660);
and_8  g07284(n6770, n3842, new_n7661);
xor_4  g07285(new_n7661, new_n7660, new_n7662);
and_8  g07286(n4921, n3627, new_n7663);
and_8  g07287(n11917, n9920, new_n7664);
and_8  g07288(n9956, n4516, new_n7665);
xnor_4 g07289(new_n7665, new_n7664, new_n7666);
xor_4  g07290(new_n7666, new_n7663, new_n7667);
xor_4  g07291(new_n7667, new_n7662, new_n7668);
or_8   g07292(new_n7640, new_n7637, new_n7669);
xnor_4 g07293(new_n7640, new_n7637, new_n7670);
or_8   g07294(new_n7644, new_n7670, new_n7671);
and_8  g07295(new_n7671, new_n7669, new_n7672);
and_8  g07296(n9637, n2564, new_n7673);
and_8  g07297(n4189, n2577, new_n7674);
and_8  g07298(n6687, n1835, new_n7675);
xnor_4 g07299(new_n7675, new_n7674, new_n7676_1);
xor_4  g07300(new_n7676_1, new_n7673, new_n7677);
xor_4  g07301(new_n7677, new_n7672, new_n7678);
xor_4  g07302(new_n7678, new_n7668, new_n7679);
nand_5 g07303(new_n7648, new_n7645, new_n7680);
and_8  g07304(new_n7647, new_n7646_1, new_n7681);
and_8  g07305(new_n7652, new_n7681, new_n7682);
nor_6  g07306(new_n7652, new_n7681, new_n7683);
or_8   g07307(new_n7683, new_n7682, new_n7684);
and_8  g07308(new_n7684, new_n7680, new_n7685);
xor_4  g07309(new_n7685, new_n7679, new_n7686);
nor_6  g07310(new_n7686, new_n7659, new_n7687);
and_8  g07311(new_n7686, new_n7659, new_n7688);
or_8   g07312(new_n7688, new_n7687, new_n7689);
nand_5 g07313(n9637, n6687, new_n7690_1);
not_8  g07314(new_n7690_1, new_n7691);
not_8  g07315(new_n7654, new_n7692);
or_8   g07316(new_n7657, new_n7692, new_n7693);
and_8  g07317(new_n7693, new_n7659, new_n7694);
nand_5 g07318(new_n7694, new_n7691, new_n7695);
nand_5 g07319(new_n4172, new_n4153, new_n7696);
xor_4  g07320(new_n7694, new_n7690_1, new_n7697);
or_8   g07321(new_n7697, new_n7696, new_n7698);
and_8  g07322(new_n7698, new_n7695, new_n7699);
xor_4  g07323(new_n7699, new_n7689, new_n7700);
not_8  g07324(new_n7700, new_n7701);
and_8  g07325(n6126, n2226, new_n7702);
and_8  g07326(n3602, n1094, new_n7703);
and_8  g07327(n10678, n3719, new_n7704);
xor_4  g07328(new_n7704, new_n7703, new_n7705);
xor_4  g07329(new_n7705, new_n7702, new_n7706);
or_8   g07330(new_n4359, new_n4180, new_n7707);
or_8   g07331(new_n4360, new_n4358, new_n7708);
and_8  g07332(new_n7708, new_n7707, new_n7709);
xor_4  g07333(new_n7709, new_n7706, new_n7710);
and_8  g07334(n10928, n10439, new_n7711);
and_8  g07335(n8595, n6986, new_n7712);
xor_4  g07336(new_n7712, new_n7711, new_n7713);
xor_4  g07337(new_n7713, new_n7710, new_n7714);
and_8  g07338(new_n4356, new_n4352, new_n7715);
or_8   g07339(new_n4362, new_n7715, new_n7716);
and_8  g07340(new_n7716, new_n7714, new_n7717);
nor_6  g07341(new_n7716, new_n7714, new_n7718);
or_8   g07342(new_n7718, new_n7717, new_n7719);
and_8  g07343(new_n4350, new_n4347, new_n7720);
nor_6  g07344(new_n4364, new_n4351, new_n7721);
or_8   g07345(new_n7721, new_n7720, new_n7722);
not_8  g07346(new_n7722, new_n7723);
or_8   g07347(new_n7723, new_n7719, new_n7724);
or_8   g07348(new_n7705, new_n7702, new_n7725);
xnor_4 g07349(new_n7705, new_n7702, new_n7726);
or_8   g07350(new_n7709, new_n7726, new_n7727);
and_8  g07351(new_n7727, new_n7725, new_n7728);
and_8  g07352(n10928, n8065, new_n7729);
and_8  g07353(n10439, n6986, new_n7730_1);
and_8  g07354(n10391, n8336, new_n7731);
xnor_4 g07355(new_n7731, new_n7730_1, new_n7732);
xor_4  g07356(new_n7732, new_n7729, new_n7733_1);
xor_4  g07357(new_n7733_1, new_n7728, new_n7734);
and_8  g07358(new_n7704, new_n7703, new_n7735);
and_8  g07359(n8595, n2226, new_n7736);
xnor_4 g07360(new_n7736, new_n7735, new_n7737);
and_8  g07361(n10678, n3602, new_n7738);
and_8  g07362(n6126, n1094, new_n7739);
and_8  g07363(n7320, n3719, new_n7740);
xnor_4 g07364(new_n7740, new_n7739, new_n7741);
xor_4  g07365(new_n7741, new_n7738, new_n7742);
xor_4  g07366(new_n7742, new_n7737, new_n7743);
xor_4  g07367(new_n7743, new_n7734, new_n7744);
nand_5 g07368(new_n7713, new_n7710, new_n7745);
and_8  g07369(new_n7712, new_n7711, new_n7746);
and_8  g07370(new_n7717, new_n7746, new_n7747);
nor_6  g07371(new_n7717, new_n7746, new_n7748);
or_8   g07372(new_n7748, new_n7747, new_n7749);
and_8  g07373(new_n7749, new_n7745, new_n7750);
or_8   g07374(new_n7750, new_n7744, new_n7751);
not_8  g07375(new_n7751, new_n7752);
and_8  g07376(new_n7750, new_n7744, new_n7753);
or_8   g07377(new_n7753, new_n7752, new_n7754);
nor_6  g07378(new_n7754, new_n7724, new_n7755);
and_8  g07379(new_n7754, new_n7724, new_n7756);
or_8   g07380(new_n7756, new_n7755, new_n7757);
and_8  g07381(n8336, n8065, new_n7758);
xor_4  g07382(new_n7723, new_n7719, new_n7759);
nor_6  g07383(new_n7759, new_n7758, new_n7760);
not_8  g07384(new_n7760, new_n7761);
nand_5 g07385(new_n4365, new_n4346, new_n7762);
not_8  g07386(new_n7762, new_n7763);
and_8  g07387(new_n7759, new_n7758, new_n7764);
or_8   g07388(new_n7764, new_n7760, new_n7765);
or_8   g07389(new_n7765, new_n7763, new_n7766);
and_8  g07390(new_n7766, new_n7761, new_n7767);
xor_4  g07391(new_n7767, new_n7757, new_n7768);
and_8  g07392(n7160, n4826, new_n7769);
and_8  g07393(n7733, n4828, new_n7770);
and_8  g07394(n12925, n2515, new_n7771);
xor_4  g07395(new_n7771, new_n7770, new_n7772);
xor_4  g07396(new_n7772, new_n7769, new_n7773);
or_8   g07397(new_n4406, new_n4205, new_n7774);
or_8   g07398(new_n4407, new_n4405, new_n7775);
and_8  g07399(new_n7775, new_n7774, new_n7776);
and_8  g07400(new_n7776, new_n7773, new_n7777);
nor_6  g07401(new_n7776, new_n7773, new_n7778);
or_8   g07402(new_n7778, new_n7777, new_n7779);
and_8  g07403(n12391, n4970, new_n7780);
and_8  g07404(n7891, n7610, new_n7781);
xor_4  g07405(new_n7781, new_n7780, new_n7782);
not_8  g07406(new_n7782, new_n7783);
or_8   g07407(new_n7783, new_n7779, new_n7784);
xor_4  g07408(new_n7776, new_n7773, new_n7785);
or_8   g07409(new_n7782, new_n7785, new_n7786);
and_8  g07410(new_n7786, new_n7784, new_n7787);
or_8   g07411(new_n4411, new_n4412, new_n7788);
and_8  g07412(new_n7788, new_n7787, new_n7789);
nor_6  g07413(new_n7788, new_n7787, new_n7790);
or_8   g07414(new_n7790, new_n7789, new_n7791);
or_8   g07415(new_n4417, new_n4399, new_n7792);
not_8  g07416(new_n4423, new_n7793);
or_8   g07417(new_n7793, new_n4420, new_n7794);
and_8  g07418(new_n7794, new_n7792, new_n7795);
or_8   g07419(new_n7795, new_n7791, new_n7796);
and_8  g07420(new_n7772, new_n7769, new_n7797);
or_8   g07421(new_n7777, new_n7797, new_n7798);
and_8  g07422(n12391, n503, new_n7799);
and_8  g07423(n7891, n4970, new_n7800);
and_8  g07424(n12069, n10965, new_n7801);
xnor_4 g07425(new_n7801, new_n7800, new_n7802);
xor_4  g07426(new_n7802, new_n7799, new_n7803);
xor_4  g07427(new_n7803, new_n7798, new_n7804);
and_8  g07428(new_n7771, new_n7770, new_n7805);
and_8  g07429(n7610, n7160, new_n7806);
xnor_4 g07430(new_n7806, new_n7805, new_n7807);
and_8  g07431(n7733, n2515, new_n7808);
and_8  g07432(n4828, n4826, new_n7809);
and_8  g07433(n12925, n1199, new_n7810);
xnor_4 g07434(new_n7810, new_n7809, new_n7811);
xor_4  g07435(new_n7811, new_n7808, new_n7812);
xor_4  g07436(new_n7812, new_n7807, new_n7813);
xor_4  g07437(new_n7813, new_n7804, new_n7814);
and_8  g07438(new_n7781, new_n7780, new_n7815);
and_8  g07439(new_n7789, new_n7815, new_n7816);
nor_6  g07440(new_n7789, new_n7815, new_n7817);
or_8   g07441(new_n7817, new_n7816, new_n7818);
and_8  g07442(new_n7818, new_n7784, new_n7819);
or_8   g07443(new_n7819, new_n7814, new_n7820);
not_8  g07444(new_n7820, new_n7821);
and_8  g07445(new_n7819, new_n7814, new_n7822);
or_8   g07446(new_n7822, new_n7821, new_n7823_1);
or_8   g07447(new_n7823_1, new_n7796, new_n7824);
xor_4  g07448(new_n7788, new_n7787, new_n7825);
xor_4  g07449(new_n4417, new_n4399, new_n7826);
and_8  g07450(new_n4423, new_n7826, new_n7827);
or_8   g07451(new_n7827, new_n4418, new_n7828);
and_8  g07452(new_n7828, new_n7825, new_n7829);
not_8  g07453(new_n7822, new_n7830);
and_8  g07454(new_n7830, new_n7820, new_n7831);
or_8   g07455(new_n7831, new_n7829, new_n7832);
and_8  g07456(new_n7832, new_n7824, new_n7833);
nand_5 g07457(n12069, n503, new_n7834);
not_8  g07458(new_n7834, new_n7835);
or_8   g07459(new_n7828, new_n7825, new_n7836);
and_8  g07460(new_n7836, new_n7796, new_n7837);
and_8  g07461(new_n7837, new_n7835, new_n7838);
and_8  g07462(new_n7795, new_n7791, new_n7839);
or_8   g07463(new_n7839, new_n7829, new_n7840);
or_8   g07464(new_n7840, new_n7834, new_n7841);
or_8   g07465(new_n7837, new_n7835, new_n7842);
and_8  g07466(new_n7842, new_n7841, new_n7843);
and_8  g07467(new_n7843, new_n4425, new_n7844);
or_8   g07468(new_n7844, new_n7838, new_n7845);
xor_4  g07469(new_n7845, new_n7833, new_n7846);
nand_5 g07470(n11222, n6359, new_n7847);
not_8  g07471(new_n7847, new_n7848);
and_8  g07472(n4086, n996, new_n7849);
not_8  g07473(new_n7849, new_n7850);
and_8  g07474(n5767, n405, new_n7851);
and_8  g07475(n8433, n5319, new_n7852);
xor_4  g07476(new_n7852, new_n7851, new_n7853);
xor_4  g07477(new_n7853, new_n7850, new_n7854);
or_8   g07478(new_n4372, new_n4371, new_n7855);
and_8  g07479(new_n4372, new_n4371, new_n7856);
or_8   g07480(new_n7856, new_n4370_1, new_n7857);
and_8  g07481(new_n7857, new_n7855, new_n7858);
xor_4  g07482(new_n7858, new_n7854, new_n7859);
and_8  g07483(n11153, n6611, new_n7860);
and_8  g07484(n5314, n217, new_n7861);
xor_4  g07485(new_n7861, new_n7860, new_n7862_1);
not_8  g07486(new_n7862_1, new_n7863);
or_8   g07487(new_n7863, new_n7859, new_n7864);
nand_5 g07488(new_n7857, new_n7855, new_n7865);
xor_4  g07489(new_n7865, new_n7854, new_n7866);
or_8   g07490(new_n7862_1, new_n7866, new_n7867);
and_8  g07491(new_n7867, new_n7864, new_n7868);
and_8  g07492(new_n4387, new_n4386, new_n7869);
or_8   g07493(new_n7869, new_n4375, new_n7870);
and_8  g07494(new_n7870, new_n7868, new_n7871);
nor_6  g07495(new_n7870, new_n7868, new_n7872);
or_8   g07496(new_n7872, new_n7871, new_n7873);
not_8  g07497(new_n4367, new_n7874);
xor_4  g07498(new_n4387, new_n4380, new_n7875);
or_8   g07499(new_n7875, new_n7874, new_n7876);
xor_4  g07500(new_n4389, new_n7874, new_n7877);
not_8  g07501(new_n4393, new_n7878);
or_8   g07502(new_n7878, new_n7877, new_n7879);
and_8  g07503(new_n7879, new_n7876, new_n7880);
or_8   g07504(new_n7880, new_n7873, new_n7881);
xor_4  g07505(new_n7870, new_n7868, new_n7882);
not_8  g07506(new_n7876, new_n7883);
and_8  g07507(new_n4393, new_n4390, new_n7884);
or_8   g07508(new_n7884, new_n7883, new_n7885);
or_8   g07509(new_n7885, new_n7882, new_n7886);
and_8  g07510(new_n7886, new_n7881, new_n7887);
and_8  g07511(new_n7887, new_n7848, new_n7888);
and_8  g07512(new_n4394, new_n4250, new_n7889);
and_8  g07513(new_n7885, new_n7882, new_n7890);
and_8  g07514(new_n7880, new_n7873, new_n7891_1);
or_8   g07515(new_n7891_1, new_n7890, new_n7892);
or_8   g07516(new_n7892, new_n7847, new_n7893);
or_8   g07517(new_n7887, new_n7848, new_n7894);
and_8  g07518(new_n7894, new_n7893, new_n7895);
and_8  g07519(new_n7895, new_n7889, new_n7896);
or_8   g07520(new_n7896, new_n7888, new_n7897);
and_8  g07521(new_n7852, new_n7851, new_n7898);
and_8  g07522(n996, n217, new_n7899);
xnor_4 g07523(new_n7899, new_n7898, new_n7900);
and_8  g07524(n5319, n405, new_n7901);
and_8  g07525(n5767, n4086, new_n7902);
and_8  g07526(n9457, n8433, new_n7903);
xnor_4 g07527(new_n7903, new_n7902, new_n7904);
xor_4  g07528(new_n7904, new_n7901, new_n7905);
nor_6  g07529(new_n7905, new_n7900, new_n7906);
and_8  g07530(new_n7905, new_n7900, new_n7907);
or_8   g07531(new_n7907, new_n7906, new_n7908);
and_8  g07532(n11153, n6359, new_n7909);
and_8  g07533(n6611, n5314, new_n7910);
and_8  g07534(n11296, n11222, new_n7911);
xnor_4 g07535(new_n7911, new_n7910, new_n7912);
xor_4  g07536(new_n7912, new_n7909, new_n7913);
nand_5 g07537(new_n7853, new_n7849, new_n7914);
or_8   g07538(new_n7865, new_n7854, new_n7915);
and_8  g07539(new_n7915, new_n7914, new_n7916);
xor_4  g07540(new_n7916, new_n7913, new_n7917);
xor_4  g07541(new_n7917, new_n7908, new_n7918);
not_8  g07542(new_n7918, new_n7919);
not_8  g07543(new_n7864, new_n7920);
and_8  g07544(new_n7861, new_n7860, new_n7921);
xor_4  g07545(new_n7871, new_n7921, new_n7922);
or_8   g07546(new_n7922, new_n7920, new_n7923);
and_8  g07547(new_n7923, new_n7919, new_n7924);
nor_6  g07548(new_n7922, new_n7920, new_n7925);
and_8  g07549(new_n7925, new_n7918, new_n7926);
or_8   g07550(new_n7926, new_n7924, new_n7927);
or_8   g07551(new_n7927, new_n7881, new_n7928);
or_8   g07552(new_n7925, new_n7918, new_n7929);
or_8   g07553(new_n7923, new_n7919, new_n7930);
and_8  g07554(new_n7930, new_n7929, new_n7931);
or_8   g07555(new_n7931, new_n7890, new_n7932);
and_8  g07556(new_n7932, new_n7928, new_n7933);
xor_4  g07557(new_n7933, new_n7897, new_n7934);
or_8   g07558(new_n7934, new_n7846, new_n7935);
and_8  g07559(new_n7845, new_n7833, new_n7936);
nor_6  g07560(new_n7845, new_n7833, new_n7937);
or_8   g07561(new_n7937, new_n7936, new_n7938);
and_8  g07562(new_n7933, new_n7897, new_n7939);
nor_6  g07563(new_n7933, new_n7897, new_n7940);
or_8   g07564(new_n7940, new_n7939, new_n7941);
or_8   g07565(new_n7941, new_n7938, new_n7942);
and_8  g07566(new_n7942, new_n7935, new_n7943);
nor_6  g07567(new_n7843, new_n4425, new_n7944);
or_8   g07568(new_n7944, new_n7844, new_n7945);
not_8  g07569(new_n7889, new_n7946_1);
xor_4  g07570(new_n7895, new_n7946_1, new_n7947);
and_8  g07571(new_n7947, new_n7945, new_n7948);
nor_6  g07572(new_n4431, new_n4395, new_n7949);
or_8   g07573(new_n7949, new_n4430, new_n7950);
xor_4  g07574(new_n7843, new_n4425, new_n7951);
xor_4  g07575(new_n7895, new_n7889, new_n7952);
or_8   g07576(new_n7952, new_n7951, new_n7953);
or_8   g07577(new_n7947, new_n7945, new_n7954);
and_8  g07578(new_n7954, new_n7953, new_n7955);
and_8  g07579(new_n7955, new_n7950, new_n7956);
or_8   g07580(new_n7956, new_n7948, new_n7957);
xor_4  g07581(new_n7957, new_n7943, new_n7958);
and_8  g07582(new_n7958, new_n7768, new_n7959);
xor_4  g07583(new_n7754, new_n7724, new_n7960);
xor_4  g07584(new_n7767, new_n7960, new_n7961);
and_8  g07585(new_n7941, new_n7938, new_n7962);
and_8  g07586(new_n7934, new_n7846, new_n7963);
or_8   g07587(new_n7963, new_n7962, new_n7964);
xor_4  g07588(new_n7957, new_n7964, new_n7965_1);
and_8  g07589(new_n7965_1, new_n7961, new_n7966_1);
or_8   g07590(new_n7966_1, new_n7959, new_n7967);
xor_4  g07591(new_n7765, new_n7762, new_n7968);
nor_6  g07592(new_n7949, new_n4430, new_n7969);
and_8  g07593(new_n7952, new_n7951, new_n7970);
or_8   g07594(new_n7970, new_n7948, new_n7971);
and_8  g07595(new_n7971, new_n7969, new_n7972);
or_8   g07596(new_n7972, new_n7956, new_n7973);
or_8   g07597(new_n7973, new_n7968, new_n7974);
not_8  g07598(new_n7968, new_n7975);
or_8   g07599(new_n7971, new_n7969, new_n7976);
or_8   g07600(new_n7955, new_n7950, new_n7977);
and_8  g07601(new_n7977, new_n7976, new_n7978);
and_8  g07602(new_n7978, new_n7975, new_n7979);
and_8  g07603(new_n7973, new_n7968, new_n7980);
or_8   g07604(new_n7980, new_n7979, new_n7981_1);
or_8   g07605(new_n4432, new_n4437, new_n7982);
not_8  g07606(new_n7982, new_n7983);
or_8   g07607(new_n4439, new_n7983, new_n7984);
or_8   g07608(new_n7984, new_n7981_1, new_n7985);
and_8  g07609(new_n7985, new_n7974, new_n7986);
xor_4  g07610(new_n7986, new_n7967, new_n7987);
or_8   g07611(new_n7987, new_n7701, new_n7988);
xor_4  g07612(new_n7697, new_n7696, new_n7989);
not_8  g07613(new_n7989, new_n7990);
nor_6  g07614(new_n4342, new_n4335, new_n7991);
or_8   g07615(new_n7991, new_n4340, new_n7992);
or_8   g07616(new_n7992, new_n4173, new_n7993);
or_8   g07617(new_n4440, new_n4345, new_n7994);
and_8  g07618(new_n7994, new_n7993, new_n7995);
and_8  g07619(new_n7995, new_n7990, new_n7996);
nor_6  g07620(new_n7980, new_n7979, new_n7997);
or_8   g07621(new_n4435, new_n4433, new_n7998);
and_8  g07622(new_n7998, new_n7982, new_n7999);
xor_4  g07623(new_n7999, new_n7997, new_n8000);
xor_4  g07624(new_n7995, new_n7990, new_n8001);
and_8  g07625(new_n8001, new_n8000, new_n8002);
or_8   g07626(new_n8002, new_n7996, new_n8003);
or_8   g07627(new_n7965_1, new_n7961, new_n8004);
or_8   g07628(new_n7958, new_n7768, new_n8005);
and_8  g07629(new_n8005, new_n8004, new_n8006);
xor_4  g07630(new_n7986, new_n8006, new_n8007);
and_8  g07631(new_n8007, new_n7700, new_n8008);
and_8  g07632(new_n7987, new_n7701, new_n8009);
or_8   g07633(new_n8009, new_n8008, new_n8010);
or_8   g07634(new_n8010, new_n8003, new_n8011);
and_8  g07635(new_n8011, new_n7988, new_n8012);
or_8   g07636(new_n7821, new_n7816, new_n8013);
nand_5 g07637(new_n7806, new_n7805, new_n8014);
or_8   g07638(new_n7812, new_n7807, new_n8015);
nand_5 g07639(new_n8015, new_n8014, new_n8016);
or_8   g07640(new_n7675, new_n7674, new_n8017);
or_8   g07641(new_n7676_1, new_n7673, new_n8018);
and_8  g07642(new_n8018, new_n8017, new_n8019);
not_8  g07643(n2577, new_n8020);
not_8  g07644(n6770, new_n8021);
or_8   g07645(new_n8021, new_n8020, new_n8022);
xor_4  g07646(new_n8022, new_n8019, new_n8023);
and_8  g07647(n9637, n4189, new_n8024);
and_8  g07648(n11917, n3627, new_n8025);
xor_4  g07649(new_n8025, new_n8024, new_n8026);
not_8  g07650(new_n8026, new_n8027);
xor_4  g07651(new_n8027, new_n8023, new_n8028_1);
or_8   g07652(new_n7801, new_n7800, new_n8029);
or_8   g07653(new_n7802, new_n7799, new_n8030);
nand_5 g07654(new_n8030, new_n8029, new_n8031);
nor_6  g07655(new_n7661, new_n7660, new_n8032);
and_8  g07656(new_n7667, new_n7662, new_n8033);
or_8   g07657(new_n8033, new_n8032, new_n8034);
xor_4  g07658(new_n8034, new_n8031, new_n8035);
xor_4  g07659(new_n8035, new_n8028_1, new_n8036);
xor_4  g07660(new_n8036, new_n8016, new_n8037);
not_8  g07661(new_n7798, new_n8038);
nand_5 g07662(new_n7803, new_n8038, new_n8039);
or_8   g07663(new_n7813, new_n7804, new_n8040);
and_8  g07664(new_n8040, new_n8039, new_n8041);
or_8   g07665(new_n7740, new_n7739, new_n8042);
or_8   g07666(new_n7741, new_n7738, new_n8043);
and_8  g07667(new_n8043, new_n8042, new_n8044);
and_8  g07668(n7523, n3719, new_n8045);
and_8  g07669(n11222, n1357, new_n8046);
xor_4  g07670(new_n8046, new_n8045, new_n8047);
and_8  g07671(n8336, n4190, new_n8048);
and_8  g07672(n7320, n3602, new_n8049);
xnor_4 g07673(new_n8049, new_n8048, new_n8050);
xor_4  g07674(new_n8050, new_n8047, new_n8051);
xor_4  g07675(new_n8051, new_n8044, new_n8052);
xor_4  g07676(new_n8052, new_n8041, new_n8053);
or_8   g07677(new_n8053, new_n8037, new_n8054);
not_8  g07678(new_n8016, new_n8055);
xor_4  g07679(new_n8036, new_n8055, new_n8056);
not_8  g07680(new_n8053, new_n8057);
or_8   g07681(new_n8057, new_n8056, new_n8058);
and_8  g07682(new_n8058, new_n8054, new_n8059);
not_8  g07683(new_n7679, new_n8060);
nor_6  g07684(new_n7685, new_n8060, new_n8061);
or_8   g07685(new_n8061, new_n7682, new_n8062);
or_8   g07686(new_n7752, new_n7747, new_n8063);
or_8   g07687(new_n8063, new_n8062, new_n8064);
nor_6  g07688(new_n8061, new_n7682, new_n8065_1);
nor_6  g07689(new_n7752, new_n7747, new_n8066);
or_8   g07690(new_n8066, new_n8065_1, new_n8067);
and_8  g07691(new_n8067, new_n8064, new_n8068);
xor_4  g07692(new_n8068, new_n8059, new_n8069);
and_8  g07693(new_n8069, new_n8013, new_n8070);
not_8  g07694(new_n8013, new_n8071);
and_8  g07695(new_n8068, new_n8059, new_n8072);
nor_6  g07696(new_n8068, new_n8059, new_n8073);
or_8   g07697(new_n8073, new_n8072, new_n8074);
and_8  g07698(new_n8074, new_n8071, new_n8075);
or_8   g07699(new_n8075, new_n8070, new_n8076);
or_8   g07700(new_n7754, new_n7724, new_n8077);
xor_4  g07701(new_n7759, new_n7758, new_n8078);
and_8  g07702(new_n8078, new_n7762, new_n8079);
or_8   g07703(new_n8079, new_n7760, new_n8080);
or_8   g07704(new_n8080, new_n7757, new_n8081);
and_8  g07705(new_n8081, new_n8077, new_n8082);
or_8   g07706(new_n7731, new_n7730_1, new_n8083);
or_8   g07707(new_n7732, new_n7729, new_n8084);
and_8  g07708(new_n8084, new_n8083, new_n8085);
and_8  g07709(n5319, n4086, new_n8086);
and_8  g07710(n10928, n10391, new_n8087);
xor_4  g07711(new_n8087, new_n8086, new_n8088);
xor_4  g07712(new_n8088, new_n8085, new_n8089);
or_8   g07713(new_n8089, new_n8082, new_n8090);
and_8  g07714(new_n7767, new_n7960, new_n8091);
or_8   g07715(new_n8091, new_n7755, new_n8092);
not_8  g07716(new_n8089, new_n8093);
or_8   g07717(new_n8093, new_n8092, new_n8094);
and_8  g07718(new_n8094, new_n8090, new_n8095);
and_8  g07719(new_n8095, new_n8076, new_n8096);
or_8   g07720(new_n8074, new_n8071, new_n8097);
or_8   g07721(new_n8069, new_n8013, new_n8098);
and_8  g07722(new_n8098, new_n8097, new_n8099);
and_8  g07723(new_n8093, new_n8092, new_n8100_1);
and_8  g07724(new_n8089, new_n8082, new_n8101);
or_8   g07725(new_n8101, new_n8100_1, new_n8102);
and_8  g07726(new_n8102, new_n8099, new_n8103);
or_8   g07727(new_n8103, new_n8096, new_n8104);
and_8  g07728(new_n7831, new_n7829, new_n8105);
or_8   g07729(new_n7936, new_n8105, new_n8106);
not_8  g07730(new_n7928, new_n8107);
or_8   g07731(new_n7939, new_n8107, new_n8108);
xor_4  g07732(new_n8108, new_n8106, new_n8109);
not_8  g07733(new_n8109, new_n8110);
xor_4  g07734(new_n8110, new_n8104, new_n8111);
and_8  g07735(n4826, n2515, new_n8112);
and_8  g07736(n12925, n6578, new_n8113);
xor_4  g07737(new_n8113, new_n8112, new_n8114);
and_8  g07738(n6359, n5314, new_n8115);
and_8  g07739(n12069, n7546, new_n8116);
xor_4  g07740(new_n8116, new_n8115, new_n8117);
xor_4  g07741(new_n8117, new_n8114, new_n8118);
or_8   g07742(new_n7903, new_n7902, new_n8119);
or_8   g07743(new_n7904, new_n7901, new_n8120);
nand_5 g07744(new_n8120, new_n8119, new_n8121);
or_8   g07745(new_n7912, new_n7909, new_n8122);
and_8  g07746(new_n8122, new_n7910, new_n8123);
and_8  g07747(n11296, n11153, new_n8124);
nand_5 g07748(new_n8124, new_n8123, new_n8125);
and_8  g07749(new_n8124, new_n7847, new_n8126);
or_8   g07750(new_n8126, new_n8123, new_n8127);
and_8  g07751(new_n8127, new_n8125, new_n8128);
xor_4  g07752(new_n8128, new_n8121, new_n8129);
xor_4  g07753(new_n8129, new_n8118, new_n8130);
and_8  g07754(new_n8130, new_n8111, new_n8131);
xor_4  g07755(new_n8109, new_n8104, new_n8132);
not_8  g07756(new_n8130, new_n8133);
and_8  g07757(new_n8133, new_n8132, new_n8134);
or_8   g07758(new_n8134, new_n8131, new_n8135);
and_8  g07759(new_n7999, new_n7997, new_n8136);
or_8   g07760(new_n8136, new_n7979, new_n8137);
and_8  g07761(new_n8137, new_n8006, new_n8138_1);
or_8   g07762(new_n8138_1, new_n7959, new_n8139);
and_8  g07763(new_n7976, new_n7953, new_n8140);
or_8   g07764(new_n8140, new_n7964, new_n8141);
and_8  g07765(new_n8141, new_n7935, new_n8142);
not_8  g07766(new_n7687, new_n8143);
or_8   g07767(new_n7699, new_n7689, new_n8144);
and_8  g07768(new_n8144, new_n8143, new_n8145);
nand_5 g07769(new_n7871, new_n7921, new_n8146);
and_8  g07770(new_n7929, new_n8146, new_n8147);
not_8  g07771(new_n7672, new_n8148);
or_8   g07772(new_n7677, new_n8148, new_n8149);
or_8   g07773(new_n7678, new_n7668, new_n8150);
and_8  g07774(new_n8150, new_n8149, new_n8151);
not_8  g07775(new_n7733_1, new_n8152);
or_8   g07776(new_n8152, new_n7728, new_n8153);
or_8   g07777(new_n7743, new_n7734, new_n8154);
and_8  g07778(new_n8154, new_n8153, new_n8155);
xor_4  g07779(new_n8155, new_n8151, new_n8156);
not_8  g07780(new_n8156, new_n8157);
and_8  g07781(new_n7899, new_n7898, new_n8158);
or_8   g07782(new_n7906, new_n8158, new_n8159);
and_8  g07783(n8595, n1094, new_n8160);
and_8  g07784(n2564, n1835, new_n8161);
xor_4  g07785(new_n8161, new_n8160, new_n8162);
xor_4  g07786(new_n8162, new_n8159, new_n8163);
or_8   g07787(new_n7810, new_n7809, new_n8164);
or_8   g07788(new_n7811, new_n7808, new_n8165);
and_8  g07789(new_n8165, new_n8164, new_n8166);
nand_5 g07790(n12391, n10965, new_n8167);
and_8  g07791(n7891, n503, new_n8168);
and_8  g07792(n9457, n405, new_n8169);
xor_4  g07793(new_n8169, new_n8168, new_n8170);
xor_4  g07794(new_n8170, new_n8167, new_n8171);
xor_4  g07795(new_n8171, new_n8166, new_n8172);
and_8  g07796(n8065, n6986, new_n8173);
and_8  g07797(n10439, n2226, new_n8174);
xor_4  g07798(new_n8174, new_n8173, new_n8175);
xor_4  g07799(new_n8175, new_n8172, new_n8176);
xor_4  g07800(new_n8176, new_n8163, new_n8177);
or_8   g07801(new_n7665, new_n7664, new_n8178);
or_8   g07802(new_n7666, new_n7663, new_n8179);
and_8  g07803(new_n8179, new_n8178, new_n8180);
and_8  g07804(n11536, n6687, new_n8181);
and_8  g07805(n6611, n996, new_n8182);
xor_4  g07806(new_n8182, new_n8181, new_n8183);
and_8  g07807(n4921, n4516, new_n8184);
and_8  g07808(n9920, n3842, new_n8185);
xor_4  g07809(new_n8185, new_n8184, new_n8186);
xor_4  g07810(new_n8186, new_n8183, new_n8187);
xor_4  g07811(new_n8187, new_n8180, new_n8188);
nand_5 g07812(n9956, n2087, new_n8189);
and_8  g07813(n7733, n1199, new_n8190);
and_8  g07814(n5767, n217, new_n8191);
xor_4  g07815(new_n8191, new_n8190, new_n8192);
and_8  g07816(n7160, n4970, new_n8193);
and_8  g07817(n7610, n4828, new_n8194);
xor_4  g07818(new_n8194, new_n8193, new_n8195);
xor_4  g07819(new_n8195, new_n8192, new_n8196);
xor_4  g07820(new_n8196, new_n8189, new_n8197);
xor_4  g07821(new_n8197, new_n8188, new_n8198);
and_8  g07822(new_n7736, new_n7735, new_n8199);
nor_6  g07823(new_n7742, new_n7737, new_n8200);
or_8   g07824(new_n8200, new_n8199, new_n8201);
and_8  g07825(n8433, n4817, new_n8202_1);
and_8  g07826(n10678, n6126, new_n8203);
xor_4  g07827(new_n8203, new_n8202_1, new_n8204);
not_8  g07828(new_n8204, new_n8205);
xor_4  g07829(new_n8205, new_n8201, new_n8206);
xor_4  g07830(new_n8206, new_n8198, new_n8207);
xor_4  g07831(new_n8207, new_n8177, new_n8208);
xor_4  g07832(new_n8208, new_n8157, new_n8209);
and_8  g07833(new_n8209, new_n8147, new_n8210);
not_8  g07834(new_n8147, new_n8211);
xor_4  g07835(new_n8208, new_n8156, new_n8212);
and_8  g07836(new_n8212, new_n8211, new_n8213);
or_8   g07837(new_n8213, new_n8210, new_n8214);
or_8   g07838(new_n8214, new_n8145, new_n8215);
nor_6  g07839(new_n7699, new_n7689, new_n8216);
or_8   g07840(new_n8216, new_n7687, new_n8217);
or_8   g07841(new_n8212, new_n8211, new_n8218);
or_8   g07842(new_n8209, new_n8147, new_n8219);
and_8  g07843(new_n8219, new_n8218, new_n8220);
or_8   g07844(new_n8220, new_n8217, new_n8221);
and_8  g07845(new_n8221, new_n8215, new_n8222);
and_8  g07846(new_n8222, new_n8142, new_n8223);
and_8  g07847(new_n7957, new_n7943, new_n8224);
or_8   g07848(new_n8224, new_n7962, new_n8225);
and_8  g07849(new_n8220, new_n8217, new_n8226);
and_8  g07850(new_n8214, new_n8145, new_n8227);
or_8   g07851(new_n8227, new_n8226, new_n8228);
and_8  g07852(new_n8228, new_n8225, new_n8229);
or_8   g07853(new_n8229, new_n8223, new_n8230);
and_8  g07854(new_n7916, new_n7913, new_n8231);
and_8  g07855(new_n7917, new_n7908, new_n8232);
or_8   g07856(new_n8232, new_n8231, new_n8233);
xor_4  g07857(new_n8233, new_n8230, new_n8234);
or_8   g07858(new_n8234, new_n8139, new_n8235);
or_8   g07859(new_n7986, new_n7967, new_n8236_1);
and_8  g07860(new_n8236_1, new_n8004, new_n8237);
not_8  g07861(new_n8233, new_n8238);
xor_4  g07862(new_n8238, new_n8230, new_n8239);
or_8   g07863(new_n8239, new_n8237, new_n8240);
and_8  g07864(new_n8240, new_n8235, new_n8241);
xor_4  g07865(new_n8241, new_n8135, new_n8242);
and_8  g07866(new_n8242, new_n8012, new_n8243);
nor_6  g07867(new_n7992, new_n4173, new_n8244);
nor_6  g07868(new_n4440, new_n4345, new_n8245);
or_8   g07869(new_n8245, new_n8244, new_n8246);
or_8   g07870(new_n8246, new_n7989, new_n8247);
xor_4  g07871(new_n7999, new_n7981_1, new_n8248);
xor_4  g07872(new_n7995, new_n7989, new_n8249);
or_8   g07873(new_n8249, new_n8248, new_n8250);
and_8  g07874(new_n8250, new_n8247, new_n8251);
or_8   g07875(new_n8007, new_n7700, new_n8252);
and_8  g07876(new_n8252, new_n7988, new_n8253);
and_8  g07877(new_n8253, new_n8251, new_n8254);
or_8   g07878(new_n8254, new_n8008, new_n8255);
or_8   g07879(new_n8133, new_n8132, new_n8256);
or_8   g07880(new_n8130, new_n8111, new_n8257);
and_8  g07881(new_n8257, new_n8256, new_n8258);
xor_4  g07882(new_n8241, new_n8258, new_n8259);
and_8  g07883(new_n8259, new_n8255, new_n8260);
or_8   g07884(new_n8260, new_n8243, n2679);
nand_5 g07885(new_n5961, new_n5945, new_n8262);
and_8  g07886(n6687, n2253, new_n8263);
and_8  g07887(n10223, n6770, new_n8264);
and_8  g07888(n9920, n2879, new_n8265);
and_8  g07889(n7265, n3627, new_n8266);
xor_4  g07890(new_n8266, new_n8265, new_n8267);
xor_4  g07891(new_n8267, new_n8264, new_n8268);
nor_6  g07892(new_n5949, new_n5924, new_n8269);
not_8  g07893(new_n5948, new_n8270);
and_8  g07894(new_n5950, new_n8270, new_n8271);
or_8   g07895(new_n8271, new_n8269, new_n8272);
xor_4  g07896(new_n8272, new_n8268, new_n8273);
and_8  g07897(n9195, n2564, new_n8274);
and_8  g07898(n4634, n4189, new_n8275);
xor_4  g07899(new_n8275, new_n8274, new_n8276_1);
not_8  g07900(new_n8276_1, new_n8277);
or_8   g07901(new_n8277, new_n8273, new_n8278);
not_8  g07902(new_n8264, new_n8279);
xor_4  g07903(new_n8267, new_n8279, new_n8280);
xor_4  g07904(new_n8272, new_n8280, new_n8281);
or_8   g07905(new_n8276_1, new_n8281, new_n8282);
and_8  g07906(new_n8282, new_n8278, new_n8283);
and_8  g07907(new_n5951, new_n5947, new_n8284);
and_8  g07908(new_n5955, new_n5952, new_n8285);
or_8   g07909(new_n8285, new_n8284, new_n8286);
xor_4  g07910(new_n8286, new_n8283, new_n8287);
and_8  g07911(new_n5956, new_n5946, new_n8288);
and_8  g07912(new_n5960, new_n5957, new_n8289);
or_8   g07913(new_n8289, new_n8288, new_n8290);
xor_4  g07914(new_n8290, new_n8287, new_n8291);
xor_4  g07915(new_n8291, new_n8263, new_n8292);
xnor_4 g07916(new_n8292, new_n8262, new_n8293);
or_8   g07917(new_n6197, new_n5962, new_n8294);
or_8   g07918(new_n6226, new_n6199, new_n8295);
and_8  g07919(new_n8295, new_n8294, new_n8296);
xor_4  g07920(new_n8296, new_n8293, new_n8297);
and_8  g07921(new_n6006, new_n5987, new_n8298);
nand_5 g07922(n12221, n8336, new_n8299);
not_8  g07923(new_n8299, new_n8300);
and_8  g07924(n9189, n2226, new_n8301);
and_8  g07925(n2024, n1094, new_n8302);
and_8  g07926(n10678, n7946, new_n8303_1);
xor_4  g07927(new_n8303_1, new_n8302, new_n8304);
and_8  g07928(new_n8304, new_n8301, new_n8305);
nor_6  g07929(new_n8304, new_n8301, new_n8306);
or_8   g07930(new_n8306, new_n8305, new_n8307);
nor_6  g07931(new_n5996, new_n5968, new_n8308);
not_8  g07932(new_n5995, new_n8309);
and_8  g07933(new_n5997, new_n8309, new_n8310);
or_8   g07934(new_n8310, new_n8308, new_n8311);
nor_6  g07935(new_n8311, new_n8307, new_n8312);
and_8  g07936(new_n8311, new_n8307, new_n8313);
or_8   g07937(new_n8313, new_n8312, new_n8314);
and_8  g07938(n12145, n10928, new_n8315);
and_8  g07939(n6986, n2522, new_n8316);
xor_4  g07940(new_n8316, new_n8315, new_n8317);
not_8  g07941(new_n8317, new_n8318);
or_8   g07942(new_n8318, new_n8314, new_n8319);
xor_4  g07943(new_n8311, new_n8307, new_n8320);
or_8   g07944(new_n8317, new_n8320, new_n8321);
and_8  g07945(new_n8321, new_n8319, new_n8322);
and_8  g07946(new_n5993, new_n5989, new_n8323);
or_8   g07947(new_n5999, new_n8323, new_n8324);
and_8  g07948(new_n8324, new_n8322, new_n8325);
nor_6  g07949(new_n8324, new_n8322, new_n8326);
or_8   g07950(new_n8326, new_n8325, new_n8327);
or_8   g07951(new_n6001, new_n5988, new_n8328);
not_8  g07952(new_n5988, new_n8329);
xor_4  g07953(new_n6001, new_n8329, new_n8330);
not_8  g07954(new_n6005, new_n8331);
or_8   g07955(new_n8331, new_n8330, new_n8332);
and_8  g07956(new_n8332, new_n8328, new_n8333);
or_8   g07957(new_n8333, new_n8327, new_n8334);
xor_4  g07958(new_n8324, new_n8322, new_n8335);
not_8  g07959(new_n8328, new_n8336_1);
and_8  g07960(new_n6005, new_n6002, new_n8337);
or_8   g07961(new_n8337, new_n8336_1, new_n8338);
or_8   g07962(new_n8338, new_n8335, new_n8339);
and_8  g07963(new_n8339, new_n8334, new_n8340);
xor_4  g07964(new_n8340, new_n8300, new_n8341);
xor_4  g07965(new_n8341, new_n8298, new_n8342);
or_8   g07966(new_n6192_1, new_n6117, new_n8343);
xor_4  g07967(new_n8343, new_n8342, new_n8344);
and_8  g07968(new_n6154, new_n6034, new_n8345);
not_8  g07969(new_n8345, new_n8346);
and_8  g07970(n12069, n5798, new_n8347);
nand_5 g07971(n7160, n5579, new_n8348);
not_8  g07972(new_n8348, new_n8349);
or_8   g07973(new_n6146, new_n6142, new_n8350);
and_8  g07974(new_n8350, new_n6143, new_n8351);
nor_6  g07975(new_n8351, new_n8349, new_n8352);
or_8   g07976(new_n8351, new_n6019, new_n8353);
and_8  g07977(new_n8353, new_n8349, new_n8354);
or_8   g07978(new_n8354, new_n8352, new_n8355);
and_8  g07979(n4828, n2498, new_n8356);
and_8  g07980(n2558, n2515, new_n8357);
xnor_4 g07981(new_n8357, new_n8356, new_n8358);
xor_4  g07982(new_n8358, new_n8355, new_n8359);
and_8  g07983(n12391, n6016, new_n8360);
and_8  g07984(n7891, n521, new_n8361);
xor_4  g07985(new_n8361, new_n8360, new_n8362);
and_8  g07986(new_n8362, new_n8359, new_n8363);
nor_6  g07987(new_n8362, new_n8359, new_n8364);
or_8   g07988(new_n8364, new_n8363, new_n8365);
not_8  g07989(new_n6141, new_n8366);
and_8  g07990(new_n6149, new_n8366, new_n8367);
or_8   g07991(new_n8367, new_n6139, new_n8368);
not_8  g07992(new_n8368, new_n8369);
or_8   g07993(new_n8369, new_n8365, new_n8370);
xor_4  g07994(new_n8362, new_n8359, new_n8371);
or_8   g07995(new_n8368, new_n8371, new_n8372);
and_8  g07996(new_n8372, new_n8370, new_n8373);
nor_6  g07997(new_n6150, new_n6133, new_n8374);
and_8  g07998(new_n6153, new_n6151, new_n8375);
or_8   g07999(new_n8375, new_n8374, new_n8376);
xor_4  g08000(new_n8376, new_n8373, new_n8377);
and_8  g08001(new_n8377, new_n8347, new_n8378);
not_8  g08002(new_n8347, new_n8379);
and_8  g08003(new_n8376, new_n8373, new_n8380);
nor_6  g08004(new_n8376, new_n8373, new_n8381);
or_8   g08005(new_n8381, new_n8380, new_n8382);
and_8  g08006(new_n8382, new_n8379, new_n8383);
or_8   g08007(new_n8383, new_n8378, new_n8384_1);
or_8   g08008(new_n8384_1, new_n8346, new_n8385);
or_8   g08009(new_n8382, new_n8379, new_n8386);
or_8   g08010(new_n8377, new_n8347, new_n8387);
and_8  g08011(new_n8387, new_n8386, new_n8388);
or_8   g08012(new_n8388, new_n8345, new_n8389);
and_8  g08013(new_n8389, new_n8385, new_n8390);
and_8  g08014(new_n6176, new_n6087, new_n8391);
and_8  g08015(n11222, n5153, new_n8392);
and_8  g08016(n3342, n996, new_n8393);
and_8  g08017(n9111, n5767, new_n8394);
and_8  g08018(n9763, n5319, new_n8395);
xor_4  g08019(new_n8395, new_n8394, new_n8396);
xor_4  g08020(new_n8396, new_n8393, new_n8397);
or_8   g08021(new_n6166, new_n6040, new_n8398_1);
and_8  g08022(new_n6166, new_n6040, new_n8399);
or_8   g08023(new_n8399, new_n6165, new_n8400);
and_8  g08024(new_n8400, new_n8398_1, new_n8401);
and_8  g08025(new_n8401, new_n8397, new_n8402);
nor_6  g08026(new_n8401, new_n8397, new_n8403);
or_8   g08027(new_n8403, new_n8402, new_n8404);
and_8  g08028(n11153, n7270, new_n8405);
and_8  g08029(n5314, n806, new_n8406);
xor_4  g08030(new_n8406, new_n8405, new_n8407);
not_8  g08031(new_n8407, new_n8408);
xor_4  g08032(new_n8408, new_n8404, new_n8409);
not_8  g08033(new_n6164, new_n8410);
and_8  g08034(new_n6168, new_n8410, new_n8411);
or_8   g08035(new_n8411, new_n6162, new_n8412);
and_8  g08036(new_n8412, new_n8409, new_n8413);
nor_6  g08037(new_n8412, new_n8409, new_n8414);
or_8   g08038(new_n8414, new_n8413, new_n8415);
nor_6  g08039(new_n6175, new_n6172, new_n8416);
nor_6  g08040(new_n8416, new_n6170, new_n8417);
or_8   g08041(new_n8417, new_n8415, new_n8418);
xor_4  g08042(new_n8412, new_n8409, new_n8419);
or_8   g08043(new_n8416, new_n6170, new_n8420);
or_8   g08044(new_n8420, new_n8419, new_n8421);
and_8  g08045(new_n8421, new_n8418, new_n8422);
and_8  g08046(new_n8422, new_n8392, new_n8423);
or_8   g08047(new_n8422, new_n8392, new_n8424);
not_8  g08048(new_n8424, new_n8425);
or_8   g08049(new_n8425, new_n8423, new_n8426);
and_8  g08050(new_n8426, new_n8391, new_n8427);
not_8  g08051(new_n8391, new_n8428);
xor_4  g08052(new_n8422, new_n8392, new_n8429);
and_8  g08053(new_n8429, new_n8428, new_n8430);
or_8   g08054(new_n8430, new_n8427, new_n8431);
and_8  g08055(new_n8431, new_n8390, new_n8432);
and_8  g08056(new_n8388, new_n8345, new_n8433_1);
and_8  g08057(new_n8384_1, new_n8346, new_n8434);
or_8   g08058(new_n8434, new_n8433_1, new_n8435);
or_8   g08059(new_n8429, new_n8428, new_n8436);
or_8   g08060(new_n8426, new_n8391, new_n8437);
and_8  g08061(new_n8437, new_n8436, new_n8438);
and_8  g08062(new_n8438, new_n8435, new_n8439);
or_8   g08063(new_n8439, new_n8432, new_n8440);
or_8   g08064(new_n6189, new_n6179, new_n8441);
xor_4  g08065(new_n8441, new_n8440, new_n8442);
xor_4  g08066(new_n8442, new_n8344, new_n8443);
xor_4  g08067(new_n8443, new_n8297, n2708);
xnor_4 g08068(new_n880, new_n879, n2818);
xnor_4 g08069(new_n2102, new_n2076, n2902);
and_8  g08070(n11407, n5305, new_n8447);
and_8  g08071(n12709, n8759, new_n8448);
and_8  g08072(n12489, n5331, new_n8449);
and_8  g08073(n10990, n7965, new_n8450);
xor_4  g08074(new_n8450, new_n8449, new_n8451);
xor_4  g08075(new_n8451, new_n8448, new_n8452);
xor_4  g08076(new_n8452, new_n8447, n3071);
xnor_4 g08077(new_n3041, new_n3037, n3124);
and_8  g08078(new_n8452, new_n8447, new_n8455);
and_8  g08079(n11407, n5964, new_n8456);
and_8  g08080(n5305, n5212, new_n8457);
xor_4  g08081(new_n8457, new_n8456, new_n8458);
or_8   g08082(new_n8458, new_n8455, new_n8459);
and_8  g08083(new_n8451, new_n8448, new_n8460);
and_8  g08084(n11728, n8759, new_n8461);
and_8  g08085(n12709, n6776, new_n8462);
xor_4  g08086(new_n8462, new_n8461, new_n8463);
xnor_4 g08087(new_n8463, new_n8460, new_n8464);
and_8  g08088(new_n8450, new_n8449, new_n8465);
and_8  g08089(n7159, n5331, new_n8466);
and_8  g08090(n12489, n8476, new_n8467);
xor_4  g08091(new_n8467, new_n8466, new_n8468);
xor_4  g08092(new_n8468, new_n8465, new_n8469);
and_8  g08093(n7965, n5760, new_n8470);
and_8  g08094(n10990, n7388, new_n8471);
xnor_4 g08095(new_n8471, new_n8470, new_n8472);
xor_4  g08096(new_n8472, new_n8469, new_n8473);
xor_4  g08097(new_n8473, new_n8464, new_n8474);
xnor_4 g08098(new_n8458, new_n8455, new_n8475);
or_8   g08099(new_n8475, new_n8474, new_n8476_1);
and_8  g08100(new_n8476_1, new_n8459, new_n8477);
not_8  g08101(new_n8447, new_n8478);
and_8  g08102(n5964, n5212, new_n8479);
and_8  g08103(new_n8479, new_n8478, new_n8480);
and_8  g08104(n11407, n1097, new_n8481);
and_8  g08105(n11877, n5305, new_n8482);
xor_4  g08106(new_n8482, new_n8481, new_n8483);
or_8   g08107(new_n8483, new_n8480, new_n8484);
or_8   g08108(new_n8482, new_n8481, new_n8485);
nand_5 g08109(new_n8485, new_n8480, new_n8486);
and_8  g08110(new_n8486, new_n8484, new_n8487);
xor_4  g08111(new_n8487, new_n8477, new_n8488);
and_8  g08112(new_n8463, new_n8460, new_n8489);
nor_6  g08113(new_n8473, new_n8464, new_n8490);
or_8   g08114(new_n8490, new_n8489, new_n8491);
not_8  g08115(new_n8448, new_n8492);
and_8  g08116(n11728, n6776, new_n8493);
nand_5 g08117(new_n8493, new_n8492, new_n8494);
and_8  g08118(n12709, n12299, new_n8495);
and_8  g08119(n8759, n6429, new_n8496);
xnor_4 g08120(new_n8496, new_n8495, new_n8497);
and_8  g08121(new_n8497, new_n8494, new_n8498);
not_8  g08122(new_n8494, new_n8499);
or_8   g08123(new_n8496, new_n8495, new_n8500);
and_8  g08124(new_n8500, new_n8499, new_n8501);
nor_6  g08125(new_n8501, new_n8498, new_n8502);
xor_4  g08126(new_n8502, new_n8491, new_n8503);
not_8  g08127(new_n8449, new_n8504);
and_8  g08128(n8476, n7159, new_n8505);
nand_5 g08129(new_n8505, new_n8504, new_n8506);
and_8  g08130(n12489, n2530, new_n8507);
and_8  g08131(n12777, n5331, new_n8508);
or_8   g08132(new_n8508, new_n8507, new_n8509);
not_8  g08133(new_n8509, new_n8510);
and_8  g08134(n12777, n2530, new_n8511);
and_8  g08135(new_n8511, new_n8449, new_n8512);
or_8   g08136(new_n8512, new_n8510, new_n8513);
and_8  g08137(new_n8513, new_n8506, new_n8514);
nor_6  g08138(new_n8510, new_n8506, new_n8515);
or_8   g08139(new_n8515, new_n8514, new_n8516);
not_8  g08140(new_n8450, new_n8517);
and_8  g08141(n7388, n5760, new_n8518);
nand_5 g08142(new_n8518, new_n8517, new_n8519);
and_8  g08143(n11892, n10990, new_n8520);
and_8  g08144(n7965, n1478, new_n8521);
xnor_4 g08145(new_n8521, new_n8520, new_n8522);
and_8  g08146(new_n8522, new_n8519, new_n8523);
not_8  g08147(new_n8519, new_n8524);
or_8   g08148(new_n8521, new_n8520, new_n8525);
and_8  g08149(new_n8525, new_n8524, new_n8526);
or_8   g08150(new_n8526, new_n8523, new_n8527);
xor_4  g08151(new_n8527, new_n8516, new_n8528);
or_8   g08152(new_n8468, new_n8465, new_n8529);
nand_5 g08153(new_n8472, new_n8469, new_n8530);
and_8  g08154(new_n8530, new_n8529, new_n8531);
xor_4  g08155(new_n8531, new_n8528, new_n8532);
xor_4  g08156(new_n8532, new_n8503, new_n8533);
xor_4  g08157(new_n8533, new_n8488, n3214);
xnor_4 g08158(new_n5788, new_n5786, n3230);
xor_4  g08159(new_n5189, new_n5136, n3272);
and_8  g08160(n5964, n4370, new_n8537);
and_8  g08161(n11407, n4312, new_n8538);
and_8  g08162(n11877, n5964, new_n8539);
or_8   g08163(new_n8539, new_n8538, new_n8540);
and_8  g08164(new_n8539, new_n8538, new_n8541);
and_8  g08165(n5212, n1097, new_n8542);
or_8   g08166(new_n8542, new_n8541, new_n8543);
and_8  g08167(new_n8543, new_n8540, new_n8544);
and_8  g08168(new_n8544, new_n8537, new_n8545);
xor_4  g08169(new_n8544, new_n8537, new_n8546);
and_8  g08170(n5212, n4312, new_n8547);
and_8  g08171(n11877, n1097, new_n8548);
and_8  g08172(n12705, n11407, new_n8549);
xor_4  g08173(new_n8549, new_n8548, new_n8550);
xor_4  g08174(new_n8550, new_n8547, new_n8551);
and_8  g08175(new_n8551, new_n8546, new_n8552);
or_8   g08176(new_n8552, new_n8545, new_n8553);
and_8  g08177(n5964, n5320, new_n8554);
and_8  g08178(n4370, n1097, new_n8555);
xnor_4 g08179(new_n8555, new_n8554, new_n8556);
xor_4  g08180(new_n8556, new_n8553, new_n8557);
and_8  g08181(n11877, n4312, new_n8558);
and_8  g08182(n12705, n5212, new_n8559);
and_8  g08183(n12025, n11407, new_n8560);
xor_4  g08184(new_n8560, new_n8559, new_n8561);
xor_4  g08185(new_n8561, new_n8558, new_n8562);
or_8   g08186(new_n8549, new_n8548, new_n8563);
and_8  g08187(new_n8549, new_n8548, new_n8564);
or_8   g08188(new_n8564, new_n8547, new_n8565);
nand_5 g08189(new_n8565, new_n8563, new_n8566);
xor_4  g08190(new_n8566, new_n8562, new_n8567);
xor_4  g08191(new_n8567, new_n8557, new_n8568);
and_8  g08192(n5320, n5305, new_n8569);
xor_4  g08193(new_n8551, new_n8546, new_n8570);
or_8   g08194(new_n8570, new_n8569, new_n8571);
not_8  g08195(new_n8569, new_n8572);
xor_4  g08196(new_n8570, new_n8572, new_n8573);
and_8  g08197(n5305, n4370, new_n8574);
and_8  g08198(new_n8482, new_n8481, new_n8575);
or_8   g08199(new_n8575, new_n8479, new_n8576);
and_8  g08200(new_n8576, new_n8485, new_n8577);
and_8  g08201(new_n8577, new_n8574, new_n8578);
xor_4  g08202(new_n8577, new_n8574, new_n8579);
xor_4  g08203(new_n8539, new_n8538, new_n8580);
xor_4  g08204(new_n8580, new_n8542, new_n8581);
and_8  g08205(new_n8581, new_n8579, new_n8582);
or_8   g08206(new_n8582, new_n8578, new_n8583);
or_8   g08207(new_n8583, new_n8573, new_n8584);
and_8  g08208(new_n8584, new_n8571, new_n8585);
and_8  g08209(new_n8585, new_n8568, new_n8586);
nor_6  g08210(new_n8561, new_n8558, new_n8587);
and_8  g08211(new_n8566, new_n8562, new_n8588);
or_8   g08212(new_n8588, new_n8587, new_n8589);
and_8  g08213(n12000, n5964, new_n8590);
and_8  g08214(n5320, n1097, new_n8591);
and_8  g08215(n9725, n5305, new_n8592);
xnor_4 g08216(new_n8592, new_n8591, new_n8593);
xor_4  g08217(new_n8593, new_n8590, new_n8594);
xor_4  g08218(new_n8594, new_n8589, new_n8595_1);
and_8  g08219(new_n8560, new_n8559, new_n8596);
and_8  g08220(n4370, n4312, new_n8597);
xor_4  g08221(new_n8597, new_n8596, new_n8598);
and_8  g08222(n12025, n5212, new_n8599);
and_8  g08223(n12705, n11877, new_n8600);
and_8  g08224(n11407, n11257, new_n8601);
xnor_4 g08225(new_n8601, new_n8600, new_n8602);
xor_4  g08226(new_n8602, new_n8599, new_n8603);
xor_4  g08227(new_n8603, new_n8598, new_n8604);
xor_4  g08228(new_n8604, new_n8595_1, new_n8605);
not_8  g08229(new_n8553, new_n8606);
or_8   g08230(new_n8556, new_n8606, new_n8607);
and_8  g08231(new_n8555, new_n8554, new_n8608);
or_8   g08232(new_n8567, new_n8557, new_n8609);
xor_4  g08233(new_n8609, new_n8608, new_n8610);
and_8  g08234(new_n8610, new_n8607, new_n8611);
xor_4  g08235(new_n8611, new_n8605, new_n8612);
xor_4  g08236(new_n8612, new_n8586, new_n8613);
and_8  g08237(n12000, n5305, new_n8614);
xor_4  g08238(new_n8585, new_n8568, new_n8615);
and_8  g08239(new_n8615, new_n8614, new_n8616);
xor_4  g08240(new_n8581, new_n8579, new_n8617);
not_8  g08241(new_n8484, new_n8618);
and_8  g08242(new_n8618, new_n8479, new_n8619);
and_8  g08243(new_n8619, new_n8617, new_n8620);
not_8  g08244(new_n8620, new_n8621);
xor_4  g08245(new_n8583, new_n8573, new_n8622);
nor_6  g08246(new_n8622, new_n8621, new_n8623);
xor_4  g08247(new_n8615, new_n8614, new_n8624);
and_8  g08248(new_n8624, new_n8623, new_n8625);
or_8   g08249(new_n8625, new_n8616, new_n8626);
xor_4  g08250(new_n8626, new_n8613, new_n8627);
not_8  g08251(new_n8627, new_n8628);
and_8  g08252(n8759, n8717, new_n8629);
and_8  g08253(n7436, n6429, new_n8630);
and_8  g08254(n12709, n9241, new_n8631);
and_8  g08255(n11728, n8276, new_n8632);
xor_4  g08256(new_n8632, new_n8631, new_n8633);
xor_4  g08257(new_n8633, new_n8630, new_n8634);
and_8  g08258(n12299, n6429, new_n8635);
and_8  g08259(n12709, n8276, new_n8636);
or_8   g08260(new_n8636, new_n8635, new_n8637);
and_8  g08261(new_n8636, new_n8635, new_n8638);
and_8  g08262(n11728, n7436, new_n8639);
or_8   g08263(new_n8639, new_n8638, new_n8640);
nand_5 g08264(new_n8640, new_n8637, new_n8641);
and_8  g08265(new_n8641, new_n8634, new_n8642);
nor_6  g08266(new_n8641, new_n8634, new_n8643);
or_8   g08267(new_n8643, new_n8642, new_n8644);
and_8  g08268(n6776, n2433, new_n8645);
and_8  g08269(n12299, n8819, new_n8646);
xor_4  g08270(new_n8646, new_n8645, new_n8647);
xor_4  g08271(new_n8647, new_n8644, new_n8648);
and_8  g08272(n8819, n6776, new_n8649);
and_8  g08273(n12709, n7436, new_n8650);
and_8  g08274(n6776, n6429, new_n8651);
or_8   g08275(new_n8651, new_n8650, new_n8652);
and_8  g08276(new_n8651, new_n8650, new_n8653);
and_8  g08277(n12299, n11728, new_n8654);
or_8   g08278(new_n8654, new_n8653, new_n8655);
and_8  g08279(new_n8655, new_n8652, new_n8656);
and_8  g08280(new_n8656, new_n8649, new_n8657);
xnor_4 g08281(new_n8656, new_n8649, new_n8658);
not_8  g08282(new_n8658, new_n8659);
xor_4  g08283(new_n8636, new_n8635, new_n8660);
xor_4  g08284(new_n8660, new_n8639, new_n8661);
and_8  g08285(new_n8661, new_n8659, new_n8662);
or_8   g08286(new_n8662, new_n8657, new_n8663);
and_8  g08287(new_n8663, new_n8648, new_n8664);
nor_6  g08288(new_n8663, new_n8648, new_n8665_1);
or_8   g08289(new_n8665_1, new_n8664, new_n8666);
not_8  g08290(n2433, new_n8667);
not_8  g08291(n8759, new_n8668);
or_8   g08292(new_n8668, new_n8667, new_n8669);
xor_4  g08293(new_n8661, new_n8658, new_n8670);
and_8  g08294(new_n8670, new_n8669, new_n8671);
nor_6  g08295(new_n8670, new_n8669, new_n8672);
or_8   g08296(new_n8672, new_n8671, new_n8673);
and_8  g08297(n8819, n8759, new_n8674);
and_8  g08298(new_n8496, new_n8495, new_n8675);
or_8   g08299(new_n8675, new_n8493, new_n8676);
and_8  g08300(new_n8676, new_n8500, new_n8677);
and_8  g08301(new_n8677, new_n8674, new_n8678);
xor_4  g08302(new_n8677, new_n8674, new_n8679);
xor_4  g08303(new_n8651, new_n8650, new_n8680);
xor_4  g08304(new_n8680, new_n8654, new_n8681);
and_8  g08305(new_n8681, new_n8679, new_n8682);
or_8   g08306(new_n8682, new_n8678, new_n8683);
nor_6  g08307(new_n8683, new_n8673, new_n8684);
or_8   g08308(new_n8684, new_n8671, new_n8685);
xor_4  g08309(new_n8685, new_n8666, new_n8686);
and_8  g08310(new_n8686, new_n8629, new_n8687);
not_8  g08311(new_n8687, new_n8688);
xor_4  g08312(new_n8681, new_n8679, new_n8689);
and_8  g08313(new_n8498, new_n8493, new_n8690);
nand_5 g08314(new_n8690, new_n8689, new_n8691);
xor_4  g08315(new_n8683, new_n8673, new_n8692);
or_8   g08316(new_n8692, new_n8691, new_n8693);
not_8  g08317(new_n8686, new_n8694);
xor_4  g08318(new_n8694, new_n8629, new_n8695);
or_8   g08319(new_n8695, new_n8693, new_n8696);
and_8  g08320(new_n8696, new_n8688, new_n8697);
or_8   g08321(new_n8685, new_n8666, new_n8698);
not_8  g08322(new_n8698, new_n8699);
nor_6  g08323(new_n8633, new_n8630, new_n8700);
nor_6  g08324(new_n8642, new_n8700, new_n8701);
and_8  g08325(n8717, n6776, new_n8702);
and_8  g08326(n12299, n2433, new_n8703);
and_8  g08327(n8759, n7730, new_n8704);
xnor_4 g08328(new_n8704, new_n8703, new_n8705);
xor_4  g08329(new_n8705, new_n8702, new_n8706);
xor_4  g08330(new_n8706, new_n8701, new_n8707);
and_8  g08331(new_n8632, new_n8631, new_n8708);
and_8  g08332(n8819, n7436, new_n8709);
xnor_4 g08333(new_n8709, new_n8708, new_n8710);
and_8  g08334(n11728, n9241, new_n8711);
and_8  g08335(n8276, n6429, new_n8712);
and_8  g08336(n12709, n10510, new_n8713);
xnor_4 g08337(new_n8713, new_n8712, new_n8714);
xor_4  g08338(new_n8714, new_n8711, new_n8715);
xor_4  g08339(new_n8715, new_n8710, new_n8716);
xor_4  g08340(new_n8716, new_n8707, new_n8717_1);
not_8  g08341(new_n8717_1, new_n8718);
and_8  g08342(new_n8647, new_n8644, new_n8719);
and_8  g08343(new_n8646, new_n8645, new_n8720);
xor_4  g08344(new_n8664, new_n8720, new_n8721);
or_8   g08345(new_n8721, new_n8719, new_n8722);
xor_4  g08346(new_n8722, new_n8718, new_n8723);
xor_4  g08347(new_n8723, new_n8699, new_n8724);
xor_4  g08348(new_n8724, new_n8697, new_n8725);
not_8  g08349(n1478, new_n8726);
or_8   g08350(new_n2748, new_n8726, new_n8727);
and_8  g08351(n5860, n5760, new_n8728);
and_8  g08352(n10990, n3986, new_n8729);
xor_4  g08353(new_n8729, new_n8728, new_n8730);
xor_4  g08354(new_n8730, new_n8727, new_n8731);
and_8  g08355(n11892, n1478, new_n8732);
and_8  g08356(n10990, n5860, new_n8733);
or_8   g08357(new_n8733, new_n8732, new_n8734);
and_8  g08358(new_n8733, new_n8732, new_n8735);
and_8  g08359(n5760, n2393, new_n8736);
or_8   g08360(new_n8736, new_n8735, new_n8737);
and_8  g08361(new_n8737, new_n8734, new_n8738);
xor_4  g08362(new_n8738, new_n8731, new_n8739);
and_8  g08363(n12947, n7388, new_n8740);
and_8  g08364(n11892, n11791, new_n8741);
xor_4  g08365(new_n8741, new_n8740, new_n8742);
not_8  g08366(new_n8742, new_n8743);
or_8   g08367(new_n8743, new_n8739, new_n8744);
nand_5 g08368(new_n8737, new_n8734, new_n8745);
xor_4  g08369(new_n8745, new_n8731, new_n8746);
or_8   g08370(new_n8742, new_n8746, new_n8747);
and_8  g08371(new_n8747, new_n8744, new_n8748);
and_8  g08372(n11791, n7388, new_n8749);
and_8  g08373(n10990, n2393, new_n8750);
and_8  g08374(n7388, n1478, new_n8751);
or_8   g08375(new_n8751, new_n8750, new_n8752);
and_8  g08376(new_n8751, new_n8750, new_n8753);
and_8  g08377(n11892, n5760, new_n8754);
or_8   g08378(new_n8754, new_n8753, new_n8755);
and_8  g08379(new_n8755, new_n8752, new_n8756);
and_8  g08380(new_n8756, new_n8749, new_n8757);
xnor_4 g08381(new_n8756, new_n8749, new_n8758);
xnor_4 g08382(new_n8733, new_n8732, new_n8759_1);
xor_4  g08383(new_n8759_1, new_n8736, new_n8760);
nor_6  g08384(new_n8760, new_n8758, new_n8761);
or_8   g08385(new_n8761, new_n8757, new_n8762);
and_8  g08386(new_n8762, new_n8748, new_n8763);
nor_6  g08387(new_n8762, new_n8748, new_n8764);
or_8   g08388(new_n8764, new_n8763, new_n8765);
and_8  g08389(n12947, n7965, new_n8766);
and_8  g08390(n11791, n7965, new_n8767);
and_8  g08391(new_n8521, new_n8520, new_n8768);
or_8   g08392(new_n8768, new_n8518, new_n8769);
and_8  g08393(new_n8769, new_n8525, new_n8770);
and_8  g08394(new_n8770, new_n8767, new_n8771);
xor_4  g08395(new_n8770, new_n8767, new_n8772);
xor_4  g08396(new_n8751, new_n8750, new_n8773);
xor_4  g08397(new_n8773, new_n8754, new_n8774);
and_8  g08398(new_n8774, new_n8772, new_n8775);
or_8   g08399(new_n8775, new_n8771, new_n8776);
nor_6  g08400(new_n8776, new_n8766, new_n8777);
and_8  g08401(new_n8760, new_n8758, new_n8778);
or_8   g08402(new_n8778, new_n8761, new_n8779);
not_8  g08403(new_n8779, new_n8780);
and_8  g08404(new_n8776, new_n8766, new_n8781);
or_8   g08405(new_n8781, new_n8777, new_n8782);
nor_6  g08406(new_n8782, new_n8780, new_n8783);
or_8   g08407(new_n8783, new_n8777, new_n8784);
or_8   g08408(new_n8784, new_n8765, new_n8785);
and_8  g08409(new_n8729, new_n8728, new_n8786);
and_8  g08410(n11791, n2393, new_n8787);
xnor_4 g08411(new_n8787, new_n8786, new_n8788);
and_8  g08412(n5760, n3986, new_n8789);
and_8  g08413(n5860, n1478, new_n8790);
and_8  g08414(n10990, n5857, new_n8791);
xnor_4 g08415(new_n8791, new_n8790, new_n8792);
xor_4  g08416(new_n8792, new_n8789, new_n8793);
nor_6  g08417(new_n8793, new_n8788, new_n8794);
and_8  g08418(new_n8793, new_n8788, new_n8795);
or_8   g08419(new_n8795, new_n8794, new_n8796);
and_8  g08420(n7388, n6441, new_n8797);
and_8  g08421(n12947, n11892, new_n8798);
and_8  g08422(n11999, n7965, new_n8799);
xnor_4 g08423(new_n8799, new_n8798, new_n8800);
xor_4  g08424(new_n8800, new_n8797, new_n8801);
not_8  g08425(new_n8730, new_n8802);
or_8   g08426(new_n8802, new_n8727, new_n8803);
or_8   g08427(new_n8745, new_n8731, new_n8804);
and_8  g08428(new_n8804, new_n8803, new_n8805);
xor_4  g08429(new_n8805, new_n8801, new_n8806);
xor_4  g08430(new_n8806, new_n8796, new_n8807);
not_8  g08431(new_n8807, new_n8808);
not_8  g08432(new_n8744, new_n8809);
and_8  g08433(new_n8741, new_n8740, new_n8810);
xor_4  g08434(new_n8763, new_n8810, new_n8811);
or_8   g08435(new_n8811, new_n8809, new_n8812);
and_8  g08436(new_n8812, new_n8808, new_n8813);
nor_6  g08437(new_n8811, new_n8809, new_n8814);
and_8  g08438(new_n8814, new_n8807, new_n8815);
or_8   g08439(new_n8815, new_n8813, new_n8816);
or_8   g08440(new_n8816, new_n8785, new_n8817);
not_8  g08441(new_n8785, new_n8818);
or_8   g08442(new_n8814, new_n8807, new_n8819_1);
or_8   g08443(new_n8812, new_n8808, new_n8820);
and_8  g08444(new_n8820, new_n8819_1, new_n8821);
or_8   g08445(new_n8821, new_n8818, new_n8822);
and_8  g08446(new_n8822, new_n8817, new_n8823);
not_8  g08447(n6441, new_n8824);
not_8  g08448(n7965, new_n8825);
or_8   g08449(new_n8825, new_n8824, new_n8826);
not_8  g08450(new_n8826, new_n8827);
xor_4  g08451(new_n8762, new_n8748, new_n8828);
nor_6  g08452(new_n8783, new_n8777, new_n8829);
or_8   g08453(new_n8829, new_n8828, new_n8830);
and_8  g08454(new_n8830, new_n8785, new_n8831);
and_8  g08455(new_n8831, new_n8827, new_n8832);
xor_4  g08456(new_n8829, new_n8765, new_n8833);
and_8  g08457(new_n8833, new_n8826, new_n8834);
xor_4  g08458(new_n8774, new_n8772, new_n8835);
and_8  g08459(new_n8523, new_n8518, new_n8836);
nand_5 g08460(new_n8836, new_n8835, new_n8837);
xor_4  g08461(new_n8782, new_n8780, new_n8838);
or_8   g08462(new_n8838, new_n8837, new_n8839);
nor_6  g08463(new_n8839, new_n8834, new_n8840);
or_8   g08464(new_n8840, new_n8832, new_n8841);
and_8  g08465(new_n8841, new_n8823, new_n8842);
nor_6  g08466(new_n8841, new_n8823, new_n8843);
or_8   g08467(new_n8843, new_n8842, new_n8844);
not_8  g08468(n12777, new_n8845);
or_8   g08469(new_n8845, new_n702, new_n8846);
and_8  g08470(n10545, n7159, new_n8847);
and_8  g08471(n12489, n7690, new_n8848);
xor_4  g08472(new_n8848, new_n8847, new_n8849);
xor_4  g08473(new_n8849, new_n8846, new_n8850);
and_8  g08474(n12489, n10545, new_n8851);
or_8   g08475(new_n8851, new_n8511, new_n8852);
and_8  g08476(new_n8851, new_n8511, new_n8853);
and_8  g08477(n12648, n7159, new_n8854);
or_8   g08478(new_n8854, new_n8853, new_n8855);
and_8  g08479(new_n8855, new_n8852, new_n8856);
xor_4  g08480(new_n8856, new_n8850, new_n8857);
and_8  g08481(n6254, n2530, new_n8858);
and_8  g08482(n11967, n8476, new_n8859);
xor_4  g08483(new_n8859, new_n8858, new_n8860);
not_8  g08484(new_n8860, new_n8861);
or_8   g08485(new_n8861, new_n8857, new_n8862);
nand_5 g08486(new_n8855, new_n8852, new_n8863);
xor_4  g08487(new_n8863, new_n8850, new_n8864);
or_8   g08488(new_n8860, new_n8864, new_n8865);
and_8  g08489(new_n8865, new_n8862, new_n8866);
and_8  g08490(n8476, n6254, new_n8867);
and_8  g08491(n12648, n12489, new_n8868);
and_8  g08492(n12777, n8476, new_n8869);
or_8   g08493(new_n8869, new_n8868, new_n8870);
and_8  g08494(new_n8869, new_n8868, new_n8871);
and_8  g08495(n7159, n2530, new_n8872);
or_8   g08496(new_n8872, new_n8871, new_n8873);
and_8  g08497(new_n8873, new_n8870, new_n8874);
and_8  g08498(new_n8874, new_n8867, new_n8875);
xnor_4 g08499(new_n8874, new_n8867, new_n8876);
xnor_4 g08500(new_n8851, new_n8511, new_n8877);
xor_4  g08501(new_n8877, new_n8854, new_n8878);
nor_6  g08502(new_n8878, new_n8876, new_n8879);
or_8   g08503(new_n8879, new_n8875, new_n8880);
and_8  g08504(new_n8880, new_n8866, new_n8881);
nor_6  g08505(new_n8880, new_n8866, new_n8882);
or_8   g08506(new_n8882, new_n8881, new_n8883);
and_8  g08507(n11967, n5331, new_n8884);
not_8  g08508(new_n8884, new_n8885);
and_8  g08509(new_n8878, new_n8876, new_n8886);
or_8   g08510(new_n8886, new_n8879, new_n8887);
and_8  g08511(new_n8887, new_n8885, new_n8888);
xor_4  g08512(new_n8878, new_n8876, new_n8889);
or_8   g08513(new_n8889, new_n8884, new_n8890);
or_8   g08514(new_n8887, new_n8885, new_n8891);
and_8  g08515(new_n8891, new_n8890, new_n8892);
and_8  g08516(n6254, n5331, new_n8893);
or_8   g08517(new_n8512, new_n8505, new_n8894);
and_8  g08518(new_n8894, new_n8509, new_n8895);
and_8  g08519(new_n8895, new_n8893, new_n8896);
xnor_4 g08520(new_n8895, new_n8893, new_n8897);
xnor_4 g08521(new_n8869, new_n8868, new_n8898);
xor_4  g08522(new_n8898, new_n8872, new_n8899);
nor_6  g08523(new_n8899, new_n8897, new_n8900);
or_8   g08524(new_n8900, new_n8896, new_n8901);
not_8  g08525(new_n8901, new_n8902);
and_8  g08526(new_n8902, new_n8892, new_n8903);
or_8   g08527(new_n8903, new_n8888, new_n8904);
or_8   g08528(new_n8904, new_n8883, new_n8905);
and_8  g08529(n5331, n1353, new_n8906);
and_8  g08530(n11967, n2530, new_n8907);
and_8  g08531(n8476, n447, new_n8908);
xnor_4 g08532(new_n8908, new_n8907, new_n8909);
xor_4  g08533(new_n8909, new_n8906, new_n8910);
not_8  g08534(new_n8849, new_n8911);
or_8   g08535(new_n8911, new_n8846, new_n8912);
or_8   g08536(new_n8863, new_n8850, new_n8913);
and_8  g08537(new_n8913, new_n8912, new_n8914);
xor_4  g08538(new_n8914, new_n8910, new_n8915);
not_8  g08539(new_n8915, new_n8916);
and_8  g08540(new_n8848, new_n8847, new_n8917);
and_8  g08541(n12648, n6254, new_n8918);
xnor_4 g08542(new_n8918, new_n8917, new_n8919);
and_8  g08543(n7690, n7159, new_n8920);
and_8  g08544(n12777, n10545, new_n8921);
and_8  g08545(n12489, n3616, new_n8922);
xnor_4 g08546(new_n8922, new_n8921, new_n8923);
xor_4  g08547(new_n8923, new_n8920, new_n8924);
xor_4  g08548(new_n8924, new_n8919, new_n8925);
xor_4  g08549(new_n8925, new_n8916, new_n8926);
not_8  g08550(new_n8926, new_n8927);
not_8  g08551(new_n8862, new_n8928);
nand_5 g08552(new_n8859, new_n8858, new_n8929);
not_8  g08553(new_n8929, new_n8930);
xor_4  g08554(new_n8881, new_n8930, new_n8931);
or_8   g08555(new_n8931, new_n8928, new_n8932);
and_8  g08556(new_n8932, new_n8927, new_n8933);
nor_6  g08557(new_n8931, new_n8928, new_n8934);
and_8  g08558(new_n8934, new_n8926, new_n8935);
or_8   g08559(new_n8935, new_n8933, new_n8936);
or_8   g08560(new_n8936, new_n8905, new_n8937);
not_8  g08561(new_n8905, new_n8938);
or_8   g08562(new_n8934, new_n8926, new_n8939);
or_8   g08563(new_n8932, new_n8927, new_n8940);
and_8  g08564(new_n8940, new_n8939, new_n8941);
or_8   g08565(new_n8941, new_n8938, new_n8942);
and_8  g08566(new_n8942, new_n8937, new_n8943);
and_8  g08567(n5331, n447, new_n8944);
not_8  g08568(new_n8883, new_n8945);
and_8  g08569(new_n8889, new_n8884, new_n8946);
or_8   g08570(new_n8946, new_n8888, new_n8947);
or_8   g08571(new_n8901, new_n8947, new_n8948);
and_8  g08572(new_n8948, new_n8890, new_n8949);
or_8   g08573(new_n8949, new_n8945, new_n8950);
and_8  g08574(new_n8950, new_n8905, new_n8951);
and_8  g08575(new_n8951, new_n8944, new_n8952);
or_8   g08576(new_n8951, new_n8944, new_n8953);
xor_4  g08577(new_n8899, new_n8897, new_n8954);
and_8  g08578(new_n8514, new_n8505, new_n8955);
and_8  g08579(new_n8955, new_n8954, new_n8956);
xor_4  g08580(new_n8901, new_n8892, new_n8957);
and_8  g08581(new_n8957, new_n8956, new_n8958);
and_8  g08582(new_n8958, new_n8953, new_n8959);
or_8   g08583(new_n8959, new_n8952, new_n8960);
and_8  g08584(new_n8960, new_n8943, new_n8961);
nor_6  g08585(new_n8960, new_n8943, new_n8962);
or_8   g08586(new_n8962, new_n8961, new_n8963);
and_8  g08587(new_n8963, new_n8844, new_n8964);
xor_4  g08588(new_n8841, new_n8823, new_n8965);
xor_4  g08589(new_n8960, new_n8943, new_n8966);
and_8  g08590(new_n8966, new_n8965, new_n8967);
or_8   g08591(new_n8967, new_n8964, new_n8968);
not_8  g08592(new_n8839, new_n8969);
xor_4  g08593(new_n8831, new_n8827, new_n8970);
or_8   g08594(new_n8970, new_n8969, new_n8971);
or_8   g08595(new_n8834, new_n8832, new_n8972);
or_8   g08596(new_n8972, new_n8839, new_n8973);
and_8  g08597(new_n8973, new_n8971, new_n8974);
xor_4  g08598(new_n8951, new_n8944, new_n8975);
or_8   g08599(new_n8975, new_n8958, new_n8976);
not_8  g08600(new_n8958, new_n8977);
not_8  g08601(new_n8944, new_n8978);
xor_4  g08602(new_n8951, new_n8978, new_n8979);
or_8   g08603(new_n8979, new_n8977, new_n8980);
and_8  g08604(new_n8980, new_n8976, new_n8981);
or_8   g08605(new_n8981, new_n8974, new_n8982);
not_8  g08606(new_n8956, new_n8983);
xor_4  g08607(new_n8901, new_n8947, new_n8984);
and_8  g08608(new_n8984, new_n8983, new_n8985);
nor_6  g08609(new_n8985, new_n8958, new_n8986);
xor_4  g08610(new_n8838, new_n8837, new_n8987);
or_8   g08611(new_n8987, new_n8986, new_n8988);
or_8   g08612(new_n8985, new_n8958, new_n8989);
xor_4  g08613(new_n8987, new_n8989, new_n8990);
xor_4  g08614(new_n8955, new_n8954, new_n8991);
xor_4  g08615(new_n8836, new_n8835, new_n8992);
and_8  g08616(new_n8992, new_n8991, new_n8993);
nor_6  g08617(new_n8527, new_n8516, new_n8994);
and_8  g08618(new_n8531, new_n8528, new_n8995);
or_8   g08619(new_n8995, new_n8994, new_n8996);
xor_4  g08620(new_n8992, new_n8991, new_n8997);
and_8  g08621(new_n8997, new_n8996, new_n8998);
or_8   g08622(new_n8998, new_n8993, new_n8999);
or_8   g08623(new_n8999, new_n8990, new_n9000);
and_8  g08624(new_n9000, new_n8988, new_n9001);
and_8  g08625(new_n8972, new_n8839, new_n9002);
and_8  g08626(new_n8970, new_n8969, new_n9003);
or_8   g08627(new_n9003, new_n9002, new_n9004);
and_8  g08628(new_n8979, new_n8977, new_n9005);
and_8  g08629(new_n8975, new_n8958, new_n9006);
or_8   g08630(new_n9006, new_n9005, new_n9007);
and_8  g08631(new_n9007, new_n9004, new_n9008);
and_8  g08632(new_n8981, new_n8974, new_n9009);
or_8   g08633(new_n9009, new_n9008, new_n9010);
or_8   g08634(new_n9010, new_n9001, new_n9011);
and_8  g08635(new_n9011, new_n8982, new_n9012);
or_8   g08636(new_n9012, new_n8968, new_n9013);
or_8   g08637(new_n8966, new_n8965, new_n9014);
or_8   g08638(new_n8963, new_n8844, new_n9015);
and_8  g08639(new_n9015, new_n9014, new_n9016);
not_8  g08640(new_n8988, new_n9017);
xor_4  g08641(new_n8987, new_n8986, new_n9018);
nor_6  g08642(new_n8998, new_n8993, new_n9019);
and_8  g08643(new_n9019, new_n9018, new_n9020);
or_8   g08644(new_n9020, new_n9017, new_n9021);
or_8   g08645(new_n9007, new_n9004, new_n9022);
and_8  g08646(new_n9022, new_n8982, new_n9023);
and_8  g08647(new_n9023, new_n9021, new_n9024);
or_8   g08648(new_n9024, new_n9008, new_n9025);
or_8   g08649(new_n9025, new_n9016, new_n9026);
and_8  g08650(new_n9026, new_n9013, new_n9027);
and_8  g08651(new_n9027, new_n8725, new_n9028);
nor_6  g08652(new_n9027, new_n8725, new_n9029);
or_8   g08653(new_n9029, new_n9028, new_n9030);
xor_4  g08654(new_n8695, new_n8693, new_n9031);
xor_4  g08655(new_n9023, new_n9001, new_n9032);
or_8   g08656(new_n9032, new_n9031, new_n9033);
or_8   g08657(new_n9023, new_n9021, new_n9034);
and_8  g08658(new_n9034, new_n9011, new_n9035);
xor_4  g08659(new_n9035, new_n9031, new_n9036);
xor_4  g08660(new_n8692, new_n8691, new_n9037);
and_8  g08661(new_n8999, new_n8990, new_n9038);
or_8   g08662(new_n9038, new_n9020, new_n9039);
and_8  g08663(new_n9039, new_n9037, new_n9040);
xor_4  g08664(new_n8690, new_n8689, new_n9041);
not_8  g08665(new_n9041, new_n9042);
nor_6  g08666(new_n8997, new_n8996, new_n9043);
or_8   g08667(new_n9043, new_n8998, new_n9044);
or_8   g08668(new_n9044, new_n9042, new_n9045);
not_8  g08669(new_n9045, new_n9046);
xor_4  g08670(new_n8997, new_n8996, new_n9047);
or_8   g08671(new_n9047, new_n9041, new_n9048);
and_8  g08672(new_n9048, new_n9045, new_n9049);
and_8  g08673(new_n8502, new_n8491, new_n9050);
and_8  g08674(new_n8532, new_n8503, new_n9051);
or_8   g08675(new_n9051, new_n9050, new_n9052);
and_8  g08676(new_n9052, new_n9049, new_n9053);
or_8   g08677(new_n9053, new_n9046, new_n9054);
not_8  g08678(new_n9037, new_n9055);
or_8   g08679(new_n9019, new_n9018, new_n9056);
and_8  g08680(new_n9056, new_n9000, new_n9057);
or_8   g08681(new_n9057, new_n9055, new_n9058);
or_8   g08682(new_n9039, new_n9037, new_n9059);
and_8  g08683(new_n9059, new_n9058, new_n9060);
and_8  g08684(new_n9060, new_n9054, new_n9061);
or_8   g08685(new_n9061, new_n9040, new_n9062);
or_8   g08686(new_n9062, new_n9036, new_n9063);
and_8  g08687(new_n9063, new_n9033, new_n9064);
or_8   g08688(new_n9064, new_n9030, new_n9065);
xor_4  g08689(new_n9027, new_n8725, new_n9066);
not_8  g08690(new_n9033, new_n9067);
not_8  g08691(new_n8693, new_n9068);
xor_4  g08692(new_n8695, new_n9068, new_n9069);
xor_4  g08693(new_n9035, new_n9069, new_n9070);
xor_4  g08694(new_n9047, new_n9042, new_n9071);
not_8  g08695(new_n9052, new_n9072);
or_8   g08696(new_n9072, new_n9071, new_n9073);
and_8  g08697(new_n9073, new_n9045, new_n9074);
and_8  g08698(new_n9057, new_n9055, new_n9075);
or_8   g08699(new_n9075, new_n9040, new_n9076);
or_8   g08700(new_n9076, new_n9074, new_n9077);
and_8  g08701(new_n9077, new_n9058, new_n9078);
and_8  g08702(new_n9078, new_n9070, new_n9079);
or_8   g08703(new_n9079, new_n9067, new_n9080_1);
or_8   g08704(new_n9080_1, new_n9066, new_n9081);
and_8  g08705(new_n9081, new_n9065, new_n9082);
nor_6  g08706(new_n9082, new_n8628, new_n9083);
xor_4  g08707(new_n9082, new_n8628, new_n9084);
xor_4  g08708(new_n8624, new_n8623, new_n9085);
xor_4  g08709(new_n9078, new_n9036, new_n9086);
or_8   g08710(new_n9086, new_n9085, new_n9087);
not_8  g08711(new_n9085, new_n9088);
xor_4  g08712(new_n9078, new_n9070, new_n9089);
and_8  g08713(new_n9089, new_n9088, new_n9090);
and_8  g08714(new_n9086, new_n9085, new_n9091);
or_8   g08715(new_n9091, new_n9090, new_n9092);
xor_4  g08716(new_n8622, new_n8621, new_n9093);
or_8   g08717(new_n9060, new_n9054, new_n9094);
and_8  g08718(new_n9094, new_n9077, new_n9095);
or_8   g08719(new_n9095, new_n9093, new_n9096);
not_8  g08720(new_n9096, new_n9097);
not_8  g08721(new_n9093, new_n9098);
and_8  g08722(new_n9076, new_n9074, new_n9099);
or_8   g08723(new_n9099, new_n9061, new_n9100);
or_8   g08724(new_n9100, new_n9098, new_n9101);
and_8  g08725(new_n9101, new_n9096, new_n9102);
xor_4  g08726(new_n8619, new_n8617, new_n9103);
or_8   g08727(new_n9052, new_n9049, new_n9104);
and_8  g08728(new_n9104, new_n9073, new_n9105);
or_8   g08729(new_n9105, new_n9103, new_n9106);
not_8  g08730(new_n9106, new_n9107);
and_8  g08731(new_n8487, new_n8477, new_n9108);
and_8  g08732(new_n8533, new_n8488, new_n9109);
or_8   g08733(new_n9109, new_n9108, new_n9110);
not_8  g08734(new_n9110, new_n9111_1);
not_8  g08735(new_n9103, new_n9112);
and_8  g08736(new_n9072, new_n9071, new_n9113);
or_8   g08737(new_n9113, new_n9053, new_n9114);
or_8   g08738(new_n9114, new_n9112, new_n9115);
and_8  g08739(new_n9115, new_n9106, new_n9116);
and_8  g08740(new_n9116, new_n9111_1, new_n9117);
or_8   g08741(new_n9117, new_n9107, new_n9118);
and_8  g08742(new_n9118, new_n9102, new_n9119);
nor_6  g08743(new_n9119, new_n9097, new_n9120);
or_8   g08744(new_n9120, new_n9092, new_n9121);
and_8  g08745(new_n9121, new_n9087, new_n9122);
and_8  g08746(new_n9122, new_n9084, new_n9123);
or_8   g08747(new_n9123, new_n9083, new_n9124);
and_8  g08748(new_n9080_1, new_n9066, new_n9125);
nor_6  g08749(new_n9125, new_n9028, new_n9126);
and_8  g08750(new_n8612, new_n8586, new_n9127);
and_8  g08751(new_n8626, new_n8613, new_n9128);
or_8   g08752(new_n9128, new_n9127, new_n9129);
or_8   g08753(new_n8601, new_n8600, new_n9130);
or_8   g08754(new_n8602, new_n8599, new_n9131);
and_8  g08755(new_n9131, new_n9130, new_n9132);
or_8   g08756(new_n8592, new_n8591, new_n9133);
or_8   g08757(new_n8593, new_n8590, new_n9134);
and_8  g08758(new_n9134, new_n9133, new_n9135);
nand_5 g08759(n9725, n5964, new_n9136);
xor_4  g08760(new_n9136, new_n9135, new_n9137_1);
xor_4  g08761(new_n9137_1, new_n9132, new_n9138);
xor_4  g08762(new_n9138, new_n9129, new_n9139);
not_8  g08763(new_n9139, new_n9140);
and_8  g08764(new_n8723, new_n8699, new_n9141);
not_8  g08765(new_n9141, new_n9142);
xor_4  g08766(new_n8723, new_n8698, new_n9143);
or_8   g08767(new_n9143, new_n8697, new_n9144);
and_8  g08768(new_n9144, new_n9142, new_n9145);
not_8  g08769(new_n8937, new_n9146);
or_8   g08770(new_n8961, new_n9146, new_n9147);
or_8   g08771(new_n9147, new_n9145, new_n9148);
xor_4  g08772(new_n8686, new_n8629, new_n9149);
and_8  g08773(new_n9149, new_n9068, new_n9150);
or_8   g08774(new_n9150, new_n8687, new_n9151);
and_8  g08775(new_n8724, new_n9151, new_n9152);
or_8   g08776(new_n9152, new_n9141, new_n9153);
nor_6  g08777(new_n8961, new_n9146, new_n9154);
or_8   g08778(new_n9154, new_n9153, new_n9155);
and_8  g08779(new_n9155, new_n9148, new_n9156);
not_8  g08780(new_n8817, new_n9157);
nor_6  g08781(new_n8842, new_n9157, new_n9158);
and_8  g08782(new_n8914, new_n8910, new_n9159);
not_8  g08783(new_n9159, new_n9160);
or_8   g08784(new_n8925, new_n8916, new_n9161);
and_8  g08785(new_n9161, new_n9160, new_n9162);
and_8  g08786(new_n8704, new_n8703, new_n9163);
or_8   g08787(new_n8704, new_n8703, new_n9164);
and_8  g08788(new_n9164, new_n8702, new_n9165);
or_8   g08789(new_n9165, new_n9163, new_n9166);
nand_5 g08790(n3986, n1478, new_n9167);
and_8  g08791(n9241, n6429, new_n9168);
and_8  g08792(n10022, n7965, new_n9169);
xor_4  g08793(new_n9169, new_n9168, new_n9170);
xor_4  g08794(new_n9170, new_n9167, new_n9171);
xnor_4 g08795(new_n9171, new_n9166, new_n9172);
xor_4  g08796(new_n9172, new_n9162, new_n9173);
or_8   g08797(new_n8922, new_n8921, new_n9174);
or_8   g08798(new_n8923, new_n8920, new_n9175);
nand_5 g08799(new_n9175, new_n9174, new_n9176);
not_8  g08800(new_n9176, new_n9177);
or_8   g08801(new_n8800, new_n8797, new_n9178);
and_8  g08802(new_n9178, new_n8798, new_n9179);
and_8  g08803(n11999, n7388, new_n9180);
nand_5 g08804(new_n9180, new_n9179, new_n9181);
and_8  g08805(new_n9180, new_n8826, new_n9182);
or_8   g08806(new_n9182, new_n9179, new_n9183);
and_8  g08807(new_n9183, new_n9181, new_n9184);
xor_4  g08808(new_n9184, new_n9177, new_n9185);
and_8  g08809(new_n8918, new_n8917, new_n9186);
nor_6  g08810(new_n8924, new_n8919, new_n9187);
or_8   g08811(new_n9187, new_n9186, new_n9188);
and_8  g08812(new_n8791, new_n8790, new_n9189_1);
or_8   g08813(new_n8791, new_n8790, new_n9190);
and_8  g08814(new_n9190, new_n8789, new_n9191);
or_8   g08815(new_n9191, new_n9189_1, new_n9192);
nand_5 g08816(n2530, n447, new_n9193);
and_8  g08817(n12777, n7690, new_n9194);
and_8  g08818(n8476, n1353, new_n9195_1);
xor_4  g08819(new_n9195_1, new_n9194, new_n9196);
xor_4  g08820(new_n9196, new_n9193, new_n9197);
xor_4  g08821(new_n9197, new_n9192, new_n9198);
xor_4  g08822(new_n9198, new_n9188, new_n9199);
or_8   g08823(new_n9199, new_n9185, new_n9200);
xor_4  g08824(new_n9184, new_n9176, new_n9201);
not_8  g08825(new_n9199, new_n9202);
or_8   g08826(new_n9202, new_n9201, new_n9203);
and_8  g08827(new_n9203, new_n9200, new_n9204);
and_8  g08828(n8759, n1198, new_n9205);
and_8  g08829(n11728, n10510, new_n9206);
xor_4  g08830(new_n9206, new_n9205, new_n9207);
and_8  g08831(n12489, n4499, new_n9208);
and_8  g08832(n10545, n6254, new_n9209);
xor_4  g08833(new_n9209, new_n9208, new_n9210);
and_8  g08834(n5331, n4436, new_n9211);
and_8  g08835(n12947, n2393, new_n9212);
xor_4  g08836(new_n9212, new_n9211, new_n9213);
xor_4  g08837(new_n9213, new_n9210, new_n9214);
xor_4  g08838(new_n9214, new_n9207, new_n9215);
and_8  g08839(n12648, n11967, new_n9216);
and_8  g08840(n7159, n3616, new_n9217);
and_8  g08841(n12709, n10644, new_n9218);
xor_4  g08842(new_n9218, new_n9217, new_n9219);
xor_4  g08843(new_n9219, new_n9216, new_n9220);
and_8  g08844(n8819, n8276, new_n9221);
and_8  g08845(n7730, n6776, new_n9222);
xor_4  g08846(new_n9222, new_n9221, new_n9223);
xor_4  g08847(new_n9223, new_n9220, new_n9224);
xor_4  g08848(new_n9224, new_n9215, new_n9225);
not_8  g08849(new_n9225, new_n9226);
or_8   g08850(new_n9226, new_n9204, new_n9227);
and_8  g08851(new_n9202, new_n9201, new_n9228);
and_8  g08852(new_n9199, new_n9185, new_n9229);
or_8   g08853(new_n9229, new_n9228, new_n9230);
or_8   g08854(new_n9225, new_n9230, new_n9231);
and_8  g08855(new_n9231, new_n9227, new_n9232);
xor_4  g08856(new_n9232, new_n9173, new_n9233);
nand_5 g08857(new_n8763, new_n8810, new_n9234);
and_8  g08858(new_n8819_1, new_n9234, new_n9235);
nand_5 g08859(n12705, n4370, new_n9236);
and_8  g08860(new_n8594, new_n8589, new_n9237);
and_8  g08861(new_n8604, new_n8595_1, new_n9238);
or_8   g08862(new_n9238, new_n9237, new_n9239);
and_8  g08863(new_n8805, new_n8801, new_n9240);
and_8  g08864(new_n8806, new_n8796, new_n9241_1);
or_8   g08865(new_n9241_1, new_n9240, new_n9242);
xor_4  g08866(new_n9242, new_n9239, new_n9243);
xor_4  g08867(new_n9243, new_n9236, new_n9244);
xor_4  g08868(new_n9244, new_n9235, new_n9245);
xor_4  g08869(new_n9245, new_n9233, new_n9246);
and_8  g08870(new_n9246, new_n9158, new_n9247);
or_8   g08871(new_n8842, new_n9157, new_n9248);
and_8  g08872(new_n9245, new_n9233, new_n9249);
nor_6  g08873(new_n9245, new_n9233, new_n9250);
or_8   g08874(new_n9250, new_n9249, new_n9251);
and_8  g08875(new_n9251, new_n9248, new_n9252);
or_8   g08876(new_n9252, new_n9247, new_n9253);
or_8   g08877(new_n9253, new_n9156, new_n9254);
and_8  g08878(new_n9154, new_n9153, new_n9255);
and_8  g08879(new_n9147, new_n9145, new_n9256);
or_8   g08880(new_n9256, new_n9255, new_n9257);
or_8   g08881(new_n9251, new_n9248, new_n9258);
or_8   g08882(new_n9246, new_n9158, new_n9259);
and_8  g08883(new_n9259, new_n9258, new_n9260);
or_8   g08884(new_n9260, new_n9257, new_n9261);
and_8  g08885(new_n9261, new_n9254, new_n9262);
xor_4  g08886(new_n9262, new_n9140, new_n9263);
and_8  g08887(new_n9013, new_n9014, new_n9264);
and_8  g08888(new_n8664, new_n8720, new_n9265);
and_8  g08889(new_n8722, new_n8718, new_n9266);
nor_6  g08890(new_n9266, new_n9265, new_n9267);
and_8  g08891(n11407, n10547, new_n9268);
and_8  g08892(n5320, n4312, new_n9269);
xor_4  g08893(new_n9269, new_n9268, new_n9270);
and_8  g08894(n12299, n8717, new_n9271);
and_8  g08895(n5857, n5760, new_n9272);
xor_4  g08896(new_n9272, new_n9271, new_n9273);
and_8  g08897(n12025, n11877, new_n9274);
and_8  g08898(n12000, n1097, new_n9275);
xor_4  g08899(new_n9275, new_n9274, new_n9276);
xor_4  g08900(new_n9276, new_n9273, new_n9277);
xor_4  g08901(new_n9277, new_n9270, new_n9278);
or_8   g08902(new_n8713, new_n8712, new_n9279);
or_8   g08903(new_n8714, new_n8711, new_n9280);
and_8  g08904(new_n9280, new_n9279, new_n9281);
and_8  g08905(n10990, n45, new_n9282);
xor_4  g08906(new_n9282, new_n9281, new_n9283);
xor_4  g08907(new_n9283, new_n9278, new_n9284);
nand_5 g08908(new_n8709, new_n8708, new_n9285);
or_8   g08909(new_n8715, new_n8710, new_n9286);
and_8  g08910(new_n9286, new_n9285, new_n9287);
and_8  g08911(n7436, n2433, new_n9288);
xor_4  g08912(new_n9288, new_n9287, new_n9289);
xor_4  g08913(new_n9289, new_n9284, new_n9290);
or_8   g08914(new_n8908, new_n8907, new_n9291);
or_8   g08915(new_n8909, new_n8906, new_n9292);
and_8  g08916(new_n9292, new_n9291, new_n9293);
or_8   g08917(new_n8642, new_n8700, new_n9294);
nand_5 g08918(new_n8706, new_n9294, new_n9295);
or_8   g08919(new_n8716, new_n8707, new_n9296);
and_8  g08920(new_n9296, new_n9295, new_n9297);
xor_4  g08921(new_n9297, new_n9293, new_n9298);
xor_4  g08922(new_n9298, new_n9290, new_n9299);
xor_4  g08923(new_n9299, new_n9267, new_n9300);
nand_5 g08924(new_n8881, new_n8930, new_n9301);
and_8  g08925(new_n8939, new_n9301, new_n9302);
and_8  g08926(new_n8787, new_n8786, new_n9303);
or_8   g08927(new_n8794, new_n9303, new_n9304);
and_8  g08928(n11892, n6441, new_n9305);
and_8  g08929(n11791, n5860, new_n9306);
xor_4  g08930(new_n9306, new_n9305, new_n9307);
and_8  g08931(n11257, n5212, new_n9308);
and_8  g08932(n6604, n5305, new_n9309);
xnor_4 g08933(new_n9309, new_n9308, new_n9310);
xor_4  g08934(new_n9310, new_n9307, new_n9311);
xor_4  g08935(new_n9311, new_n9304, new_n9312);
xor_4  g08936(new_n9312, new_n9302, new_n9313);
not_8  g08937(new_n9313, new_n9314);
xor_4  g08938(new_n9314, new_n9300, new_n9315);
or_8   g08939(new_n8597, new_n8596, new_n9316);
nand_5 g08940(new_n8603, new_n8598, new_n9317);
and_8  g08941(new_n9317, new_n9316, new_n9318);
not_8  g08942(new_n8608, new_n9319);
or_8   g08943(new_n8609, new_n9319, new_n9320);
or_8   g08944(new_n8611, new_n8605, new_n9321);
and_8  g08945(new_n9321, new_n9320, new_n9322);
xor_4  g08946(new_n9322, new_n9318, new_n9323);
not_8  g08947(new_n9323, new_n9324);
or_8   g08948(new_n9324, new_n9315, new_n9325);
xor_4  g08949(new_n9313, new_n9300, new_n9326);
or_8   g08950(new_n9323, new_n9326, new_n9327);
and_8  g08951(new_n9327, new_n9325, new_n9328);
and_8  g08952(new_n9328, new_n9264, new_n9329);
nor_6  g08953(new_n9328, new_n9264, new_n9330);
or_8   g08954(new_n9330, new_n9329, new_n9331);
or_8   g08955(new_n9331, new_n9263, new_n9332);
xor_4  g08956(new_n9262, new_n9139, new_n9333);
xor_4  g08957(new_n9328, new_n9264, new_n9334);
or_8   g08958(new_n9334, new_n9333, new_n9335);
and_8  g08959(new_n9335, new_n9332, new_n9336);
xor_4  g08960(new_n9336, new_n9126, new_n9337);
and_8  g08961(new_n9337, new_n9124, new_n9338);
or_8   g08962(new_n9082, new_n8628, new_n9339);
xor_4  g08963(new_n9082, new_n8627, new_n9340);
or_8   g08964(new_n9089, new_n9088, new_n9341);
and_8  g08965(new_n9341, new_n9087, new_n9342);
or_8   g08966(new_n9119, new_n9097, new_n9343);
and_8  g08967(new_n9343, new_n9342, new_n9344);
or_8   g08968(new_n9344, new_n9090, new_n9345);
or_8   g08969(new_n9345, new_n9340, new_n9346);
and_8  g08970(new_n9346, new_n9339, new_n9347);
or_8   g08971(new_n9125, new_n9028, new_n9348);
xor_4  g08972(new_n9336, new_n9348, new_n9349);
and_8  g08973(new_n9349, new_n9347, new_n9350);
or_8   g08974(new_n9350, new_n9338, n3287);
xor_4  g08975(new_n9120, new_n9342, n3339);
xnor_4 g08976(new_n4052, new_n4051, n3456);
nand_5 g08977(n6687, n4005, new_n9354);
and_8  g08978(n12720, n6770, new_n9355);
and_8  g08979(n9920, n2509, new_n9356);
and_8  g08980(n6038, n3627, new_n9357);
xor_4  g08981(new_n9357, new_n9356, new_n9358);
xnor_4 g08982(new_n9358, new_n9355, new_n9359);
and_8  g08983(n9920, n6038, new_n9360);
and_8  g08984(n12720, n4189, new_n9361);
or_8   g08985(new_n9361, new_n9360, new_n9362);
and_8  g08986(n6770, n2509, new_n9363);
xnor_4 g08987(new_n9361, new_n9360, new_n9364);
or_8   g08988(new_n9364, new_n9363, new_n9365);
and_8  g08989(new_n9365, new_n9362, new_n9366);
xor_4  g08990(new_n9366, new_n9359, new_n9367);
and_8  g08991(n2564, n2508, new_n9368);
and_8  g08992(n6770, n6038, new_n9369);
and_8  g08993(n4189, n2509, new_n9370);
or_8   g08994(new_n9370, new_n9369, new_n9371);
and_8  g08995(n12720, n2564, new_n9372);
nor_6  g08996(new_n9370, new_n9369, new_n9373);
and_8  g08997(new_n9370, new_n9369, new_n9374);
or_8   g08998(new_n9374, new_n9373, new_n9375);
or_8   g08999(new_n9375, new_n9372, new_n9376);
and_8  g09000(new_n9376, new_n9371, new_n9377);
and_8  g09001(new_n9377, new_n9368, new_n9378);
nor_6  g09002(new_n9364, new_n9363, new_n9379);
and_8  g09003(new_n9364, new_n9363, new_n9380);
or_8   g09004(new_n9380, new_n9379, new_n9381);
xor_4  g09005(new_n9377, new_n9368, new_n9382);
and_8  g09006(new_n9382, new_n9381, new_n9383);
or_8   g09007(new_n9383, new_n9378, new_n9384);
and_8  g09008(n2585, n2564, new_n9385);
and_8  g09009(n4189, n2508, new_n9386);
xor_4  g09010(new_n9386, new_n9385, new_n9387_1);
nor_6  g09011(new_n9387_1, new_n9384, new_n9388);
and_8  g09012(new_n9387_1, new_n9384, new_n9389);
or_8   g09013(new_n9389, new_n9388, new_n9390);
xor_4  g09014(new_n9390, new_n9367, new_n9391);
and_8  g09015(n6687, n2585, new_n9392);
and_8  g09016(n6687, n2508, new_n9393);
and_8  g09017(new_n9361, new_n377, new_n9394);
and_8  g09018(n6038, n4189, new_n9395);
and_8  g09019(n12720, n6687, new_n9396);
or_8   g09020(new_n9396, new_n9395, new_n9397);
and_8  g09021(n2564, n2509, new_n9398);
and_8  g09022(new_n9398, new_n9397, new_n9399);
or_8   g09023(new_n9399, new_n9394, new_n9400_1);
and_8  g09024(new_n9400_1, new_n9393, new_n9401);
xor_4  g09025(new_n9400_1, new_n9393, new_n9402);
xnor_4 g09026(new_n9375, new_n9372, new_n9403);
and_8  g09027(new_n9403, new_n9402, new_n9404);
or_8   g09028(new_n9404, new_n9401, new_n9405);
nor_6  g09029(new_n9405, new_n9392, new_n9406);
xnor_4 g09030(new_n9382, new_n9381, new_n9407);
xor_4  g09031(new_n9405, new_n9392, new_n9408);
and_8  g09032(new_n9408, new_n9407, new_n9409);
or_8   g09033(new_n9409, new_n9406, new_n9410);
xor_4  g09034(new_n9410, new_n9391, new_n9411);
or_8   g09035(new_n9411, new_n9354, new_n9412);
not_8  g09036(new_n9412, new_n9413);
xnor_4 g09037(new_n9403, new_n9402, new_n9414);
not_8  g09038(new_n9394, new_n9415);
nand_5 g09039(new_n9397, new_n9415, new_n9416);
not_8  g09040(new_n9416, new_n9417);
and_8  g09041(n6687, n2509, new_n9418);
and_8  g09042(n6038, n2564, new_n9419);
nand_5 g09043(new_n9419, new_n9418, new_n9420);
or_8   g09044(new_n9420, new_n9417, new_n9421);
or_8   g09045(new_n9421, new_n9414, new_n9422);
xor_4  g09046(new_n9408, new_n9407, new_n9423);
or_8   g09047(new_n9423, new_n9422, new_n9424);
not_8  g09048(new_n9424, new_n9425);
not_8  g09049(new_n9354, new_n9426);
not_8  g09050(new_n9367, new_n9427);
xor_4  g09051(new_n9390, new_n9427, new_n9428);
or_8   g09052(new_n9410, new_n9428, new_n9429);
nor_6  g09053(new_n9409, new_n9406, new_n9430);
or_8   g09054(new_n9430, new_n9391, new_n9431);
and_8  g09055(new_n9431, new_n9429, new_n9432);
xor_4  g09056(new_n9432, new_n9426, new_n9433);
and_8  g09057(new_n9433, new_n9425, new_n9434);
or_8   g09058(new_n9434, new_n9413, new_n9435);
not_8  g09059(new_n9429, new_n9436);
nor_6  g09060(new_n9358, new_n9355, new_n9437);
nor_6  g09061(new_n9366, new_n9359, new_n9438);
or_8   g09062(new_n9438, new_n9437, new_n9439);
and_8  g09063(n4005, n2564, new_n9440);
and_8  g09064(n4189, n2585, new_n9441);
and_8  g09065(n12706, n6687, new_n9442);
xnor_4 g09066(new_n9442, new_n9441, new_n9443);
xor_4  g09067(new_n9443, new_n9440, new_n9444);
xor_4  g09068(new_n9444, new_n9439, new_n9445);
and_8  g09069(new_n9357, new_n9356, new_n9446);
and_8  g09070(n6770, n2508, new_n9447);
xor_4  g09071(new_n9447, new_n9446, new_n9448);
and_8  g09072(n3627, n2509, new_n9449);
and_8  g09073(n12720, n9920, new_n9450);
and_8  g09074(n6038, n4516, new_n9451);
xnor_4 g09075(new_n9451, new_n9450, new_n9452);
xor_4  g09076(new_n9452, new_n9449, new_n9453);
xor_4  g09077(new_n9453, new_n9448, new_n9454);
xor_4  g09078(new_n9454, new_n9445, new_n9455);
not_8  g09079(new_n9389, new_n9456);
nand_5 g09080(new_n9386, new_n9385, new_n9457_1);
not_8  g09081(new_n9457_1, new_n9458);
or_8   g09082(new_n9390, new_n9367, new_n9459);
xor_4  g09083(new_n9459, new_n9458, new_n9460);
and_8  g09084(new_n9460, new_n9456, new_n9461);
or_8   g09085(new_n9461, new_n9455, new_n9462);
and_8  g09086(new_n9454, new_n9445, new_n9463);
nor_6  g09087(new_n9454, new_n9445, new_n9464);
or_8   g09088(new_n9464, new_n9463, new_n9465);
xor_4  g09089(new_n9459, new_n9457_1, new_n9466);
or_8   g09090(new_n9466, new_n9389, new_n9467);
or_8   g09091(new_n9467, new_n9465, new_n9468);
and_8  g09092(new_n9468, new_n9462, new_n9469);
xor_4  g09093(new_n9469, new_n9436, new_n9470);
xor_4  g09094(new_n9470, new_n9435, new_n9471);
and_8  g09095(n8336, n5105, new_n9472);
and_8  g09096(n10928, n7500, new_n9473);
and_8  g09097(n8336, n1209, new_n9474);
and_8  g09098(n7354, n6986, new_n9475);
or_8   g09099(new_n9475, new_n9474, new_n9476);
and_8  g09100(new_n9476, new_n9473, new_n9477);
and_8  g09101(new_n9475, new_n9474, new_n9478);
or_8   g09102(new_n9478, new_n9477, new_n9479);
xor_4  g09103(new_n9479, new_n9472, new_n9480);
and_8  g09104(n7500, n6986, new_n9481);
and_8  g09105(n7354, n2226, new_n9482);
and_8  g09106(n10928, n1209, new_n9483);
xor_4  g09107(new_n9483, new_n9482, new_n9484);
xor_4  g09108(new_n9484, new_n9481, new_n9485);
xnor_4 g09109(new_n9485, new_n9480, new_n9486);
xnor_4 g09110(new_n9475, new_n9474, new_n9487);
and_8  g09111(n10928, n7354, new_n9488);
and_8  g09112(n8336, n7500, new_n9489);
and_8  g09113(new_n9489, new_n9488, new_n9490);
nand_5 g09114(new_n9490, new_n9487, new_n9491);
or_8   g09115(new_n9491, new_n9486, new_n9492);
and_8  g09116(n8336, n4141, new_n9493);
and_8  g09117(new_n9479, new_n9472, new_n9494);
and_8  g09118(new_n9485, new_n9480, new_n9495);
or_8   g09119(new_n9495, new_n9494, new_n9496);
xnor_4 g09120(new_n9496, new_n9493, new_n9497);
and_8  g09121(n10928, n5105, new_n9498);
or_8   g09122(new_n9483, new_n9482, new_n9499);
and_8  g09123(new_n9483, new_n9482, new_n9500);
or_8   g09124(new_n9500, new_n9481, new_n9501);
and_8  g09125(new_n9501, new_n9499, new_n9502);
xor_4  g09126(new_n9502, new_n9498, new_n9503);
and_8  g09127(n6986, n1209, new_n9504);
and_8  g09128(n7354, n1094, new_n9505);
and_8  g09129(n7500, n2226, new_n9506);
xnor_4 g09130(new_n9506, new_n9505, new_n9507);
xnor_4 g09131(new_n9507, new_n9504, new_n9508);
xor_4  g09132(new_n9508, new_n9503, new_n9509);
xor_4  g09133(new_n9509, new_n9497, new_n9510);
nor_6  g09134(new_n9510, new_n9492, new_n9511);
and_8  g09135(n8336, n4928, new_n9512);
not_8  g09136(new_n9512, new_n9513);
and_8  g09137(n2226, n1209, new_n9514);
or_8   g09138(new_n9506, new_n9505, new_n9515);
or_8   g09139(new_n9507, new_n9504, new_n9516);
and_8  g09140(new_n9516, new_n9515, new_n9517);
and_8  g09141(new_n9517, new_n9514, new_n9518);
nor_6  g09142(new_n9517, new_n9514, new_n9519);
or_8   g09143(new_n9519, new_n9518, new_n9520);
and_8  g09144(n7500, n1094, new_n9521);
and_8  g09145(n10678, n7354, new_n9522);
xor_4  g09146(new_n9522, new_n9521, new_n9523);
not_8  g09147(new_n9523, new_n9524);
xor_4  g09148(new_n9524, new_n9520, new_n9525);
and_8  g09149(n10928, n4141, new_n9526);
and_8  g09150(n6986, n5105, new_n9527);
xor_4  g09151(new_n9527, new_n9526, new_n9528);
xor_4  g09152(new_n9528, new_n9525, new_n9529);
and_8  g09153(new_n9502, new_n9498, new_n9530);
and_8  g09154(new_n9508, new_n9503, new_n9531);
or_8   g09155(new_n9531, new_n9530, new_n9532);
and_8  g09156(new_n9532, new_n9529, new_n9533);
xor_4  g09157(new_n9523, new_n9520, new_n9534);
xor_4  g09158(new_n9528, new_n9534, new_n9535);
not_8  g09159(new_n9532, new_n9536);
and_8  g09160(new_n9536, new_n9535, new_n9537);
or_8   g09161(new_n9537, new_n9533, new_n9538);
or_8   g09162(new_n9496, new_n9493, new_n9539);
or_8   g09163(new_n9509, new_n9497, new_n9540);
and_8  g09164(new_n9540, new_n9539, new_n9541);
xor_4  g09165(new_n9541, new_n9538, new_n9542);
and_8  g09166(new_n9542, new_n9513, new_n9543);
nor_6  g09167(new_n9542, new_n9513, new_n9544);
or_8   g09168(new_n9544, new_n9543, new_n9545);
nor_6  g09169(new_n9545, new_n9511, new_n9546);
and_8  g09170(new_n9545, new_n9511, new_n9547);
or_8   g09171(new_n9547, new_n9546, new_n9548);
and_8  g09172(n11222, n7294, new_n9549);
and_8  g09173(n11222, n1980, new_n9550);
and_8  g09174(n8028, n5314, new_n9551);
and_8  g09175(new_n9551, new_n9550, new_n9552);
or_8   g09176(new_n9551, new_n9550, new_n9553);
and_8  g09177(n11153, n10848, new_n9554);
and_8  g09178(new_n9554, new_n9553, new_n9555);
or_8   g09179(new_n9555, new_n9552, new_n9556);
xor_4  g09180(new_n9556, new_n9549, new_n9557);
and_8  g09181(n10848, n5314, new_n9558);
and_8  g09182(n8028, n996, new_n9559);
and_8  g09183(n11153, n1980, new_n9560);
xor_4  g09184(new_n9560, new_n9559, new_n9561);
xor_4  g09185(new_n9561, new_n9558, new_n9562);
and_8  g09186(new_n9562, new_n9557, new_n9563);
nor_6  g09187(new_n9562, new_n9557, new_n9564);
or_8   g09188(new_n9564, new_n9563, new_n9565);
xnor_4 g09189(new_n9551, new_n9550, new_n9566);
and_8  g09190(n11153, n8028, new_n9567);
and_8  g09191(n11222, n10848, new_n9568);
and_8  g09192(new_n9568, new_n9567, new_n9569);
nand_5 g09193(new_n9569, new_n9566, new_n9570);
nor_6  g09194(new_n9570, new_n9565, new_n9571_1);
not_8  g09195(new_n9571_1, new_n9572);
and_8  g09196(new_n9556, new_n9549, new_n9573);
or_8   g09197(new_n9563, new_n9573, new_n9574);
nand_5 g09198(n12704, n11222, new_n9575);
not_8  g09199(new_n9575, new_n9576);
and_8  g09200(n11153, n7294, new_n9577);
or_8   g09201(new_n9560, new_n9559, new_n9578_1);
and_8  g09202(new_n9560, new_n9559, new_n9579);
or_8   g09203(new_n9579, new_n9558, new_n9580);
and_8  g09204(new_n9580, new_n9578_1, new_n9581);
xor_4  g09205(new_n9581, new_n9577, new_n9582);
and_8  g09206(n10848, n996, new_n9583_1);
and_8  g09207(n5314, n1980, new_n9584);
and_8  g09208(n8028, n5767, new_n9585);
xor_4  g09209(new_n9585, new_n9584, new_n9586);
xor_4  g09210(new_n9586, new_n9583_1, new_n9587);
and_8  g09211(new_n9587, new_n9582, new_n9588);
nor_6  g09212(new_n9587, new_n9582, new_n9589);
or_8   g09213(new_n9589, new_n9588, new_n9590);
xor_4  g09214(new_n9590, new_n9576, new_n9591);
xor_4  g09215(new_n9591, new_n9574, new_n9592);
or_8   g09216(new_n9592, new_n9572, new_n9593);
nand_5 g09217(n11222, n5814, new_n9594);
and_8  g09218(n1980, n996, new_n9595);
and_8  g09219(n8028, n5319, new_n9596);
and_8  g09220(n10848, n5767, new_n9597);
xor_4  g09221(new_n9597, new_n9596, new_n9598);
and_8  g09222(new_n9598, new_n9595, new_n9599);
nor_6  g09223(new_n9598, new_n9595, new_n9600);
or_8   g09224(new_n9600, new_n9599, new_n9601);
or_8   g09225(new_n9585, new_n9584, new_n9602);
and_8  g09226(new_n9585, new_n9584, new_n9603);
or_8   g09227(new_n9603, new_n9583_1, new_n9604);
and_8  g09228(new_n9604, new_n9602, new_n9605);
xor_4  g09229(new_n9605, new_n9601, new_n9606);
and_8  g09230(n12704, n11153, new_n9607);
and_8  g09231(n7294, n5314, new_n9608);
xor_4  g09232(new_n9608, new_n9607, new_n9609);
not_8  g09233(new_n9609, new_n9610);
or_8   g09234(new_n9610, new_n9606, new_n9611);
nand_5 g09235(new_n9604, new_n9602, new_n9612);
or_8   g09236(new_n9612, new_n9601, new_n9613);
xor_4  g09237(new_n9598, new_n9595, new_n9614);
or_8   g09238(new_n9605, new_n9614, new_n9615);
and_8  g09239(new_n9615, new_n9613, new_n9616);
or_8   g09240(new_n9609, new_n9616, new_n9617);
and_8  g09241(new_n9617, new_n9611, new_n9618);
and_8  g09242(new_n9581, new_n9577, new_n9619);
or_8   g09243(new_n9588, new_n9619, new_n9620);
and_8  g09244(new_n9620, new_n9618, new_n9621);
nor_6  g09245(new_n9620, new_n9618, new_n9622);
or_8   g09246(new_n9622, new_n9621, new_n9623);
and_8  g09247(new_n9590, new_n9575, new_n9624);
not_8  g09248(new_n9574, new_n9625);
xor_4  g09249(new_n9590, new_n9575, new_n9626);
and_8  g09250(new_n9626, new_n9625, new_n9627);
or_8   g09251(new_n9627, new_n9624, new_n9628);
or_8   g09252(new_n9628, new_n9623, new_n9629);
xor_4  g09253(new_n9620, new_n9618, new_n9630);
not_8  g09254(new_n9624, new_n9631);
or_8   g09255(new_n9591, new_n9574, new_n9632);
and_8  g09256(new_n9632, new_n9631, new_n9633);
or_8   g09257(new_n9633, new_n9630, new_n9634);
and_8  g09258(new_n9634, new_n9629, new_n9635);
xor_4  g09259(new_n9635, new_n9594, new_n9636);
or_8   g09260(new_n9636, new_n9593, new_n9637_1);
xor_4  g09261(new_n9626, new_n9574, new_n9638);
and_8  g09262(new_n9638, new_n9571_1, new_n9639);
not_8  g09263(new_n9594, new_n9640_1);
xor_4  g09264(new_n9635, new_n9640_1, new_n9641);
or_8   g09265(new_n9641, new_n9639, new_n9642);
and_8  g09266(new_n9642, new_n9637_1, new_n9643);
and_8  g09267(n12069, n2802, new_n9644);
and_8  g09268(n7891, n1564, new_n9645);
and_8  g09269(n12069, n533, new_n9646);
or_8   g09270(new_n9646, new_n9645, new_n9647);
and_8  g09271(n12391, n1512, new_n9648);
and_8  g09272(new_n9648, new_n9647, new_n9649);
and_8  g09273(new_n9646, new_n9645, new_n9650);
or_8   g09274(new_n9650, new_n9649, new_n9651);
xor_4  g09275(new_n9651, new_n9644, new_n9652);
and_8  g09276(n7891, n1512, new_n9653);
and_8  g09277(n7160, n1564, new_n9654);
and_8  g09278(n12391, n533, new_n9655);
nor_6  g09279(new_n9655, new_n9654, new_n9656);
and_8  g09280(new_n9655, new_n9654, new_n9657);
or_8   g09281(new_n9657, new_n9656, new_n9658);
nor_6  g09282(new_n9658, new_n9653, new_n9659);
and_8  g09283(new_n9658, new_n9653, new_n9660);
or_8   g09284(new_n9660, new_n9659, new_n9661);
and_8  g09285(new_n9661, new_n9652, new_n9662);
nor_6  g09286(new_n9661, new_n9652, new_n9663);
or_8   g09287(new_n9663, new_n9662, new_n9664);
xnor_4 g09288(new_n9646, new_n9645, new_n9665);
and_8  g09289(n12391, n1564, new_n9666);
and_8  g09290(n12069, n1512, new_n9667);
and_8  g09291(new_n9667, new_n9666, new_n9668);
nand_5 g09292(new_n9668, new_n9665, new_n9669);
nor_6  g09293(new_n9669, new_n9664, new_n9670);
not_8  g09294(new_n9670, new_n9671);
and_8  g09295(n12069, n6806, new_n9672);
and_8  g09296(n12391, n2802, new_n9673);
not_8  g09297(new_n9673, new_n9674);
or_8   g09298(new_n9659, new_n9656, new_n9675);
or_8   g09299(new_n9675, new_n9674, new_n9676);
or_8   g09300(new_n9655, new_n9654, new_n9677);
or_8   g09301(new_n9658, new_n9653, new_n9678);
and_8  g09302(new_n9678, new_n9677, new_n9679);
or_8   g09303(new_n9679, new_n9673, new_n9680);
and_8  g09304(new_n9680, new_n9676, new_n9681);
and_8  g09305(n7891, n533, new_n9682);
and_8  g09306(n4828, n1564, new_n9683);
and_8  g09307(n7160, n1512, new_n9684);
xor_4  g09308(new_n9684, new_n9683, new_n9685);
xor_4  g09309(new_n9685, new_n9682, new_n9686);
and_8  g09310(new_n9686, new_n9681, new_n9687);
and_8  g09311(new_n9679, new_n9673, new_n9688);
and_8  g09312(new_n9675, new_n9674, new_n9689);
or_8   g09313(new_n9689, new_n9688, new_n9690);
not_8  g09314(new_n9682, new_n9691);
xor_4  g09315(new_n9685, new_n9691, new_n9692);
and_8  g09316(new_n9692, new_n9690, new_n9693);
or_8   g09317(new_n9693, new_n9687, new_n9694);
xor_4  g09318(new_n9694, new_n9672, new_n9695);
and_8  g09319(new_n9651, new_n9644, new_n9696);
or_8   g09320(new_n9662, new_n9696, new_n9697);
xor_4  g09321(new_n9697, new_n9695, new_n9698);
or_8   g09322(new_n9698, new_n9671, new_n9699);
not_8  g09323(new_n9699, new_n9700);
nand_5 g09324(n12069, n5069, new_n9701);
not_8  g09325(new_n9701, new_n9702);
and_8  g09326(n7160, n533, new_n9703);
and_8  g09327(n2515, n1564, new_n9704);
and_8  g09328(n4828, n1512, new_n9705);
xor_4  g09329(new_n9705, new_n9704, new_n9706_1);
and_8  g09330(new_n9706_1, new_n9703, new_n9707);
nor_6  g09331(new_n9706_1, new_n9703, new_n9708);
or_8   g09332(new_n9708, new_n9707, new_n9709);
nor_6  g09333(new_n9684, new_n9683, new_n9710);
and_8  g09334(new_n9685, new_n9691, new_n9711);
or_8   g09335(new_n9711, new_n9710, new_n9712);
nor_6  g09336(new_n9712, new_n9709, new_n9713);
and_8  g09337(new_n9712, new_n9709, new_n9714);
or_8   g09338(new_n9714, new_n9713, new_n9715);
and_8  g09339(n7891, n2802, new_n9716);
and_8  g09340(n12391, n6806, new_n9717);
xor_4  g09341(new_n9717, new_n9716, new_n9718);
not_8  g09342(new_n9718, new_n9719);
or_8   g09343(new_n9719, new_n9715, new_n9720);
nor_6  g09344(new_n9714, new_n9713, new_n9721);
or_8   g09345(new_n9718, new_n9721, new_n9722);
and_8  g09346(new_n9722, new_n9720, new_n9723);
or_8   g09347(new_n9687, new_n9688, new_n9724);
and_8  g09348(new_n9724, new_n9723, new_n9725_1);
nor_6  g09349(new_n9724, new_n9723, new_n9726);
or_8   g09350(new_n9726, new_n9725_1, new_n9727);
not_8  g09351(new_n9672, new_n9728);
and_8  g09352(new_n9694, new_n9728, new_n9729);
xor_4  g09353(new_n9694, new_n9728, new_n9730);
not_8  g09354(new_n9697, new_n9731);
and_8  g09355(new_n9731, new_n9730, new_n9732);
or_8   g09356(new_n9732, new_n9729, new_n9733);
or_8   g09357(new_n9733, new_n9727, new_n9734);
xor_4  g09358(new_n9724, new_n9723, new_n9735);
nor_6  g09359(new_n9693, new_n9687, new_n9736);
or_8   g09360(new_n9736, new_n9672, new_n9737);
or_8   g09361(new_n9697, new_n9695, new_n9738);
and_8  g09362(new_n9738, new_n9737, new_n9739);
or_8   g09363(new_n9739, new_n9735, new_n9740);
and_8  g09364(new_n9740, new_n9734, new_n9741);
or_8   g09365(new_n9741, new_n9702, new_n9742);
and_8  g09366(new_n9739, new_n9735, new_n9743);
and_8  g09367(new_n9733, new_n9727, new_n9744);
or_8   g09368(new_n9744, new_n9743, new_n9745);
or_8   g09369(new_n9745, new_n9701, new_n9746);
and_8  g09370(new_n9746, new_n9742, new_n9747);
xor_4  g09371(new_n9747, new_n9700, new_n9748);
or_8   g09372(new_n9748, new_n9643, new_n9749);
and_8  g09373(new_n9641, new_n9639, new_n9750);
and_8  g09374(new_n9636, new_n9593, new_n9751);
or_8   g09375(new_n9751, new_n9750, new_n9752);
xor_4  g09376(new_n9747, new_n9699, new_n9753);
or_8   g09377(new_n9753, new_n9752, new_n9754);
and_8  g09378(new_n9754, new_n9749, new_n9755);
or_8   g09379(new_n9638, new_n9571_1, new_n9756_1);
and_8  g09380(new_n9756_1, new_n9593, new_n9757);
and_8  g09381(new_n9669, new_n9664, new_n9758);
or_8   g09382(new_n9758, new_n9670, new_n9759);
and_8  g09383(new_n9570, new_n9565, new_n9760);
or_8   g09384(new_n9760, new_n9571_1, new_n9761);
and_8  g09385(new_n9761, new_n9759, new_n9762);
not_8  g09386(new_n9762, new_n9763_1);
not_8  g09387(new_n9648, new_n9764);
or_8   g09388(new_n9764, new_n380, new_n9765);
and_8  g09389(new_n9765, new_n9665, new_n9766);
not_8  g09390(new_n380, new_n9767_1);
and_8  g09391(new_n9649, new_n9767_1, new_n9768);
or_8   g09392(new_n9768, new_n9766, new_n9769);
not_8  g09393(new_n9554, new_n9770);
or_8   g09394(new_n9770, new_n379, new_n9771);
and_8  g09395(new_n9771, new_n9566, new_n9772);
nor_6  g09396(new_n9770, new_n379, new_n9773);
and_8  g09397(new_n9773, new_n9553, new_n9774);
or_8   g09398(new_n9774, new_n9772, new_n9775);
nor_6  g09399(new_n9775, new_n9769, new_n9776);
and_8  g09400(new_n380, new_n379, new_n9777);
xor_4  g09401(new_n9568, new_n9567, new_n9778);
or_8   g09402(new_n9778, new_n9777, new_n9779);
xor_4  g09403(new_n9778, new_n9777, new_n9780);
not_8  g09404(new_n9780, new_n9781);
xor_4  g09405(new_n9667, new_n9666, new_n9782);
or_8   g09406(new_n9782, new_n9781, new_n9783);
and_8  g09407(new_n9783, new_n9779, new_n9784);
xor_4  g09408(new_n9775, new_n9769, new_n9785);
and_8  g09409(new_n9785, new_n9784, new_n9786);
or_8   g09410(new_n9786, new_n9776, new_n9787);
xor_4  g09411(new_n9669, new_n9664, new_n9788);
xor_4  g09412(new_n9570, new_n9565, new_n9789);
and_8  g09413(new_n9789, new_n9788, new_n9790);
or_8   g09414(new_n9790, new_n9762, new_n9791);
or_8   g09415(new_n9791, new_n9787, new_n9792);
and_8  g09416(new_n9792, new_n9763_1, new_n9793);
nor_6  g09417(new_n9793, new_n9757, new_n9794);
not_8  g09418(new_n9794, new_n9795);
xor_4  g09419(new_n9698, new_n9671, new_n9796);
and_8  g09420(new_n9793, new_n9757, new_n9797);
or_8   g09421(new_n9797, new_n9794, new_n9798);
or_8   g09422(new_n9798, new_n9796, new_n9799);
and_8  g09423(new_n9799, new_n9795, new_n9800);
xor_4  g09424(new_n9800, new_n9755, new_n9801);
and_8  g09425(new_n9801, new_n9548, new_n9802);
not_8  g09426(new_n9802, new_n9803);
nor_6  g09427(new_n9801, new_n9548, new_n9804);
or_8   g09428(new_n9804, new_n9802, new_n9805);
xor_4  g09429(new_n9510, new_n9492, new_n9806);
not_8  g09430(new_n9806, new_n9807);
xor_4  g09431(new_n9698, new_n9670, new_n9808);
xor_4  g09432(new_n9793, new_n9757, new_n9809);
or_8   g09433(new_n9809, new_n9808, new_n9810);
and_8  g09434(new_n9810, new_n9799, new_n9811);
or_8   g09435(new_n9811, new_n9807, new_n9812);
and_8  g09436(new_n9809, new_n9808, new_n9813);
and_8  g09437(new_n9798, new_n9796, new_n9814);
or_8   g09438(new_n9814, new_n9813, new_n9815);
and_8  g09439(new_n9815, new_n9806, new_n9816);
and_8  g09440(new_n9811, new_n9807, new_n9817);
or_8   g09441(new_n9817, new_n9816, new_n9818);
xnor_4 g09442(new_n9491, new_n9486, new_n9819);
xor_4  g09443(new_n9791, new_n9787, new_n9820_1);
nor_6  g09444(new_n9820_1, new_n9819, new_n9821);
xor_4  g09445(new_n9820_1, new_n9819, new_n9822);
xor_4  g09446(new_n9785, new_n9784, new_n9823);
not_8  g09447(new_n378, new_n9824);
nand_5 g09448(new_n9473, new_n9824, new_n9825);
or_8   g09449(new_n9825, new_n9476, new_n9826);
not_8  g09450(new_n9825, new_n9827);
or_8   g09451(new_n9827, new_n9487, new_n9828);
and_8  g09452(new_n9828, new_n9826, new_n9829);
not_8  g09453(new_n9829, new_n9830);
or_8   g09454(new_n9830, new_n9823, new_n9831);
xor_4  g09455(new_n9829, new_n9823, new_n9832);
xor_4  g09456(new_n9782, new_n9780, new_n9833);
xor_4  g09457(new_n9489, new_n9488, new_n9834);
and_8  g09458(new_n9834, new_n9833, new_n9835);
and_8  g09459(new_n381_1, new_n378, new_n9836);
xor_4  g09460(new_n9834, new_n9833, new_n9837);
and_8  g09461(new_n9837, new_n9836, new_n9838);
or_8   g09462(new_n9838, new_n9835, new_n9839);
or_8   g09463(new_n9839, new_n9832, new_n9840);
and_8  g09464(new_n9840, new_n9831, new_n9841);
and_8  g09465(new_n9841, new_n9822, new_n9842);
or_8   g09466(new_n9842, new_n9821, new_n9843);
not_8  g09467(new_n9843, new_n9844);
or_8   g09468(new_n9844, new_n9818, new_n9845);
and_8  g09469(new_n9845, new_n9812, new_n9846);
or_8   g09470(new_n9846, new_n9805, new_n9847);
and_8  g09471(new_n9847, new_n9803, new_n9848);
nor_6  g09472(new_n9537, new_n9533, new_n9849);
and_8  g09473(new_n9541, new_n9849, new_n9850);
nor_6  g09474(new_n9524, new_n9520, new_n9851);
or_8   g09475(new_n9851, new_n9518, new_n9852);
and_8  g09476(n10928, n4928, new_n9853);
and_8  g09477(n6986, n4141, new_n9854);
and_8  g09478(n8336, n8236, new_n9855);
xnor_4 g09479(new_n9855, new_n9854, new_n9856);
xor_4  g09480(new_n9856, new_n9853, new_n9857);
xor_4  g09481(new_n9857, new_n9852, new_n9858);
and_8  g09482(new_n9522, new_n9521, new_n9859);
and_8  g09483(n5105, n2226, new_n9860);
xnor_4 g09484(new_n9860, new_n9859, new_n9861);
and_8  g09485(n10678, n7500, new_n9862);
and_8  g09486(n7354, n7320, new_n9863);
and_8  g09487(n1209, n1094, new_n9864);
xnor_4 g09488(new_n9864, new_n9863, new_n9865);
xor_4  g09489(new_n9865, new_n9862, new_n9866);
xor_4  g09490(new_n9866, new_n9861, new_n9867);
xor_4  g09491(new_n9867, new_n9858, new_n9868);
nand_5 g09492(new_n9528, new_n9525, new_n9869);
nand_5 g09493(new_n9527, new_n9526, new_n9870);
not_8  g09494(new_n9870, new_n9871);
and_8  g09495(new_n9533, new_n9871, new_n9872);
or_8   g09496(new_n9536, new_n9535, new_n9873);
and_8  g09497(new_n9873, new_n9870, new_n9874);
or_8   g09498(new_n9874, new_n9872, new_n9875);
and_8  g09499(new_n9875, new_n9869, new_n9876);
xor_4  g09500(new_n9876, new_n9868, new_n9877);
xor_4  g09501(new_n9877, new_n9850, new_n9878);
not_8  g09502(new_n9543, new_n9879);
or_8   g09503(new_n9545, new_n9511, new_n9880);
and_8  g09504(new_n9880, new_n9879, new_n9881);
and_8  g09505(new_n9881, new_n9878, new_n9882);
nor_6  g09506(new_n9881, new_n9878, new_n9883);
nor_6  g09507(new_n9883, new_n9882, new_n9884);
not_8  g09508(new_n9613, new_n9885);
or_8   g09509(new_n9885, new_n9599, new_n9886);
and_8  g09510(n11153, n5814, new_n9887);
and_8  g09511(n12704, n5314, new_n9888);
and_8  g09512(n11222, n4903, new_n9889);
xnor_4 g09513(new_n9889, new_n9888, new_n9890);
xor_4  g09514(new_n9890, new_n9887, new_n9891);
xor_4  g09515(new_n9891, new_n9886, new_n9892);
and_8  g09516(new_n9597, new_n9596, new_n9893);
and_8  g09517(n7294, n996, new_n9894);
xor_4  g09518(new_n9894, new_n9893, new_n9895);
and_8  g09519(n10848, n5319, new_n9896);
not_8  g09520(new_n9896, new_n9897);
and_8  g09521(n5767, n1980, new_n9898);
and_8  g09522(n9457, n8028, new_n9899);
xnor_4 g09523(new_n9899, new_n9898, new_n9900);
xor_4  g09524(new_n9900, new_n9897, new_n9901);
xor_4  g09525(new_n9901, new_n9895, new_n9902);
xor_4  g09526(new_n9902, new_n9892, new_n9903);
nand_5 g09527(new_n9608, new_n9607, new_n9904);
xor_4  g09528(new_n9621, new_n9904, new_n9905);
and_8  g09529(new_n9905, new_n9611, new_n9906);
nor_6  g09530(new_n9906, new_n9903, new_n9907);
and_8  g09531(new_n9906, new_n9903, new_n9908);
or_8   g09532(new_n9908, new_n9907, new_n9909);
or_8   g09533(new_n9909, new_n9629, new_n9910);
not_8  g09534(new_n9910, new_n9911);
and_8  g09535(new_n9909, new_n9629, new_n9912);
or_8   g09536(new_n9912, new_n9911, new_n9913);
nand_5 g09537(new_n9635, new_n9640_1, new_n9914);
and_8  g09538(new_n9637_1, new_n9914, new_n9915);
nor_6  g09539(new_n9915, new_n9913, new_n9916);
and_8  g09540(new_n9915, new_n9913, new_n9917);
or_8   g09541(new_n9917, new_n9916, new_n9918);
not_8  g09542(new_n9720, new_n9919);
and_8  g09543(new_n9717, new_n9716, new_n9920_1);
xor_4  g09544(new_n9725_1, new_n9920_1, new_n9921);
or_8   g09545(new_n9921, new_n9919, new_n9922);
and_8  g09546(new_n9705, new_n9704, new_n9923);
and_8  g09547(n7160, n2802, new_n9924);
xnor_4 g09548(new_n9924, new_n9923, new_n9925);
and_8  g09549(n2515, n1512, new_n9926);
and_8  g09550(n1564, n1199, new_n9927);
and_8  g09551(n4828, n533, new_n9928);
xnor_4 g09552(new_n9928, new_n9927, new_n9929);
xor_4  g09553(new_n9929, new_n9926, new_n9930);
xnor_4 g09554(new_n9930, new_n9925, new_n9931);
nor_6  g09555(new_n9713, new_n9707, new_n9932);
and_8  g09556(n12391, n5069, new_n9933);
and_8  g09557(n7891, n6806, new_n9934);
and_8  g09558(n12069, n12044, new_n9935);
xnor_4 g09559(new_n9935, new_n9934, new_n9936);
xor_4  g09560(new_n9936, new_n9933, new_n9937);
xor_4  g09561(new_n9937, new_n9932, new_n9938_1);
nor_6  g09562(new_n9938_1, new_n9931, new_n9939);
and_8  g09563(new_n9938_1, new_n9931, new_n9940);
or_8   g09564(new_n9940, new_n9939, new_n9941);
xor_4  g09565(new_n9941, new_n9922, new_n9942);
and_8  g09566(new_n9942, new_n9743, new_n9943);
and_8  g09567(new_n9941, new_n9922, new_n9944);
nor_6  g09568(new_n9941, new_n9922, new_n9945);
or_8   g09569(new_n9945, new_n9944, new_n9946);
and_8  g09570(new_n9946, new_n9734, new_n9947);
or_8   g09571(new_n9947, new_n9943, new_n9948);
and_8  g09572(new_n9745, new_n9701, new_n9949);
or_8   g09573(new_n9949, new_n9699, new_n9950);
and_8  g09574(new_n9950, new_n9746, new_n9951);
xor_4  g09575(new_n9951, new_n9948, new_n9952);
and_8  g09576(new_n9753, new_n9752, new_n9953);
and_8  g09577(new_n9748, new_n9643, new_n9954);
or_8   g09578(new_n9954, new_n9953, new_n9955);
or_8   g09579(new_n9800, new_n9955, new_n9956_1);
and_8  g09580(new_n9956_1, new_n9749, new_n9957);
or_8   g09581(new_n9957, new_n9952, new_n9958);
nor_6  g09582(new_n9951, new_n9948, new_n9959);
and_8  g09583(new_n9951, new_n9948, new_n9960);
or_8   g09584(new_n9960, new_n9959, new_n9961);
or_8   g09585(new_n9813, new_n9794, new_n9962);
and_8  g09586(new_n9962, new_n9755, new_n9963);
or_8   g09587(new_n9963, new_n9953, new_n9964);
or_8   g09588(new_n9964, new_n9961, new_n9965);
and_8  g09589(new_n9965, new_n9958, new_n9966);
and_8  g09590(new_n9966, new_n9918, new_n9967);
nor_6  g09591(new_n9966, new_n9918, new_n9968);
or_8   g09592(new_n9968, new_n9967, new_n9969);
or_8   g09593(new_n9969, new_n9884, new_n9970);
or_8   g09594(new_n9883, new_n9882, new_n9971);
xor_4  g09595(new_n9966, new_n9918, new_n9972);
or_8   g09596(new_n9972, new_n9971, new_n9973);
and_8  g09597(new_n9973, new_n9970, new_n9974);
and_8  g09598(new_n9974, new_n9848, new_n9975);
nor_6  g09599(new_n9846, new_n9805, new_n9976);
or_8   g09600(new_n9976, new_n9802, new_n9977);
and_8  g09601(new_n9972, new_n9971, new_n9978);
and_8  g09602(new_n9969, new_n9884, new_n9979);
or_8   g09603(new_n9979, new_n9978, new_n9980);
and_8  g09604(new_n9980, new_n9977, new_n9981);
or_8   g09605(new_n9981, new_n9975, new_n9982);
or_8   g09606(new_n9982, new_n9471, new_n9983);
xor_4  g09607(new_n9433, new_n9425, new_n9984);
xor_4  g09608(new_n9423, new_n9422, new_n9985);
or_8   g09609(new_n9815, new_n9806, new_n9986);
and_8  g09610(new_n9986, new_n9812, new_n9987);
or_8   g09611(new_n9843, new_n9987, new_n9988);
and_8  g09612(new_n9988, new_n9845, new_n9989);
or_8   g09613(new_n9989, new_n9985, new_n9990);
xor_4  g09614(new_n9421, new_n9414, new_n9991);
not_8  g09615(new_n9991, new_n9992);
nor_6  g09616(new_n9841, new_n9822, new_n9993);
or_8   g09617(new_n9993, new_n9842, new_n9994);
and_8  g09618(new_n9994, new_n9992, new_n9995);
not_8  g09619(new_n9995, new_n9996);
not_8  g09620(new_n9842, new_n9997);
or_8   g09621(new_n9841, new_n9822, new_n9998);
and_8  g09622(new_n9998, new_n9997, new_n9999);
and_8  g09623(new_n9999, new_n9991, new_n10000);
or_8   g09624(new_n10000, new_n9995, new_n10001);
xor_4  g09625(new_n9839, new_n9832, new_n10002);
not_8  g09626(new_n377, new_n10003);
and_8  g09627(new_n9398, new_n10003, new_n10004);
or_8   g09628(new_n10004, new_n9417, new_n10005);
nand_5 g09629(new_n10004, new_n9397, new_n10006);
nand_5 g09630(new_n10006, new_n10005, new_n10007);
nand_5 g09631(new_n10007, new_n10002, new_n10008);
not_8  g09632(new_n10007, new_n10009);
xor_4  g09633(new_n10009, new_n10002, new_n10010);
and_8  g09634(new_n382, new_n377, new_n10011);
xor_4  g09635(new_n9419, new_n9418, new_n10012);
or_8   g09636(new_n10012, new_n10011, new_n10013);
xor_4  g09637(new_n9837, new_n9836, new_n10014);
xnor_4 g09638(new_n10012, new_n10011, new_n10015);
or_8   g09639(new_n10015, new_n10014, new_n10016);
and_8  g09640(new_n10016, new_n10013, new_n10017);
or_8   g09641(new_n10017, new_n10010, new_n10018);
and_8  g09642(new_n10018, new_n10008, new_n10019);
or_8   g09643(new_n10019, new_n10001, new_n10020);
and_8  g09644(new_n10020, new_n9996, new_n10021);
not_8  g09645(new_n9985, new_n10022_1);
and_8  g09646(new_n9843, new_n9987, new_n10023);
and_8  g09647(new_n9844, new_n9818, new_n10024);
or_8   g09648(new_n10024, new_n10023, new_n10025);
and_8  g09649(new_n10025, new_n10022_1, new_n10026);
and_8  g09650(new_n9989, new_n9985, new_n10027);
or_8   g09651(new_n10027, new_n10026, new_n10028);
or_8   g09652(new_n10028, new_n10021, new_n10029);
and_8  g09653(new_n10029, new_n9990, new_n10030);
or_8   g09654(new_n10030, new_n9984, new_n10031);
xor_4  g09655(new_n9846, new_n9805, new_n10032);
not_8  g09656(new_n9984, new_n10033);
xor_4  g09657(new_n10030, new_n10033, new_n10034);
or_8   g09658(new_n10034, new_n10032, new_n10035);
and_8  g09659(new_n10035, new_n10031, new_n10036);
not_8  g09660(new_n9471, new_n10037);
or_8   g09661(new_n9980, new_n9977, new_n10038);
or_8   g09662(new_n9974, new_n9848, new_n10039);
and_8  g09663(new_n10039, new_n10038, new_n10040);
and_8  g09664(new_n10040, new_n10037, new_n10041);
and_8  g09665(new_n9982, new_n9471, new_n10042);
or_8   g09666(new_n10042, new_n10041, new_n10043);
or_8   g09667(new_n10043, new_n10036, new_n10044);
and_8  g09668(new_n10044, new_n9983, new_n10045);
not_8  g09669(new_n9958, new_n10046);
or_8   g09670(new_n9967, new_n10046, new_n10047);
or_8   g09671(new_n9975, new_n9978, new_n10048);
or_8   g09672(new_n10048, new_n10047, new_n10049);
not_8  g09673(new_n10047, new_n10050);
and_8  g09674(new_n10038, new_n9970, new_n10051);
or_8   g09675(new_n10051, new_n10050, new_n10052);
and_8  g09676(new_n10052, new_n10049, new_n10053);
and_8  g09677(new_n9877, new_n9850, new_n10054);
or_8   g09678(new_n9882, new_n10054, new_n10055);
and_8  g09679(new_n9725_1, new_n9920_1, new_n10056);
nor_6  g09680(new_n9944, new_n10056, new_n10057);
nand_5 g09681(new_n9894, new_n9893, new_n10058);
nand_5 g09682(new_n9901, new_n9895, new_n10059);
and_8  g09683(new_n10059, new_n10058, new_n10060);
and_8  g09684(new_n9928, new_n9927, new_n10061);
or_8   g09685(new_n9928, new_n9927, new_n10062);
and_8  g09686(new_n10062, new_n9926, new_n10063);
or_8   g09687(new_n10063, new_n10061, new_n10064);
xor_4  g09688(new_n10064, new_n10060, new_n10065);
and_8  g09689(n8028, n4817, new_n10066);
and_8  g09690(n7523, n7354, new_n10067);
xor_4  g09691(new_n10067, new_n10066, new_n10068);
and_8  g09692(n10848, n9457, new_n10069);
and_8  g09693(n11222, n1906, new_n10070);
xor_4  g09694(new_n10070, new_n10069, new_n10071);
and_8  g09695(n6986, n4928, new_n10072);
and_8  g09696(n4141, n2226, new_n10073);
xor_4  g09697(new_n10073, new_n10072, new_n10074);
xnor_4 g09698(new_n10074, new_n10071, new_n10075);
xor_4  g09699(new_n10075, new_n10068, new_n10076);
and_8  g09700(new_n9451, new_n9450, new_n10077);
or_8   g09701(new_n9451, new_n9450, new_n10078);
and_8  g09702(new_n10078, new_n9449, new_n10079);
or_8   g09703(new_n10079, new_n10077, new_n10080);
nand_5 g09704(n4516, n2509, new_n10081);
and_8  g09705(n12704, n996, new_n10082);
and_8  g09706(n12720, n3627, new_n10083);
xor_4  g09707(new_n10083, new_n10082, new_n10084);
xor_4  g09708(new_n10084, new_n10081, new_n10085);
xor_4  g09709(new_n10085, new_n10080, new_n10086);
xor_4  g09710(new_n10086, new_n10076, new_n10087);
nand_5 g09711(n2515, n533, new_n10088);
and_8  g09712(n1512, n1199, new_n10089);
and_8  g09713(n12391, n12044, new_n10090);
xor_4  g09714(new_n10090, new_n10089, new_n10091);
xor_4  g09715(new_n10091, new_n10088, new_n10092);
xor_4  g09716(new_n10092, new_n10087, new_n10093);
xor_4  g09717(new_n10093, new_n10065, new_n10094);
not_8  g09718(new_n9891, new_n10095);
or_8   g09719(new_n10095, new_n9886, new_n10096);
or_8   g09720(new_n9902, new_n9892, new_n10097);
and_8  g09721(new_n10097, new_n10096, new_n10098);
or_8   g09722(new_n9899, new_n9898, new_n10099);
or_8   g09723(new_n9900, new_n9896, new_n10100);
and_8  g09724(new_n10100, new_n10099, new_n10101);
and_8  g09725(n12069, n5694, new_n10102);
and_8  g09726(n11153, n4903, new_n10103);
xor_4  g09727(new_n10103, new_n10102, new_n10104);
and_8  g09728(n7294, n5767, new_n10105);
and_8  g09729(n8336, n783, new_n10106);
xor_4  g09730(new_n10106, new_n10105, new_n10107);
xnor_4 g09731(new_n10107, new_n10104, new_n10108);
xor_4  g09732(new_n10108, new_n10101, new_n10109);
and_8  g09733(n4189, n4005, new_n10110);
and_8  g09734(n5814, n5314, new_n10111);
xor_4  g09735(new_n10111, new_n10110, new_n10112);
xor_4  g09736(new_n10112, new_n10109, new_n10113);
xor_4  g09737(new_n10113, new_n10098, new_n10114);
xor_4  g09738(new_n10114, new_n10094, new_n10115);
xor_4  g09739(new_n10115, new_n10057, new_n10116);
xor_4  g09740(new_n10116, new_n10055, new_n10117);
not_8  g09741(new_n10117, new_n10118);
or_8   g09742(new_n9959, new_n9943, new_n10119);
not_8  g09743(new_n10119, new_n10120);
or_8   g09744(new_n9915, new_n9913, new_n10121);
and_8  g09745(new_n10121, new_n9910, new_n10122);
and_8  g09746(new_n9444, new_n9439, new_n10123);
or_8   g09747(new_n9463, new_n10123, new_n10124);
or_8   g09748(new_n9442, new_n9441, new_n10125);
or_8   g09749(new_n9443, new_n9440, new_n10126);
and_8  g09750(new_n10126, new_n10125, new_n10127);
xor_4  g09751(new_n10127, new_n10124, new_n10128);
or_8   g09752(new_n9889, new_n9888, new_n10129);
or_8   g09753(new_n9890, new_n9887, new_n10130);
and_8  g09754(new_n10130, new_n10129, new_n10131);
or_8   g09755(new_n9935, new_n9934, new_n10132);
or_8   g09756(new_n9936, new_n9933, new_n10133);
and_8  g09757(new_n10133, new_n10132, new_n10134);
xor_4  g09758(new_n10134, new_n10131, new_n10135);
xor_4  g09759(new_n10135, new_n10128, new_n10136);
or_8   g09760(new_n10136, new_n10122, new_n10137);
or_8   g09761(new_n9916, new_n9911, new_n10138);
not_8  g09762(new_n10136, new_n10139);
or_8   g09763(new_n10139, new_n10138, new_n10140);
and_8  g09764(new_n10140, new_n10137, new_n10141);
and_8  g09765(new_n9469, new_n9436, new_n10142);
not_8  g09766(new_n10142, new_n10143);
xor_4  g09767(new_n9432, new_n9354, new_n10144);
or_8   g09768(new_n10144, new_n9424, new_n10145);
and_8  g09769(new_n10145, new_n9412, new_n10146);
xor_4  g09770(new_n9469, new_n9429, new_n10147);
or_8   g09771(new_n10147, new_n10146, new_n10148);
and_8  g09772(new_n10148, new_n10143, new_n10149);
and_8  g09773(new_n9937, new_n9932, new_n10150);
or_8   g09774(new_n9940, new_n10150, new_n10151);
and_8  g09775(n6578, n1564, new_n10152);
xor_4  g09776(new_n10152, new_n10151, new_n10153);
or_8   g09777(new_n10153, new_n10149, new_n10154);
and_8  g09778(new_n9470, new_n9435, new_n10155);
or_8   g09779(new_n10155, new_n10142, new_n10156);
not_8  g09780(new_n10153, new_n10157);
or_8   g09781(new_n10157, new_n10156, new_n10158);
and_8  g09782(new_n10158, new_n10154, new_n10159);
xor_4  g09783(new_n10159, new_n10141, new_n10160);
not_8  g09784(new_n9904, new_n10161);
nand_5 g09785(new_n9621, new_n10161, new_n10162);
or_8   g09786(new_n9906, new_n9903, new_n10163);
and_8  g09787(new_n10163, new_n10162, new_n10164);
nand_5 g09788(new_n9860, new_n9859, new_n10165);
or_8   g09789(new_n9866, new_n9861, new_n10166);
and_8  g09790(new_n10166, new_n10165, new_n10167);
or_8   g09791(new_n9855, new_n9854, new_n10168);
or_8   g09792(new_n9856, new_n9853, new_n10169);
and_8  g09793(new_n10169, new_n10168, new_n10170);
nand_5 g09794(n5319, n1980, new_n10171);
and_8  g09795(n9920, n2508, new_n10172);
and_8  g09796(n10678, n1209, new_n10173);
xor_4  g09797(new_n10173, new_n10172, new_n10174_1);
xor_4  g09798(new_n10174_1, new_n10171, new_n10175);
xnor_4 g09799(new_n10175, new_n10170, new_n10176);
xor_4  g09800(new_n10176, new_n10167, new_n10177);
xor_4  g09801(new_n10177, new_n10164, new_n10178);
not_8  g09802(new_n9852, new_n10179);
and_8  g09803(new_n9857, new_n10179, new_n10180);
nor_6  g09804(new_n9867, new_n9858, new_n10181);
or_8   g09805(new_n10181, new_n10180, new_n10182);
or_8   g09806(new_n9864, new_n9863, new_n10183);
or_8   g09807(new_n9865, new_n9862, new_n10184);
and_8  g09808(new_n10184, new_n10183, new_n10185);
nand_5 g09809(n4828, n2802, new_n10186);
and_8  g09810(n10928, n8236, new_n10187);
and_8  g09811(n5105, n1094, new_n10188);
xor_4  g09812(new_n10188, new_n10187, new_n10189);
xor_4  g09813(new_n10189, new_n10186, new_n10190);
xor_4  g09814(new_n10190, new_n10185, new_n10191);
xor_4  g09815(new_n10191, new_n10182, new_n10192);
xor_4  g09816(new_n10192, new_n10178, new_n10193);
nand_5 g09817(new_n9924, new_n9923, new_n10194);
or_8   g09818(new_n9930, new_n9925, new_n10195);
and_8  g09819(new_n10195, new_n10194, new_n10196);
and_8  g09820(n7891, n5069, new_n10197);
and_8  g09821(n6038, n2087, new_n10198);
xor_4  g09822(new_n10198, new_n10197, new_n10199);
xor_4  g09823(new_n10199, new_n10196, new_n10200);
and_8  g09824(n7160, n6806, new_n10201);
and_8  g09825(n6687, n615, new_n10202);
xor_4  g09826(new_n10202, new_n10201, new_n10203);
xor_4  g09827(new_n10203, new_n10200, new_n10204);
xor_4  g09828(new_n10204, new_n10193, new_n10205);
or_8   g09829(new_n9459, new_n9457_1, new_n10206);
and_8  g09830(new_n9462, new_n10206, new_n10207);
not_8  g09831(new_n10207, new_n10208);
not_8  g09832(new_n9872, new_n10209);
or_8   g09833(new_n9876, new_n9868, new_n10210);
and_8  g09834(new_n10210, new_n10209, new_n10211);
or_8   g09835(new_n9447, new_n9446, new_n10212);
nand_5 g09836(new_n9453, new_n9448, new_n10213);
and_8  g09837(new_n10213, new_n10212, new_n10214);
nand_5 g09838(n7500, n7320, new_n10215);
and_8  g09839(n12706, n2564, new_n10216);
and_8  g09840(n6770, n2585, new_n10217_1);
xor_4  g09841(new_n10217_1, new_n10216, new_n10218);
xor_4  g09842(new_n10218, new_n10215, new_n10219);
xor_4  g09843(new_n10219, new_n10214, new_n10220);
xor_4  g09844(new_n10220, new_n10211, new_n10221);
or_8   g09845(new_n10221, new_n10208, new_n10222);
not_8  g09846(new_n10220, new_n10223_1);
xor_4  g09847(new_n10223_1, new_n10211, new_n10224);
or_8   g09848(new_n10224, new_n10207, new_n10225);
and_8  g09849(new_n10225, new_n10222, new_n10226);
and_8  g09850(new_n10226, new_n10205, new_n10227);
not_8  g09851(new_n10204, new_n10228);
xor_4  g09852(new_n10228, new_n10193, new_n10229);
and_8  g09853(new_n10224, new_n10207, new_n10230);
and_8  g09854(new_n10221, new_n10208, new_n10231);
or_8   g09855(new_n10231, new_n10230, new_n10232);
and_8  g09856(new_n10232, new_n10229, new_n10233);
or_8   g09857(new_n10233, new_n10227, new_n10234);
or_8   g09858(new_n10234, new_n10160, new_n10235);
nor_6  g09859(new_n10159, new_n10141, new_n10236);
and_8  g09860(new_n10159, new_n10141, new_n10237);
or_8   g09861(new_n10237, new_n10236, new_n10238);
or_8   g09862(new_n10232, new_n10229, new_n10239);
or_8   g09863(new_n10226, new_n10205, new_n10240);
and_8  g09864(new_n10240, new_n10239, new_n10241);
or_8   g09865(new_n10241, new_n10238, new_n10242);
and_8  g09866(new_n10242, new_n10235, new_n10243);
and_8  g09867(new_n10243, new_n10120, new_n10244);
and_8  g09868(new_n10241, new_n10238, new_n10245);
and_8  g09869(new_n10234, new_n10160, new_n10246);
or_8   g09870(new_n10246, new_n10245, new_n10247);
and_8  g09871(new_n10247, new_n10119, new_n10248);
or_8   g09872(new_n10248, new_n10244, new_n10249);
and_8  g09873(new_n10249, new_n10118, new_n10250);
or_8   g09874(new_n10247, new_n10119, new_n10251);
or_8   g09875(new_n10243, new_n10120, new_n10252);
and_8  g09876(new_n10252, new_n10251, new_n10253);
and_8  g09877(new_n10253, new_n10117, new_n10254);
or_8   g09878(new_n10254, new_n10250, new_n10255);
or_8   g09879(new_n10255, new_n10053, new_n10256);
and_8  g09880(new_n10051, new_n10050, new_n10257);
and_8  g09881(new_n10048, new_n10047, new_n10258);
or_8   g09882(new_n10258, new_n10257, new_n10259);
or_8   g09883(new_n10253, new_n10117, new_n10260);
or_8   g09884(new_n10249, new_n10118, new_n10261);
and_8  g09885(new_n10261, new_n10260, new_n10262);
or_8   g09886(new_n10262, new_n10259, new_n10263);
and_8  g09887(new_n10263, new_n10256, new_n10264);
xor_4  g09888(new_n10264, new_n10045, n3654);
xnor_4 g09889(new_n10034, new_n10032, n3661);
and_8  g09890(n7456, n5305, new_n10267);
and_8  g09891(n5964, n3932, new_n10268);
and_8  g09892(n1798, n1097, new_n10269);
and_8  g09893(n12591, n5305, new_n10270);
or_8   g09894(new_n10270, new_n10269, new_n10271);
and_8  g09895(new_n10271, new_n10268, new_n10272);
and_8  g09896(new_n10270, new_n10269, new_n10273);
or_8   g09897(new_n10273, new_n10272, new_n10274);
xor_4  g09898(new_n10274, new_n10267, new_n10275);
and_8  g09899(n3932, n1097, new_n10276);
and_8  g09900(n4312, n1798, new_n10277);
and_8  g09901(n12591, n5964, new_n10278_1);
xnor_4 g09902(new_n10278_1, new_n10277, new_n10279);
xnor_4 g09903(new_n10279, new_n10276, new_n10280);
xnor_4 g09904(new_n10280, new_n10275, new_n10281);
and_8  g09905(new_n6414, new_n6413, new_n10282);
xnor_4 g09906(new_n10270, new_n10269, new_n10283);
nand_5 g09907(new_n10283, new_n10282, new_n10284);
nor_6  g09908(new_n10284, new_n10281, new_n10285);
and_8  g09909(n11662, n5305, new_n10286);
and_8  g09910(n7456, n5964, new_n10287);
nand_5 g09911(n4312, n3932, new_n10288);
and_8  g09912(n12591, n1097, new_n10289);
and_8  g09913(n12705, n1798, new_n10290);
nor_6  g09914(new_n10290, new_n10289, new_n10291);
and_8  g09915(new_n10290, new_n10289, new_n10292);
or_8   g09916(new_n10292, new_n10291, new_n10293);
xor_4  g09917(new_n10293, new_n10288, new_n10294);
xor_4  g09918(new_n10294, new_n10287, new_n10295);
or_8   g09919(new_n10278_1, new_n10277, new_n10296);
or_8   g09920(new_n10279, new_n10276, new_n10297);
and_8  g09921(new_n10297, new_n10296, new_n10298);
xor_4  g09922(new_n10298, new_n10295, new_n10299);
xor_4  g09923(new_n10299, new_n10286, new_n10300);
and_8  g09924(new_n10274, new_n10267, new_n10301);
and_8  g09925(new_n10280, new_n10275, new_n10302);
or_8   g09926(new_n10302, new_n10301, new_n10303);
xor_4  g09927(new_n10303, new_n10300, new_n10304);
xor_4  g09928(new_n10304, new_n10285, new_n10305);
not_8  g09929(new_n10305, new_n10306);
xor_4  g09930(new_n10284, new_n10281, new_n10307);
not_8  g09931(new_n10307, new_n10308);
and_8  g09932(n11023, n8759, new_n10309);
and_8  g09933(n8759, n3022, new_n10310);
and_8  g09934(n12299, n6703, new_n10311);
or_8   g09935(new_n10311, new_n10310, new_n10312);
and_8  g09936(n12299, n3022, new_n10313);
nand_5 g09937(new_n10313, new_n6407, new_n10314);
not_8  g09938(new_n10314, new_n10315);
and_8  g09939(n9640, n6776, new_n10316);
or_8   g09940(new_n10316, new_n10315, new_n10317);
and_8  g09941(new_n10317, new_n10312, new_n10318);
xor_4  g09942(new_n10318, new_n10309, new_n10319);
and_8  g09943(n12299, n9640, new_n10320);
and_8  g09944(n6776, n3022, new_n10321);
and_8  g09945(n7436, n6703, new_n10322);
xor_4  g09946(new_n10322, new_n10321, new_n10323);
xor_4  g09947(new_n10323, new_n10320, new_n10324);
xor_4  g09948(new_n10324, new_n10319, new_n10325);
not_8  g09949(new_n6407, new_n10326);
nand_5 g09950(new_n10316, new_n10326, new_n10327_1);
nand_5 g09951(new_n10314, new_n10312, new_n10328);
nand_5 g09952(new_n10328, new_n10327_1, new_n10329);
not_8  g09953(new_n10329, new_n10330);
and_8  g09954(new_n10330, new_n10316, new_n10331);
xnor_4 g09955(new_n10331, new_n10325, new_n10332);
and_8  g09956(n11922, n5331, new_n10333);
and_8  g09957(n2530, n1067, new_n10334);
and_8  g09958(n8665, n8476, new_n10335);
and_8  g09959(n12648, n5645, new_n10336);
xor_4  g09960(new_n10336, new_n10335, new_n10337);
xor_4  g09961(new_n10337, new_n10334, new_n10338);
xor_4  g09962(new_n10338, new_n10333, new_n10339);
not_8  g09963(new_n10339, new_n10340);
and_8  g09964(n8665, n5331, new_n10341);
and_8  g09965(n5645, n2530, new_n10342);
or_8   g09966(new_n10342, new_n10341, new_n10343);
and_8  g09967(n8476, n1067, new_n10344);
and_8  g09968(n8665, n2530, new_n10345);
and_8  g09969(new_n10345, new_n6408, new_n10346);
or_8   g09970(new_n10346, new_n10344, new_n10347);
nand_5 g09971(new_n10347, new_n10343, new_n10348);
xor_4  g09972(new_n10348, new_n10340, new_n10349);
and_8  g09973(new_n6428, new_n6427, new_n10350);
not_8  g09974(new_n10346, new_n10351);
nand_5 g09975(new_n10351, new_n10343, new_n10352);
and_8  g09976(new_n10352, new_n10350, new_n10353);
xor_4  g09977(new_n10353, new_n10349, new_n10354);
and_8  g09978(n7965, n2749, new_n10355);
and_8  g09979(n7965, n3754, new_n10356);
and_8  g09980(n11892, n11876, new_n10357);
or_8   g09981(new_n10357, new_n10356, new_n10358);
and_8  g09982(n11892, n3754, new_n10359);
and_8  g09983(new_n10359, new_n6409, new_n10360);
and_8  g09984(n10898, n7388, new_n10361);
or_8   g09985(new_n10361, new_n10360, new_n10362);
and_8  g09986(new_n10362, new_n10358, new_n10363);
xor_4  g09987(new_n10363, new_n10355, new_n10364);
and_8  g09988(n11892, n10898, new_n10365);
and_8  g09989(n7388, n3754, new_n10366);
and_8  g09990(n11876, n2393, new_n10367);
nor_6  g09991(new_n10367, new_n10366, new_n10368);
and_8  g09992(new_n10367, new_n10366, new_n10369);
or_8   g09993(new_n10369, new_n10368, new_n10370);
xnor_4 g09994(new_n10370, new_n10365, new_n10371);
and_8  g09995(new_n10371, new_n10364, new_n10372);
nor_6  g09996(new_n10371, new_n10364, new_n10373);
or_8   g09997(new_n10373, new_n10372, new_n10374);
not_8  g09998(new_n10361, new_n10375);
or_8   g09999(new_n10375, new_n6409, new_n10376);
not_8  g10000(new_n10358, new_n10377);
or_8   g10001(new_n10360, new_n10377, new_n10378);
and_8  g10002(new_n10378, new_n10376, new_n10379);
not_8  g10003(new_n10379, new_n10380);
or_8   g10004(new_n10380, new_n10375, new_n10381);
xor_4  g10005(new_n10381, new_n10374, new_n10382);
xor_4  g10006(new_n10382, new_n10354, new_n10383);
or_8   g10007(new_n10376, new_n10377, new_n10384);
and_8  g10008(new_n10384, new_n10380, new_n10385);
and_8  g10009(new_n6425, new_n6422, new_n10386);
and_8  g10010(new_n6429_1, new_n6426, new_n10387);
or_8   g10011(new_n10387, new_n10386, new_n10388);
nor_6  g10012(new_n10388, new_n10385, new_n10389);
xor_4  g10013(new_n10388, new_n10385, new_n10390);
not_8  g10014(new_n6408, new_n10391_1);
nand_5 g10015(new_n10344, new_n10391_1, new_n10392);
or_8   g10016(new_n10392, new_n10343, new_n10393);
not_8  g10017(new_n10392, new_n10394);
or_8   g10018(new_n10394, new_n10352, new_n10395);
and_8  g10019(new_n10395, new_n10393, new_n10396);
and_8  g10020(new_n10396, new_n10390, new_n10397);
or_8   g10021(new_n10397, new_n10389, new_n10398);
or_8   g10022(new_n10398, new_n10383, new_n10399);
not_8  g10023(new_n10348, new_n10400);
xor_4  g10024(new_n10400, new_n10340, new_n10401);
xor_4  g10025(new_n10353, new_n10401, new_n10402);
xor_4  g10026(new_n10382, new_n10402, new_n10403);
nor_6  g10027(new_n10397, new_n10389, new_n10404);
or_8   g10028(new_n10404, new_n10403, new_n10405);
and_8  g10029(new_n10405, new_n10399, new_n10406);
nor_6  g10030(new_n10406, new_n10332, new_n10407);
and_8  g10031(new_n10406, new_n10332, new_n10408);
or_8   g10032(new_n10408, new_n10407, new_n10409);
not_8  g10033(new_n10327_1, new_n10410);
nand_5 g10034(new_n10410, new_n10312, new_n10411);
and_8  g10035(new_n10411, new_n10329, new_n10412);
and_8  g10036(new_n6420, new_n6417, new_n10413);
and_8  g10037(new_n6430, new_n6421, new_n10414);
or_8   g10038(new_n10414, new_n10413, new_n10415);
nor_6  g10039(new_n10415, new_n10412, new_n10416);
xor_4  g10040(new_n10396, new_n10390, new_n10417);
xor_4  g10041(new_n10415, new_n10412, new_n10418);
and_8  g10042(new_n10418, new_n10417, new_n10419);
nor_6  g10043(new_n10419, new_n10416, new_n10420);
xor_4  g10044(new_n10420, new_n10409, new_n10421);
or_8   g10045(new_n10421, new_n10308, new_n10422);
nor_6  g10046(new_n10408, new_n10407, new_n10423);
xor_4  g10047(new_n10420, new_n10423, new_n10424);
and_8  g10048(new_n10424, new_n10307, new_n10425);
and_8  g10049(new_n10421, new_n10308, new_n10426);
or_8   g10050(new_n10426, new_n10425, new_n10427);
xor_4  g10051(new_n10418, new_n10417, new_n10428);
not_8  g10052(new_n6406, new_n10429);
and_8  g10053(new_n10268, new_n10429, new_n10430);
not_8  g10054(new_n10430, new_n10431);
or_8   g10055(new_n10431, new_n10271, new_n10432);
or_8   g10056(new_n10430, new_n10283, new_n10433);
and_8  g10057(new_n10433, new_n10432, new_n10434);
and_8  g10058(new_n10434, new_n10428, new_n10435);
nand_5 g10059(new_n6415, new_n6412, new_n10436);
nand_5 g10060(new_n6431_1, new_n6416, new_n10437);
and_8  g10061(new_n10437, new_n10436, new_n10438);
xor_4  g10062(new_n10434, new_n10428, new_n10439_1);
and_8  g10063(new_n10439_1, new_n10438, new_n10440);
or_8   g10064(new_n10440, new_n10435, new_n10441);
or_8   g10065(new_n10441, new_n10427, new_n10442);
and_8  g10066(new_n10442, new_n10422, new_n10443);
and_8  g10067(new_n10443, new_n10306, new_n10444);
or_8   g10068(new_n10424, new_n10307, new_n10445);
and_8  g10069(new_n10445, new_n10422, new_n10446);
not_8  g10070(new_n10435, new_n10447);
not_8  g10071(new_n10438, new_n10448);
nor_6  g10072(new_n10418, new_n10417, new_n10449);
or_8   g10073(new_n10449, new_n10419, new_n10450);
xor_4  g10074(new_n10434, new_n10450, new_n10451_1);
or_8   g10075(new_n10451_1, new_n10448, new_n10452);
and_8  g10076(new_n10452, new_n10447, new_n10453);
and_8  g10077(new_n10453, new_n10446, new_n10454);
or_8   g10078(new_n10454, new_n10425, new_n10455);
and_8  g10079(new_n10455, new_n10305, new_n10456);
or_8   g10080(new_n10456, new_n10444, new_n10457);
and_8  g10081(new_n10331, new_n10325, new_n10458);
nand_5 g10082(n10451, n8759, new_n10459);
and_8  g10083(n11023, n6776, new_n10460);
or_8   g10084(new_n10322, new_n10321, new_n10461);
and_8  g10085(new_n10322, new_n10321, new_n10462);
or_8   g10086(new_n10462, new_n10320, new_n10463);
and_8  g10087(new_n10463, new_n10461, new_n10464);
xor_4  g10088(new_n10464, new_n10460, new_n10465);
and_8  g10089(n9640, n7436, new_n10466);
and_8  g10090(n8276, n6703, new_n10467);
xor_4  g10091(new_n10467, new_n10313, new_n10468);
xor_4  g10092(new_n10468, new_n10466, new_n10469);
xnor_4 g10093(new_n10469, new_n10465, new_n10470);
xor_4  g10094(new_n10470, new_n10459, new_n10471);
and_8  g10095(new_n10318, new_n10309, new_n10472);
and_8  g10096(new_n10324, new_n10319, new_n10473);
or_8   g10097(new_n10473, new_n10472, new_n10474);
xor_4  g10098(new_n10474, new_n10471, new_n10475);
xor_4  g10099(new_n10475, new_n10458, new_n10476_1);
nor_6  g10100(new_n10381, new_n10374, new_n10477);
and_8  g10101(n7965, n159, new_n10478);
and_8  g10102(new_n10363, new_n10355, new_n10479);
or_8   g10103(new_n10372, new_n10479, new_n10480);
and_8  g10104(new_n10480, new_n10478, new_n10481);
nor_6  g10105(new_n10480, new_n10478, new_n10482);
or_8   g10106(new_n10482, new_n10481, new_n10483);
and_8  g10107(n7388, n2749, new_n10484);
or_8   g10108(new_n10367, new_n10366, new_n10485);
or_8   g10109(new_n10370, new_n10365, new_n10486);
and_8  g10110(new_n10486, new_n10485, new_n10487);
and_8  g10111(new_n10487, new_n10484, new_n10488);
nor_6  g10112(new_n10487, new_n10484, new_n10489);
or_8   g10113(new_n10489, new_n10488, new_n10490);
not_8  g10114(new_n10359, new_n10491);
and_8  g10115(n11876, n5860, new_n10492);
and_8  g10116(n10898, n2393, new_n10493);
xor_4  g10117(new_n10493, new_n10492, new_n10494);
xor_4  g10118(new_n10494, new_n10491, new_n10495);
xor_4  g10119(new_n10495, new_n10490, new_n10496);
not_8  g10120(new_n10496, new_n10497);
xor_4  g10121(new_n10497, new_n10483, new_n10498);
xor_4  g10122(new_n10498, new_n10477, new_n10499);
nand_5 g10123(new_n10353, new_n10349, new_n10500);
not_8  g10124(new_n10500, new_n10501);
and_8  g10125(n5331, n2551, new_n10502);
not_8  g10126(new_n10502, new_n10503);
and_8  g10127(n11922, n8476, new_n10504);
or_8   g10128(new_n10336, new_n10335, new_n10505);
and_8  g10129(new_n10336, new_n10335, new_n10506);
or_8   g10130(new_n10506, new_n10334, new_n10507);
and_8  g10131(new_n10507, new_n10505, new_n10508);
xor_4  g10132(new_n10508, new_n10504, new_n10509);
and_8  g10133(n12648, n1067, new_n10510_1);
and_8  g10134(n10545, n5645, new_n10511);
xor_4  g10135(new_n10511, new_n10345, new_n10512);
xor_4  g10136(new_n10512, new_n10510_1, new_n10513);
and_8  g10137(new_n10513, new_n10509, new_n10514);
nor_6  g10138(new_n10513, new_n10509, new_n10515);
or_8   g10139(new_n10515, new_n10514, new_n10516);
xor_4  g10140(new_n10516, new_n10503, new_n10517);
and_8  g10141(new_n10338, new_n10333, new_n10518);
and_8  g10142(new_n10400, new_n10339, new_n10519);
or_8   g10143(new_n10519, new_n10518, new_n10520);
xor_4  g10144(new_n10520, new_n10517, new_n10521);
xor_4  g10145(new_n10521, new_n10501, new_n10522);
xor_4  g10146(new_n10522, new_n10499, new_n10523);
and_8  g10147(new_n10381, new_n10374, new_n10524);
or_8   g10148(new_n10524, new_n10477, new_n10525);
and_8  g10149(new_n10525, new_n10402, new_n10526);
and_8  g10150(new_n10398, new_n10383, new_n10527);
or_8   g10151(new_n10527, new_n10526, new_n10528);
and_8  g10152(new_n10528, new_n10523, new_n10529);
and_8  g10153(new_n10522, new_n10499, new_n10530);
nor_6  g10154(new_n10522, new_n10499, new_n10531);
or_8   g10155(new_n10531, new_n10530, new_n10532);
not_8  g10156(new_n10528, new_n10533);
and_8  g10157(new_n10533, new_n10532, new_n10534);
or_8   g10158(new_n10534, new_n10529, new_n10535);
and_8  g10159(new_n10535, new_n10476_1, new_n10536);
not_8  g10160(new_n10476_1, new_n10537);
or_8   g10161(new_n10533, new_n10532, new_n10538);
or_8   g10162(new_n10528, new_n10523, new_n10539);
and_8  g10163(new_n10539, new_n10538, new_n10540);
and_8  g10164(new_n10540, new_n10537, new_n10541);
or_8   g10165(new_n10541, new_n10536, new_n10542);
nor_6  g10166(new_n10420, new_n10409, new_n10543);
or_8   g10167(new_n10543, new_n10408, new_n10544);
not_8  g10168(new_n10544, new_n10545_1);
xor_4  g10169(new_n10545_1, new_n10542, new_n10546);
xor_4  g10170(new_n10546, new_n10457, n3677);
xor_4  g10171(new_n9116, new_n9110, n3849);
xor_4  g10172(new_n6402, new_n6401, n4088);
xor_4  g10173(new_n1151, new_n1059, n4155);
xor_4  g10174(new_n3049, new_n3045, n4159);
xor_4  g10175(new_n6392, new_n6233, n4226);
nand_5 g10176(n12591, n4312, new_n10553);
or_8   g10177(new_n10290, new_n10289, new_n10554);
and_8  g10178(n4312, n3932, new_n10555);
or_8   g10179(new_n10293, new_n10555, new_n10556);
and_8  g10180(new_n10556, new_n10554, new_n10557);
xor_4  g10181(new_n10557, new_n10553, new_n10558);
and_8  g10182(n12705, n3932, new_n10559);
and_8  g10183(n12025, n1798, new_n10560);
xor_4  g10184(new_n10560, new_n10559, new_n10561);
xor_4  g10185(new_n10561, new_n10558, new_n10562);
and_8  g10186(n11662, n5964, new_n10563);
and_8  g10187(n7456, n1097, new_n10564);
xnor_4 g10188(new_n10564, new_n10563, new_n10565);
and_8  g10189(new_n10565, new_n10562, new_n10566);
nor_6  g10190(new_n10565, new_n10562, new_n10567);
or_8   g10191(new_n10567, new_n10566, new_n10568);
and_8  g10192(new_n10294, new_n10287, new_n10569);
and_8  g10193(new_n10298, new_n10295, new_n10570);
nor_6  g10194(new_n10570, new_n10569, new_n10571);
xor_4  g10195(new_n10571, new_n10568, new_n10572);
and_8  g10196(new_n10299, new_n10286, new_n10573);
and_8  g10197(new_n10303, new_n10300, new_n10574);
or_8   g10198(new_n10574, new_n10573, new_n10575);
and_8  g10199(new_n10575, new_n10572, new_n10576);
not_8  g10200(new_n10553, new_n10577);
or_8   g10201(new_n10557, new_n10577, new_n10578);
or_8   g10202(new_n10561, new_n10558, new_n10579);
and_8  g10203(new_n10579, new_n10578, new_n10580);
and_8  g10204(n10327, n5964, new_n10581);
and_8  g10205(n11662, n1097, new_n10582);
and_8  g10206(n9583, n5305, new_n10583);
xnor_4 g10207(new_n10583, new_n10582, new_n10584);
xnor_4 g10208(new_n10584, new_n10581, new_n10585);
xor_4  g10209(new_n10585, new_n10580, new_n10586);
and_8  g10210(new_n10560, new_n10559, new_n10587);
and_8  g10211(n7456, n4312, new_n10588);
xor_4  g10212(new_n10588, new_n10587, new_n10589_1);
and_8  g10213(n12025, n3932, new_n10590);
and_8  g10214(n12705, n12591, new_n10591);
and_8  g10215(n11257, n1798, new_n10592);
xnor_4 g10216(new_n10592, new_n10591, new_n10593);
xor_4  g10217(new_n10593, new_n10590, new_n10594);
xor_4  g10218(new_n10594, new_n10589_1, new_n10595);
xor_4  g10219(new_n10595, new_n10586, new_n10596);
not_8  g10220(new_n10567, new_n10597);
nand_5 g10221(new_n10564, new_n10563, new_n10598);
not_8  g10222(new_n10598, new_n10599);
nor_6  g10223(new_n10571, new_n10568, new_n10600);
and_8  g10224(new_n10600, new_n10599, new_n10601);
or_8   g10225(new_n10571, new_n10568, new_n10602);
and_8  g10226(new_n10602, new_n10598, new_n10603);
or_8   g10227(new_n10603, new_n10601, new_n10604);
and_8  g10228(new_n10604, new_n10597, new_n10605);
xor_4  g10229(new_n10605, new_n10596, new_n10606);
xor_4  g10230(new_n10606, new_n10576, new_n10607);
nand_5 g10231(n10327, n5305, new_n10608);
not_8  g10232(new_n10608, new_n10609);
xor_4  g10233(new_n10575, new_n10572, new_n10610);
or_8   g10234(new_n10610, new_n10609, new_n10611);
and_8  g10235(new_n10304, new_n10285, new_n10612);
xor_4  g10236(new_n10610, new_n10608, new_n10613);
or_8   g10237(new_n10613, new_n10612, new_n10614);
and_8  g10238(new_n10614, new_n10611, new_n10615);
xor_4  g10239(new_n10615, new_n10607, new_n10616);
not_8  g10240(new_n10616, new_n10617);
and_8  g10241(new_n10464, new_n10460, new_n10618);
and_8  g10242(new_n10469, new_n10465, new_n10619);
or_8   g10243(new_n10619, new_n10618, new_n10620);
and_8  g10244(n10451, n6776, new_n10621);
and_8  g10245(n12299, n11023, new_n10622);
xnor_4 g10246(new_n10622, new_n10621, new_n10623);
xor_4  g10247(new_n10623, new_n10620, new_n10624);
and_8  g10248(n7436, n3022, new_n10625);
and_8  g10249(n9640, n8276, new_n10626);
and_8  g10250(n9241, n6703, new_n10627);
xor_4  g10251(new_n10627, new_n10626, new_n10628);
xor_4  g10252(new_n10628, new_n10625, new_n10629);
or_8   g10253(new_n10467, new_n10313, new_n10630);
and_8  g10254(new_n10467, new_n10313, new_n10631);
or_8   g10255(new_n10631, new_n10466, new_n10632);
nand_5 g10256(new_n10632, new_n10630, new_n10633);
xor_4  g10257(new_n10633, new_n10629, new_n10634);
xor_4  g10258(new_n10634, new_n10624, new_n10635);
nor_6  g10259(new_n10470, new_n10459, new_n10636);
and_8  g10260(new_n10474, new_n10471, new_n10637);
or_8   g10261(new_n10637, new_n10636, new_n10638);
and_8  g10262(new_n10638, new_n10635, new_n10639);
nor_6  g10263(new_n10628, new_n10625, new_n10640);
and_8  g10264(new_n10633, new_n10629, new_n10641);
or_8   g10265(new_n10641, new_n10640, new_n10642);
and_8  g10266(n10278, n6776, new_n10643);
and_8  g10267(n12299, n10451, new_n10644_1);
and_8  g10268(n11423, n8759, new_n10645);
xnor_4 g10269(new_n10645, new_n10644_1, new_n10646);
xor_4  g10270(new_n10646, new_n10643, new_n10647);
xnor_4 g10271(new_n10647, new_n10642, new_n10648);
and_8  g10272(new_n10627, new_n10626, new_n10649);
and_8  g10273(n11023, n7436, new_n10650);
xnor_4 g10274(new_n10650, new_n10649, new_n10651);
and_8  g10275(n9640, n9241, new_n10652);
and_8  g10276(n8276, n3022, new_n10653);
and_8  g10277(n10510, n6703, new_n10654);
xnor_4 g10278(new_n10654, new_n10653, new_n10655);
xor_4  g10279(new_n10655, new_n10652, new_n10656);
xor_4  g10280(new_n10656, new_n10651, new_n10657);
xor_4  g10281(new_n10657, new_n10648, new_n10658);
not_8  g10282(new_n10620, new_n10659);
or_8   g10283(new_n10623, new_n10659, new_n10660);
and_8  g10284(new_n10622, new_n10621, new_n10661);
or_8   g10285(new_n10634, new_n10624, new_n10662);
xor_4  g10286(new_n10662, new_n10661, new_n10663);
and_8  g10287(new_n10663, new_n10660, new_n10664);
xor_4  g10288(new_n10664, new_n10658, new_n10665);
xor_4  g10289(new_n10665, new_n10639, new_n10666);
nand_5 g10290(n10278, n8759, new_n10667);
not_8  g10291(new_n10667, new_n10668);
xor_4  g10292(new_n10638, new_n10635, new_n10669);
and_8  g10293(new_n10669, new_n10668, new_n10670);
and_8  g10294(new_n10475, new_n10458, new_n10671);
xor_4  g10295(new_n10669, new_n10668, new_n10672);
and_8  g10296(new_n10672, new_n10671, new_n10673);
or_8   g10297(new_n10673, new_n10670, new_n10674);
and_8  g10298(new_n10674, new_n10666, new_n10675);
nor_6  g10299(new_n10674, new_n10666, new_n10676);
or_8   g10300(new_n10676, new_n10675, new_n10677);
and_8  g10301(n12648, n8665, new_n10678_1);
and_8  g10302(n10545, n1067, new_n10679);
and_8  g10303(n7690, n5645, new_n10680);
xor_4  g10304(new_n10680, new_n10679, new_n10681);
and_8  g10305(new_n10681, new_n10678_1, new_n10682);
nor_6  g10306(new_n10681, new_n10678_1, new_n10683);
or_8   g10307(new_n10683, new_n10682, new_n10684);
or_8   g10308(new_n10511, new_n10345, new_n10685_1);
and_8  g10309(new_n10511, new_n10345, new_n10686);
or_8   g10310(new_n10686, new_n10510_1, new_n10687);
and_8  g10311(new_n10687, new_n10685_1, new_n10688);
xor_4  g10312(new_n10688, new_n10684, new_n10689);
and_8  g10313(n8476, n2551, new_n10690);
and_8  g10314(n11922, n2530, new_n10691);
xor_4  g10315(new_n10691, new_n10690, new_n10692);
not_8  g10316(new_n10692, new_n10693);
or_8   g10317(new_n10693, new_n10689, new_n10694);
nand_5 g10318(new_n10687, new_n10685_1, new_n10695_1);
or_8   g10319(new_n10695_1, new_n10684, new_n10696);
xor_4  g10320(new_n10681, new_n10678_1, new_n10697);
or_8   g10321(new_n10688, new_n10697, new_n10698);
and_8  g10322(new_n10698, new_n10696, new_n10699);
or_8   g10323(new_n10692, new_n10699, new_n10700);
and_8  g10324(new_n10700, new_n10694, new_n10701);
and_8  g10325(new_n10508, new_n10504, new_n10702);
or_8   g10326(new_n10514, new_n10702, new_n10703);
xor_4  g10327(new_n10703, new_n10701, new_n10704);
nor_6  g10328(new_n10516, new_n10503, new_n10705);
and_8  g10329(new_n10520, new_n10517, new_n10706);
or_8   g10330(new_n10706, new_n10705, new_n10707);
and_8  g10331(new_n10707, new_n10704, new_n10708);
not_8  g10332(new_n10708, new_n10709);
and_8  g10333(new_n10680, new_n10679, new_n10710);
and_8  g10334(n12648, n11922, new_n10711);
xor_4  g10335(new_n10711, new_n10710, new_n10712);
not_8  g10336(new_n10712, new_n10713);
nand_5 g10337(n7690, n1067, new_n10714);
not_8  g10338(new_n10714, new_n10715);
and_8  g10339(n10545, n8665, new_n10716);
and_8  g10340(n5645, n3616, new_n10717);
xnor_4 g10341(new_n10717, new_n10716, new_n10718);
xor_4  g10342(new_n10718, new_n10715, new_n10719);
or_8   g10343(new_n10719, new_n10713, new_n10720);
xor_4  g10344(new_n10718, new_n10714, new_n10721);
or_8   g10345(new_n10721, new_n10712, new_n10722);
and_8  g10346(new_n10722, new_n10720, new_n10723);
and_8  g10347(new_n10688, new_n10697, new_n10724);
or_8   g10348(new_n10724, new_n10682, new_n10725);
and_8  g10349(n12826, n8476, new_n10726);
and_8  g10350(n2551, n2530, new_n10727);
and_8  g10351(n5331, n4094, new_n10728);
xnor_4 g10352(new_n10728, new_n10727, new_n10729);
nor_6  g10353(new_n10729, new_n10726, new_n10730);
and_8  g10354(new_n10729, new_n10726, new_n10731);
or_8   g10355(new_n10731, new_n10730, new_n10732);
nor_6  g10356(new_n10732, new_n10725, new_n10733);
and_8  g10357(new_n10732, new_n10725, new_n10734);
or_8   g10358(new_n10734, new_n10733, new_n10735);
xor_4  g10359(new_n10735, new_n10723, new_n10736);
and_8  g10360(new_n10691, new_n10690, new_n10737);
and_8  g10361(new_n10703, new_n10701, new_n10738);
and_8  g10362(new_n10738, new_n10737, new_n10739);
nor_6  g10363(new_n10738, new_n10737, new_n10740);
or_8   g10364(new_n10740, new_n10739, new_n10741);
and_8  g10365(new_n10741, new_n10694, new_n10742);
nor_6  g10366(new_n10742, new_n10736, new_n10743);
and_8  g10367(new_n10742, new_n10736, new_n10744);
or_8   g10368(new_n10744, new_n10743, new_n10745);
xor_4  g10369(new_n10745, new_n10709, new_n10746);
nand_5 g10370(n12826, n5331, new_n10747);
not_8  g10371(new_n10747, new_n10748);
xor_4  g10372(new_n10707, new_n10704, new_n10749);
or_8   g10373(new_n10749, new_n10748, new_n10750);
and_8  g10374(new_n10521, new_n10501, new_n10751);
xor_4  g10375(new_n10749, new_n10747, new_n10752);
or_8   g10376(new_n10752, new_n10751, new_n10753);
and_8  g10377(new_n10753, new_n10750, new_n10754);
and_8  g10378(new_n10754, new_n10746, new_n10755);
xor_4  g10379(new_n10745, new_n10708, new_n10756);
not_8  g10380(new_n10750, new_n10757);
not_8  g10381(new_n10521, new_n10758);
or_8   g10382(new_n10758, new_n10500, new_n10759);
xor_4  g10383(new_n10749, new_n10748, new_n10760);
and_8  g10384(new_n10760, new_n10759, new_n10761);
or_8   g10385(new_n10761, new_n10757, new_n10762);
and_8  g10386(new_n10762, new_n10756, new_n10763);
or_8   g10387(new_n10763, new_n10755, new_n10764);
and_8  g10388(n7965, n1510, new_n10765);
nor_6  g10389(new_n10495, new_n10490, new_n10766);
or_8   g10390(new_n10766, new_n10488, new_n10767);
and_8  g10391(n7388, n159, new_n10768);
and_8  g10392(n11892, n2749, new_n10769);
xor_4  g10393(new_n10769, new_n10768, new_n10770);
xor_4  g10394(new_n10770, new_n10767, new_n10771);
and_8  g10395(n3754, n2393, new_n10772);
and_8  g10396(n10898, n5860, new_n10773);
and_8  g10397(n11876, n3986, new_n10774);
xor_4  g10398(new_n10774, new_n10773, new_n10775);
xor_4  g10399(new_n10775, new_n10772, new_n10776);
not_8  g10400(new_n10776, new_n10777);
nor_6  g10401(new_n10493, new_n10492, new_n10778);
and_8  g10402(new_n10494, new_n10491, new_n10779);
or_8   g10403(new_n10779, new_n10778, new_n10780);
xor_4  g10404(new_n10780, new_n10777, new_n10781);
not_8  g10405(new_n10781, new_n10782);
and_8  g10406(new_n10782, new_n10771, new_n10783);
nor_6  g10407(new_n10770, new_n10767, new_n10784);
and_8  g10408(new_n10770, new_n10767, new_n10785);
or_8   g10409(new_n10785, new_n10784, new_n10786);
and_8  g10410(new_n10781, new_n10786, new_n10787);
or_8   g10411(new_n10787, new_n10783, new_n10788);
xor_4  g10412(new_n10480, new_n10478, new_n10789_1);
and_8  g10413(new_n10496, new_n10789_1, new_n10790);
or_8   g10414(new_n10790, new_n10481, new_n10791);
and_8  g10415(new_n10791, new_n10788, new_n10792);
or_8   g10416(new_n10781, new_n10786, new_n10793);
or_8   g10417(new_n10782, new_n10771, new_n10794);
and_8  g10418(new_n10794, new_n10793, new_n10795);
not_8  g10419(new_n10481, new_n10796);
or_8   g10420(new_n10497, new_n10483, new_n10797);
and_8  g10421(new_n10797, new_n10796, new_n10798);
and_8  g10422(new_n10798, new_n10795, new_n10799);
nor_6  g10423(new_n10799, new_n10792, new_n10800);
and_8  g10424(new_n10800, new_n10765, new_n10801);
and_8  g10425(new_n10498, new_n10477, new_n10802);
not_8  g10426(new_n10765, new_n10803);
or_8   g10427(new_n10799, new_n10792, new_n10804);
or_8   g10428(new_n10804, new_n10803, new_n10805);
or_8   g10429(new_n10800, new_n10765, new_n10806);
and_8  g10430(new_n10806, new_n10805, new_n10807);
and_8  g10431(new_n10807, new_n10802, new_n10808);
nor_6  g10432(new_n10808, new_n10801, new_n10809);
not_8  g10433(new_n10792, new_n10810);
and_8  g10434(new_n10769, new_n10768, new_n10811);
or_8   g10435(new_n10783, new_n10784, new_n10812);
xor_4  g10436(new_n10812, new_n10811, new_n10813);
and_8  g10437(n7388, n1510, new_n10814);
and_8  g10438(n11892, n159, new_n10815);
and_8  g10439(n12247, n7965, new_n10816);
xnor_4 g10440(new_n10816, new_n10815, new_n10817);
xor_4  g10441(new_n10817, new_n10814, new_n10818);
nand_5 g10442(new_n10775, new_n10772, new_n10819);
or_8   g10443(new_n10780, new_n10777, new_n10820);
and_8  g10444(new_n10820, new_n10819, new_n10821);
xor_4  g10445(new_n10821, new_n10818, new_n10822);
and_8  g10446(new_n10774, new_n10773, new_n10823);
and_8  g10447(n2749, n2393, new_n10824);
xnor_4 g10448(new_n10824, new_n10823, new_n10825);
and_8  g10449(n10898, n3986, new_n10826);
and_8  g10450(n11876, n5857, new_n10827);
and_8  g10451(n5860, n3754, new_n10828);
xnor_4 g10452(new_n10828, new_n10827, new_n10829);
xor_4  g10453(new_n10829, new_n10826, new_n10830);
nor_6  g10454(new_n10830, new_n10825, new_n10831);
and_8  g10455(new_n10830, new_n10825, new_n10832);
or_8   g10456(new_n10832, new_n10831, new_n10833);
xor_4  g10457(new_n10833, new_n10822, new_n10834);
or_8   g10458(new_n10834, new_n10813, new_n10835);
not_8  g10459(new_n10811, new_n10836);
xor_4  g10460(new_n10812, new_n10836, new_n10837);
not_8  g10461(new_n10834, new_n10838);
or_8   g10462(new_n10838, new_n10837, new_n10839);
and_8  g10463(new_n10839, new_n10835, new_n10840);
xor_4  g10464(new_n10840, new_n10810, new_n10841);
or_8   g10465(new_n10841, new_n10809, new_n10842);
or_8   g10466(new_n10808, new_n10801, new_n10843);
xor_4  g10467(new_n10840, new_n10792, new_n10844);
or_8   g10468(new_n10844, new_n10843, new_n10845);
and_8  g10469(new_n10845, new_n10842, new_n10846);
xor_4  g10470(new_n10846, new_n10764, new_n10847);
xor_4  g10471(new_n10807, new_n10802, new_n10848_1);
and_8  g10472(new_n10752, new_n10751, new_n10849);
or_8   g10473(new_n10849, new_n10761, new_n10850);
or_8   g10474(new_n10850, new_n10848_1, new_n10851_1);
or_8   g10475(new_n10522, new_n10499, new_n10852);
and_8  g10476(new_n10538, new_n10852, new_n10853);
not_8  g10477(new_n10802, new_n10854);
xor_4  g10478(new_n10807, new_n10854, new_n10855);
or_8   g10479(new_n10760, new_n10759, new_n10856);
and_8  g10480(new_n10856, new_n10753, new_n10857);
and_8  g10481(new_n10857, new_n10855, new_n10858);
and_8  g10482(new_n10850, new_n10848_1, new_n10859);
or_8   g10483(new_n10859, new_n10858, new_n10860);
or_8   g10484(new_n10860, new_n10853, new_n10861);
and_8  g10485(new_n10861, new_n10851_1, new_n10862);
or_8   g10486(new_n10862, new_n10847, new_n10863);
or_8   g10487(new_n10762, new_n10756, new_n10864);
or_8   g10488(new_n10754, new_n10746, new_n10865);
and_8  g10489(new_n10865, new_n10864, new_n10866);
xor_4  g10490(new_n10846, new_n10866, new_n10867);
or_8   g10491(new_n10529, new_n10531, new_n10868);
or_8   g10492(new_n10857, new_n10855, new_n10869);
and_8  g10493(new_n10869, new_n10851_1, new_n10870);
and_8  g10494(new_n10870, new_n10868, new_n10871);
or_8   g10495(new_n10871, new_n10858, new_n10872);
or_8   g10496(new_n10872, new_n10867, new_n10873);
and_8  g10497(new_n10873, new_n10863, new_n10874);
and_8  g10498(new_n10874, new_n10677, new_n10875);
xor_4  g10499(new_n10674, new_n10666, new_n10876);
and_8  g10500(new_n10872, new_n10867, new_n10877);
and_8  g10501(new_n10862, new_n10847, new_n10878);
or_8   g10502(new_n10878, new_n10877, new_n10879);
and_8  g10503(new_n10879, new_n10876, new_n10880);
or_8   g10504(new_n10880, new_n10875, new_n10881);
nor_6  g10505(new_n10672, new_n10671, new_n10882);
or_8   g10506(new_n10882, new_n10673, new_n10883);
or_8   g10507(new_n10870, new_n10868, new_n10884);
and_8  g10508(new_n10884, new_n10861, new_n10885);
and_8  g10509(new_n10885, new_n10883, new_n10886);
or_8   g10510(new_n10540, new_n10537, new_n10887);
or_8   g10511(new_n10544, new_n10542, new_n10888);
and_8  g10512(new_n10888, new_n10887, new_n10889);
xor_4  g10513(new_n10672, new_n10671, new_n10890);
and_8  g10514(new_n10860, new_n10853, new_n10891);
or_8   g10515(new_n10891, new_n10871, new_n10892);
or_8   g10516(new_n10892, new_n10890, new_n10893);
or_8   g10517(new_n10885, new_n10883, new_n10894);
and_8  g10518(new_n10894, new_n10893, new_n10895);
and_8  g10519(new_n10895, new_n10889, new_n10896);
nor_6  g10520(new_n10896, new_n10886, new_n10897);
or_8   g10521(new_n10897, new_n10881, new_n10898_1);
or_8   g10522(new_n10879, new_n10876, new_n10899);
or_8   g10523(new_n10874, new_n10677, new_n10900);
and_8  g10524(new_n10900, new_n10899, new_n10901);
or_8   g10525(new_n10896, new_n10886, new_n10902);
or_8   g10526(new_n10902, new_n10901, new_n10903);
and_8  g10527(new_n10903, new_n10898_1, new_n10904);
and_8  g10528(new_n10904, new_n10617, new_n10905);
and_8  g10529(new_n10902, new_n10901, new_n10906);
and_8  g10530(new_n10897, new_n10881, new_n10907);
or_8   g10531(new_n10907, new_n10906, new_n10908);
or_8   g10532(new_n10908, new_n10616, new_n10909);
or_8   g10533(new_n10904, new_n10617, new_n10910);
and_8  g10534(new_n10910, new_n10909, new_n10911);
xor_4  g10535(new_n10613, new_n10612, new_n10912);
xor_4  g10536(new_n10895, new_n10889, new_n10913_1);
and_8  g10537(new_n10913_1, new_n10912, new_n10914);
not_8  g10538(new_n10912, new_n10915);
or_8   g10539(new_n10535, new_n10476_1, new_n10916);
and_8  g10540(new_n10916, new_n10887, new_n10917);
and_8  g10541(new_n10545_1, new_n10917, new_n10918);
or_8   g10542(new_n10918, new_n10536, new_n10919);
xor_4  g10543(new_n10895, new_n10919, new_n10920);
or_8   g10544(new_n10920, new_n10915, new_n10921);
or_8   g10545(new_n10913_1, new_n10912, new_n10922);
and_8  g10546(new_n10922, new_n10921, new_n10923);
or_8   g10547(new_n10443, new_n10306, new_n10924);
or_8   g10548(new_n10546, new_n10457, new_n10925);
and_8  g10549(new_n10925, new_n10924, new_n10926);
and_8  g10550(new_n10926, new_n10923, new_n10927);
or_8   g10551(new_n10927, new_n10914, new_n10928_1);
and_8  g10552(new_n10928_1, new_n10911, new_n10929);
nor_6  g10553(new_n10929, new_n10905, new_n10930);
and_8  g10554(new_n10665, new_n10639, new_n10931);
or_8   g10555(new_n10675, new_n10931, new_n10932);
or_8   g10556(new_n10906, new_n10875, new_n10933);
or_8   g10557(new_n10588, new_n10587, new_n10934);
nand_5 g10558(new_n10594, new_n10589_1, new_n10935);
and_8  g10559(new_n10935, new_n10934, new_n10936);
and_8  g10560(n11662, n4312, new_n10937);
xor_4  g10561(new_n10937, new_n10936, new_n10938);
nand_5 g10562(new_n10650, new_n10649, new_n10939);
or_8   g10563(new_n10656, new_n10651, new_n10940);
and_8  g10564(new_n10940, new_n10939, new_n10941);
and_8  g10565(n12299, n10278, new_n10942);
xor_4  g10566(new_n10942, new_n10941, new_n10943);
or_8   g10567(new_n10645, new_n10644_1, new_n10944);
or_8   g10568(new_n10646, new_n10643, new_n10945);
and_8  g10569(new_n10945, new_n10944, new_n10946);
and_8  g10570(n10451, n7436, new_n10947);
and_8  g10571(n9241, n3022, new_n10948);
xor_4  g10572(new_n10948, new_n10947, new_n10949_1);
and_8  g10573(n11257, n3932, new_n10950);
and_8  g10574(n10327, n1097, new_n10951);
xor_4  g10575(new_n10951, new_n10950, new_n10952);
xor_4  g10576(new_n10952, new_n10949_1, new_n10953);
xor_4  g10577(new_n10953, new_n10946, new_n10954);
or_8   g10578(new_n10828, new_n10827, new_n10955);
or_8   g10579(new_n10829, new_n10826, new_n10956);
and_8  g10580(new_n10956, new_n10955, new_n10957);
and_8  g10581(n2393, n159, new_n10958);
and_8  g10582(n5860, n2749, new_n10959);
xor_4  g10583(new_n10959, new_n10958, new_n10960);
xnor_4 g10584(new_n10960, new_n10957, new_n10961);
xor_4  g10585(new_n10961, new_n10954, new_n10962);
xor_4  g10586(new_n10962, new_n10943, new_n10963);
xor_4  g10587(new_n10963, new_n10938, new_n10964);
or_8   g10588(new_n10745, new_n10709, new_n10965_1);
and_8  g10589(new_n10864, new_n10965_1, new_n10966);
xor_4  g10590(new_n10966, new_n10964, new_n10967);
not_8  g10591(new_n10967, new_n10968);
nor_6  g10592(new_n10812, new_n10836, new_n10969);
not_8  g10593(new_n10835, new_n10970);
or_8   g10594(new_n10970, new_n10969, new_n10971);
or_8   g10595(new_n10817, new_n10814, new_n10972);
nand_5 g10596(new_n10972, new_n10815, new_n10973);
nand_5 g10597(n12247, n7388, new_n10974);
nor_6  g10598(new_n10974, new_n10973, new_n10975);
or_8   g10599(new_n10974, new_n10765, new_n10976);
and_8  g10600(new_n10976, new_n10973, new_n10977);
or_8   g10601(new_n10977, new_n10975, new_n10978);
nand_5 g10602(n10898, n5857, new_n10979);
and_8  g10603(n12591, n12025, new_n10980);
and_8  g10604(n11876, n45, new_n10981);
xor_4  g10605(new_n10981, new_n10980, new_n10982);
xor_4  g10606(new_n10982, new_n10979, new_n10983);
xor_4  g10607(new_n10983, new_n10978, new_n10984);
not_8  g10608(new_n10984, new_n10985);
xor_4  g10609(new_n10985, new_n10971, new_n10986);
or_8   g10610(new_n10654, new_n10653, new_n10987);
or_8   g10611(new_n10655, new_n10652, new_n10988);
and_8  g10612(new_n10988, new_n10987, new_n10989);
and_8  g10613(n12705, n7456, new_n10990_1);
and_8  g10614(n11023, n8276, new_n10991);
xor_4  g10615(new_n10991, new_n10990_1, new_n10992);
xor_4  g10616(new_n10992, new_n10989, new_n10993);
and_8  g10617(n9583, n5964, new_n10994);
and_8  g10618(n12511, n7965, new_n10995);
xor_4  g10619(new_n10995, new_n10994, new_n10996);
xor_4  g10620(new_n10996, new_n10993, new_n10997);
not_8  g10621(new_n10997, new_n10998);
not_8  g10622(new_n10661, new_n10999);
or_8   g10623(new_n10662, new_n10999, new_n11000);
or_8   g10624(new_n10664, new_n10658, new_n11001);
and_8  g10625(new_n11001, new_n11000, new_n11002);
nand_5 g10626(new_n10647, new_n10642, new_n11003);
or_8   g10627(new_n10657, new_n10648, new_n11004);
and_8  g10628(new_n11004, new_n11003, new_n11005);
not_8  g10629(new_n11005, new_n11006);
xor_4  g10630(new_n11006, new_n11002, new_n11007);
or_8   g10631(new_n11007, new_n10998, new_n11008);
xor_4  g10632(new_n11005, new_n11002, new_n11009);
or_8   g10633(new_n11009, new_n10997, new_n11010);
and_8  g10634(new_n11010, new_n11008, new_n11011);
or_8   g10635(new_n11011, new_n10986, new_n11012);
xor_4  g10636(new_n10984, new_n10971, new_n11013);
and_8  g10637(new_n11009, new_n10997, new_n11014);
and_8  g10638(new_n11007, new_n10998, new_n11015);
or_8   g10639(new_n11015, new_n11014, new_n11016);
or_8   g10640(new_n11016, new_n11013, new_n11017);
and_8  g10641(new_n11017, new_n11012, new_n11018);
xor_4  g10642(new_n10834, new_n10837, new_n11019);
or_8   g10643(new_n11019, new_n10810, new_n11020);
not_8  g10644(new_n11020, new_n11021);
and_8  g10645(new_n10844, new_n10843, new_n11022);
or_8   g10646(new_n11022, new_n11021, new_n11023_1);
not_8  g10647(new_n10739, new_n11024);
or_8   g10648(new_n10742, new_n10736, new_n11025);
and_8  g10649(new_n11025, new_n11024, new_n11026);
nor_6  g10650(new_n10585, new_n10580, new_n11027);
and_8  g10651(new_n10595, new_n10586, new_n11028);
or_8   g10652(new_n11028, new_n11027, new_n11029);
not_8  g10653(new_n11029, new_n11030);
and_8  g10654(new_n11030, new_n11026, new_n11031);
nor_6  g10655(new_n11030, new_n11026, new_n11032);
or_8   g10656(new_n11032, new_n11031, new_n11033);
and_8  g10657(n3986, n3754, new_n11034);
and_8  g10658(n11423, n6776, new_n11035);
xor_4  g10659(new_n11035, new_n11034, new_n11036);
and_8  g10660(n8759, n2278, new_n11037);
and_8  g10661(n10510, n9640, new_n11038);
xor_4  g10662(new_n11038, new_n11037, new_n11039);
xnor_4 g10663(new_n11039, new_n11036, new_n11040);
and_8  g10664(n8476, n4094, new_n11041);
and_8  g10665(n5305, n753, new_n11042);
xor_4  g10666(new_n11042, new_n11041, new_n11043);
and_8  g10667(n3616, n1067, new_n11044);
and_8  g10668(n10644, n6703, new_n11045);
xor_4  g10669(new_n11045, new_n11044, new_n11046);
xor_4  g10670(new_n11046, new_n11043, new_n11047);
xor_4  g10671(new_n11047, new_n11040, new_n11048);
or_8   g10672(new_n10583, new_n10582, new_n11049);
or_8   g10673(new_n10584, new_n10581, new_n11050);
and_8  g10674(new_n11050, new_n11049, new_n11051);
or_8   g10675(new_n10592, new_n10591, new_n11052);
or_8   g10676(new_n10593, new_n10590, new_n11053);
and_8  g10677(new_n11053, new_n11052, new_n11054);
xor_4  g10678(new_n11054, new_n11051, new_n11055);
xor_4  g10679(new_n11055, new_n11048, new_n11056);
xor_4  g10680(new_n11056, new_n11033, new_n11057);
not_8  g10681(new_n10601, new_n11058);
or_8   g10682(new_n10605, new_n10596, new_n11059);
and_8  g10683(new_n11059, new_n11058, new_n11060);
and_8  g10684(new_n10821, new_n10818, new_n11061);
and_8  g10685(new_n10833, new_n10822, new_n11062);
or_8   g10686(new_n11062, new_n11061, new_n11063);
and_8  g10687(new_n10824, new_n10823, new_n11064);
nor_6  g10688(new_n10831, new_n11064, new_n11065);
or_8   g10689(new_n10717, new_n10716, new_n11066);
or_8   g10690(new_n10718, new_n10715, new_n11067);
and_8  g10691(new_n11067, new_n11066, new_n11068);
and_8  g10692(n10547, n1798, new_n11069);
and_8  g10693(n8665, n7690, new_n11070);
xnor_4 g10694(new_n11070, new_n11069, new_n11071);
and_8  g10695(n12826, n2530, new_n11072);
and_8  g10696(n11892, n1510, new_n11073);
xor_4  g10697(new_n11073, new_n11072, new_n11074);
xor_4  g10698(new_n11074, new_n11071, new_n11075);
xor_4  g10699(new_n11075, new_n11068, new_n11076);
and_8  g10700(new_n11076, new_n11065, new_n11077);
or_8   g10701(new_n10831, new_n11064, new_n11078);
not_8  g10702(new_n11074, new_n11079);
xor_4  g10703(new_n11079, new_n11071, new_n11080);
xor_4  g10704(new_n11080, new_n11068, new_n11081);
and_8  g10705(new_n11081, new_n11078, new_n11082);
or_8   g10706(new_n11082, new_n11077, new_n11083);
xor_4  g10707(new_n11083, new_n11063, new_n11084);
nand_5 g10708(n11922, n10545, new_n11085);
not_8  g10709(new_n10733, new_n11086);
or_8   g10710(new_n10735, new_n10723, new_n11087);
and_8  g10711(new_n11087, new_n11086, new_n11088);
xor_4  g10712(new_n11088, new_n11085, new_n11089);
nand_5 g10713(new_n10711, new_n10710, new_n11090);
not_8  g10714(new_n11090, new_n11091);
and_8  g10715(new_n10721, new_n10712, new_n11092);
or_8   g10716(new_n11092, new_n11091, new_n11093);
nor_6  g10717(new_n10728, new_n10727, new_n11094);
or_8   g10718(new_n10730, new_n11094, new_n11095);
and_8  g10719(new_n11095, new_n11093, new_n11096);
and_8  g10720(new_n10720, new_n11090, new_n11097);
not_8  g10721(new_n11095, new_n11098);
and_8  g10722(new_n11098, new_n11097, new_n11099);
or_8   g10723(new_n11099, new_n11096, new_n11100);
or_8   g10724(new_n702, new_n6663, new_n11101);
and_8  g10725(n10685, n5331, new_n11102);
and_8  g10726(n5645, n4499, new_n11103);
xor_4  g10727(new_n11103, new_n11102, new_n11104);
xor_4  g10728(new_n11104, new_n11101, new_n11105);
xor_4  g10729(new_n11105, new_n11100, new_n11106);
and_8  g10730(new_n11106, new_n11089, new_n11107);
not_8  g10731(new_n11085, new_n11108);
xor_4  g10732(new_n11088, new_n11108, new_n11109);
not_8  g10733(new_n11105, new_n11110);
xor_4  g10734(new_n11110, new_n11100, new_n11111);
and_8  g10735(new_n11111, new_n11109, new_n11112);
or_8   g10736(new_n11112, new_n11107, new_n11113);
or_8   g10737(new_n11113, new_n11084, new_n11114);
nor_6  g10738(new_n11082, new_n11077, new_n11115);
xor_4  g10739(new_n11115, new_n11063, new_n11116);
or_8   g10740(new_n11111, new_n11109, new_n11117);
or_8   g10741(new_n11106, new_n11089, new_n11118);
and_8  g10742(new_n11118, new_n11117, new_n11119);
or_8   g10743(new_n11119, new_n11116, new_n11120);
and_8  g10744(new_n11120, new_n11114, new_n11121);
xor_4  g10745(new_n11121, new_n11060, new_n11122);
and_8  g10746(new_n11122, new_n11057, new_n11123);
not_8  g10747(new_n11056, new_n11124);
xor_4  g10748(new_n11124, new_n11033, new_n11125);
and_8  g10749(new_n11121, new_n11060, new_n11126);
nor_6  g10750(new_n11121, new_n11060, new_n11127);
or_8   g10751(new_n11127, new_n11126, new_n11128);
and_8  g10752(new_n11128, new_n11125, new_n11129);
or_8   g10753(new_n11129, new_n11123, new_n11130);
or_8   g10754(new_n11130, new_n11023_1, new_n11131);
and_8  g10755(new_n10842, new_n11020, new_n11132);
or_8   g10756(new_n11128, new_n11125, new_n11133);
or_8   g10757(new_n11122, new_n11057, new_n11134);
and_8  g10758(new_n11134, new_n11133, new_n11135);
or_8   g10759(new_n11135, new_n11132, new_n11136);
and_8  g10760(new_n11136, new_n11131, new_n11137);
and_8  g10761(new_n11137, new_n11018, new_n11138);
nor_6  g10762(new_n11137, new_n11018, new_n11139);
or_8   g10763(new_n11139, new_n11138, new_n11140);
or_8   g10764(new_n11140, new_n10968, new_n11141);
xor_4  g10765(new_n11137, new_n11018, new_n11142);
or_8   g10766(new_n11142, new_n10967, new_n11143);
and_8  g10767(new_n11143, new_n11141, new_n11144);
and_8  g10768(new_n10606, new_n10576, new_n11145);
and_8  g10769(new_n10615, new_n10607, new_n11146);
or_8   g10770(new_n11146, new_n11145, new_n11147);
nor_6  g10771(new_n10846, new_n10866, new_n11148);
or_8   g10772(new_n10877, new_n11148, new_n11149);
or_8   g10773(new_n11149, new_n11147, new_n11150);
nor_6  g10774(new_n11146, new_n11145, new_n11151);
or_8   g10775(new_n10846, new_n10866, new_n11152);
and_8  g10776(new_n10863, new_n11152, new_n11153_1);
or_8   g10777(new_n11153_1, new_n11151, new_n11154);
and_8  g10778(new_n11154, new_n11150, new_n11155);
and_8  g10779(new_n11155, new_n11144, new_n11156);
and_8  g10780(new_n11142, new_n10967, new_n11157);
and_8  g10781(new_n11140, new_n10968, new_n11158);
or_8   g10782(new_n11158, new_n11157, new_n11159);
and_8  g10783(new_n11153_1, new_n11151, new_n11160);
and_8  g10784(new_n11149, new_n11147, new_n11161);
or_8   g10785(new_n11161, new_n11160, new_n11162);
and_8  g10786(new_n11162, new_n11159, new_n11163);
or_8   g10787(new_n11163, new_n11156, new_n11164);
or_8   g10788(new_n11164, new_n10933, new_n11165);
and_8  g10789(new_n10898_1, new_n10899, new_n11166);
or_8   g10790(new_n11162, new_n11159, new_n11167);
or_8   g10791(new_n11155, new_n11144, new_n11168);
and_8  g10792(new_n11168, new_n11167, new_n11169);
or_8   g10793(new_n11169, new_n11166, new_n11170);
and_8  g10794(new_n11170, new_n11165, new_n11171);
xor_4  g10795(new_n11171, new_n10932, new_n11172);
or_8   g10796(new_n11172, new_n10930, new_n11173);
or_8   g10797(new_n10929, new_n10905, new_n11174);
not_8  g10798(new_n10932, new_n11175);
xor_4  g10799(new_n11171, new_n11175, new_n11176);
or_8   g10800(new_n11176, new_n11174, new_n11177);
and_8  g10801(new_n11177, new_n11173, n4230);
xnor_4 g10802(new_n6224, new_n6222, n4300);
xnor_4 g10803(new_n3788, new_n3787, n4326);
nand_5 g10804(new_n1265, new_n1260, new_n11181);
and_8  g10805(n6687, n5320, new_n11182);
and_8  g10806(new_n1253, new_n1246, new_n11183);
and_8  g10807(new_n1259, new_n1254, new_n11184);
or_8   g10808(new_n11184, new_n11183, new_n11185);
xor_4  g10809(new_n11185, new_n11182, new_n11186);
nand_5 g10810(n4370, n2564, new_n11187);
not_8  g10811(new_n11187, new_n11188);
or_8   g10812(new_n1257, new_n1256, new_n11189);
or_8   g10813(new_n1258, new_n1255, new_n11190);
and_8  g10814(new_n11190, new_n11189, new_n11191);
xor_4  g10815(new_n11191, new_n11188, new_n11192);
not_8  g10816(new_n11192, new_n11193);
and_8  g10817(n6770, n5212, new_n11194);
and_8  g10818(n11877, n4189, new_n11195);
and_8  g10819(n11407, n9920, new_n11196);
xnor_4 g10820(new_n11196, new_n11195, new_n11197);
xor_4  g10821(new_n11197, new_n11194, new_n11198);
xor_4  g10822(new_n11198, new_n11193, new_n11199);
xor_4  g10823(new_n11199, new_n11186, new_n11200);
not_8  g10824(new_n11200, new_n11201);
xor_4  g10825(new_n11201, new_n11181, new_n11202);
not_8  g10826(new_n11202, new_n11203);
and_8  g10827(new_n1364, new_n1362, new_n11204);
nand_5 g10828(n8336, n2433, new_n11205);
and_8  g10829(n10928, n8819, new_n11206);
or_8   g10830(new_n1356, new_n1355, new_n11207);
and_8  g10831(new_n1356, new_n1355, new_n11208);
or_8   g10832(new_n11208, new_n1354, new_n11209);
and_8  g10833(new_n11209, new_n11207, new_n11210);
xnor_4 g10834(new_n11210, new_n11206, new_n11211);
and_8  g10835(n11728, n2226, new_n11212);
and_8  g10836(n12709, n1094, new_n11213);
xor_4  g10837(new_n11213, new_n1292, new_n11214);
xor_4  g10838(new_n11214, new_n11212, new_n11215);
xor_4  g10839(new_n11215, new_n11211, new_n11216_1);
nor_6  g10840(new_n11216_1, new_n11205, new_n11217);
and_8  g10841(new_n11216_1, new_n11205, new_n11218);
or_8   g10842(new_n11218, new_n11217, new_n11219);
and_8  g10843(new_n1358, new_n1353_1, new_n11220);
and_8  g10844(new_n1361, new_n1359, new_n11221);
or_8   g10845(new_n11221, new_n11220, new_n11222_1);
not_8  g10846(new_n11222_1, new_n11223);
xor_4  g10847(new_n11223, new_n11219, new_n11224);
xor_4  g10848(new_n11224, new_n11204, new_n11225);
and_8  g10849(new_n1426, new_n1365, new_n11226);
or_8   g10850(new_n1300, new_n1288, new_n11227);
xor_4  g10851(new_n1300, new_n1287, new_n11228);
xor_4  g10852(new_n1421, new_n1327, new_n11229);
or_8   g10853(new_n11229, new_n11228, new_n11230);
and_8  g10854(new_n11230, new_n11227, new_n11231);
and_8  g10855(new_n11231, new_n1427, new_n11232);
or_8   g10856(new_n11232, new_n11226, new_n11233);
and_8  g10857(new_n11233, new_n11225, new_n11234);
and_8  g10858(new_n11224, new_n11204, new_n11235);
nor_6  g10859(new_n11224, new_n11204, new_n11236);
or_8   g10860(new_n11236, new_n11235, new_n11237);
nor_6  g10861(new_n1364, new_n1362, new_n11238);
or_8   g10862(new_n11204, new_n11238, new_n11239);
xor_4  g10863(new_n1423, new_n1420, new_n11240);
or_8   g10864(new_n11240, new_n11239, new_n11241);
xor_4  g10865(new_n11240, new_n1365, new_n11242);
or_8   g10866(new_n1430, new_n11242, new_n11243);
and_8  g10867(new_n11243, new_n11241, new_n11244);
and_8  g10868(new_n11244, new_n11237, new_n11245);
or_8   g10869(new_n11245, new_n11234, new_n11246);
nand_5 g10870(n12069, n11967, new_n11247);
not_8  g10871(new_n11247, new_n11248);
and_8  g10872(n12391, n6254, new_n11249);
or_8   g10873(new_n1374, new_n1373, new_n11250);
or_8   g10874(new_n1377, new_n1372, new_n11251);
and_8  g10875(new_n11251, new_n11250, new_n11252);
xor_4  g10876(new_n11252, new_n11249, new_n11253);
and_8  g10877(n7160, n7159, new_n11254);
and_8  g10878(n12777, n7891, new_n11255);
and_8  g10879(n12489, n4828, new_n11256);
xor_4  g10880(new_n11256, new_n11255, new_n11257_1);
xor_4  g10881(new_n11257_1, new_n11254, new_n11258);
xor_4  g10882(new_n11258, new_n11253, new_n11259);
xor_4  g10883(new_n11259, new_n11248, new_n11260);
or_8   g10884(new_n1382, new_n1369, new_n11261);
xor_4  g10885(new_n11261, new_n11260, new_n11262);
xor_4  g10886(new_n11262, new_n1387, new_n11263);
and_8  g10887(n12947, n11222, new_n11264);
and_8  g10888(n11791, n11153, new_n11265);
or_8   g10889(new_n1398, new_n1397, new_n11266);
or_8   g10890(new_n1401, new_n1396, new_n11267);
and_8  g10891(new_n11267, new_n11266, new_n11268);
xor_4  g10892(new_n11268, new_n11265, new_n11269);
and_8  g10893(n5760, n996, new_n11270);
and_8  g10894(n5314, n1478, new_n11271);
and_8  g10895(n10990, n5767, new_n11272);
xor_4  g10896(new_n11272, new_n11271, new_n11273);
xor_4  g10897(new_n11273, new_n11270, new_n11274);
xor_4  g10898(new_n11274, new_n11269, new_n11275);
xor_4  g10899(new_n11275, new_n11264, new_n11276);
or_8   g10900(new_n1403, new_n1393, new_n11277);
and_8  g10901(new_n11277, new_n11276, new_n11278);
and_8  g10902(new_n11275, new_n11264, new_n11279);
nor_6  g10903(new_n11275, new_n11264, new_n11280);
or_8   g10904(new_n11280, new_n11279, new_n11281);
not_8  g10905(new_n11277, new_n11282);
and_8  g10906(new_n11282, new_n11281, new_n11283);
or_8   g10907(new_n11283, new_n11278, new_n11284);
and_8  g10908(new_n11284, new_n1407, new_n11285);
or_8   g10909(new_n11282, new_n11281, new_n11286);
or_8   g10910(new_n11277, new_n11276, new_n11287);
and_8  g10911(new_n11287, new_n11286, new_n11288);
and_8  g10912(new_n11288, new_n1416, new_n11289);
or_8   g10913(new_n11289, new_n11285, new_n11290);
or_8   g10914(new_n1424, new_n1419, new_n11291);
or_8   g10915(new_n11291, new_n11290, new_n11292);
nor_6  g10916(new_n11289, new_n11285, new_n11293);
nor_6  g10917(new_n1424, new_n1419, new_n11294);
or_8   g10918(new_n11294, new_n11293, new_n11295);
and_8  g10919(new_n11295, new_n11292, new_n11296_1);
xor_4  g10920(new_n11296_1, new_n11263, new_n11297);
or_8   g10921(new_n11297, new_n11246, new_n11298);
or_8   g10922(new_n11244, new_n11237, new_n11299);
or_8   g10923(new_n11233, new_n11225, new_n11300);
and_8  g10924(new_n11300, new_n11299, new_n11301);
xor_4  g10925(new_n11262, new_n1414, new_n11302);
xor_4  g10926(new_n11296_1, new_n11302, new_n11303);
or_8   g10927(new_n11303, new_n11301, new_n11304);
and_8  g10928(new_n11304, new_n11298, new_n11305);
xor_4  g10929(new_n11305, new_n11203, new_n11306);
not_8  g10930(new_n1351, new_n11307);
or_8   g10931(new_n11307, new_n1266, new_n11308);
or_8   g10932(new_n1431, new_n1352, new_n11309);
and_8  g10933(new_n11309, new_n11308, new_n11310);
xor_4  g10934(new_n11310, new_n11306, n4333);
and_8  g10935(n11877, n11757, new_n11312);
and_8  g10936(n5240, n5212, new_n11313);
and_8  g10937(n11821, n11407, new_n11314);
xor_4  g10938(new_n11314, new_n11313, new_n11315);
xor_4  g10939(new_n11315, new_n11312, new_n11316);
and_8  g10940(n11407, n5240, new_n11317);
and_8  g10941(n11877, n3172, new_n11318);
or_8   g10942(new_n11318, new_n11317, new_n11319);
and_8  g10943(n11757, n5212, new_n11320);
xnor_4 g10944(new_n11318, new_n11317, new_n11321);
or_8   g10945(new_n11321, new_n11320, new_n11322);
and_8  g10946(new_n11322, new_n11319, new_n11323);
xor_4  g10947(new_n11323, new_n11316, new_n11324);
and_8  g10948(n5320, n1333, new_n11325);
and_8  g10949(n4370, n3172, new_n11326_1);
xor_4  g10950(new_n11326_1, new_n11325, new_n11327);
xor_4  g10951(new_n11327, new_n11324, new_n11328);
and_8  g10952(n4370, n1333, new_n11329);
and_8  g10953(n11877, n1333, new_n11330);
and_8  g10954(n11757, n11407, new_n11331);
or_8   g10955(new_n11331, new_n11330, new_n11332);
and_8  g10956(n5212, n3172, new_n11333);
xnor_4 g10957(new_n11331, new_n11330, new_n11334);
or_8   g10958(new_n11334, new_n11333, new_n11335);
and_8  g10959(new_n11335, new_n11332, new_n11336);
and_8  g10960(new_n11336, new_n11329, new_n11337);
xor_4  g10961(new_n11336, new_n11329, new_n11338);
xnor_4 g10962(new_n11321, new_n11320, new_n11339);
and_8  g10963(new_n11339, new_n11338, new_n11340);
or_8   g10964(new_n11340, new_n11337, new_n11341);
xor_4  g10965(new_n11341, new_n11328, new_n11342);
and_8  g10966(n7862, n5320, new_n11343);
not_8  g10967(new_n11343, new_n11344);
nor_6  g10968(new_n11339, new_n11338, new_n11345);
or_8   g10969(new_n11345, new_n11340, new_n11346);
nand_5 g10970(new_n11346, new_n11344, new_n11347);
xor_4  g10971(new_n11346, new_n11343, new_n11348);
and_8  g10972(n7862, n4370, new_n11349);
and_8  g10973(n11407, n3172, new_n11350);
and_8  g10974(n11877, n7862, new_n11351);
or_8   g10975(new_n11351, new_n11350, new_n11352);
and_8  g10976(n11407, n7862, new_n11353);
and_8  g10977(new_n11353, new_n11318, new_n11354);
and_8  g10978(n5212, n1333, new_n11355);
or_8   g10979(new_n11355, new_n11354, new_n11356);
and_8  g10980(new_n11356, new_n11352, new_n11357);
and_8  g10981(new_n11357, new_n11349, new_n11358);
xor_4  g10982(new_n11357, new_n11349, new_n11359);
xnor_4 g10983(new_n11334, new_n11333, new_n11360);
and_8  g10984(new_n11360, new_n11359, new_n11361);
or_8   g10985(new_n11361, new_n11358, new_n11362);
or_8   g10986(new_n11362, new_n11348, new_n11363);
and_8  g10987(new_n11363, new_n11347, new_n11364);
and_8  g10988(new_n11364, new_n11342, new_n11365);
and_8  g10989(new_n11327, new_n11324, new_n11366);
and_8  g10990(new_n11326_1, new_n11325, new_n11367);
and_8  g10991(new_n11341, new_n11328, new_n11368);
xor_4  g10992(new_n11368, new_n11367, new_n11369);
nor_6  g10993(new_n11369, new_n11366, new_n11370);
and_8  g10994(new_n11314, new_n11313, new_n11371);
and_8  g10995(n11757, n4370, new_n11372);
xor_4  g10996(new_n11372, new_n11371, new_n11373);
and_8  g10997(n11821, n5212, new_n11374);
and_8  g10998(n11877, n5240, new_n11375);
and_8  g10999(n11407, n9080, new_n11376);
xnor_4 g11000(new_n11376, new_n11375, new_n11377);
xor_4  g11001(new_n11377, new_n11374, new_n11378);
xor_4  g11002(new_n11378, new_n11373, new_n11379);
or_8   g11003(new_n11315, new_n11312, new_n11380);
not_8  g11004(new_n11316, new_n11381);
or_8   g11005(new_n11323, new_n11381, new_n11382);
and_8  g11006(new_n11382, new_n11380, new_n11383);
and_8  g11007(n12000, n1333, new_n11384);
and_8  g11008(n5320, n3172, new_n11385);
and_8  g11009(n9725, n7862, new_n11386);
xnor_4 g11010(new_n11386, new_n11385, new_n11387);
xnor_4 g11011(new_n11387, new_n11384, new_n11388);
xor_4  g11012(new_n11388, new_n11383, new_n11389);
xor_4  g11013(new_n11389, new_n11379, new_n11390);
xor_4  g11014(new_n11390, new_n11370, new_n11391);
xor_4  g11015(new_n11391, new_n11365, new_n11392);
not_8  g11016(new_n11392, new_n11393);
and_8  g11017(n12000, n7862, new_n11394);
xor_4  g11018(new_n11364, new_n11342, new_n11395);
nor_6  g11019(new_n11395, new_n11394, new_n11396);
xnor_4 g11020(new_n11360, new_n11359, new_n11397);
not_8  g11021(new_n11352, new_n11398);
or_8   g11022(new_n11354, new_n11398, new_n11399);
and_8  g11023(n11407, n1333, new_n11400);
and_8  g11024(n7862, n5212, new_n11401);
and_8  g11025(new_n11401, new_n11400, new_n11402);
and_8  g11026(new_n11402, new_n11399, new_n11403);
not_8  g11027(new_n11403, new_n11404);
or_8   g11028(new_n11404, new_n11397, new_n11405);
xor_4  g11029(new_n11362, new_n11348, new_n11406);
nor_6  g11030(new_n11406, new_n11405, new_n11407_1);
and_8  g11031(new_n11395, new_n11394, new_n11408);
or_8   g11032(new_n11408, new_n11396, new_n11409);
nor_6  g11033(new_n11409, new_n11407_1, new_n11410);
or_8   g11034(new_n11410, new_n11396, new_n11411);
xor_4  g11035(new_n11411, new_n11393, new_n11412);
and_8  g11036(n8819, n6877, new_n11413);
and_8  g11037(n12709, n2464, new_n11414);
and_8  g11038(n6877, n6429, new_n11415);
and_8  g11039(new_n11415, new_n11414, new_n11416);
or_8   g11040(new_n11415, new_n11414, new_n11417);
and_8  g11041(n11728, n9400, new_n11418);
and_8  g11042(new_n11418, new_n11417, new_n11419);
or_8   g11043(new_n11419, new_n11416, new_n11420);
xor_4  g11044(new_n11420, new_n11413, new_n11421);
and_8  g11045(n11728, n2464, new_n11422);
and_8  g11046(n12709, n11311, new_n11423_1);
and_8  g11047(n9400, n6429, new_n11424);
xor_4  g11048(new_n11424, new_n11423_1, new_n11425);
xor_4  g11049(new_n11425, new_n11422, new_n11426);
xnor_4 g11050(new_n11426, new_n11421, new_n11427);
xnor_4 g11051(new_n11415, new_n11414, new_n11428);
and_8  g11052(n12709, n9400, new_n11429);
and_8  g11053(n11728, n6877, new_n11430);
and_8  g11054(new_n11430, new_n11429, new_n11431);
nand_5 g11055(new_n11431, new_n11428, new_n11432);
nor_6  g11056(new_n11432, new_n11427, new_n11433);
not_8  g11057(n6877, new_n11434);
or_8   g11058(new_n11434, new_n8667, new_n11435);
and_8  g11059(n9400, n8819, new_n11436);
or_8   g11060(new_n11424, new_n11423_1, new_n11437);
and_8  g11061(new_n11424, new_n11423_1, new_n11438);
or_8   g11062(new_n11438, new_n11422, new_n11439);
and_8  g11063(new_n11439, new_n11437, new_n11440);
xnor_4 g11064(new_n11440, new_n11436, new_n11441);
nand_5 g11065(n11728, n11311, new_n11442);
and_8  g11066(n6429, n2464, new_n11443);
and_8  g11067(n12709, n4187, new_n11444);
xnor_4 g11068(new_n11444, new_n11443, new_n11445);
xor_4  g11069(new_n11445, new_n11442, new_n11446);
xor_4  g11070(new_n11446, new_n11441, new_n11447);
xor_4  g11071(new_n11447, new_n11435, new_n11448);
and_8  g11072(new_n11420, new_n11413, new_n11449);
and_8  g11073(new_n11426, new_n11421, new_n11450);
or_8   g11074(new_n11450, new_n11449, new_n11451);
xor_4  g11075(new_n11451, new_n11448, new_n11452);
and_8  g11076(new_n11452, new_n11433, new_n11453);
and_8  g11077(n8717, n6877, new_n11454);
and_8  g11078(n11311, n6429, new_n11455);
and_8  g11079(n12709, n4203, new_n11456);
and_8  g11080(n11728, n4187, new_n11457);
xor_4  g11081(new_n11457, new_n11456, new_n11458);
xor_4  g11082(new_n11458, new_n11455, new_n11459);
or_8   g11083(new_n11444, new_n11443, new_n11460);
not_8  g11084(new_n11442, new_n11461);
or_8   g11085(new_n11445, new_n11461, new_n11462);
and_8  g11086(new_n11462, new_n11460, new_n11463);
xor_4  g11087(new_n11463, new_n11459, new_n11464);
and_8  g11088(n9400, n2433, new_n11465);
and_8  g11089(n8819, n2464, new_n11466);
xor_4  g11090(new_n11466, new_n11465, new_n11467);
xor_4  g11091(new_n11467, new_n11464, new_n11468);
and_8  g11092(new_n11440, new_n11436, new_n11469);
not_8  g11093(new_n11441, new_n11470);
and_8  g11094(new_n11446, new_n11470, new_n11471);
or_8   g11095(new_n11471, new_n11469, new_n11472);
xor_4  g11096(new_n11472, new_n11468, new_n11473);
nor_6  g11097(new_n11447, new_n11435, new_n11474);
and_8  g11098(new_n11451, new_n11448, new_n11475);
or_8   g11099(new_n11475, new_n11474, new_n11476);
xor_4  g11100(new_n11476, new_n11473, new_n11477);
not_8  g11101(new_n11477, new_n11478_1);
xor_4  g11102(new_n11478_1, new_n11454, new_n11479);
xor_4  g11103(new_n11479, new_n11453, new_n11480);
nor_6  g11104(new_n11452, new_n11433, new_n11481);
or_8   g11105(new_n11481, new_n11453, new_n11482);
xor_4  g11106(new_n11432, new_n11427, new_n11483);
not_8  g11107(new_n11483, new_n11484);
and_8  g11108(n12489, n4805, new_n11485);
and_8  g11109(n10990, n7236, new_n11486);
and_8  g11110(new_n11486, new_n11485, new_n11487);
and_8  g11111(n12489, n11478, new_n11488);
and_8  g11112(n7159, n4805, new_n11489);
xor_4  g11113(new_n11489, new_n11488, new_n11490);
or_8   g11114(new_n11490, new_n11487, new_n11491);
xor_4  g11115(new_n11490, new_n11487, new_n11492);
not_8  g11116(new_n11492, new_n11493);
and_8  g11117(n10990, n3992, new_n11494);
and_8  g11118(n7236, n5760, new_n11495);
xor_4  g11119(new_n11495, new_n11494, new_n11496);
or_8   g11120(new_n11496, new_n11493, new_n11497);
and_8  g11121(new_n11497, new_n11491, new_n11498);
and_8  g11122(n10990, n8384, new_n11499);
and_8  g11123(n7236, n1478, new_n11500);
and_8  g11124(new_n11500, new_n11499, new_n11501);
not_8  g11125(n10990, new_n11502);
or_8   g11126(new_n11502, new_n3576, new_n11503);
and_8  g11127(n5760, n3992, new_n11504);
and_8  g11128(new_n11504, new_n11503, new_n11505);
or_8   g11129(new_n11500, new_n11499, new_n11506);
nor_6  g11130(new_n11506, new_n11505, new_n11507);
or_8   g11131(new_n11507, new_n11501, new_n11508);
and_8  g11132(new_n11506, new_n11505, new_n11509);
nor_6  g11133(new_n11509, new_n11508, new_n11510);
nor_6  g11134(new_n11510, new_n11498, new_n11511);
xor_4  g11135(new_n11510, new_n11498, new_n11512);
not_8  g11136(new_n11485, new_n11513);
and_8  g11137(n11478, n7159, new_n11514);
and_8  g11138(new_n11514, new_n11513, new_n11515);
and_8  g11139(n12489, n5283, new_n11516);
and_8  g11140(n12777, n4805, new_n11517);
xor_4  g11141(new_n11517, new_n11516, new_n11518);
nor_6  g11142(new_n11518, new_n11515, new_n11519);
or_8   g11143(new_n11517, new_n11516, new_n11520);
and_8  g11144(new_n11520, new_n11515, new_n11521);
or_8   g11145(new_n11521, new_n11519, new_n11522);
and_8  g11146(new_n11522, new_n11512, new_n11523);
nor_6  g11147(new_n11523, new_n11511, new_n11524);
and_8  g11148(n6254, n4805, new_n11525);
and_8  g11149(new_n11517, new_n11516, new_n11526);
and_8  g11150(new_n11520, new_n11514, new_n11527);
or_8   g11151(new_n11527, new_n11526, new_n11528);
xor_4  g11152(new_n11528, new_n11525, new_n11529);
and_8  g11153(n7159, n5283, new_n11530);
and_8  g11154(n12489, n137, new_n11531);
and_8  g11155(n12777, n11478, new_n11532);
nor_6  g11156(new_n11532, new_n11531, new_n11533);
and_8  g11157(new_n11532, new_n11531, new_n11534);
or_8   g11158(new_n11534, new_n11533, new_n11535);
nor_6  g11159(new_n11535, new_n11530, new_n11536_1);
and_8  g11160(new_n11535, new_n11530, new_n11537);
or_8   g11161(new_n11537, new_n11536_1, new_n11538);
and_8  g11162(new_n11538, new_n11529, new_n11539);
nor_6  g11163(new_n11538, new_n11529, new_n11540);
or_8   g11164(new_n11540, new_n11539, new_n11541);
nand_5 g11165(new_n11489, new_n11488, new_n11542);
or_8   g11166(new_n11518, new_n11542, new_n11543);
nor_6  g11167(new_n11543, new_n11541, new_n11544);
and_8  g11168(new_n11543, new_n11541, new_n11545);
or_8   g11169(new_n11545, new_n11544, new_n11546);
and_8  g11170(n11791, n7236, new_n11547);
or_8   g11171(new_n11504, new_n11501, new_n11548);
and_8  g11172(new_n11548, new_n11506, new_n11549);
xor_4  g11173(new_n11549, new_n11547, new_n11550);
and_8  g11174(n8384, n5760, new_n11551);
and_8  g11175(n10990, n6358, new_n11552);
and_8  g11176(n3992, n1478, new_n11553);
nor_6  g11177(new_n11553, new_n11552, new_n11554);
and_8  g11178(new_n11553, new_n11552, new_n11555);
or_8   g11179(new_n11555, new_n11554, new_n11556);
nor_6  g11180(new_n11556, new_n11551, new_n11557);
and_8  g11181(new_n11556, new_n11551, new_n11558);
or_8   g11182(new_n11558, new_n11557, new_n11559);
xor_4  g11183(new_n11559, new_n11550, new_n11560);
and_8  g11184(new_n11508, new_n11504, new_n11561);
and_8  g11185(new_n11561, new_n11560, new_n11562);
nor_6  g11186(new_n11561, new_n11560, new_n11563);
or_8   g11187(new_n11563, new_n11562, new_n11564);
and_8  g11188(new_n11564, new_n11546, new_n11565);
nor_6  g11189(new_n11564, new_n11546, new_n11566);
or_8   g11190(new_n11566, new_n11565, new_n11567);
xor_4  g11191(new_n11567, new_n11524, new_n11568);
or_8   g11192(new_n11568, new_n11484, new_n11569);
xor_4  g11193(new_n11568, new_n11483, new_n11570);
xor_4  g11194(new_n11522, new_n11512, new_n11571);
nand_5 g11195(n12709, n6877, new_n11572);
nand_5 g11196(new_n11572, new_n11418, new_n11573);
and_8  g11197(new_n11573, new_n11428, new_n11574);
not_8  g11198(new_n11573, new_n11575);
and_8  g11199(new_n11575, new_n11417, new_n11576);
or_8   g11200(new_n11576, new_n11574, new_n11577);
or_8   g11201(new_n11577, new_n11571, new_n11578);
and_8  g11202(new_n11510, new_n11498, new_n11579);
or_8   g11203(new_n11579, new_n11511, new_n11580);
xor_4  g11204(new_n11522, new_n11580, new_n11581);
xor_4  g11205(new_n11577, new_n11581, new_n11582);
xor_4  g11206(new_n11496, new_n11492, new_n11583);
xor_4  g11207(new_n11430, new_n11429, new_n11584);
and_8  g11208(new_n11584, new_n11583, new_n11585);
not_8  g11209(new_n11572, new_n11586);
xor_4  g11210(new_n11486, new_n11485, new_n11587);
and_8  g11211(new_n11587, new_n11586, new_n11588);
xor_4  g11212(new_n11584, new_n11583, new_n11589);
and_8  g11213(new_n11589, new_n11588, new_n11590);
or_8   g11214(new_n11590, new_n11585, new_n11591);
not_8  g11215(new_n11591, new_n11592);
or_8   g11216(new_n11592, new_n11582, new_n11593);
and_8  g11217(new_n11593, new_n11578, new_n11594);
or_8   g11218(new_n11594, new_n11570, new_n11595);
and_8  g11219(new_n11595, new_n11569, new_n11596);
and_8  g11220(new_n11596, new_n11482, new_n11597);
not_8  g11221(new_n11482, new_n11598);
not_8  g11222(new_n11569, new_n11599);
xor_4  g11223(new_n11568, new_n11484, new_n11600);
not_8  g11224(new_n11578, new_n11601);
xor_4  g11225(new_n11577, new_n11571, new_n11602);
and_8  g11226(new_n11591, new_n11602, new_n11603);
or_8   g11227(new_n11603, new_n11601, new_n11604);
and_8  g11228(new_n11604, new_n11600, new_n11605);
or_8   g11229(new_n11605, new_n11599, new_n11606);
or_8   g11230(new_n11606, new_n11598, new_n11607);
or_8   g11231(new_n11596, new_n11482, new_n11608);
and_8  g11232(new_n11608, new_n11607, new_n11609);
and_8  g11233(n7159, n137, new_n11610);
and_8  g11234(n12777, n5283, new_n11611);
and_8  g11235(n12489, n6294, new_n11612);
xnor_4 g11236(new_n11612, new_n11611, new_n11613);
nor_6  g11237(new_n11613, new_n11610, new_n11614);
and_8  g11238(new_n11613, new_n11610, new_n11615);
or_8   g11239(new_n11615, new_n11614, new_n11616);
and_8  g11240(n11478, n6254, new_n11617);
or_8   g11241(new_n11532, new_n11531, new_n11618);
or_8   g11242(new_n11535, new_n11530, new_n11619);
and_8  g11243(new_n11619, new_n11618, new_n11620);
xor_4  g11244(new_n11620, new_n11617, new_n11621);
and_8  g11245(new_n11621, new_n11616, new_n11622);
nor_6  g11246(new_n11621, new_n11616, new_n11623);
or_8   g11247(new_n11623, new_n11622, new_n11624);
and_8  g11248(n11967, n4805, new_n11625);
and_8  g11249(new_n11528, new_n11525, new_n11626);
or_8   g11250(new_n11539, new_n11626, new_n11627);
xor_4  g11251(new_n11627, new_n11625, new_n11628);
and_8  g11252(new_n11628, new_n11624, new_n11629);
nor_6  g11253(new_n11628, new_n11624, new_n11630);
or_8   g11254(new_n11630, new_n11629, new_n11631);
xor_4  g11255(new_n11631, new_n11544, new_n11632);
not_8  g11256(new_n11562, new_n11633);
and_8  g11257(n6358, n5760, new_n11634);
and_8  g11258(n8384, n1478, new_n11635);
and_8  g11259(n10990, n5198, new_n11636);
xnor_4 g11260(new_n11636, new_n11635, new_n11637);
nor_6  g11261(new_n11637, new_n11634, new_n11638);
and_8  g11262(new_n11637, new_n11634, new_n11639);
or_8   g11263(new_n11639, new_n11638, new_n11640);
and_8  g11264(n11791, n3992, new_n11641);
or_8   g11265(new_n11553, new_n11552, new_n11642);
or_8   g11266(new_n11556, new_n11551, new_n11643);
and_8  g11267(new_n11643, new_n11642, new_n11644);
xor_4  g11268(new_n11644, new_n11641, new_n11645);
and_8  g11269(new_n11645, new_n11640, new_n11646);
nor_6  g11270(new_n11645, new_n11640, new_n11647);
or_8   g11271(new_n11647, new_n11646, new_n11648);
and_8  g11272(n12947, n7236, new_n11649);
and_8  g11273(new_n11549, new_n11547, new_n11650);
and_8  g11274(new_n11559, new_n11550, new_n11651);
or_8   g11275(new_n11651, new_n11650, new_n11652);
xor_4  g11276(new_n11652, new_n11649, new_n11653);
xor_4  g11277(new_n11653, new_n11648, new_n11654);
or_8   g11278(new_n11654, new_n11633, new_n11655);
and_8  g11279(new_n11653, new_n11648, new_n11656);
nor_6  g11280(new_n11653, new_n11648, new_n11657);
or_8   g11281(new_n11657, new_n11656, new_n11658);
or_8   g11282(new_n11658, new_n11562, new_n11659);
and_8  g11283(new_n11659, new_n11655, new_n11660);
and_8  g11284(new_n11660, new_n11632, new_n11661);
nor_6  g11285(new_n11660, new_n11632, new_n11662_1);
or_8   g11286(new_n11662_1, new_n11661, new_n11663);
or_8   g11287(new_n11567, new_n11524, new_n11664);
not_8  g11288(new_n11664, new_n11665);
or_8   g11289(new_n11665, new_n11565, new_n11666);
xor_4  g11290(new_n11666, new_n11663, new_n11667);
not_8  g11291(new_n11667, new_n11668);
and_8  g11292(new_n11668, new_n11609, new_n11669);
or_8   g11293(new_n11669, new_n11597, new_n11670);
and_8  g11294(new_n11670, new_n11480, new_n11671);
not_8  g11295(new_n11655, new_n11672);
and_8  g11296(n7236, n6441, new_n11673);
and_8  g11297(new_n11644, new_n11641, new_n11674);
or_8   g11298(new_n11646, new_n11674, new_n11675);
and_8  g11299(n12947, n3992, new_n11676);
and_8  g11300(n11791, n8384, new_n11677);
xor_4  g11301(new_n11677, new_n11676, new_n11678);
and_8  g11302(new_n11678, new_n11675, new_n11679);
nor_6  g11303(new_n11678, new_n11675, new_n11680);
or_8   g11304(new_n11680, new_n11679, new_n11681);
and_8  g11305(n6358, n1478, new_n11682);
and_8  g11306(n5760, n5198, new_n11683);
and_8  g11307(n10990, n1471, new_n11684);
xor_4  g11308(new_n11684, new_n11683, new_n11685);
xor_4  g11309(new_n11685, new_n11682, new_n11686);
not_8  g11310(new_n11686, new_n11687);
nor_6  g11311(new_n11636, new_n11635, new_n11688);
or_8   g11312(new_n11638, new_n11688, new_n11689);
xor_4  g11313(new_n11689, new_n11687, new_n11690);
xor_4  g11314(new_n11690, new_n11681, new_n11691);
nor_6  g11315(new_n11652, new_n11649, new_n11692);
or_8   g11316(new_n11656, new_n11692, new_n11693);
or_8   g11317(new_n11693, new_n11691, new_n11694);
xor_4  g11318(new_n11689, new_n11686, new_n11695);
xor_4  g11319(new_n11695, new_n11681, new_n11696);
not_8  g11320(new_n11693, new_n11697);
or_8   g11321(new_n11697, new_n11696, new_n11698);
and_8  g11322(new_n11698, new_n11694, new_n11699);
xor_4  g11323(new_n11699, new_n11673, new_n11700);
xor_4  g11324(new_n11700, new_n11672, new_n11701);
and_8  g11325(new_n11631, new_n11544, new_n11702);
not_8  g11326(n447, new_n11703);
or_8   g11327(new_n3601, new_n11703, new_n11704);
and_8  g11328(new_n11620, new_n11617, new_n11705);
or_8   g11329(new_n11622, new_n11705, new_n11706);
and_8  g11330(n11967, n11478, new_n11707_1);
and_8  g11331(n6254, n5283, new_n11708);
xor_4  g11332(new_n11708, new_n11707_1, new_n11709);
and_8  g11333(new_n11709, new_n11706, new_n11710);
nor_6  g11334(new_n11709, new_n11706, new_n11711);
or_8   g11335(new_n11711, new_n11710, new_n11712);
and_8  g11336(n12777, n137, new_n11713);
and_8  g11337(n7159, n6294, new_n11714);
and_8  g11338(n12489, n6797, new_n11715);
xor_4  g11339(new_n11715, new_n11714, new_n11716);
xor_4  g11340(new_n11716, new_n11713, new_n11717);
nor_6  g11341(new_n11612, new_n11611, new_n11718);
or_8   g11342(new_n11614, new_n11718, new_n11719);
xor_4  g11343(new_n11719, new_n11717, new_n11720);
xor_4  g11344(new_n11720, new_n11712, new_n11721);
nor_6  g11345(new_n11627, new_n11625, new_n11722);
or_8   g11346(new_n11629, new_n11722, new_n11723);
not_8  g11347(new_n11723, new_n11724);
and_8  g11348(new_n11724, new_n11721, new_n11725);
not_8  g11349(new_n11717, new_n11726);
xor_4  g11350(new_n11719, new_n11726, new_n11727);
xor_4  g11351(new_n11727, new_n11712, new_n11728_1);
and_8  g11352(new_n11723, new_n11728_1, new_n11729);
or_8   g11353(new_n11729, new_n11725, new_n11730);
or_8   g11354(new_n11730, new_n11704, new_n11731);
not_8  g11355(new_n11704, new_n11732);
or_8   g11356(new_n11723, new_n11728_1, new_n11733);
or_8   g11357(new_n11724, new_n11721, new_n11734);
and_8  g11358(new_n11734, new_n11733, new_n11735);
or_8   g11359(new_n11735, new_n11732, new_n11736);
and_8  g11360(new_n11736, new_n11731, new_n11737);
and_8  g11361(new_n11737, new_n11702, new_n11738);
nor_6  g11362(new_n11737, new_n11702, new_n11739);
or_8   g11363(new_n11739, new_n11738, new_n11740);
not_8  g11364(new_n11661, new_n11741);
or_8   g11365(new_n11666, new_n11663, new_n11742);
and_8  g11366(new_n11742, new_n11741, new_n11743);
and_8  g11367(new_n11743, new_n11740, new_n11744);
xor_4  g11368(new_n11737, new_n11702, new_n11745);
xor_4  g11369(new_n11660, new_n11632, new_n11746);
nor_6  g11370(new_n11665, new_n11565, new_n11747);
and_8  g11371(new_n11747, new_n11746, new_n11748);
or_8   g11372(new_n11748, new_n11661, new_n11749);
and_8  g11373(new_n11749, new_n11745, new_n11750);
or_8   g11374(new_n11750, new_n11744, new_n11751);
xor_4  g11375(new_n11751, new_n11701, new_n11752);
not_8  g11376(new_n11453, new_n11753);
xor_4  g11377(new_n11479, new_n11753, new_n11754);
and_8  g11378(new_n11606, new_n11598, new_n11755_1);
or_8   g11379(new_n11755_1, new_n11597, new_n11756);
or_8   g11380(new_n11667, new_n11756, new_n11757_1);
and_8  g11381(new_n11757_1, new_n11607, new_n11758);
or_8   g11382(new_n11758, new_n11754, new_n11759);
or_8   g11383(new_n11670, new_n11480, new_n11760);
and_8  g11384(new_n11760, new_n11759, new_n11761);
and_8  g11385(new_n11761, new_n11752, new_n11762);
or_8   g11386(new_n11762, new_n11671, new_n11763);
and_8  g11387(new_n11476, new_n11473, new_n11764);
and_8  g11388(new_n11467, new_n11464, new_n11765);
and_8  g11389(new_n11466, new_n11465, new_n11766);
and_8  g11390(new_n11472, new_n11468, new_n11767);
xor_4  g11391(new_n11767, new_n11766, new_n11768);
or_8   g11392(new_n11768, new_n11765, new_n11769);
and_8  g11393(new_n11458, new_n11455, new_n11770);
and_8  g11394(new_n11463, new_n11459, new_n11771);
or_8   g11395(new_n11771, new_n11770, new_n11772);
and_8  g11396(n9400, n8717, new_n11773);
and_8  g11397(n2464, n2433, new_n11774);
and_8  g11398(n7730, n6877, new_n11775);
xnor_4 g11399(new_n11775, new_n11774, new_n11776);
xnor_4 g11400(new_n11776, new_n11773, new_n11777);
xor_4  g11401(new_n11777, new_n11772, new_n11778);
and_8  g11402(new_n11457, new_n11456, new_n11779);
and_8  g11403(n11311, n8819, new_n11780_1);
xnor_4 g11404(new_n11780_1, new_n11779, new_n11781);
and_8  g11405(n11728, n4203, new_n11782);
and_8  g11406(n6429, n4187, new_n11783);
and_8  g11407(n12753, n12709, new_n11784);
xnor_4 g11408(new_n11784, new_n11783, new_n11785);
xor_4  g11409(new_n11785, new_n11782, new_n11786);
xor_4  g11410(new_n11786, new_n11781, new_n11787);
xor_4  g11411(new_n11787, new_n11778, new_n11788);
and_8  g11412(new_n11788, new_n11769, new_n11789);
nor_6  g11413(new_n11788, new_n11769, new_n11790);
or_8   g11414(new_n11790, new_n11789, new_n11791_1);
xor_4  g11415(new_n11791_1, new_n11764, new_n11792);
and_8  g11416(new_n11477, new_n11454, new_n11793);
not_8  g11417(new_n11793, new_n11794);
or_8   g11418(new_n11479, new_n11753, new_n11795);
and_8  g11419(new_n11795, new_n11794, new_n11796);
xor_4  g11420(new_n11796, new_n11792, new_n11797);
and_8  g11421(n11478, n447, new_n11798);
and_8  g11422(n11967, n5283, new_n11799);
and_8  g11423(n4805, n1353, new_n11800);
xnor_4 g11424(new_n11800, new_n11799, new_n11801);
xor_4  g11425(new_n11801, new_n11798, new_n11802);
and_8  g11426(new_n11716, new_n11713, new_n11803);
nor_6  g11427(new_n11719, new_n11726, new_n11804);
or_8   g11428(new_n11804, new_n11803, new_n11805);
xor_4  g11429(new_n11805, new_n11802, new_n11806);
and_8  g11430(new_n11715, new_n11714, new_n11807);
and_8  g11431(n6254, n137, new_n11808);
xnor_4 g11432(new_n11808, new_n11807, new_n11809);
and_8  g11433(n7159, n6797, new_n11810);
and_8  g11434(n12777, n6294, new_n11811);
and_8  g11435(n12489, n3146, new_n11812);
xnor_4 g11436(new_n11812, new_n11811, new_n11813);
xor_4  g11437(new_n11813, new_n11810, new_n11814);
xor_4  g11438(new_n11814, new_n11809, new_n11815);
xor_4  g11439(new_n11815, new_n11806, new_n11816);
nand_5 g11440(new_n11708, new_n11707_1, new_n11817);
or_8   g11441(new_n11720, new_n11712, new_n11818);
or_8   g11442(new_n11818, new_n11817, new_n11819);
not_8  g11443(new_n11817, new_n11820);
xor_4  g11444(new_n11709, new_n11706, new_n11821_1);
and_8  g11445(new_n11727, new_n11821_1, new_n11822);
or_8   g11446(new_n11822, new_n11820, new_n11823);
and_8  g11447(new_n11823, new_n11819, new_n11824);
nor_6  g11448(new_n11824, new_n11710, new_n11825);
or_8   g11449(new_n11825, new_n11816, new_n11826);
not_8  g11450(new_n11802, new_n11827);
xor_4  g11451(new_n11805, new_n11827, new_n11828);
xor_4  g11452(new_n11815, new_n11828, new_n11829);
or_8   g11453(new_n11824, new_n11710, new_n11830);
or_8   g11454(new_n11830, new_n11829, new_n11831);
and_8  g11455(new_n11831, new_n11826, new_n11832);
xor_4  g11456(new_n11832, new_n11725, new_n11833);
and_8  g11457(new_n11735, new_n11732, new_n11834);
or_8   g11458(new_n11738, new_n11834, new_n11835);
and_8  g11459(new_n11835, new_n11833, new_n11836);
xor_4  g11460(new_n11832, new_n11733, new_n11837);
nor_6  g11461(new_n11738, new_n11834, new_n11838);
and_8  g11462(new_n11838, new_n11837, new_n11839);
or_8   g11463(new_n11839, new_n11836, new_n11840);
nand_5 g11464(new_n11685, new_n11682, new_n11841);
or_8   g11465(new_n11689, new_n11687, new_n11842);
and_8  g11466(new_n11842, new_n11841, new_n11843);
and_8  g11467(n6441, n3992, new_n11844);
and_8  g11468(n12947, n8384, new_n11845);
and_8  g11469(n11999, n7236, new_n11846);
xnor_4 g11470(new_n11846, new_n11845, new_n11847);
xor_4  g11471(new_n11847, new_n11844, new_n11848);
not_8  g11472(new_n11848, new_n11849);
xor_4  g11473(new_n11849, new_n11843, new_n11850);
and_8  g11474(new_n11684, new_n11683, new_n11851);
and_8  g11475(n11791, n6358, new_n11852);
xnor_4 g11476(new_n11852, new_n11851, new_n11853);
and_8  g11477(n5760, n1471, new_n11854);
and_8  g11478(n5198, n1478, new_n11855);
and_8  g11479(n10990, n7646, new_n11856);
xnor_4 g11480(new_n11856, new_n11855, new_n11857);
xor_4  g11481(new_n11857, new_n11854, new_n11858);
xor_4  g11482(new_n11858, new_n11853, new_n11859);
xor_4  g11483(new_n11859, new_n11850, new_n11860);
nand_5 g11484(new_n11677, new_n11676, new_n11861);
or_8   g11485(new_n11695, new_n11681, new_n11862);
or_8   g11486(new_n11862, new_n11861, new_n11863);
not_8  g11487(new_n11861, new_n11864);
xor_4  g11488(new_n11678, new_n11675, new_n11865);
and_8  g11489(new_n11690, new_n11865, new_n11866);
or_8   g11490(new_n11866, new_n11864, new_n11867);
and_8  g11491(new_n11867, new_n11863, new_n11868);
nor_6  g11492(new_n11868, new_n11679, new_n11869);
or_8   g11493(new_n11869, new_n11860, new_n11870);
xor_4  g11494(new_n11848, new_n11843, new_n11871);
xor_4  g11495(new_n11859, new_n11871, new_n11872);
or_8   g11496(new_n11868, new_n11679, new_n11873);
or_8   g11497(new_n11873, new_n11872, new_n11874);
and_8  g11498(new_n11874, new_n11870, new_n11875);
xor_4  g11499(new_n11875, new_n11694, new_n11876_1);
not_8  g11500(new_n11673, new_n11877_1);
xor_4  g11501(new_n11697, new_n11691, new_n11878);
or_8   g11502(new_n11878, new_n11877_1, new_n11879);
xor_4  g11503(new_n11699, new_n11877_1, new_n11880);
or_8   g11504(new_n11880, new_n11655, new_n11881);
and_8  g11505(new_n11881, new_n11879, new_n11882);
and_8  g11506(new_n11882, new_n11876_1, new_n11883);
not_8  g11507(new_n11694, new_n11884);
xor_4  g11508(new_n11875, new_n11884, new_n11885);
not_8  g11509(new_n11879, new_n11886);
and_8  g11510(new_n11700, new_n11672, new_n11887);
or_8   g11511(new_n11887, new_n11886, new_n11888);
and_8  g11512(new_n11888, new_n11885, new_n11889);
or_8   g11513(new_n11889, new_n11883, new_n11890);
or_8   g11514(new_n11890, new_n11840, new_n11891);
or_8   g11515(new_n11838, new_n11837, new_n11892_1);
or_8   g11516(new_n11835, new_n11833, new_n11893);
and_8  g11517(new_n11893, new_n11892_1, new_n11894);
or_8   g11518(new_n11888, new_n11885, new_n11895);
or_8   g11519(new_n11882, new_n11876_1, new_n11896);
and_8  g11520(new_n11896, new_n11895, new_n11897);
or_8   g11521(new_n11897, new_n11894, new_n11898);
and_8  g11522(new_n11898, new_n11891, new_n11899);
or_8   g11523(new_n11749, new_n11745, new_n11900);
or_8   g11524(new_n11751, new_n11701, new_n11901);
and_8  g11525(new_n11901, new_n11900, new_n11902);
xor_4  g11526(new_n11902, new_n11899, new_n11903);
or_8   g11527(new_n11903, new_n11797, new_n11904);
not_8  g11528(new_n11764, new_n11905);
xor_4  g11529(new_n11791_1, new_n11905, new_n11906);
xor_4  g11530(new_n11796, new_n11906, new_n11907);
and_8  g11531(new_n11902, new_n11899, new_n11908);
nor_6  g11532(new_n11902, new_n11899, new_n11909);
or_8   g11533(new_n11909, new_n11908, new_n11910);
or_8   g11534(new_n11910, new_n11907, new_n11911);
and_8  g11535(new_n11911, new_n11904, new_n11912);
and_8  g11536(new_n11912, new_n11763, new_n11913);
not_8  g11537(new_n11701, new_n11914);
xor_4  g11538(new_n11751, new_n11914, new_n11915);
and_8  g11539(new_n11758, new_n11754, new_n11916);
or_8   g11540(new_n11916, new_n11671, new_n11917_1);
or_8   g11541(new_n11917_1, new_n11915, new_n11918);
and_8  g11542(new_n11918, new_n11759, new_n11919_1);
and_8  g11543(new_n11910, new_n11907, new_n11920);
and_8  g11544(new_n11903, new_n11797, new_n11921);
or_8   g11545(new_n11921, new_n11920, new_n11922_1);
and_8  g11546(new_n11922_1, new_n11919_1, new_n11923);
or_8   g11547(new_n11923, new_n11913, new_n11924);
or_8   g11548(new_n11924, new_n11412, new_n11925);
not_8  g11549(new_n11412, new_n11926);
or_8   g11550(new_n11922_1, new_n11919_1, new_n11927);
or_8   g11551(new_n11912, new_n11763, new_n11928);
and_8  g11552(new_n11928, new_n11927, new_n11929);
and_8  g11553(new_n11929, new_n11926, new_n11930);
and_8  g11554(new_n11924, new_n11412, new_n11931);
or_8   g11555(new_n11931, new_n11930, new_n11932);
xor_4  g11556(new_n11409, new_n11407_1, new_n11933);
not_8  g11557(new_n11933, new_n11934);
xor_4  g11558(new_n11406, new_n11405, new_n11935);
and_8  g11559(new_n11667, new_n11756, new_n11936);
or_8   g11560(new_n11936, new_n11669, new_n11937);
or_8   g11561(new_n11937, new_n11935, new_n11938);
not_8  g11562(new_n11935, new_n11939);
or_8   g11563(new_n11668, new_n11609, new_n11940);
and_8  g11564(new_n11940, new_n11757_1, new_n11941);
and_8  g11565(new_n11941, new_n11939, new_n11942);
and_8  g11566(new_n11937, new_n11935, new_n11943);
or_8   g11567(new_n11943, new_n11942, new_n11944);
xor_4  g11568(new_n11404, new_n11397, new_n11945);
not_8  g11569(new_n11945, new_n11946);
xor_4  g11570(new_n11594, new_n11600, new_n11947);
and_8  g11571(new_n11947, new_n11946, new_n11948);
not_8  g11572(new_n11948, new_n11949);
xor_4  g11573(new_n11592, new_n11582, new_n11950);
not_8  g11574(new_n11353, new_n11951);
and_8  g11575(new_n11355, new_n11951, new_n11952);
nand_5 g11576(new_n11952, new_n11398, new_n11953);
or_8   g11577(new_n11952, new_n11399, new_n11954);
and_8  g11578(new_n11954, new_n11953, new_n11955);
not_8  g11579(new_n11955, new_n11956);
or_8   g11580(new_n11956, new_n11950, new_n11957);
xor_4  g11581(new_n11955, new_n11950, new_n11958);
xor_4  g11582(new_n11587, new_n11586, new_n11959);
and_8  g11583(new_n11959, new_n11353, new_n11960);
xor_4  g11584(new_n11401, new_n11400, new_n11961);
or_8   g11585(new_n11961, new_n11960, new_n11962);
xor_4  g11586(new_n11589, new_n11588, new_n11963);
xnor_4 g11587(new_n11961, new_n11960, new_n11964);
or_8   g11588(new_n11964, new_n11963, new_n11965);
and_8  g11589(new_n11965, new_n11962, new_n11966);
or_8   g11590(new_n11966, new_n11958, new_n11967_1);
and_8  g11591(new_n11967_1, new_n11957, new_n11968);
xor_4  g11592(new_n11594, new_n11570, new_n11969);
and_8  g11593(new_n11969, new_n11945, new_n11970);
or_8   g11594(new_n11970, new_n11948, new_n11971);
or_8   g11595(new_n11971, new_n11968, new_n11972);
and_8  g11596(new_n11972, new_n11949, new_n11973);
or_8   g11597(new_n11973, new_n11944, new_n11974);
and_8  g11598(new_n11974, new_n11938, new_n11975);
or_8   g11599(new_n11975, new_n11934, new_n11976);
xor_4  g11600(new_n11761, new_n11915, new_n11977);
xor_4  g11601(new_n11975, new_n11933, new_n11978);
or_8   g11602(new_n11978, new_n11977, new_n11979);
and_8  g11603(new_n11979, new_n11976, new_n11980);
or_8   g11604(new_n11980, new_n11932, new_n11981);
and_8  g11605(new_n11981, new_n11925, new_n11982);
and_8  g11606(new_n11904, new_n11919_1, new_n11983);
or_8   g11607(new_n11983, new_n11921, new_n11984);
nand_5 g11608(new_n11391, new_n11365, new_n11985);
or_8   g11609(new_n11411, new_n11393, new_n11986);
and_8  g11610(new_n11986, new_n11985, new_n11987);
nand_5 g11611(new_n11826, new_n11819, new_n11988);
not_8  g11612(new_n11988, new_n11989);
or_8   g11613(new_n11846, new_n11845, new_n11990);
or_8   g11614(new_n11847, new_n11844, new_n11991);
and_8  g11615(new_n11991, new_n11990, new_n11992);
nand_5 g11616(n4805, n4436, new_n11993);
and_8  g11617(n8384, n6441, new_n11994);
and_8  g11618(n11791, n5198, new_n11995);
xor_4  g11619(new_n11995, new_n11994, new_n11996);
xor_4  g11620(new_n11996, new_n11993, new_n11997);
xor_4  g11621(new_n11997, new_n11992, new_n11998);
and_8  g11622(n7159, n3146, new_n11999_1);
and_8  g11623(n11967, n137, new_n12000_1);
xor_4  g11624(new_n12000_1, new_n11999_1, new_n12001);
and_8  g11625(n6294, n6254, new_n12002);
and_8  g11626(n12947, n6358, new_n12003);
xor_4  g11627(new_n12003, new_n12002, new_n12004);
and_8  g11628(n11407, n6826, new_n12005_1);
and_8  g11629(n7862, n6604, new_n12006);
xor_4  g11630(new_n12006, new_n12005_1, new_n12007);
xor_4  g11631(new_n12007, new_n12004, new_n12008);
xor_4  g11632(new_n12008, new_n12001, new_n12009);
xor_4  g11633(new_n12009, new_n11998, new_n12010);
and_8  g11634(n6429, n4203, new_n12011);
nand_5 g11635(new_n11808, new_n11807, new_n12012);
or_8   g11636(new_n11814, new_n11809, new_n12013);
and_8  g11637(new_n12013, new_n12012, new_n12014_1);
xor_4  g11638(new_n12014_1, new_n12011, new_n12015);
xor_4  g11639(new_n12015, new_n12010, new_n12016);
or_8   g11640(new_n11805, new_n11827, new_n12017);
or_8   g11641(new_n11815, new_n11806, new_n12018);
and_8  g11642(new_n12018, new_n12017, new_n12019);
not_8  g11643(new_n12019, new_n12020_1);
nand_5 g11644(new_n11848, new_n11843, new_n12021);
or_8   g11645(new_n11859, new_n11850, new_n12022);
and_8  g11646(new_n12022, new_n12021, new_n12023);
and_8  g11647(n11478, n1353, new_n12024);
or_8   g11648(new_n11801, new_n11798, new_n12025_1);
and_8  g11649(new_n12025_1, new_n11799, new_n12026);
nand_5 g11650(new_n12026, new_n12024, new_n12027);
and_8  g11651(new_n12024, new_n11704, new_n12028);
or_8   g11652(new_n12028, new_n12026, new_n12029);
and_8  g11653(new_n12029, new_n12027, new_n12030);
and_8  g11654(new_n11812, new_n11811, new_n12031);
or_8   g11655(new_n11812, new_n11811, new_n12032);
and_8  g11656(new_n12032, new_n11810, new_n12033);
or_8   g11657(new_n12033, new_n12031, new_n12034);
xor_4  g11658(new_n12034, new_n12030, new_n12035);
xor_4  g11659(new_n12035, new_n12023, new_n12036);
xor_4  g11660(new_n12036, new_n12020_1, new_n12037);
or_8   g11661(new_n12037, new_n12016, new_n12038);
not_8  g11662(new_n12016, new_n12039);
xor_4  g11663(new_n12036, new_n12019, new_n12040);
or_8   g11664(new_n12040, new_n12039, new_n12041);
and_8  g11665(new_n12041, new_n12038, new_n12042);
nand_5 g11666(new_n11368, new_n11367, new_n12043);
or_8   g11667(new_n11390, new_n11370, new_n12044_1);
and_8  g11668(new_n12044_1, new_n12043, new_n12045);
and_8  g11669(n12777, n6797, new_n12046);
xor_4  g11670(new_n12046, new_n12045, new_n12047);
and_8  g11671(new_n12047, new_n12042, new_n12048);
nor_6  g11672(new_n12047, new_n12042, new_n12049);
or_8   g11673(new_n12049, new_n12048, new_n12050);
or_8   g11674(new_n12050, new_n11989, new_n12051);
and_8  g11675(new_n12050, new_n11989, new_n12052);
not_8  g11676(new_n12052, new_n12053);
and_8  g11677(new_n12053, new_n12051, new_n12054);
and_8  g11678(new_n12054, new_n11987, new_n12055);
not_8  g11679(new_n11985, new_n12056);
nor_6  g11680(new_n11411, new_n11393, new_n12057);
or_8   g11681(new_n12057, new_n12056, new_n12058);
not_8  g11682(new_n12051, new_n12059);
or_8   g11683(new_n12052, new_n12059, new_n12060);
and_8  g11684(new_n12060, new_n12058, new_n12061);
or_8   g11685(new_n12061, new_n12055, new_n12062);
or_8   g11686(new_n12062, new_n11984, new_n12063);
or_8   g11687(new_n11920, new_n11763, new_n12064);
and_8  g11688(new_n12064, new_n11911, new_n12065);
or_8   g11689(new_n12060, new_n12058, new_n12066);
or_8   g11690(new_n12054, new_n11987, new_n12067);
and_8  g11691(new_n12067, new_n12066, new_n12068);
or_8   g11692(new_n12068, new_n12065, new_n12069_1);
and_8  g11693(new_n12069_1, new_n12063, new_n12070);
or_8   g11694(new_n11791_1, new_n11905, new_n12071);
or_8   g11695(new_n11796, new_n11792, new_n12072);
and_8  g11696(new_n12072, new_n12071, new_n12073);
and_8  g11697(new_n11832, new_n11725, new_n12074);
or_8   g11698(new_n11836, new_n12074, new_n12075);
and_8  g11699(new_n12075, new_n12073, new_n12076_1);
not_8  g11700(new_n12071, new_n12077);
xnor_4 g11701(new_n11478_1, new_n11454, new_n12078);
and_8  g11702(new_n12078, new_n11453, new_n12079);
or_8   g11703(new_n12079, new_n11793, new_n12080);
and_8  g11704(new_n12080, new_n11906, new_n12081);
or_8   g11705(new_n12081, new_n12077, new_n12082);
nor_6  g11706(new_n11836, new_n12074, new_n12083);
and_8  g11707(new_n12083, new_n12082, new_n12084);
or_8   g11708(new_n12084, new_n12076_1, new_n12085);
nand_5 g11709(new_n11875, new_n11884, new_n12086);
and_8  g11710(new_n11896, new_n12086, new_n12087);
and_8  g11711(new_n11777, new_n11772, new_n12088);
and_8  g11712(new_n11787, new_n11778, new_n12089);
or_8   g11713(new_n12089, new_n12088, new_n12090);
or_8   g11714(new_n11775, new_n11774, new_n12091);
or_8   g11715(new_n11776, new_n11773, new_n12092);
and_8  g11716(new_n12092, new_n12091, new_n12093);
and_8  g11717(n5283, n447, new_n12094);
and_8  g11718(n11999, n3992, new_n12095);
xor_4  g11719(new_n12095, new_n12094, new_n12096);
xnor_4 g11720(new_n12096, new_n12093, new_n12097);
xor_4  g11721(new_n12097, new_n12090, new_n12098);
and_8  g11722(n7646, n5760, new_n12099);
and_8  g11723(n10990, n4722, new_n12100);
xor_4  g11724(new_n12100, new_n12099, new_n12101);
xor_4  g11725(new_n12101, new_n12098, new_n12102);
xor_4  g11726(new_n12102, new_n12087, new_n12103);
xor_4  g11727(new_n12103, new_n12085, new_n12104);
and_8  g11728(new_n11897, new_n11894, new_n12105);
or_8   g11729(new_n11908, new_n12105, new_n12106);
and_8  g11730(new_n11767, new_n11766, new_n12107);
or_8   g11731(new_n11789, new_n12107, new_n12108);
nor_6  g11732(new_n11388, new_n11383, new_n12109);
and_8  g11733(new_n11389, new_n11379, new_n12110);
nor_6  g11734(new_n12110, new_n12109, new_n12111_1);
or_8   g11735(new_n11784, new_n11783, new_n12112);
or_8   g11736(new_n11785, new_n11782, new_n12113);
and_8  g11737(new_n12113, new_n12112, new_n12114);
nand_5 g11738(n12000, n3172, new_n12115);
and_8  g11739(n9725, n1333, new_n12116);
and_8  g11740(n12709, n10174, new_n12117);
xor_4  g11741(new_n12117, new_n12116, new_n12118);
xor_4  g11742(new_n12118, new_n12115, new_n12119);
xor_4  g11743(new_n12119, new_n12114, new_n12120);
nand_5 g11744(new_n11780_1, new_n11779, new_n12121);
or_8   g11745(new_n11786, new_n11781, new_n12122);
and_8  g11746(new_n12122, new_n12121, new_n12123);
or_8   g11747(new_n11856, new_n11855, new_n12124);
or_8   g11748(new_n11857, new_n11854, new_n12125);
and_8  g11749(new_n12125, new_n12124, new_n12126);
and_8  g11750(n6877, n1198, new_n12127);
and_8  g11751(n12753, n11728, new_n12128);
xor_4  g11752(new_n12128, new_n12127, new_n12129);
xor_4  g11753(new_n12129, new_n12126, new_n12130);
xor_4  g11754(new_n12130, new_n12123, new_n12131);
xor_4  g11755(new_n12131, new_n12120, new_n12132);
xor_4  g11756(new_n12132, new_n12111_1, new_n12133);
nand_5 g11757(n12489, n4938, new_n12134);
or_8   g11758(new_n11386, new_n11385, new_n12135);
or_8   g11759(new_n11387, new_n11384, new_n12136);
and_8  g11760(new_n12136, new_n12135, new_n12137);
and_8  g11761(n11757, n5320, new_n12138);
and_8  g11762(n9080, n5212, new_n12139);
xnor_4 g11763(new_n12139, new_n12138, new_n12140);
and_8  g11764(n11877, n11821, new_n12141);
and_8  g11765(n5240, n4370, new_n12142);
xor_4  g11766(new_n12142, new_n12141, new_n12143);
xor_4  g11767(new_n12143, new_n12140, new_n12144);
xor_4  g11768(new_n12144, new_n12137, new_n12145_1);
and_8  g11769(n9400, n7730, new_n12146);
and_8  g11770(n11311, n2433, new_n12147);
xor_4  g11771(new_n12147, new_n12146, new_n12148);
not_8  g11772(new_n12148, new_n12149);
xor_4  g11773(new_n12149, new_n12145_1, new_n12150);
or_8   g11774(new_n11376, new_n11375, new_n12151);
or_8   g11775(new_n11377, new_n11374, new_n12152);
nand_5 g11776(new_n12152, new_n12151, new_n12153);
nor_6  g11777(new_n11372, new_n11371, new_n12154);
and_8  g11778(new_n11378, new_n11373, new_n12155);
or_8   g11779(new_n12155, new_n12154, new_n12156);
xor_4  g11780(new_n12156, new_n12153, new_n12157);
xor_4  g11781(new_n12157, new_n12150, new_n12158);
xor_4  g11782(new_n12158, new_n12134, new_n12159);
xor_4  g11783(new_n12159, new_n12133, new_n12160);
or_8   g11784(new_n12160, new_n12108, new_n12161);
not_8  g11785(new_n12108, new_n12162);
and_8  g11786(new_n12159, new_n12133, new_n12163);
nor_6  g11787(new_n12159, new_n12133, new_n12164);
or_8   g11788(new_n12164, new_n12163, new_n12165);
or_8   g11789(new_n12165, new_n12162, new_n12166);
and_8  g11790(new_n12166, new_n12161, new_n12167);
and_8  g11791(new_n11870, new_n11863, new_n12168);
and_8  g11792(n8819, n4187, new_n12169);
and_8  g11793(n1478, n1471, new_n12170);
xor_4  g11794(new_n12170, new_n12169, new_n12171);
and_8  g11795(n8717, n2464, new_n12172);
and_8  g11796(n10022, n7236, new_n12173);
xor_4  g11797(new_n12173, new_n12172, new_n12174);
xnor_4 g11798(new_n12174, new_n12171, new_n12175);
nand_5 g11799(new_n11852, new_n11851, new_n12176);
or_8   g11800(new_n11858, new_n11853, new_n12177);
and_8  g11801(new_n12177, new_n12176, new_n12178);
xor_4  g11802(new_n12178, new_n12175, new_n12179);
xor_4  g11803(new_n12179, new_n12168, new_n12180);
or_8   g11804(new_n12180, new_n12167, new_n12181);
and_8  g11805(new_n12165, new_n12162, new_n12182);
and_8  g11806(new_n12160, new_n12108, new_n12183);
or_8   g11807(new_n12183, new_n12182, new_n12184);
not_8  g11808(new_n12180, new_n12185);
or_8   g11809(new_n12185, new_n12184, new_n12186);
and_8  g11810(new_n12186, new_n12181, new_n12187);
xor_4  g11811(new_n12187, new_n12106, new_n12188);
or_8   g11812(new_n12188, new_n12104, new_n12189);
and_8  g11813(new_n12103, new_n12085, new_n12190);
nor_6  g11814(new_n12103, new_n12085, new_n12191);
or_8   g11815(new_n12191, new_n12190, new_n12192);
nor_6  g11816(new_n11908, new_n12105, new_n12193);
xor_4  g11817(new_n12187, new_n12193, new_n12194);
or_8   g11818(new_n12194, new_n12192, new_n12195);
and_8  g11819(new_n12195, new_n12189, new_n12196);
xor_4  g11820(new_n12196, new_n12070, new_n12197);
xor_4  g11821(new_n12197, new_n11982, n4378);
xor_4  g11822(new_n4044, new_n3954, n4397);
xor_4  g11823(new_n4326_1, new_n4134, n4553);
xor_4  g11824(new_n875, new_n866, n4686);
xnor_4 g11825(new_n10019, new_n10001, n4689);
xor_4  g11826(new_n5187, new_n5182, n4733);
xnor_4 g11827(new_n2096_1, new_n2089, n4757);
xnor_4 g11828(new_n5178, new_n5176, n4971);
xnor_4 g11829(new_n6920, new_n6918, n5030);
xnor_4 g11830(new_n3043, new_n3008, n5034);
xnor_4 g11831(new_n3035, new_n3027, n5094);
and_8  g11832(new_n11191, new_n11188, new_n12209);
not_8  g11833(new_n11198, new_n12210);
and_8  g11834(new_n12210, new_n11192, new_n12211);
or_8   g11835(new_n12211, new_n12209, new_n12212);
and_8  g11836(n5320, n2564, new_n12213);
and_8  g11837(n4370, n4189, new_n12214);
xor_4  g11838(new_n12214, new_n12213, new_n12215);
and_8  g11839(new_n12215, new_n12212, new_n12216);
nor_6  g11840(new_n12215, new_n12212, new_n12217);
or_8   g11841(new_n12217, new_n12216, new_n12218);
and_8  g11842(n11877, n6770, new_n12219);
or_8   g11843(new_n11196, new_n11195, new_n12220);
or_8   g11844(new_n11197, new_n11194, new_n12221_1);
and_8  g11845(new_n12221_1, new_n12220, new_n12222);
xor_4  g11846(new_n12222, new_n12219, new_n12223);
and_8  g11847(n9920, n5212, new_n12224);
and_8  g11848(n11407, n3627, new_n12225);
xor_4  g11849(new_n12225, new_n12224, new_n12226);
xor_4  g11850(new_n12226, new_n12223, new_n12227);
not_8  g11851(new_n12227, new_n12228);
or_8   g11852(new_n12228, new_n12218, new_n12229);
xor_4  g11853(new_n12215, new_n12212, new_n12230);
or_8   g11854(new_n12227, new_n12230, new_n12231);
and_8  g11855(new_n12231, new_n12229, new_n12232);
and_8  g11856(new_n11185, new_n11182, new_n12233);
and_8  g11857(new_n11199, new_n11186, new_n12234);
or_8   g11858(new_n12234, new_n12233, new_n12235);
and_8  g11859(new_n12235, new_n12232, new_n12236);
and_8  g11860(new_n12222, new_n12219, new_n12237);
and_8  g11861(new_n12226, new_n12223, new_n12238);
or_8   g11862(new_n12238, new_n12237, new_n12239);
and_8  g11863(n12000, n2564, new_n12240);
and_8  g11864(n5320, n4189, new_n12241);
and_8  g11865(n9725, n6687, new_n12242);
xnor_4 g11866(new_n12242, new_n12241, new_n12243);
xor_4  g11867(new_n12243, new_n12240, new_n12244);
xor_4  g11868(new_n12244, new_n12239, new_n12245);
and_8  g11869(new_n12225, new_n12224, new_n12246);
and_8  g11870(n6770, n4370, new_n12247_1);
xnor_4 g11871(new_n12247_1, new_n12246, new_n12248);
and_8  g11872(n5212, n3627, new_n12249);
and_8  g11873(n11877, n9920, new_n12250);
and_8  g11874(n11407, n4516, new_n12251);
xnor_4 g11875(new_n12251, new_n12250, new_n12252);
xor_4  g11876(new_n12252, new_n12249, new_n12253);
xor_4  g11877(new_n12253, new_n12248, new_n12254);
or_8   g11878(new_n12254, new_n12245, new_n12255);
not_8  g11879(new_n12255, new_n12256);
and_8  g11880(new_n12254, new_n12245, new_n12257);
or_8   g11881(new_n12257, new_n12256, new_n12258);
nand_5 g11882(new_n12214, new_n12213, new_n12259);
or_8   g11883(new_n12229, new_n12259, new_n12260);
not_8  g11884(new_n12259, new_n12261);
and_8  g11885(new_n12227, new_n12230, new_n12262);
or_8   g11886(new_n12262, new_n12261, new_n12263);
and_8  g11887(new_n12263, new_n12260, new_n12264);
or_8   g11888(new_n12264, new_n12216, new_n12265);
or_8   g11889(new_n12265, new_n12258, new_n12266);
xor_4  g11890(new_n12254, new_n12245, new_n12267);
not_8  g11891(new_n12216, new_n12268);
and_8  g11892(new_n12262, new_n12261, new_n12269);
and_8  g11893(new_n12229, new_n12259, new_n12270);
or_8   g11894(new_n12270, new_n12269, new_n12271);
and_8  g11895(new_n12271, new_n12268, new_n12272);
or_8   g11896(new_n12272, new_n12267, new_n12273);
and_8  g11897(new_n12273, new_n12266, new_n12274);
xor_4  g11898(new_n12274, new_n12236, new_n12275);
nand_5 g11899(n12000, n6687, new_n12276);
not_8  g11900(new_n12276, new_n12277);
xor_4  g11901(new_n12235, new_n12232, new_n12278);
and_8  g11902(new_n12278, new_n12277, new_n12279);
not_8  g11903(new_n11181, new_n12280);
and_8  g11904(new_n11200, new_n12280, new_n12281);
and_8  g11905(new_n12228, new_n12218, new_n12282);
or_8   g11906(new_n12282, new_n12262, new_n12283);
xor_4  g11907(new_n12235, new_n12283, new_n12284);
or_8   g11908(new_n12284, new_n12276, new_n12285);
or_8   g11909(new_n12278, new_n12277, new_n12286);
and_8  g11910(new_n12286, new_n12285, new_n12287);
and_8  g11911(new_n12287, new_n12281, new_n12288);
or_8   g11912(new_n12288, new_n12279, new_n12289);
xor_4  g11913(new_n12289, new_n12275, new_n12290);
and_8  g11914(n8717, n8336, new_n12291);
and_8  g11915(n6429, n2226, new_n12292);
and_8  g11916(n11728, n1094, new_n12293);
and_8  g11917(n12709, n10678, new_n12294);
xor_4  g11918(new_n12294, new_n12293, new_n12295);
xor_4  g11919(new_n12295, new_n12292, new_n12296);
or_8   g11920(new_n11213, new_n1292, new_n12297);
and_8  g11921(new_n11213, new_n1292, new_n12298);
or_8   g11922(new_n12298, new_n11212, new_n12299_1);
and_8  g11923(new_n12299_1, new_n12297, new_n12300);
xor_4  g11924(new_n12300, new_n12296, new_n12301);
and_8  g11925(n10928, n2433, new_n12302);
and_8  g11926(n8819, n6986, new_n12303);
xor_4  g11927(new_n12303, new_n12302, new_n12304);
xor_4  g11928(new_n12304, new_n12301, new_n12305);
and_8  g11929(new_n11210, new_n11206, new_n12306);
not_8  g11930(new_n11211, new_n12307);
and_8  g11931(new_n11215, new_n12307, new_n12308);
or_8   g11932(new_n12308, new_n12306, new_n12309);
xor_4  g11933(new_n12309, new_n12305, new_n12310);
nor_6  g11934(new_n11223, new_n11219, new_n12311);
or_8   g11935(new_n12311, new_n11217, new_n12312);
xor_4  g11936(new_n12312, new_n12310, new_n12313);
and_8  g11937(new_n12313, new_n12291, new_n12314);
xor_4  g11938(new_n12313, new_n12291, new_n12315);
and_8  g11939(new_n12315, new_n11235, new_n12316);
or_8   g11940(new_n12316, new_n12314, new_n12317);
and_8  g11941(new_n12312, new_n12310, new_n12318);
and_8  g11942(new_n12295, new_n12292, new_n12319);
and_8  g11943(new_n12300, new_n12296, new_n12320);
nor_6  g11944(new_n12320, new_n12319, new_n12321);
and_8  g11945(n10928, n8717, new_n12322);
and_8  g11946(n6986, n2433, new_n12323);
and_8  g11947(n8336, n7730, new_n12324);
xnor_4 g11948(new_n12324, new_n12323, new_n12325);
xor_4  g11949(new_n12325, new_n12322, new_n12326);
xnor_4 g11950(new_n12326, new_n12321, new_n12327);
and_8  g11951(new_n12294, new_n12293, new_n12328);
and_8  g11952(n8819, n2226, new_n12329);
xnor_4 g11953(new_n12329, new_n12328, new_n12330);
and_8  g11954(n11728, n10678, new_n12331);
and_8  g11955(n6429, n1094, new_n12332);
and_8  g11956(n12709, n7320, new_n12333);
xnor_4 g11957(new_n12333, new_n12332, new_n12334);
xor_4  g11958(new_n12334, new_n12331, new_n12335);
xor_4  g11959(new_n12335, new_n12330, new_n12336);
xor_4  g11960(new_n12336, new_n12327, new_n12337);
nand_5 g11961(new_n12304, new_n12301, new_n12338);
nand_5 g11962(new_n12303, new_n12302, new_n12339);
and_8  g11963(new_n12309, new_n12305, new_n12340);
xor_4  g11964(new_n12340, new_n12339, new_n12341);
and_8  g11965(new_n12341, new_n12338, new_n12342);
xor_4  g11966(new_n12342, new_n12337, new_n12343);
xor_4  g11967(new_n12343, new_n12318, new_n12344);
xor_4  g11968(new_n12344, new_n12317, new_n12345);
not_8  g11969(new_n11235, new_n12346);
not_8  g11970(new_n12291, new_n12347);
xor_4  g11971(new_n12313, new_n12347, new_n12348);
or_8   g11972(new_n12348, new_n12346, new_n12349);
or_8   g11973(new_n12315, new_n11235, new_n12350);
and_8  g11974(new_n12350, new_n12349, new_n12351);
and_8  g11975(new_n11303, new_n11301, new_n12352);
or_8   g11976(new_n12352, new_n11234, new_n12353);
or_8   g11977(new_n12353, new_n12351, new_n12354);
and_8  g11978(n11222, n6441, new_n12355);
not_8  g11979(new_n12355, new_n12356);
and_8  g11980(new_n11268, new_n11265, new_n12357);
and_8  g11981(new_n11274, new_n11269, new_n12358);
or_8   g11982(new_n12358, new_n12357, new_n12359);
and_8  g11983(n12947, n11153, new_n12360);
and_8  g11984(n11791, n5314, new_n12361);
xor_4  g11985(new_n12361, new_n12360, new_n12362);
xor_4  g11986(new_n12362, new_n12359, new_n12363);
and_8  g11987(n1478, n996, new_n12364);
and_8  g11988(n10990, n5319, new_n12365);
and_8  g11989(n5767, n5760, new_n12366);
xor_4  g11990(new_n12366, new_n12365, new_n12367);
xor_4  g11991(new_n12367, new_n12364, new_n12368);
not_8  g11992(new_n12368, new_n12369);
or_8   g11993(new_n11272, new_n11271, new_n12370);
and_8  g11994(new_n11272, new_n11271, new_n12371);
or_8   g11995(new_n12371, new_n11270, new_n12372);
nand_5 g11996(new_n12372, new_n12370, new_n12373);
xor_4  g11997(new_n12373, new_n12369, new_n12374);
xor_4  g11998(new_n12374, new_n12363, new_n12375);
or_8   g11999(new_n11278, new_n11279, new_n12376);
and_8  g12000(new_n12376, new_n12375, new_n12377);
nor_6  g12001(new_n12376, new_n12375, new_n12378);
or_8   g12002(new_n12378, new_n12377, new_n12379);
or_8   g12003(new_n12379, new_n12356, new_n12380);
xor_4  g12004(new_n12376, new_n12375, new_n12381);
or_8   g12005(new_n12381, new_n12355, new_n12382);
and_8  g12006(new_n12382, new_n12380, new_n12383);
xor_4  g12007(new_n12383, new_n11289, new_n12384);
and_8  g12008(new_n11262, new_n1414, new_n12385);
and_8  g12009(n12069, n447, new_n12386);
and_8  g12010(n12777, n7160, new_n12387);
and_8  g12011(n7159, n4828, new_n12388);
and_8  g12012(n12489, n2515, new_n12389);
xor_4  g12013(new_n12389, new_n12388, new_n12390);
xor_4  g12014(new_n12390, new_n12387, new_n12391_1);
or_8   g12015(new_n11256, new_n11255, new_n12392);
and_8  g12016(new_n11256, new_n11255, new_n12393);
or_8   g12017(new_n12393, new_n11254, new_n12394);
and_8  g12018(new_n12394, new_n12392, new_n12395);
and_8  g12019(new_n12395, new_n12391_1, new_n12396);
nor_6  g12020(new_n12395, new_n12391_1, new_n12397);
or_8   g12021(new_n12397, new_n12396, new_n12398);
and_8  g12022(n12391, n11967, new_n12399);
and_8  g12023(n7891, n6254, new_n12400);
xor_4  g12024(new_n12400, new_n12399, new_n12401);
not_8  g12025(new_n12401, new_n12402);
or_8   g12026(new_n12402, new_n12398, new_n12403);
xor_4  g12027(new_n12395, new_n12391_1, new_n12404);
or_8   g12028(new_n12401, new_n12404, new_n12405);
and_8  g12029(new_n12405, new_n12403, new_n12406);
and_8  g12030(new_n11252, new_n11249, new_n12407);
and_8  g12031(new_n11258, new_n11253, new_n12408);
or_8   g12032(new_n12408, new_n12407, new_n12409);
xor_4  g12033(new_n12409, new_n12406, new_n12410);
not_8  g12034(new_n12410, new_n12411);
and_8  g12035(new_n11259, new_n11248, new_n12412);
not_8  g12036(new_n12412, new_n12413);
xor_4  g12037(new_n11259, new_n11247, new_n12414);
not_8  g12038(new_n11261, new_n12415);
or_8   g12039(new_n12415, new_n12414, new_n12416);
and_8  g12040(new_n12416, new_n12413, new_n12417);
or_8   g12041(new_n12417, new_n12411, new_n12418);
and_8  g12042(new_n11261, new_n11260, new_n12419);
or_8   g12043(new_n12419, new_n12412, new_n12420);
or_8   g12044(new_n12420, new_n12410, new_n12421);
and_8  g12045(new_n12421, new_n12418, new_n12422);
and_8  g12046(new_n12422, new_n12386, new_n12423);
not_8  g12047(new_n12386, new_n12424);
and_8  g12048(new_n12420, new_n12410, new_n12425);
and_8  g12049(new_n12417, new_n12411, new_n12426);
or_8   g12050(new_n12426, new_n12425, new_n12427);
and_8  g12051(new_n12427, new_n12424, new_n12428);
or_8   g12052(new_n12428, new_n12423, new_n12429);
xor_4  g12053(new_n12429, new_n12385, new_n12430);
and_8  g12054(new_n11294, new_n11293, new_n12431);
and_8  g12055(new_n11291, new_n11290, new_n12432);
or_8   g12056(new_n12432, new_n12431, new_n12433);
or_8   g12057(new_n12433, new_n11263, new_n12434);
and_8  g12058(new_n12434, new_n11292, new_n12435);
or_8   g12059(new_n12435, new_n12430, new_n12436);
and_8  g12060(new_n12429, new_n12385, new_n12437);
nor_6  g12061(new_n12429, new_n12385, new_n12438);
or_8   g12062(new_n12438, new_n12437, new_n12439);
and_8  g12063(new_n11296_1, new_n11302, new_n12440);
or_8   g12064(new_n12440, new_n12431, new_n12441);
or_8   g12065(new_n12441, new_n12439, new_n12442);
and_8  g12066(new_n12442, new_n12436, new_n12443);
xor_4  g12067(new_n12443, new_n12384, new_n12444_1);
and_8  g12068(new_n12348, new_n12346, new_n12445);
or_8   g12069(new_n12445, new_n12316, new_n12446);
and_8  g12070(new_n11298, new_n11299, new_n12447);
and_8  g12071(new_n12447, new_n12446, new_n12448);
and_8  g12072(new_n12353, new_n12351, new_n12449);
or_8   g12073(new_n12449, new_n12448, new_n12450);
or_8   g12074(new_n12450, new_n12444_1, new_n12451);
and_8  g12075(new_n12451, new_n12354, new_n12452);
or_8   g12076(new_n12452, new_n12345, new_n12453);
not_8  g12077(new_n12345, new_n12454);
and_8  g12078(new_n12383, new_n11289, new_n12455);
nor_6  g12079(new_n12383, new_n11289, new_n12456);
or_8   g12080(new_n12456, new_n12455, new_n12457);
xor_4  g12081(new_n12443, new_n12457, new_n12458);
or_8   g12082(new_n12447, new_n12446, new_n12459);
and_8  g12083(new_n12459, new_n12354, new_n12460);
and_8  g12084(new_n12460, new_n12458, new_n12461);
or_8   g12085(new_n12461, new_n12448, new_n12462);
or_8   g12086(new_n12462, new_n12454, new_n12463);
and_8  g12087(new_n12463, new_n12453, new_n12464);
nand_5 g12088(new_n12367, new_n12364, new_n12465);
or_8   g12089(new_n12373, new_n12369, new_n12466);
and_8  g12090(new_n12466, new_n12465, new_n12467);
and_8  g12091(n11153, n6441, new_n12468);
and_8  g12092(n12947, n5314, new_n12469);
and_8  g12093(n11999, n11222, new_n12470);
xnor_4 g12094(new_n12470, new_n12469, new_n12471);
xor_4  g12095(new_n12471, new_n12468, new_n12472);
xnor_4 g12096(new_n12472, new_n12467, new_n12473);
and_8  g12097(new_n12366, new_n12365, new_n12474);
and_8  g12098(n11791, n996, new_n12475);
xor_4  g12099(new_n12475, new_n12474, new_n12476);
nand_5 g12100(n5760, n5319, new_n12477);
and_8  g12101(n5767, n1478, new_n12478);
and_8  g12102(n10990, n9457, new_n12479);
xnor_4 g12103(new_n12479, new_n12478, new_n12480);
xor_4  g12104(new_n12480, new_n12477, new_n12481);
xor_4  g12105(new_n12481, new_n12476, new_n12482);
xor_4  g12106(new_n12482, new_n12473, new_n12483);
nand_5 g12107(new_n12362, new_n12359, new_n12484);
nand_5 g12108(new_n12361, new_n12360, new_n12485);
and_8  g12109(new_n12374, new_n12363, new_n12486);
xor_4  g12110(new_n12486, new_n12485, new_n12487);
and_8  g12111(new_n12487, new_n12484, new_n12488);
xor_4  g12112(new_n12488, new_n12483, new_n12489_1);
nor_6  g12113(new_n12489_1, new_n12377, new_n12490);
and_8  g12114(new_n12489_1, new_n12377, new_n12491);
or_8   g12115(new_n12491, new_n12490, new_n12492);
not_8  g12116(new_n12492, new_n12493);
not_8  g12117(new_n12380, new_n12494);
or_8   g12118(new_n12455, new_n12494, new_n12495);
xor_4  g12119(new_n12495, new_n12493, new_n12496);
and_8  g12120(new_n12390, new_n12387, new_n12497);
or_8   g12121(new_n12396, new_n12497, new_n12498);
not_8  g12122(new_n12498, new_n12499);
and_8  g12123(n12391, n447, new_n12500);
and_8  g12124(n11967, n7891, new_n12501);
and_8  g12125(n12069, n1353, new_n12502);
xnor_4 g12126(new_n12502, new_n12501, new_n12503);
xor_4  g12127(new_n12503, new_n12500, new_n12504);
xor_4  g12128(new_n12504, new_n12499, new_n12505);
and_8  g12129(new_n12389, new_n12388, new_n12506);
and_8  g12130(n7160, n6254, new_n12507);
xor_4  g12131(new_n12507, new_n12506, new_n12508);
nand_5 g12132(n7159, n2515, new_n12509);
not_8  g12133(new_n12509, new_n12510);
and_8  g12134(n12777, n4828, new_n12511_1);
and_8  g12135(n12489, n1199, new_n12512);
xor_4  g12136(new_n12512, new_n12511_1, new_n12513);
xor_4  g12137(new_n12513, new_n12510, new_n12514);
xor_4  g12138(new_n12514, new_n12508, new_n12515);
xor_4  g12139(new_n12515, new_n12505, new_n12516);
not_8  g12140(new_n12403, new_n12517);
and_8  g12141(new_n12400, new_n12399, new_n12518);
and_8  g12142(new_n12409, new_n12406, new_n12519);
xor_4  g12143(new_n12519, new_n12518, new_n12520);
or_8   g12144(new_n12520, new_n12517, new_n12521);
xor_4  g12145(new_n12521, new_n12516, new_n12522);
xor_4  g12146(new_n12522, new_n12425, new_n12523);
nor_6  g12147(new_n12438, new_n12428, new_n12524);
xor_4  g12148(new_n12524, new_n12523, new_n12525);
and_8  g12149(new_n12525, new_n12496, new_n12526);
nor_6  g12150(new_n12455, new_n12494, new_n12527);
and_8  g12151(new_n12527, new_n12492, new_n12528);
and_8  g12152(new_n12495, new_n12493, new_n12529);
or_8   g12153(new_n12529, new_n12528, new_n12530);
nor_6  g12154(new_n12524, new_n12523, new_n12531);
and_8  g12155(new_n12524, new_n12523, new_n12532);
or_8   g12156(new_n12532, new_n12531, new_n12533);
and_8  g12157(new_n12533, new_n12530, new_n12534);
or_8   g12158(new_n12534, new_n12526, new_n12535);
not_8  g12159(new_n12436, new_n12536);
and_8  g12160(new_n12443, new_n12384, new_n12537);
nor_6  g12161(new_n12537, new_n12536, new_n12538);
xor_4  g12162(new_n12538, new_n12535, new_n12539);
xor_4  g12163(new_n12539, new_n12464, new_n12540);
or_8   g12164(new_n12540, new_n12290, new_n12541);
not_8  g12165(new_n12290, new_n12542);
and_8  g12166(new_n12462, new_n12454, new_n12543);
and_8  g12167(new_n12452, new_n12345, new_n12544);
or_8   g12168(new_n12544, new_n12543, new_n12545);
xor_4  g12169(new_n12539, new_n12545, new_n12546);
or_8   g12170(new_n12546, new_n12542, new_n12547);
and_8  g12171(new_n12547, new_n12541, new_n12548);
xor_4  g12172(new_n12287, new_n12281, new_n12549);
nand_5 g12173(new_n11305, new_n11202, new_n12550);
not_8  g12174(new_n12550, new_n12551);
nor_6  g12175(new_n11310, new_n11306, new_n12552);
or_8   g12176(new_n12552, new_n12551, new_n12553);
or_8   g12177(new_n12553, new_n12549, new_n12554);
or_8   g12178(new_n11310, new_n11306, new_n12555);
and_8  g12179(new_n12555, new_n12550, new_n12556);
xor_4  g12180(new_n12556, new_n12549, new_n12557);
xor_4  g12181(new_n12460, new_n12458, new_n12558);
not_8  g12182(new_n12558, new_n12559);
or_8   g12183(new_n12559, new_n12557, new_n12560);
and_8  g12184(new_n12560, new_n12554, new_n12561);
xor_4  g12185(new_n12561, new_n12548, n5132);
xor_4  g12186(new_n11959, new_n11353, n5191);
or_8   g12187(new_n3802, new_n3373, new_n12564);
or_8   g12188(new_n3947, new_n3942, new_n12565);
or_8   g12189(new_n12565, new_n3804, new_n12566);
and_8  g12190(new_n12566, new_n12564, new_n12567);
or_8   g12191(new_n3942, new_n3944, new_n12568);
or_8   g12192(new_n3345, new_n3319, new_n12569);
or_8   g12193(new_n3372, new_n3349, new_n12570);
and_8  g12194(new_n12570, new_n12569, new_n12571);
not_8  g12195(new_n3341, new_n12572);
nand_5 g12196(new_n3342_1, new_n12572, new_n12573);
or_8   g12197(new_n3344, new_n3338, new_n12574);
and_8  g12198(new_n12574, new_n12573, new_n12575);
and_8  g12199(n11478, n10965, new_n12576);
nand_5 g12200(new_n3816, new_n3815, new_n12577);
or_8   g12201(new_n3822, new_n3817, new_n12578);
and_8  g12202(new_n12578, new_n12577, new_n12579);
and_8  g12203(n8433, n4722, new_n12580);
and_8  g12204(n8065, n2464, new_n12581);
and_8  g12205(n7646, n405, new_n12582);
xor_4  g12206(new_n12582, new_n12581, new_n12583);
xor_4  g12207(new_n12583, new_n12580, new_n12584);
xor_4  g12208(new_n12584, new_n12579, new_n12585);
xor_4  g12209(new_n12585, new_n12576, new_n12586);
xor_4  g12210(new_n12586, new_n12575, new_n12587);
not_8  g12211(new_n3887, new_n12588);
and_8  g12212(new_n12588, new_n3885, new_n12589);
or_8   g12213(new_n3898, new_n12589, new_n12590);
and_8  g12214(new_n3851, new_n3850, new_n12591_1);
nor_6  g12215(new_n3857, new_n3852, new_n12592);
or_8   g12216(new_n12592, new_n12591_1, new_n12593);
nand_5 g12217(new_n3890, new_n3889, new_n12594);
or_8   g12218(new_n3896, new_n3891, new_n12595);
and_8  g12219(new_n12595, new_n12594, new_n12596);
xor_4  g12220(new_n12596, new_n12593, new_n12597);
and_8  g12221(n8384, n6359, new_n12598);
and_8  g12222(n7546, n4805, new_n12599);
xor_4  g12223(new_n12599, new_n12598, new_n12600);
and_8  g12224(n12925, n4938, new_n12601);
and_8  g12225(n11536, n7862, new_n12602);
xor_4  g12226(new_n12602, new_n12601, new_n12603);
and_8  g12227(new_n3894, new_n3893, new_n12604);
or_8   g12228(new_n3894, new_n3893, new_n12605);
and_8  g12229(new_n12605, new_n3892, new_n12606);
or_8   g12230(new_n12606, new_n12604, new_n12607);
xor_4  g12231(new_n12607, new_n12603, new_n12608);
xnor_4 g12232(new_n12608, new_n12600, new_n12609);
xor_4  g12233(new_n12609, new_n12597, new_n12610);
nor_6  g12234(new_n12610, new_n12590, new_n12611);
and_8  g12235(new_n12610, new_n12590, new_n12612);
or_8   g12236(new_n12612, new_n12611, new_n12613);
not_8  g12237(new_n3845, new_n12614);
or_8   g12238(new_n3848, new_n12614, new_n12615);
or_8   g12239(new_n3858, new_n3849_1, new_n12616);
and_8  g12240(new_n12616, new_n12615, new_n12617);
or_8   g12241(new_n3883, new_n3882, new_n12618);
or_8   g12242(new_n3884, new_n3881, new_n12619);
and_8  g12243(new_n12619, new_n12618, new_n12620);
and_8  g12244(n9956, n6826, new_n12621);
and_8  g12245(n6797, n4826, new_n12622);
xor_4  g12246(new_n12622, new_n12621, new_n12623);
and_8  g12247(n7610, n6294, new_n12624);
and_8  g12248(n6611, n6358, new_n12625);
xor_4  g12249(new_n12625, new_n12624, new_n12626);
xor_4  g12250(new_n12626, new_n12623, new_n12627);
xor_4  g12251(new_n12627, new_n12620, new_n12628);
nand_5 g12252(n7733, n3146, new_n12629);
or_8   g12253(new_n3843, new_n3842_1, new_n12630);
or_8   g12254(new_n3844, new_n3841, new_n12631);
and_8  g12255(new_n12631, new_n12630, new_n12632);
xor_4  g12256(new_n12632, new_n12629, new_n12633);
xor_4  g12257(new_n12633, new_n12628, new_n12634);
and_8  g12258(n5198, n217, new_n12635);
and_8  g12259(n5283, n503, new_n12636);
xor_4  g12260(new_n12636, new_n12635, new_n12637);
and_8  g12261(n4970, n137, new_n12638);
and_8  g12262(n11296, n3992, new_n12639);
xnor_4 g12263(new_n12639, new_n12638, new_n12640);
xor_4  g12264(new_n12640, new_n12637, new_n12641);
and_8  g12265(new_n3855, new_n3854, new_n12642);
or_8   g12266(new_n3855, new_n3854, new_n12643);
and_8  g12267(new_n12643, new_n3853, new_n12644);
or_8   g12268(new_n12644, new_n12642, new_n12645);
and_8  g12269(n11311, n10439, new_n12646);
and_8  g12270(n6126, n4203, new_n12647);
xor_4  g12271(new_n12647, new_n12646, new_n12648_1);
xor_4  g12272(new_n12648_1, new_n12645, new_n12649);
xor_4  g12273(new_n12649, new_n12641, new_n12650);
xor_4  g12274(new_n12650, new_n12634, new_n12651);
xor_4  g12275(new_n12651, new_n12617, new_n12652);
not_8  g12276(new_n12652, new_n12653);
and_8  g12277(new_n12653, new_n12613, new_n12654);
xor_4  g12278(new_n12610, new_n12590, new_n12655);
and_8  g12279(new_n12652, new_n12655, new_n12656);
or_8   g12280(new_n12656, new_n12654, new_n12657);
and_8  g12281(new_n3444, new_n3827, new_n12658);
and_8  g12282(new_n3829, new_n3833, new_n12659);
or_8   g12283(new_n12659, new_n12658, new_n12660);
and_8  g12284(new_n3720, new_n3861, new_n12661);
or_8   g12285(new_n3870, new_n12661, new_n12662);
or_8   g12286(new_n12662, new_n12660, new_n12663);
nor_6  g12287(new_n12659, new_n12658, new_n12664);
nor_6  g12288(new_n3870, new_n12661, new_n12665);
or_8   g12289(new_n12665, new_n12664, new_n12666);
and_8  g12290(new_n12666, new_n12663, new_n12667);
and_8  g12291(new_n12667, new_n12657, new_n12668);
nor_6  g12292(new_n12667, new_n12657, new_n12669);
or_8   g12293(new_n12669, new_n12668, new_n12670);
or_8   g12294(new_n12670, new_n12587, new_n12671);
not_8  g12295(new_n12586, new_n12672);
xor_4  g12296(new_n12672, new_n12575, new_n12673);
xor_4  g12297(new_n12667, new_n12657, new_n12674);
or_8   g12298(new_n12674, new_n12673, new_n12675);
and_8  g12299(new_n12675, new_n12671, new_n12676);
and_8  g12300(new_n12676, new_n12571, new_n12677);
or_8   g12301(new_n3347, new_n3318, new_n12678);
and_8  g12302(new_n12569, new_n12678, new_n12679);
and_8  g12303(new_n3375, new_n3365, new_n12680);
or_8   g12304(new_n12680, new_n3368, new_n12681);
and_8  g12305(new_n12681, new_n12679, new_n12682);
or_8   g12306(new_n12682, new_n3348, new_n12683);
and_8  g12307(new_n12674, new_n12673, new_n12684);
and_8  g12308(new_n12670, new_n12587, new_n12685);
or_8   g12309(new_n12685, new_n12684, new_n12686);
and_8  g12310(new_n12686, new_n12683, new_n12687);
or_8   g12311(new_n12687, new_n12677, new_n12688);
nor_6  g12312(new_n3835, new_n3831, new_n12689);
nor_6  g12313(new_n3456_1, new_n3837, new_n12690);
and_8  g12314(new_n12690, new_n12689, new_n12691);
or_8   g12315(new_n12691, new_n3835, new_n12692);
and_8  g12316(new_n3813, new_n3810, new_n12693);
and_8  g12317(new_n3824, new_n3814, new_n12694);
or_8   g12318(new_n12694, new_n12693, new_n12695);
and_8  g12319(n4086, n1471, new_n12696);
not_8  g12320(new_n12696, new_n12697);
and_8  g12321(n10391, n9400, new_n12698);
or_8   g12322(new_n3809, new_n3806, new_n12699);
and_8  g12323(new_n12699, new_n3807, new_n12700);
and_8  g12324(new_n12700, new_n12698, new_n12701);
and_8  g12325(new_n12698, new_n3425, new_n12702);
nor_6  g12326(new_n12702, new_n12700, new_n12703);
nor_6  g12327(new_n12703, new_n12701, new_n12704_1);
nand_5 g12328(n11757, n2577, new_n12705_1);
and_8  g12329(n9637, n3172, new_n12706_1);
and_8  g12330(n5240, n3842, new_n12707);
xor_4  g12331(new_n12707, new_n12706_1, new_n12708);
xor_4  g12332(new_n12708, new_n12705_1, new_n12709_1);
and_8  g12333(new_n3325, new_n3324, new_n12710);
or_8   g12334(new_n3325, new_n3324, new_n12711);
and_8  g12335(new_n12711, new_n3323, new_n12712);
or_8   g12336(new_n12712, new_n12710, new_n12713);
xor_4  g12337(new_n12713, new_n12709_1, new_n12714);
xor_4  g12338(new_n12714, new_n12704_1, new_n12715);
xor_4  g12339(new_n12715, new_n12697, new_n12716);
and_8  g12340(n7236, n1357, new_n12717);
nand_5 g12341(new_n3330, new_n3329, new_n12718);
or_8   g12342(new_n3336, new_n3331, new_n12719);
and_8  g12343(new_n12719, new_n12718, new_n12720_1);
xor_4  g12344(new_n12720_1, new_n12717, new_n12721);
not_8  g12345(new_n12721, new_n12722);
and_8  g12346(new_n12722, new_n12716, new_n12723);
xor_4  g12347(new_n12715, new_n12696, new_n12724);
and_8  g12348(new_n12721, new_n12724, new_n12725);
or_8   g12349(new_n12725, new_n12723, new_n12726);
xor_4  g12350(new_n12726, new_n12695, new_n12727);
and_8  g12351(n1835, n1333, new_n12728);
and_8  g12352(n11917, n11821, new_n12729);
xnor_4 g12353(new_n12729, new_n12728, new_n12730);
and_8  g12354(n12753, n3602, new_n12731);
and_8  g12355(n8595, n4187, new_n12732);
xor_4  g12356(new_n12732, new_n12731, new_n12733);
and_8  g12357(n6877, n4190, new_n12734);
and_8  g12358(n10174, n3719, new_n12735);
xor_4  g12359(new_n12735, new_n12734, new_n12736);
xor_4  g12360(new_n12736, new_n12733, new_n12737);
xor_4  g12361(new_n12737, new_n12730, new_n12738);
or_8   g12362(new_n3820, new_n3819, new_n12739);
or_8   g12363(new_n3821, new_n3818, new_n12740);
and_8  g12364(new_n12740, new_n12739, new_n12741);
and_8  g12365(n9080, n4921, new_n12742);
xor_4  g12366(new_n12742, new_n12741, new_n12743);
xor_4  g12367(new_n12743, new_n12738, new_n12744);
and_8  g12368(new_n3327, new_n3322, new_n12745);
and_8  g12369(new_n3337, new_n3328, new_n12746);
or_8   g12370(new_n12746, new_n12745, new_n12747);
xor_4  g12371(new_n12747, new_n12744, new_n12748);
not_8  g12372(new_n12748, new_n12749);
and_8  g12373(new_n12749, new_n12727, new_n12750);
not_8  g12374(new_n12695, new_n12751);
xor_4  g12375(new_n12726, new_n12751, new_n12752);
and_8  g12376(new_n12748, new_n12752, new_n12753_1);
or_8   g12377(new_n12753_1, new_n12750, new_n12754);
and_8  g12378(new_n3913, new_n3900, new_n12755);
or_8   g12379(new_n12755, new_n3905, new_n12756);
not_8  g12380(new_n12756, new_n12757);
and_8  g12381(new_n12757, new_n12754, new_n12758);
nor_6  g12382(new_n12753_1, new_n12750, new_n12759);
and_8  g12383(new_n12756, new_n12759, new_n12760);
or_8   g12384(new_n12760, new_n12758, new_n12761);
and_8  g12385(new_n12761, new_n12692, new_n12762);
not_8  g12386(new_n3835, new_n12763);
or_8   g12387(new_n3838, new_n3836, new_n12764);
and_8  g12388(new_n12764, new_n12763, new_n12765);
or_8   g12389(new_n12756, new_n12759, new_n12766);
or_8   g12390(new_n12757, new_n12754, new_n12767);
and_8  g12391(new_n12767, new_n12766, new_n12768);
and_8  g12392(new_n12768, new_n12765, new_n12769);
or_8   g12393(new_n12769, new_n12762, new_n12770);
not_8  g12394(new_n3873, new_n12771);
or_8   g12395(new_n3879, new_n12771, new_n12772);
or_8   g12396(new_n12772, new_n12770, new_n12773);
or_8   g12397(new_n12768, new_n12765, new_n12774);
or_8   g12398(new_n12761, new_n12692, new_n12775);
and_8  g12399(new_n12775, new_n12774, new_n12776);
nor_6  g12400(new_n3879, new_n12771, new_n12777_1);
or_8   g12401(new_n12777_1, new_n12776, new_n12778);
and_8  g12402(new_n12778, new_n12773, new_n12779);
xor_4  g12403(new_n12779, new_n12688, new_n12780);
and_8  g12404(new_n3927, new_n3924, new_n12781);
or_8   g12405(new_n3933, new_n12781, new_n12782);
nand_5 g12406(new_n3915, new_n3697, new_n12783);
and_8  g12407(new_n3926, new_n12783, new_n12784);
or_8   g12408(new_n3334, new_n3333, new_n12785);
or_8   g12409(new_n3335, new_n3332, new_n12786);
nand_5 g12410(new_n12786, new_n12785, new_n12787);
xor_4  g12411(new_n12787, new_n12784, new_n12788);
xor_4  g12412(new_n12788, new_n12782, new_n12789);
or_8   g12413(new_n12789, new_n12780, new_n12790);
nor_6  g12414(new_n12779, new_n12688, new_n12791);
and_8  g12415(new_n12779, new_n12688, new_n12792);
or_8   g12416(new_n12792, new_n12791, new_n12793);
nor_6  g12417(new_n12788, new_n12782, new_n12794);
and_8  g12418(new_n12788, new_n12782, new_n12795);
or_8   g12419(new_n12795, new_n12794, new_n12796);
or_8   g12420(new_n12796, new_n12793, new_n12797);
and_8  g12421(new_n12797, new_n12790, new_n12798);
and_8  g12422(new_n12798, new_n12568, new_n12799);
or_8   g12423(new_n3946, new_n3945, new_n12800);
and_8  g12424(new_n12800, new_n3938, new_n12801);
and_8  g12425(new_n12796, new_n12793, new_n12802);
and_8  g12426(new_n12789, new_n12780, new_n12803);
or_8   g12427(new_n12803, new_n12802, new_n12804);
and_8  g12428(new_n12804, new_n12801, new_n12805);
or_8   g12429(new_n12805, new_n12799, new_n12806);
xor_4  g12430(new_n12806, new_n12567, n5257);
xnor_4 g12431(new_n11966, new_n11958, n5411);
xnor_4 g12432(new_n3790, new_n3782, n5435);
xor_4  g12433(new_n6411, new_n6406, n5641);
xnor_4 g12434(new_n9118, new_n9102, n5670);
xor_4  g12435(new_n5180, new_n5391, n5693);
xnor_4 g12436(new_n1349, new_n1338, n5934);
xnor_4 g12437(new_n11971, new_n11968, n6089);
and_8  g12438(new_n8290, new_n8287, new_n12815);
nand_5 g12439(new_n8267, new_n8264, new_n12816);
or_8   g12440(new_n8272, new_n8280, new_n12817);
and_8  g12441(new_n12817, new_n12816, new_n12818);
and_8  g12442(n2564, n2253, new_n12819);
and_8  g12443(n9195, n4189, new_n12820);
and_8  g12444(n6687, n3865, new_n12821);
xnor_4 g12445(new_n12821, new_n12820, new_n12822);
xor_4  g12446(new_n12822, new_n12819, new_n12823);
xor_4  g12447(new_n12823, new_n12818, new_n12824);
and_8  g12448(new_n8266, new_n8265, new_n12825);
and_8  g12449(n6770, n4634, new_n12826_1);
xor_4  g12450(new_n12826_1, new_n12825, new_n12827);
and_8  g12451(n3627, n2879, new_n12828);
and_8  g12452(n10223, n9920, new_n12829);
and_8  g12453(n7265, n4516, new_n12830);
xnor_4 g12454(new_n12830, new_n12829, new_n12831);
xor_4  g12455(new_n12831, new_n12828, new_n12832);
xor_4  g12456(new_n12832, new_n12827, new_n12833);
xor_4  g12457(new_n12833, new_n12824, new_n12834);
not_8  g12458(new_n12834, new_n12835);
not_8  g12459(new_n8278, new_n12836);
and_8  g12460(new_n8275, new_n8274, new_n12837);
and_8  g12461(new_n8286, new_n8283, new_n12838);
xor_4  g12462(new_n12838, new_n12837, new_n12839);
or_8   g12463(new_n12839, new_n12836, new_n12840);
xor_4  g12464(new_n12840, new_n12835, new_n12841);
xor_4  g12465(new_n12841, new_n12815, new_n12842);
not_8  g12466(new_n12842, new_n12843);
nor_6  g12467(new_n8291, new_n8263, new_n12844);
and_8  g12468(new_n8292, new_n8262, new_n12845);
or_8   g12469(new_n12845, new_n12844, new_n12846);
xor_4  g12470(new_n12846, new_n12843, new_n12847);
not_8  g12471(new_n8342, new_n12848);
and_8  g12472(new_n6196, new_n6186, new_n12849);
or_8   g12473(new_n12849, new_n12848, new_n12850);
xor_4  g12474(new_n8343, new_n12848, new_n12851);
not_8  g12475(new_n8441, new_n12852);
xor_4  g12476(new_n12852, new_n8440, new_n12853);
or_8   g12477(new_n12853, new_n12851, new_n12854);
and_8  g12478(new_n12854, new_n12850, new_n12855);
and_8  g12479(new_n8340, new_n8300, new_n12856);
and_8  g12480(new_n8341, new_n8298, new_n12857);
or_8   g12481(new_n12857, new_n12856, new_n12858);
nor_6  g12482(new_n8312, new_n8305, new_n12859);
and_8  g12483(n12221, n10928, new_n12860);
and_8  g12484(n12145, n6986, new_n12861);
and_8  g12485(n10217, n8336, new_n12862);
xnor_4 g12486(new_n12862, new_n12861, new_n12863);
xor_4  g12487(new_n12863, new_n12860, new_n12864);
xor_4  g12488(new_n12864, new_n12859, new_n12865);
and_8  g12489(new_n8303_1, new_n8302, new_n12866);
and_8  g12490(n2522, n2226, new_n12867);
xor_4  g12491(new_n12867, new_n12866, new_n12868);
nand_5 g12492(n10678, n2024, new_n12869);
not_8  g12493(new_n12869, new_n12870);
and_8  g12494(n9189, n1094, new_n12871);
and_8  g12495(n7946, n7320, new_n12872);
xnor_4 g12496(new_n12872, new_n12871, new_n12873);
xor_4  g12497(new_n12873, new_n12870, new_n12874);
xor_4  g12498(new_n12874, new_n12868, new_n12875);
xor_4  g12499(new_n12875, new_n12865, new_n12876);
nand_5 g12500(new_n8316, new_n8315, new_n12877);
xor_4  g12501(new_n8325, new_n12877, new_n12878);
and_8  g12502(new_n12878, new_n8319, new_n12879);
or_8   g12503(new_n12879, new_n12876, new_n12880);
not_8  g12504(new_n12880, new_n12881);
and_8  g12505(new_n12879, new_n12876, new_n12882);
or_8   g12506(new_n12882, new_n12881, new_n12883);
or_8   g12507(new_n12883, new_n8334, new_n12884);
not_8  g12508(new_n8334, new_n12885);
xor_4  g12509(new_n12879, new_n12876, new_n12886);
or_8   g12510(new_n12886, new_n12885, new_n12887);
and_8  g12511(new_n12887, new_n12884, new_n12888);
xor_4  g12512(new_n12888, new_n12858, new_n12889);
not_8  g12513(new_n8380, new_n12890);
and_8  g12514(new_n8357, new_n8356, new_n12891);
and_8  g12515(n7160, n521, new_n12892);
xnor_4 g12516(new_n12892, new_n12891, new_n12893);
and_8  g12517(n2515, n2498, new_n12894);
and_8  g12518(n2558, n1199, new_n12895);
and_8  g12519(n5579, n4828, new_n12896);
nor_6  g12520(new_n12896, new_n12895, new_n12897);
and_8  g12521(new_n12896, new_n12895, new_n12898);
or_8   g12522(new_n12898, new_n12897, new_n12899);
xor_4  g12523(new_n12899, new_n12894, new_n12900);
xnor_4 g12524(new_n12900, new_n12893, new_n12901);
nand_5 g12525(new_n8353, new_n8349, new_n12902);
or_8   g12526(new_n8358, new_n8355, new_n12903);
and_8  g12527(new_n12903, new_n12902, new_n12904);
and_8  g12528(n12391, n5798, new_n12905);
and_8  g12529(n7891, n6016, new_n12906);
and_8  g12530(n12069, n2347, new_n12907);
xnor_4 g12531(new_n12907, new_n12906, new_n12908);
xor_4  g12532(new_n12908, new_n12905, new_n12909);
xor_4  g12533(new_n12909, new_n12904, new_n12910);
xor_4  g12534(new_n12910, new_n12901, new_n12911);
not_8  g12535(new_n8363, new_n12912);
and_8  g12536(new_n8361, new_n8360, new_n12913);
not_8  g12537(new_n12913, new_n12914);
nor_6  g12538(new_n8370, new_n12914, new_n12915);
and_8  g12539(new_n8370, new_n12914, new_n12916);
or_8   g12540(new_n12916, new_n12915, new_n12917);
and_8  g12541(new_n12917, new_n12912, new_n12918);
nor_6  g12542(new_n12918, new_n12911, new_n12919);
and_8  g12543(new_n12918, new_n12911, new_n12920);
or_8   g12544(new_n12920, new_n12919, new_n12921);
or_8   g12545(new_n12921, new_n12890, new_n12922);
xor_4  g12546(new_n12918, new_n12911, new_n12923);
or_8   g12547(new_n12923, new_n8380, new_n12924);
and_8  g12548(new_n12924, new_n12922, new_n12925_1);
or_8   g12549(new_n8433_1, new_n8378, new_n12926);
and_8  g12550(new_n12926, new_n12925_1, new_n12927);
and_8  g12551(new_n12923, new_n8380, new_n12928);
and_8  g12552(new_n12921, new_n12890, new_n12929);
or_8   g12553(new_n12929, new_n12928, new_n12930);
and_8  g12554(new_n8385, new_n8386, new_n12931);
and_8  g12555(new_n12931, new_n12930, new_n12932);
or_8   g12556(new_n12932, new_n12927, new_n12933);
and_8  g12557(new_n8396, new_n8393, new_n12934);
or_8   g12558(new_n8402, new_n12934, new_n12935);
and_8  g12559(n11153, n5153, new_n12936);
and_8  g12560(n7270, n5314, new_n12937);
and_8  g12561(n11222, n2507, new_n12938);
xnor_4 g12562(new_n12938, new_n12937, new_n12939);
xor_4  g12563(new_n12939, new_n12936, new_n12940);
xor_4  g12564(new_n12940, new_n12935, new_n12941);
and_8  g12565(new_n8395, new_n8394, new_n12942);
and_8  g12566(n996, n806, new_n12943);
xnor_4 g12567(new_n12943, new_n12942, new_n12944);
and_8  g12568(n9111, n5319, new_n12945);
and_8  g12569(n5767, n3342, new_n12946);
and_8  g12570(n9763, n9457, new_n12947_1);
xnor_4 g12571(new_n12947_1, new_n12946, new_n12948);
xor_4  g12572(new_n12948, new_n12945, new_n12949);
xor_4  g12573(new_n12949, new_n12944, new_n12950);
xor_4  g12574(new_n12950, new_n12941, new_n12951);
nor_6  g12575(new_n8408, new_n8404, new_n12952);
and_8  g12576(new_n8406, new_n8405, new_n12953);
xor_4  g12577(new_n8413, new_n12953, new_n12954);
or_8   g12578(new_n12954, new_n12952, new_n12955);
xor_4  g12579(new_n12955, new_n12951, new_n12956);
or_8   g12580(new_n12956, new_n8418, new_n12957);
not_8  g12581(new_n8418, new_n12958);
not_8  g12582(new_n12951, new_n12959);
xor_4  g12583(new_n12955, new_n12959, new_n12960);
or_8   g12584(new_n12960, new_n12958, new_n12961);
and_8  g12585(new_n12961, new_n12957, new_n12962);
and_8  g12586(new_n8437, new_n8424, new_n12963);
and_8  g12587(new_n12963, new_n12962, new_n12964);
and_8  g12588(new_n12960, new_n12958, new_n12965);
and_8  g12589(new_n12956, new_n8418, new_n12966);
or_8   g12590(new_n12966, new_n12965, new_n12967);
or_8   g12591(new_n8430, new_n8425, new_n12968);
and_8  g12592(new_n12968, new_n12967, new_n12969);
or_8   g12593(new_n12969, new_n12964, new_n12970);
and_8  g12594(new_n12970, new_n12933, new_n12971);
or_8   g12595(new_n12931, new_n12930, new_n12972);
or_8   g12596(new_n12926, new_n12925_1, new_n12973);
and_8  g12597(new_n12973, new_n12972, new_n12974);
or_8   g12598(new_n12968, new_n12967, new_n12975);
or_8   g12599(new_n12963, new_n12962, new_n12976);
and_8  g12600(new_n12976, new_n12975, new_n12977);
and_8  g12601(new_n12977, new_n12974, new_n12978);
or_8   g12602(new_n12978, new_n12971, new_n12979);
or_8   g12603(new_n8438, new_n8435, new_n12980);
or_8   g12604(new_n8441, new_n8440, new_n12981);
and_8  g12605(new_n12981, new_n12980, new_n12982);
xor_4  g12606(new_n12982, new_n12979, new_n12983);
or_8   g12607(new_n12983, new_n12889, new_n12984);
not_8  g12608(new_n12889, new_n12985);
or_8   g12609(new_n12977, new_n12974, new_n12986);
or_8   g12610(new_n12970, new_n12933, new_n12987);
and_8  g12611(new_n12987, new_n12986, new_n12988);
xor_4  g12612(new_n12982, new_n12988, new_n12989);
or_8   g12613(new_n12989, new_n12985, new_n12990);
and_8  g12614(new_n12990, new_n12984, new_n12991);
and_8  g12615(new_n12991, new_n12855, new_n12992);
and_8  g12616(new_n8343, new_n8342, new_n12993);
and_8  g12617(new_n8442, new_n8344, new_n12994);
or_8   g12618(new_n12994, new_n12993, new_n12995);
and_8  g12619(new_n12989, new_n12985, new_n12996);
and_8  g12620(new_n12983, new_n12889, new_n12997);
or_8   g12621(new_n12997, new_n12996, new_n12998);
and_8  g12622(new_n12998, new_n12995, new_n12999);
or_8   g12623(new_n12999, new_n12992, new_n13000);
or_8   g12624(new_n13000, new_n12847, new_n13001);
and_8  g12625(new_n8296, new_n8293, new_n13002);
and_8  g12626(new_n8443, new_n8297, new_n13003);
or_8   g12627(new_n13003, new_n13002, new_n13004);
not_8  g12628(new_n12847, new_n13005);
or_8   g12629(new_n12998, new_n12995, new_n13006);
or_8   g12630(new_n12991, new_n12855, new_n13007);
and_8  g12631(new_n13007, new_n13006, new_n13008);
and_8  g12632(new_n13008, new_n13005, new_n13009);
and_8  g12633(new_n13000, new_n12847, new_n13010);
or_8   g12634(new_n13010, new_n13009, new_n13011);
or_8   g12635(new_n13011, new_n13004, new_n13012);
and_8  g12636(new_n13012, new_n13001, new_n13013);
or_8   g12637(new_n12992, new_n12996, new_n13014);
and_8  g12638(new_n12982, new_n12988, new_n13015);
nor_6  g12639(new_n13015, new_n12971, new_n13016);
not_8  g12640(new_n12877, new_n13017);
nand_5 g12641(new_n8325, new_n13017, new_n13018);
and_8  g12642(new_n12880, new_n13018, new_n13019);
and_8  g12643(new_n12823, new_n12818, new_n13020);
and_8  g12644(new_n12833, new_n12824, new_n13021);
or_8   g12645(new_n13021, new_n13020, new_n13022);
nand_5 g12646(n2522, n1094, new_n13023);
or_8   g12647(new_n12938, new_n12937, new_n13024);
or_8   g12648(new_n12939, new_n12936, new_n13025);
and_8  g12649(new_n13025, new_n13024, new_n13026);
xor_4  g12650(new_n13026, new_n13023, new_n13027);
xor_4  g12651(new_n13027, new_n13022, new_n13028);
and_8  g12652(new_n13028, new_n13019, new_n13029);
nor_6  g12653(new_n13028, new_n13019, new_n13030);
or_8   g12654(new_n13030, new_n13029, new_n13031);
and_8  g12655(new_n12864, new_n12859, new_n13032);
and_8  g12656(new_n12875, new_n12865, new_n13033);
or_8   g12657(new_n13033, new_n13032, new_n13034);
and_8  g12658(n10678, n9189, new_n13035);
xor_4  g12659(new_n13035, new_n13034, new_n13036);
or_8   g12660(new_n12872, new_n12871, new_n13037);
or_8   g12661(new_n12873, new_n12870, new_n13038);
and_8  g12662(new_n13038, new_n13037, new_n13039);
and_8  g12663(n7946, n7523, new_n13040);
and_8  g12664(n10223, n3627, new_n13041);
and_8  g12665(n3865, n2564, new_n13042);
xor_4  g12666(new_n13042, new_n13041, new_n13043);
xor_4  g12667(new_n13043, new_n13040, new_n13044);
xor_4  g12668(new_n13044, new_n13039, new_n13045);
and_8  g12669(n12221, n6986, new_n13046);
and_8  g12670(n8336, n7823, new_n13047);
xor_4  g12671(new_n13047, new_n13046, new_n13048);
xor_4  g12672(new_n13048, new_n13045, new_n13049);
nor_6  g12673(new_n12830, new_n12829, new_n13050);
nor_6  g12674(new_n12831, new_n12828, new_n13051);
or_8   g12675(new_n13051, new_n13050, new_n13052);
or_8   g12676(new_n12867, new_n12866, new_n13053);
not_8  g12677(new_n13053, new_n13054);
and_8  g12678(new_n12874, new_n12868, new_n13055);
or_8   g12679(new_n13055, new_n13054, new_n13056);
or_8   g12680(new_n13056, new_n13052, new_n13057);
not_8  g12681(new_n13052, new_n13058);
not_8  g12682(new_n12868, new_n13059);
xor_4  g12683(new_n12873, new_n12869, new_n13060);
or_8   g12684(new_n13060, new_n13059, new_n13061);
and_8  g12685(new_n13061, new_n13053, new_n13062);
or_8   g12686(new_n13062, new_n13058, new_n13063);
and_8  g12687(new_n13063, new_n13057, new_n13064);
or_8   g12688(new_n12907, new_n12906, new_n13065);
or_8   g12689(new_n12908, new_n12905, new_n13066);
and_8  g12690(new_n13066, new_n13065, new_n13067);
nand_5 g12691(n6687, n2512, new_n13068);
or_8   g12692(new_n12896, new_n12895, new_n13069);
and_8  g12693(new_n13069, new_n12894, new_n13070);
or_8   g12694(new_n13070, new_n12898, new_n13071);
xor_4  g12695(new_n13071, new_n13068, new_n13072);
xor_4  g12696(new_n13072, new_n13067, new_n13073);
not_8  g12697(new_n13073, new_n13074);
xor_4  g12698(new_n13074, new_n13064, new_n13075);
and_8  g12699(new_n13075, new_n13049, new_n13076);
not_8  g12700(new_n13049, new_n13077);
xor_4  g12701(new_n13073, new_n13064, new_n13078);
and_8  g12702(new_n13078, new_n13077, new_n13079);
or_8   g12703(new_n13079, new_n13076, new_n13080);
and_8  g12704(n11153, n2507, new_n13081);
and_8  g12705(n7270, n996, new_n13082);
xor_4  g12706(new_n13082, new_n13081, new_n13083);
and_8  g12707(n7160, n6016, new_n13084);
and_8  g12708(n5767, n806, new_n13085);
xor_4  g12709(new_n13085, new_n13084, new_n13086);
xnor_4 g12710(new_n13086, new_n13083, new_n13087);
and_8  g12711(n4828, n521, new_n13088);
and_8  g12712(n5579, n2515, new_n13089);
xor_4  g12713(new_n13089, new_n13088, new_n13090);
and_8  g12714(n12069, n1576, new_n13091);
and_8  g12715(n5314, n5153, new_n13092);
xnor_4 g12716(new_n13092, new_n13091, new_n13093);
xor_4  g12717(new_n13093, new_n13090, new_n13094);
xor_4  g12718(new_n13094, new_n13087, new_n13095);
and_8  g12719(new_n12821, new_n12820, new_n13096);
or_8   g12720(new_n12821, new_n12820, new_n13097);
and_8  g12721(new_n13097, new_n12819, new_n13098);
or_8   g12722(new_n13098, new_n13096, new_n13099);
not_8  g12723(n2879, new_n13100);
not_8  g12724(n4516, new_n13101);
or_8   g12725(new_n13101, new_n13100, new_n13102);
and_8  g12726(n4189, n2253, new_n13103);
and_8  g12727(n9920, n4634, new_n13104);
xor_4  g12728(new_n13104, new_n13103, new_n13105);
xor_4  g12729(new_n13105, new_n13102, new_n13106);
xor_4  g12730(new_n13106, new_n13099, new_n13107);
not_8  g12731(new_n13107, new_n13108);
xor_4  g12732(new_n13108, new_n13095, new_n13109);
nor_6  g12733(new_n12826_1, new_n12825, new_n13110);
and_8  g12734(new_n12832, new_n12827, new_n13111);
or_8   g12735(new_n13111, new_n13110, new_n13112);
and_8  g12736(new_n12943, new_n12942, new_n13113);
nor_6  g12737(new_n12949, new_n12944, new_n13114);
or_8   g12738(new_n13114, new_n13113, new_n13115);
xor_4  g12739(new_n13115, new_n13112, new_n13116);
and_8  g12740(new_n13116, new_n13109, new_n13117);
xor_4  g12741(new_n13107, new_n13095, new_n13118);
nor_6  g12742(new_n13111, new_n13110, new_n13119);
xor_4  g12743(new_n13115, new_n13119, new_n13120);
and_8  g12744(new_n13120, new_n13118, new_n13121);
or_8   g12745(new_n13121, new_n13117, new_n13122);
or_8   g12746(new_n13122, new_n13080, new_n13123);
or_8   g12747(new_n13078, new_n13077, new_n13124);
or_8   g12748(new_n13075, new_n13049, new_n13125);
and_8  g12749(new_n13125, new_n13124, new_n13126);
nor_6  g12750(new_n13121, new_n13117, new_n13127);
or_8   g12751(new_n13127, new_n13126, new_n13128);
and_8  g12752(new_n13128, new_n13123, new_n13129);
or_8   g12753(new_n13129, new_n13036, new_n13130);
not_8  g12754(new_n13036, new_n13131);
and_8  g12755(new_n13127, new_n13126, new_n13132);
and_8  g12756(new_n13122, new_n13080, new_n13133);
or_8   g12757(new_n13133, new_n13132, new_n13134);
or_8   g12758(new_n13134, new_n13131, new_n13135);
and_8  g12759(new_n13135, new_n13130, new_n13136);
xor_4  g12760(new_n13136, new_n13031, new_n13137);
and_8  g12761(new_n8413, new_n12953, new_n13138);
and_8  g12762(new_n12955, new_n12959, new_n13139);
nor_6  g12763(new_n13139, new_n13138, new_n13140);
and_8  g12764(n12145, n2226, new_n13141);
and_8  g12765(new_n12862, new_n12861, new_n13142);
or_8   g12766(new_n12862, new_n12861, new_n13143);
and_8  g12767(new_n13143, new_n12860, new_n13144);
or_8   g12768(new_n13144, new_n13142, new_n13145);
and_8  g12769(n9195, n6770, new_n13146);
and_8  g12770(n11222, n6431, new_n13147);
xor_4  g12771(new_n13147, new_n13146, new_n13148);
and_8  g12772(n10928, n10217, new_n13149);
and_8  g12773(n7320, n2024, new_n13150);
xor_4  g12774(new_n13150, new_n13149, new_n13151);
xor_4  g12775(new_n13151, new_n13148, new_n13152);
and_8  g12776(n5319, n3342, new_n13153);
and_8  g12777(n9457, n9111, new_n13154);
and_8  g12778(n9763, n4817, new_n13155);
xor_4  g12779(new_n13155, new_n13154, new_n13156);
xor_4  g12780(new_n13156, new_n13153, new_n13157);
xor_4  g12781(new_n13157, new_n13152, new_n13158);
xor_4  g12782(new_n13158, new_n13145, new_n13159);
xor_4  g12783(new_n13159, new_n13141, new_n13160);
xor_4  g12784(new_n13160, new_n13140, new_n13161);
or_8   g12785(new_n13161, new_n13137, new_n13162);
not_8  g12786(new_n13031, new_n13163);
xor_4  g12787(new_n13136, new_n13163, new_n13164);
not_8  g12788(new_n13161, new_n13165);
or_8   g12789(new_n13165, new_n13164, new_n13166);
and_8  g12790(new_n13166, new_n13162, new_n13167);
and_8  g12791(new_n12886, new_n12885, new_n13168);
and_8  g12792(new_n12888, new_n12858, new_n13169);
or_8   g12793(new_n13169, new_n13168, new_n13170);
or_8   g12794(new_n12919, new_n12915, new_n13171);
and_8  g12795(new_n12838, new_n12837, new_n13172);
and_8  g12796(new_n12840, new_n12835, new_n13173);
nor_6  g12797(new_n13173, new_n13172, new_n13174);
not_8  g12798(new_n12940, new_n13175);
or_8   g12799(new_n13175, new_n12935, new_n13176);
or_8   g12800(new_n12950, new_n12941, new_n13177);
and_8  g12801(new_n13177, new_n13176, new_n13178);
nand_5 g12802(new_n12892, new_n12891, new_n13179);
or_8   g12803(new_n12900, new_n12893, new_n13180);
and_8  g12804(new_n13180, new_n13179, new_n13181);
nand_5 g12805(n7891, n5798, new_n13182);
xor_4  g12806(new_n13182, new_n13181, new_n13183);
and_8  g12807(n12391, n2347, new_n13184);
and_8  g12808(n7265, n2087, new_n13185);
xor_4  g12809(new_n13185, new_n13184, new_n13186);
xor_4  g12810(new_n13186, new_n13183, new_n13187);
or_8   g12811(new_n13187, new_n13178, new_n13188);
nor_6  g12812(new_n13175, new_n12935, new_n13189);
nor_6  g12813(new_n12950, new_n12941, new_n13190);
or_8   g12814(new_n13190, new_n13189, new_n13191);
not_8  g12815(new_n13186, new_n13192);
xor_4  g12816(new_n13192, new_n13183, new_n13193);
or_8   g12817(new_n13193, new_n13191, new_n13194);
and_8  g12818(new_n13194, new_n13188, new_n13195);
and_8  g12819(n2498, n1199, new_n13196);
and_8  g12820(n6578, n2558, new_n13197);
xor_4  g12821(new_n13197, new_n13196, new_n13198);
xor_4  g12822(new_n13198, new_n13195, new_n13199);
and_8  g12823(new_n13199, new_n13174, new_n13200);
or_8   g12824(new_n13173, new_n13172, new_n13201);
not_8  g12825(new_n13198, new_n13202);
xor_4  g12826(new_n13202, new_n13195, new_n13203);
and_8  g12827(new_n13203, new_n13201, new_n13204);
or_8   g12828(new_n13204, new_n13200, new_n13205);
and_8  g12829(new_n13205, new_n13171, new_n13206);
nor_6  g12830(new_n12919, new_n12915, new_n13207);
or_8   g12831(new_n13203, new_n13201, new_n13208);
or_8   g12832(new_n13199, new_n13174, new_n13209);
and_8  g12833(new_n13209, new_n13208, new_n13210);
and_8  g12834(new_n13210, new_n13207, new_n13211);
or_8   g12835(new_n13211, new_n13206, new_n13212);
xor_4  g12836(new_n13212, new_n13170, new_n13213);
and_8  g12837(new_n13213, new_n13167, new_n13214);
and_8  g12838(new_n13165, new_n13164, new_n13215);
and_8  g12839(new_n13161, new_n13137, new_n13216);
or_8   g12840(new_n13216, new_n13215, new_n13217);
nor_6  g12841(new_n13212, new_n13170, new_n13218);
and_8  g12842(new_n13212, new_n13170, new_n13219);
or_8   g12843(new_n13219, new_n13218, new_n13220);
and_8  g12844(new_n13220, new_n13217, new_n13221);
or_8   g12845(new_n13221, new_n13214, new_n13222);
or_8   g12846(new_n12964, new_n12965, new_n13223);
or_8   g12847(new_n12947_1, new_n12946, new_n13224);
or_8   g12848(new_n12948, new_n12945, new_n13225);
and_8  g12849(new_n13225, new_n13224, new_n13226);
and_8  g12850(new_n12909, new_n12904, new_n13227);
and_8  g12851(new_n12910, new_n12901, new_n13228);
or_8   g12852(new_n13228, new_n13227, new_n13229);
xor_4  g12853(new_n13229, new_n13226, new_n13230);
xor_4  g12854(new_n13230, new_n13223, new_n13231);
and_8  g12855(new_n13231, new_n13222, new_n13232);
or_8   g12856(new_n13220, new_n13217, new_n13233);
or_8   g12857(new_n13213, new_n13167, new_n13234);
and_8  g12858(new_n13234, new_n13233, new_n13235);
and_8  g12859(new_n12975, new_n12957, new_n13236);
xor_4  g12860(new_n13230, new_n13236, new_n13237);
and_8  g12861(new_n13237, new_n13235, new_n13238);
or_8   g12862(new_n13238, new_n13232, new_n13239);
and_8  g12863(new_n13239, new_n13016, new_n13240);
or_8   g12864(new_n13015, new_n12971, new_n13241);
or_8   g12865(new_n13237, new_n13235, new_n13242);
or_8   g12866(new_n13231, new_n13222, new_n13243);
and_8  g12867(new_n13243, new_n13242, new_n13244);
and_8  g12868(new_n13244, new_n13241, new_n13245);
or_8   g12869(new_n13245, new_n13240, new_n13246);
and_8  g12870(new_n12841, new_n12815, new_n13247);
nor_6  g12871(new_n12846, new_n12843, new_n13248);
nor_6  g12872(new_n13248, new_n13247, new_n13249);
and_8  g12873(new_n12972, new_n12922, new_n13250);
not_8  g12874(new_n13250, new_n13251);
or_8   g12875(new_n13251, new_n13249, new_n13252);
or_8   g12876(new_n13248, new_n13247, new_n13253);
or_8   g12877(new_n13250, new_n13253, new_n13254);
and_8  g12878(new_n13254, new_n13252, new_n13255);
xor_4  g12879(new_n13255, new_n13246, new_n13256);
or_8   g12880(new_n13256, new_n13014, new_n13257);
and_8  g12881(new_n13006, new_n12984, new_n13258);
and_8  g12882(new_n13255, new_n13246, new_n13259);
nor_6  g12883(new_n13255, new_n13246, new_n13260);
or_8   g12884(new_n13260, new_n13259, new_n13261);
or_8   g12885(new_n13261, new_n13258, new_n13262);
and_8  g12886(new_n13262, new_n13257, new_n13263);
xor_4  g12887(new_n13263, new_n13013, n6192);
xor_4  g12888(new_n888, new_n860, n6273);
xor_4  g12889(new_n8001, new_n8248, n6445);
xnor_4 g12890(new_n10028, new_n10021, n6645);
xnor_4 g12891(new_n8475, new_n8474, n6689);
xor_4  g12892(new_n1340, new_n1339, n6742);
xor_4  g12893(new_n2111, new_n2062, n6809);
xor_4  g12894(new_n7111, new_n7247, n6822);
xnor_4 g12895(new_n11964, new_n11963, n6860);
xnor_4 g12896(new_n10017, new_n10010, n7193);
xor_4  g12897(new_n8253, new_n8251, n7568);
xnor_4 g12898(new_n1347, new_n1346, n7676);
and_8  g12899(new_n899, new_n483, new_n13276);
and_8  g12900(new_n1053, new_n910, new_n13277);
or_8   g12901(new_n13277, new_n13276, new_n13278);
and_8  g12902(new_n1047, new_n1049, new_n13279);
not_8  g12903(new_n1034, new_n13280);
or_8   g12904(new_n1040, new_n13280, new_n13281);
nand_5 g12905(n9241, n1209, new_n13282);
and_8  g12906(new_n1016, new_n991, new_n13283);
nor_6  g12907(new_n1028, new_n13283, new_n13284);
and_8  g12908(new_n1013, new_n1012, new_n13285);
or_8   g12909(new_n1019, new_n13285, new_n13286);
xnor_4 g12910(new_n445, new_n442, new_n13287);
or_8   g12911(new_n13287, new_n441, new_n13288);
or_8   g12912(new_n456, new_n447_1, new_n13289);
nand_5 g12913(new_n13289, new_n13288, new_n13290);
not_8  g12914(new_n13290, new_n13291);
nand_5 g12915(new_n449, new_n448, new_n13292);
or_8   g12916(new_n455, new_n450, new_n13293);
and_8  g12917(new_n13293, new_n13292, new_n13294);
nand_5 g12918(n12705, n2508, new_n13295);
and_8  g12919(new_n444, new_n443, new_n13296);
or_8   g12920(new_n444, new_n443, new_n13297);
and_8  g12921(new_n13297, new_n442, new_n13298);
or_8   g12922(new_n13298, new_n13296, new_n13299);
xor_4  g12923(new_n13299, new_n13295, new_n13300);
and_8  g12924(n3986, n1980, new_n13301);
and_8  g12925(n10848, n5857, new_n13302);
xor_4  g12926(new_n13302, new_n13301, new_n13303);
and_8  g12927(n11257, n2509, new_n13304);
and_8  g12928(n4005, n1097, new_n13305);
xor_4  g12929(new_n13305, new_n13304, new_n13306);
xor_4  g12930(new_n13306, new_n13303, new_n13307);
xor_4  g12931(new_n13307, new_n13300, new_n13308);
xor_4  g12932(new_n13308, new_n13294, new_n13309);
not_8  g12933(new_n13309, new_n13310);
and_8  g12934(n8028, n45, new_n13311);
or_8   g12935(new_n917, new_n916, new_n13312);
or_8   g12936(new_n918, new_n915, new_n13313);
and_8  g12937(new_n13313, new_n13312, new_n13314);
xor_4  g12938(new_n13314, new_n13311, new_n13315);
and_8  g12939(new_n926, new_n925, new_n13316);
or_8   g12940(new_n926, new_n925, new_n13317);
and_8  g12941(new_n13317, new_n924, new_n13318);
or_8   g12942(new_n13318, new_n13316, new_n13319);
xor_4  g12943(new_n13319, new_n13315, new_n13320);
nand_5 g12944(n4312, n2585, new_n13321);
or_8   g12945(new_n453, new_n452, new_n13322);
or_8   g12946(new_n454, new_n451, new_n13323);
and_8  g12947(new_n13323, new_n13322, new_n13324);
nand_5 g12948(n10644, n7354, new_n13325);
and_8  g12949(n12706, n5964, new_n13326);
and_8  g12950(n12720, n12025, new_n13327);
xor_4  g12951(new_n13327, new_n13326, new_n13328);
xor_4  g12952(new_n13328, new_n13325, new_n13329);
xor_4  g12953(new_n13329, new_n13324, new_n13330);
xor_4  g12954(new_n13330, new_n13321, new_n13331);
and_8  g12955(new_n13331, new_n13320, new_n13332);
nor_6  g12956(new_n13331, new_n13320, new_n13333);
or_8   g12957(new_n13333, new_n13332, new_n13334);
not_8  g12958(new_n13334, new_n13335);
xor_4  g12959(new_n13335, new_n13310, new_n13336);
xor_4  g12960(new_n13336, new_n13291, new_n13337);
and_8  g12961(n7436, n4141, new_n13338);
nand_5 g12962(new_n922, new_n921, new_n13339);
or_8   g12963(new_n928, new_n923, new_n13340);
and_8  g12964(new_n13340, new_n13339, new_n13341);
xor_4  g12965(new_n13341, new_n13338, new_n13342);
xor_4  g12966(new_n13342, new_n13337, new_n13343);
xor_4  g12967(new_n13343, new_n13286, new_n13344);
not_8  g12968(new_n13344, new_n13345);
and_8  g12969(new_n13345, new_n13284, new_n13346);
or_8   g12970(new_n1028, new_n13283, new_n13347);
and_8  g12971(new_n13344, new_n13347, new_n13348);
or_8   g12972(new_n13348, new_n13346, new_n13349);
and_8  g12973(new_n13349, new_n13282, new_n13350);
not_8  g12974(new_n13282, new_n13351);
or_8   g12975(new_n13344, new_n13347, new_n13352);
or_8   g12976(new_n13345, new_n13284, new_n13353);
and_8  g12977(new_n13353, new_n13352, new_n13354);
and_8  g12978(new_n13354, new_n13351, new_n13355);
or_8   g12979(new_n13355, new_n13350, new_n13356);
xor_4  g12980(new_n13356, new_n13281, new_n13357);
and_8  g12981(n10547, n6038, new_n13358);
or_8   g12982(new_n960, new_n959, new_n13359);
or_8   g12983(new_n961, new_n958, new_n13360);
and_8  g12984(new_n13360, new_n13359, new_n13361);
xor_4  g12985(new_n13361, new_n13358, new_n13362);
or_8   g12986(new_n969, new_n968, new_n13363);
or_8   g12987(new_n970, new_n967, new_n13364);
and_8  g12988(new_n13364, new_n13363, new_n13365);
nand_5 g12989(n12044, n8476, new_n13366);
and_8  g12990(n11892, n5814, new_n13367);
and_8  g12991(n3616, n1512, new_n13368);
xor_4  g12992(new_n13368, new_n13367, new_n13369);
xor_4  g12993(new_n13369, new_n13366, new_n13370);
xor_4  g12994(new_n13370, new_n13365, new_n13371);
xor_4  g12995(new_n13371, new_n13362, new_n13372);
and_8  g12996(n12299, n4928, new_n13373);
or_8   g12997(new_n1006, new_n1005, new_n13374);
or_8   g12998(new_n1007, new_n1004, new_n13375);
and_8  g12999(new_n13375, new_n13374, new_n13376);
xor_4  g13000(new_n13376, new_n13373, new_n13377);
and_8  g13001(n5069, n2530, new_n13378);
and_8  g13002(n10545, n2802, new_n13379);
xor_4  g13003(new_n13379, new_n13378, new_n13380);
xor_4  g13004(new_n13380, new_n13377, new_n13381);
xor_4  g13005(new_n13381, new_n13372, new_n13382);
nand_5 g13006(new_n962, new_n957, new_n13383);
or_8   g13007(new_n972, new_n963, new_n13384);
and_8  g13008(new_n13384, new_n13383, new_n13385);
nand_5 g13009(new_n1002, new_n1001, new_n13386);
or_8   g13010(new_n1008, new_n1003, new_n13387);
and_8  g13011(new_n13387, new_n13386, new_n13388);
and_8  g13012(new_n965, new_n964, new_n13389);
nor_6  g13013(new_n971, new_n966, new_n13390);
or_8   g13014(new_n13390, new_n13389, new_n13391);
nand_5 g13015(n7690, n533, new_n13392);
xor_4  g13016(new_n13392, new_n13391, new_n13393);
xor_4  g13017(new_n13393, new_n13388, new_n13394);
or_8   g13018(new_n13394, new_n13385, new_n13395);
not_8  g13019(new_n13383, new_n13396);
or_8   g13020(new_n973, new_n13396, new_n13397);
not_8  g13021(new_n13388, new_n13398);
xor_4  g13022(new_n13393, new_n13398, new_n13399);
or_8   g13023(new_n13399, new_n13397, new_n13400);
and_8  g13024(new_n13400, new_n13395, new_n13401);
nor_6  g13025(new_n13401, new_n13382, new_n13402);
and_8  g13026(new_n13401, new_n13382, new_n13403);
or_8   g13027(new_n13403, new_n13402, new_n13404);
and_8  g13028(n12704, n2393, new_n13405);
and_8  g13029(n7294, n5860, new_n13406);
xor_4  g13030(new_n13406, new_n13405, new_n13407);
and_8  g13031(n12648, n6806, new_n13408);
and_8  g13032(n4499, n1564, new_n13409);
xor_4  g13033(new_n13409, new_n13408, new_n13410);
xor_4  g13034(new_n13410, new_n13407, new_n13411);
or_8   g13035(new_n997, new_n996_1, new_n13412);
or_8   g13036(new_n998, new_n995, new_n13413);
and_8  g13037(new_n13413, new_n13412, new_n13414);
and_8  g13038(n5694, n5331, new_n13415);
and_8  g13039(n7388, n4903, new_n13416);
xor_4  g13040(new_n13416, new_n13415, new_n13417);
xor_4  g13041(new_n13417, new_n13414, new_n13418);
xor_4  g13042(new_n13418, new_n13411, new_n13419);
and_8  g13043(n8276, n5105, new_n13420);
and_8  g13044(n5305, n615, new_n13421);
xor_4  g13045(new_n13421, new_n13420, new_n13422);
xor_4  g13046(new_n13422, new_n13419, new_n13423);
not_8  g13047(new_n13423, new_n13424);
and_8  g13048(new_n13424, new_n13404, new_n13425);
xor_4  g13049(new_n13401, new_n13382, new_n13426);
and_8  g13050(new_n13423, new_n13426, new_n13427);
or_8   g13051(new_n13427, new_n13425, new_n13428);
and_8  g13052(new_n550, new_n932, new_n13429);
or_8   g13053(new_n935, new_n13429, new_n13430);
and_8  g13054(new_n788, new_n977, new_n13431);
or_8   g13055(new_n980, new_n13431, new_n13432);
xor_4  g13056(new_n13432, new_n13430, new_n13433);
or_8   g13057(new_n13433, new_n13428, new_n13434);
or_8   g13058(new_n13423, new_n13426, new_n13435);
or_8   g13059(new_n13424, new_n13404, new_n13436);
and_8  g13060(new_n13436, new_n13435, new_n13437);
not_8  g13061(new_n13432, new_n13438);
xor_4  g13062(new_n13438, new_n13430, new_n13439);
or_8   g13063(new_n13439, new_n13437, new_n13440);
and_8  g13064(new_n13440, new_n13434, new_n13441);
and_8  g13065(n8759, n783, new_n13442);
and_8  g13066(n10510, n7500, new_n13443);
xor_4  g13067(new_n13443, new_n13442, new_n13444);
not_8  g13068(new_n461, new_n13445);
or_8   g13069(new_n464, new_n457, new_n13446);
and_8  g13070(new_n13446, new_n13445, new_n13447);
nand_5 g13071(new_n999, new_n994, new_n13448);
not_8  g13072(new_n1000, new_n13449);
or_8   g13073(new_n1009, new_n13449, new_n13450);
nand_5 g13074(new_n13450, new_n13448, new_n13451);
not_8  g13075(new_n13451, new_n13452);
and_8  g13076(new_n13452, new_n13447, new_n13453);
nor_6  g13077(new_n13452, new_n13447, new_n13454);
or_8   g13078(new_n13454, new_n13453, new_n13455);
xor_4  g13079(new_n13455, new_n13444, new_n13456);
or_8   g13080(new_n13456, new_n13441, new_n13457);
and_8  g13081(new_n13439, new_n13437, new_n13458);
and_8  g13082(new_n13433, new_n13428, new_n13459);
or_8   g13083(new_n13459, new_n13458, new_n13460);
not_8  g13084(new_n13444, new_n13461);
xor_4  g13085(new_n13455, new_n13461, new_n13462);
or_8   g13086(new_n13462, new_n13460, new_n13463);
and_8  g13087(new_n13463, new_n13457, new_n13464);
not_8  g13088(new_n985, new_n13465);
or_8   g13089(new_n989, new_n1031, new_n13466);
and_8  g13090(new_n13466, new_n13465, new_n13467);
nand_5 g13091(n7965, n1906, new_n13468);
not_8  g13092(new_n13468, new_n13469);
xor_4  g13093(new_n13469, new_n13467, new_n13470);
and_8  g13094(new_n13470, new_n13464, new_n13471);
and_8  g13095(new_n13462, new_n13460, new_n13472);
and_8  g13096(new_n13456, new_n13441, new_n13473);
or_8   g13097(new_n13473, new_n13472, new_n13474);
xor_4  g13098(new_n13468, new_n13467, new_n13475);
and_8  g13099(new_n13475, new_n13474, new_n13476);
or_8   g13100(new_n13476, new_n13471, new_n13477);
and_8  g13101(new_n465, new_n438, new_n13478);
and_8  g13102(new_n482, new_n466, new_n13479);
or_8   g13103(new_n13479, new_n13478, new_n13480);
not_8  g13104(new_n949, new_n13481);
or_8   g13105(new_n953, new_n950, new_n13482);
and_8  g13106(new_n13482, new_n13481, new_n13483);
and_8  g13107(new_n919, new_n914, new_n13484);
and_8  g13108(new_n936, new_n920, new_n13485);
or_8   g13109(new_n13485, new_n13484, new_n13486);
and_8  g13110(n8236, n6776, new_n13487);
xor_4  g13111(new_n13487, new_n13486, new_n13488);
xor_4  g13112(new_n13488, new_n13483, new_n13489);
or_8   g13113(new_n13489, new_n13480, new_n13490);
nor_6  g13114(new_n13479, new_n13478, new_n13491);
not_8  g13115(new_n13488, new_n13492);
xor_4  g13116(new_n13492, new_n13483, new_n13493);
or_8   g13117(new_n13493, new_n13491, new_n13494);
and_8  g13118(new_n13494, new_n13490, new_n13495);
xor_4  g13119(new_n13495, new_n13477, new_n13496);
and_8  g13120(new_n13496, new_n13357, new_n13497);
nor_6  g13121(new_n13356, new_n13281, new_n13498);
and_8  g13122(new_n13356, new_n13281, new_n13499);
or_8   g13123(new_n13499, new_n13498, new_n13500);
nor_6  g13124(new_n13495, new_n13477, new_n13501);
and_8  g13125(new_n13495, new_n13477, new_n13502);
or_8   g13126(new_n13502, new_n13501, new_n13503);
and_8  g13127(new_n13503, new_n13500, new_n13504);
or_8   g13128(new_n13504, new_n13497, new_n13505);
or_8   g13129(new_n13505, new_n13279, new_n13506);
and_8  g13130(new_n1051, new_n1050, new_n13507);
or_8   g13131(new_n13507, new_n1043, new_n13508);
or_8   g13132(new_n13503, new_n13500, new_n13509);
or_8   g13133(new_n13496, new_n13357, new_n13510);
and_8  g13134(new_n13510, new_n13509, new_n13511);
or_8   g13135(new_n13511, new_n13508, new_n13512);
and_8  g13136(new_n13512, new_n13506, new_n13513);
xor_4  g13137(new_n13513, new_n13278, n7966);
nor_6  g13138(new_n13010, new_n13009, new_n13515);
xor_4  g13139(new_n13515, new_n13004, n7981);
and_8  g13140(new_n12546, new_n12542, new_n13517);
and_8  g13141(new_n12540, new_n12290, new_n13518);
or_8   g13142(new_n13518, new_n13517, new_n13519);
or_8   g13143(new_n12561, new_n13519, new_n13520);
and_8  g13144(new_n13520, new_n12541, new_n13521);
and_8  g13145(new_n12539, new_n12464, new_n13522);
or_8   g13146(new_n13522, new_n12544, new_n13523);
or_8   g13147(new_n12533, new_n12530, new_n13524);
or_8   g13148(new_n12538, new_n12535, new_n13525);
and_8  g13149(new_n13525, new_n13524, new_n13526);
and_8  g13150(new_n12522, new_n12425, new_n13527);
or_8   g13151(new_n12532, new_n13527, new_n13528);
and_8  g13152(new_n12273, new_n12260, new_n13529);
and_8  g13153(new_n12512, new_n12511_1, new_n13530);
or_8   g13154(new_n12512, new_n12511_1, new_n13531);
and_8  g13155(new_n13531, new_n12510, new_n13532);
or_8   g13156(new_n13532, new_n13530, new_n13533);
nand_5 g13157(n8717, n6986, new_n13534);
and_8  g13158(n11222, n10022, new_n13535);
and_8  g13159(n12391, n1353, new_n13536);
xor_4  g13160(new_n13536, new_n13535, new_n13537);
xor_4  g13161(new_n13537, new_n13534, new_n13538);
xor_4  g13162(new_n13538, new_n13533, new_n13539);
xor_4  g13163(new_n13539, new_n13529, new_n13540);
xnor_4 g13164(new_n13540, new_n13528, new_n13541);
xor_4  g13165(new_n13541, new_n13526, new_n13542);
and_8  g13166(new_n12519, new_n12518, new_n13543);
and_8  g13167(new_n12521, new_n12516, new_n13544);
or_8   g13168(new_n13544, new_n13543, new_n13545);
nand_5 g13169(new_n12504, new_n12499, new_n13546);
not_8  g13170(new_n12505, new_n13547);
or_8   g13171(new_n12515, new_n13547, new_n13548);
and_8  g13172(new_n13548, new_n13546, new_n13549);
and_8  g13173(n12069, n4436, new_n13550);
and_8  g13174(n11999, n11153, new_n13551);
xor_4  g13175(new_n13551, new_n13550, new_n13552);
and_8  g13176(n7159, n1199, new_n13553);
and_8  g13177(n11967, n7160, new_n13554);
xnor_4 g13178(new_n13554, new_n13553, new_n13555);
xor_4  g13179(new_n13555, new_n13552, new_n13556);
and_8  g13180(new_n12502, new_n12501, new_n13557);
or_8   g13181(new_n12502, new_n12501, new_n13558);
and_8  g13182(new_n13558, new_n12500, new_n13559);
or_8   g13183(new_n13559, new_n13557, new_n13560);
and_8  g13184(n6254, n4828, new_n13561);
and_8  g13185(n11407, n2087, new_n13562);
xor_4  g13186(new_n13562, new_n13561, new_n13563);
xor_4  g13187(new_n13563, new_n13560, new_n13564);
xor_4  g13188(new_n13564, new_n13556, new_n13565);
xor_4  g13189(new_n13565, new_n13549, new_n13566);
xor_4  g13190(new_n13566, new_n13545, new_n13567);
and_8  g13191(new_n12472, new_n12467, new_n13568);
not_8  g13192(new_n13568, new_n13569);
or_8   g13193(new_n12482, new_n12473, new_n13570);
and_8  g13194(new_n13570, new_n13569, new_n13571);
and_8  g13195(n12489, n6578, new_n13572);
and_8  g13196(n12947, n996, new_n13573);
and_8  g13197(n9457, n5760, new_n13574);
xor_4  g13198(new_n13574, new_n13573, new_n13575);
xor_4  g13199(new_n13575, new_n13572, new_n13576);
xor_4  g13200(new_n13576, new_n13571, new_n13577);
and_8  g13201(new_n12507, new_n12506, new_n13578);
and_8  g13202(new_n12514, new_n12508, new_n13579);
or_8   g13203(new_n13579, new_n13578, new_n13580);
and_8  g13204(n7891, n447, new_n13581);
xor_4  g13205(new_n13581, new_n13580, new_n13582);
and_8  g13206(n12777, n2515, new_n13583);
or_8   g13207(new_n12479, new_n12478, new_n13584);
not_8  g13208(new_n12477, new_n13585);
or_8   g13209(new_n12480, new_n13585, new_n13586);
and_8  g13210(new_n13586, new_n13584, new_n13587);
or_8   g13211(new_n12470, new_n12469, new_n13588);
or_8   g13212(new_n12471, new_n12468, new_n13589);
and_8  g13213(new_n13589, new_n13588, new_n13590);
xor_4  g13214(new_n13590, new_n13587, new_n13591);
xor_4  g13215(new_n13591, new_n13583, new_n13592);
xor_4  g13216(new_n13592, new_n13582, new_n13593);
and_8  g13217(n6441, n5314, new_n13594);
and_8  g13218(n11791, n5767, new_n13595);
xor_4  g13219(new_n13595, new_n13594, new_n13596);
and_8  g13220(new_n12475, new_n12474, new_n13597);
and_8  g13221(new_n12481, new_n12476, new_n13598);
or_8   g13222(new_n13598, new_n13597, new_n13599);
nand_5 g13223(n6687, n6604, new_n13600);
xor_4  g13224(new_n13600, new_n13599, new_n13601);
xor_4  g13225(new_n13601, new_n13596, new_n13602);
xor_4  g13226(new_n13602, new_n13593, new_n13603);
xor_4  g13227(new_n13603, new_n13577, new_n13604);
and_8  g13228(new_n13604, new_n13567, new_n13605);
nor_6  g13229(new_n13604, new_n13567, new_n13606);
or_8   g13230(new_n13606, new_n13605, new_n13607);
not_8  g13231(new_n12339, new_n13608);
and_8  g13232(new_n12340, new_n13608, new_n13609);
nor_6  g13233(new_n12342, new_n12337, new_n13610);
or_8   g13234(new_n13610, new_n13609, new_n13611);
nand_5 g13235(new_n12326, new_n12321, new_n13612);
or_8   g13236(new_n12336, new_n12327, new_n13613);
and_8  g13237(new_n13613, new_n13612, new_n13614);
and_8  g13238(n10678, n6429, new_n13615);
xor_4  g13239(new_n13615, new_n13614, new_n13616);
nand_5 g13240(new_n12329, new_n12328, new_n13617);
or_8   g13241(new_n12335, new_n12330, new_n13618);
and_8  g13242(new_n13618, new_n13617, new_n13619);
and_8  g13243(n2433, n2226, new_n13620);
and_8  g13244(n8819, n1094, new_n13621);
and_8  g13245(n10928, n7730, new_n13622);
xor_4  g13246(new_n13622, new_n13621, new_n13623);
xor_4  g13247(new_n13623, new_n13620, new_n13624);
xor_4  g13248(new_n13624, new_n13619, new_n13625);
xor_4  g13249(new_n13625, new_n13616, new_n13626);
xor_4  g13250(new_n13626, new_n13611, new_n13627);
and_8  g13251(new_n13627, new_n13607, new_n13628);
xor_4  g13252(new_n13604, new_n13567, new_n13629);
not_8  g13253(new_n13611, new_n13630);
xor_4  g13254(new_n13626, new_n13630, new_n13631);
and_8  g13255(new_n13631, new_n13629, new_n13632);
or_8   g13256(new_n13632, new_n13628, new_n13633);
not_8  g13257(new_n12485, new_n13634);
nand_5 g13258(new_n12486, new_n13634, new_n13635);
or_8   g13259(new_n12488, new_n12483, new_n13636);
nand_5 g13260(new_n13636, new_n13635, new_n13637);
not_8  g13261(new_n12235, new_n13638);
or_8   g13262(new_n13638, new_n12283, new_n13639);
xor_4  g13263(new_n12272, new_n12258, new_n13640);
or_8   g13264(new_n13640, new_n13639, new_n13641);
not_8  g13265(new_n13641, new_n13642);
and_8  g13266(new_n12289, new_n12275, new_n13643);
or_8   g13267(new_n13643, new_n13642, new_n13644);
or_8   g13268(new_n13644, new_n13637, new_n13645);
not_8  g13269(new_n13637, new_n13646);
xor_4  g13270(new_n12274, new_n13639, new_n13647);
or_8   g13271(new_n11201, new_n11181, new_n13648);
and_8  g13272(new_n12284, new_n12276, new_n13649);
or_8   g13273(new_n13649, new_n12279, new_n13650);
or_8   g13274(new_n13650, new_n13648, new_n13651);
and_8  g13275(new_n13651, new_n12285, new_n13652);
or_8   g13276(new_n13652, new_n13647, new_n13653);
and_8  g13277(new_n13653, new_n13641, new_n13654);
or_8   g13278(new_n13654, new_n13646, new_n13655);
and_8  g13279(new_n13655, new_n13645, new_n13656);
and_8  g13280(new_n13656, new_n13633, new_n13657);
nor_6  g13281(new_n13656, new_n13633, new_n13658);
or_8   g13282(new_n13658, new_n13657, new_n13659);
nor_6  g13283(new_n12529, new_n12491, new_n13660);
and_8  g13284(new_n12343, new_n12318, new_n13661);
and_8  g13285(new_n12344, new_n12317, new_n13662);
or_8   g13286(new_n13662, new_n13661, new_n13663);
not_8  g13287(new_n12239, new_n13664);
nand_5 g13288(new_n12244, new_n13664, new_n13665);
nand_5 g13289(new_n12255, new_n13665, new_n13666);
and_8  g13290(new_n12242, new_n12241, new_n13667);
or_8   g13291(new_n12242, new_n12241, new_n13668);
and_8  g13292(new_n13668, new_n12240, new_n13669);
or_8   g13293(new_n13669, new_n13667, new_n13670);
and_8  g13294(n12709, n7523, new_n13671);
and_8  g13295(n12000, n4189, new_n13672);
xor_4  g13296(new_n13672, new_n13671, new_n13673);
xor_4  g13297(new_n13673, new_n13670, new_n13674);
and_8  g13298(n9725, n2564, new_n13675);
and_8  g13299(n9920, n4370, new_n13676);
xor_4  g13300(new_n13676, new_n13675, new_n13677);
and_8  g13301(n5212, n4516, new_n13678);
and_8  g13302(n6770, n5320, new_n13679);
and_8  g13303(n5319, n1478, new_n13680);
xor_4  g13304(new_n13680, new_n13679, new_n13681);
xor_4  g13305(new_n13681, new_n13678, new_n13682);
xor_4  g13306(new_n13682, new_n13677, new_n13683);
and_8  g13307(n11728, n7320, new_n13684);
or_8   g13308(new_n12333, new_n12332, new_n13685);
or_8   g13309(new_n12334, new_n12331, new_n13686);
and_8  g13310(new_n13686, new_n13685, new_n13687);
xor_4  g13311(new_n13687, new_n13684, new_n13688);
xor_4  g13312(new_n13688, new_n13683, new_n13689);
xor_4  g13313(new_n13689, new_n13674, new_n13690);
and_8  g13314(new_n12251, new_n12250, new_n13691);
or_8   g13315(new_n12251, new_n12250, new_n13692);
and_8  g13316(new_n13692, new_n12249, new_n13693);
or_8   g13317(new_n13693, new_n13691, new_n13694);
nand_5 g13318(n10990, n4817, new_n13695);
and_8  g13319(n11877, n3627, new_n13696);
and_8  g13320(n8336, n1198, new_n13697);
xor_4  g13321(new_n13697, new_n13696, new_n13698);
xor_4  g13322(new_n13698, new_n13695, new_n13699);
xor_4  g13323(new_n13699, new_n13694, new_n13700);
and_8  g13324(new_n12247_1, new_n12246, new_n13701);
nor_6  g13325(new_n12253, new_n12248, new_n13702);
or_8   g13326(new_n13702, new_n13701, new_n13703);
or_8   g13327(new_n12324, new_n12323, new_n13704);
or_8   g13328(new_n12325, new_n12322, new_n13705);
and_8  g13329(new_n13705, new_n13704, new_n13706);
xor_4  g13330(new_n13706, new_n13703, new_n13707);
xor_4  g13331(new_n13707, new_n13700, new_n13708);
xor_4  g13332(new_n13708, new_n13690, new_n13709);
xor_4  g13333(new_n13709, new_n13666, new_n13710);
not_8  g13334(new_n13710, new_n13711);
or_8   g13335(new_n13711, new_n13663, new_n13712);
not_8  g13336(new_n13661, new_n13713);
not_8  g13337(new_n12314, new_n13714);
and_8  g13338(new_n12349, new_n13714, new_n13715);
not_8  g13339(new_n12343, new_n13716);
xor_4  g13340(new_n13716, new_n12318, new_n13717);
or_8   g13341(new_n13717, new_n13715, new_n13718);
and_8  g13342(new_n13718, new_n13713, new_n13719);
or_8   g13343(new_n13710, new_n13719, new_n13720);
and_8  g13344(new_n13720, new_n13712, new_n13721);
xor_4  g13345(new_n13721, new_n13660, new_n13722);
and_8  g13346(new_n13722, new_n13659, new_n13723);
xor_4  g13347(new_n13656, new_n13633, new_n13724);
or_8   g13348(new_n12529, new_n12491, new_n13725);
xor_4  g13349(new_n13721, new_n13725, new_n13726);
and_8  g13350(new_n13726, new_n13724, new_n13727);
or_8   g13351(new_n13727, new_n13723, new_n13728);
or_8   g13352(new_n13728, new_n13542, new_n13729);
xor_4  g13353(new_n13540, new_n13528, new_n13730);
xor_4  g13354(new_n13730, new_n13526, new_n13731);
or_8   g13355(new_n13726, new_n13724, new_n13732);
or_8   g13356(new_n13722, new_n13659, new_n13733);
and_8  g13357(new_n13733, new_n13732, new_n13734);
or_8   g13358(new_n13734, new_n13731, new_n13735);
and_8  g13359(new_n13735, new_n13729, new_n13736);
xor_4  g13360(new_n13736, new_n13523, new_n13737);
and_8  g13361(new_n13737, new_n13521, new_n13738);
not_8  g13362(new_n12549, new_n13739);
and_8  g13363(new_n12556, new_n13739, new_n13740);
xor_4  g13364(new_n12556, new_n13739, new_n13741);
and_8  g13365(new_n12558, new_n13741, new_n13742);
or_8   g13366(new_n13742, new_n13740, new_n13743);
and_8  g13367(new_n13743, new_n12548, new_n13744);
or_8   g13368(new_n13744, new_n13517, new_n13745);
nor_6  g13369(new_n13522, new_n12544, new_n13746);
xor_4  g13370(new_n13736, new_n13746, new_n13747);
and_8  g13371(new_n13747, new_n13745, new_n13748);
or_8   g13372(new_n13748, new_n13738, n8100);
xnor_4 g13373(new_n10015, new_n10014, n8138);
xnor_4 g13374(new_n6218, new_n6217, n8202);
xor_4  g13375(new_n3783, new_n3774, n8303);
xnor_4 g13376(new_n3033, new_n3032, n8398);
xnor_4 g13377(new_n4331, new_n4330, n9137);
xnor_4 g13378(new_n7253, new_n7243, n9387);
xnor_4 g13379(new_n11978, new_n11977, n9571);
xor_4  g13380(new_n897, new_n890, n9578);
xor_4  g13381(new_n1163, new_n1161, n9706);
xnor_4 g13382(new_n4333_1, new_n4325, n9756);
and_8  g13383(new_n6906, new_n6517, new_n13760);
and_8  g13384(new_n6924, new_n6907, new_n13761);
or_8   g13385(new_n13761, new_n13760, new_n13762);
and_8  g13386(n12826, n7891, new_n13763);
nand_5 g13387(new_n6554, new_n6593, new_n13764);
not_8  g13388(new_n6598, new_n13765);
and_8  g13389(new_n13765, new_n13764, new_n13766);
xor_4  g13390(new_n13766, new_n13763, new_n13767);
or_8   g13391(new_n6865, new_n6618, new_n13768);
or_8   g13392(new_n6905, new_n6868, new_n13769);
and_8  g13393(new_n13769, new_n13768, new_n13770);
nand_5 g13394(n8336, n2278, new_n13771);
not_8  g13395(new_n13771, new_n13772);
nor_6  g13396(new_n6503, new_n6500, new_n13773);
or_8   g13397(new_n6515, new_n6510, new_n13774);
and_8  g13398(new_n13774, new_n13773, new_n13775);
or_8   g13399(new_n13775, new_n6503, new_n13776);
or_8   g13400(new_n13776, new_n13772, new_n13777);
not_8  g13401(new_n6503, new_n13778);
or_8   g13402(new_n6516, new_n6504, new_n13779);
and_8  g13403(new_n13779, new_n13778, new_n13780);
or_8   g13404(new_n13780, new_n13771, new_n13781);
and_8  g13405(new_n13781, new_n13777, new_n13782);
not_8  g13406(new_n6702, new_n13783);
and_8  g13407(new_n6717, new_n6703_1, new_n13784);
or_8   g13408(new_n13784, new_n13783, new_n13785);
nand_5 g13409(new_n6483, new_n6482, new_n13786);
or_8   g13410(new_n6489, new_n6484, new_n13787);
nand_5 g13411(new_n13787, new_n13786, new_n13788);
not_8  g13412(new_n13788, new_n13789);
not_8  g13413(new_n6577, new_n13790);
nor_6  g13414(new_n13790, new_n6572, new_n13791);
or_8   g13415(new_n6589, new_n13791, new_n13792);
nand_5 g13416(n11662, n6770, new_n13793);
and_8  g13417(n10451, n2226, new_n13794);
and_8  g13418(n5319, n3754, new_n13795);
xor_4  g13419(new_n13795, new_n13794, new_n13796);
xor_4  g13420(new_n13796, new_n13793, new_n13797);
nor_6  g13421(new_n6585, new_n6584, new_n13798);
and_8  g13422(new_n6586, new_n6583, new_n13799);
or_8   g13423(new_n13799, new_n13798, new_n13800);
not_8  g13424(new_n13800, new_n13801);
xor_4  g13425(new_n13801, new_n13797, new_n13802);
and_8  g13426(new_n6487, new_n6486, new_n13803);
or_8   g13427(new_n6487, new_n6486, new_n13804);
and_8  g13428(new_n13804, new_n6485, new_n13805);
or_8   g13429(new_n13805, new_n13803, new_n13806);
and_8  g13430(n10278, n6986, new_n13807);
and_8  g13431(n10678, n3022, new_n13808);
xnor_4 g13432(new_n13808, new_n13807, new_n13809);
xor_4  g13433(new_n13809, new_n13806, new_n13810);
not_8  g13434(new_n13810, new_n13811);
and_8  g13435(new_n13811, new_n13802, new_n13812);
xor_4  g13436(new_n13800, new_n13797, new_n13813);
and_8  g13437(new_n13810, new_n13813, new_n13814);
or_8   g13438(new_n13814, new_n13812, new_n13815);
and_8  g13439(new_n6580, new_n6579, new_n13816);
nor_6  g13440(new_n6587, new_n6581, new_n13817);
or_8   g13441(new_n13817, new_n13816, new_n13818);
nor_6  g13442(new_n6575, new_n6574, new_n13819);
nor_6  g13443(new_n6576, new_n6573, new_n13820);
or_8   g13444(new_n13820, new_n13819, new_n13821);
not_8  g13445(new_n13821, new_n13822);
xor_4  g13446(new_n13822, new_n13818, new_n13823);
or_8   g13447(new_n13823, new_n13815, new_n13824);
or_8   g13448(new_n13810, new_n13813, new_n13825);
or_8   g13449(new_n13811, new_n13802, new_n13826);
and_8  g13450(new_n13826, new_n13825, new_n13827);
xor_4  g13451(new_n13821, new_n13818, new_n13828);
or_8   g13452(new_n13828, new_n13827, new_n13829);
and_8  g13453(new_n13829, new_n13824, new_n13830);
and_8  g13454(new_n13830, new_n13792, new_n13831);
or_8   g13455(new_n13790, new_n6572, new_n13832);
or_8   g13456(new_n6588, new_n6578_1, new_n13833);
and_8  g13457(new_n13833, new_n13832, new_n13834);
and_8  g13458(new_n13828, new_n13827, new_n13835);
and_8  g13459(new_n13823, new_n13815, new_n13836);
or_8   g13460(new_n13836, new_n13835, new_n13837);
and_8  g13461(new_n13837, new_n13834, new_n13838);
or_8   g13462(new_n13838, new_n13831, new_n13839);
xor_4  g13463(new_n13839, new_n13789, new_n13840);
or_8   g13464(new_n6478, new_n6477, new_n13841);
or_8   g13465(new_n6479, new_n6476, new_n13842);
and_8  g13466(new_n13842, new_n13841, new_n13843);
and_8  g13467(n8665, n2515, new_n13844);
and_8  g13468(n10898, n9457, new_n13845);
and_8  g13469(n12511, n11222, new_n13846);
xor_4  g13470(new_n13846, new_n13845, new_n13847);
xor_4  g13471(new_n13847, new_n13844, new_n13848);
xor_4  g13472(new_n13848, new_n13843, new_n13849);
and_8  g13473(new_n13849, new_n13840, new_n13850);
xor_4  g13474(new_n13839, new_n13788, new_n13851);
not_8  g13475(new_n13849, new_n13852);
and_8  g13476(new_n13852, new_n13851, new_n13853);
or_8   g13477(new_n13853, new_n13850, new_n13854);
nand_5 g13478(n12391, n4094, new_n13855);
not_8  g13479(new_n13855, new_n13856);
not_8  g13480(new_n6475, new_n13857);
and_8  g13481(new_n6480, new_n13857, new_n13858);
nor_6  g13482(new_n6490, new_n6481, new_n13859);
or_8   g13483(new_n13859, new_n13858, new_n13860);
and_8  g13484(n4516, n3932, new_n13861);
and_8  g13485(n7523, n6703, new_n13862);
xnor_4 g13486(new_n13862, new_n13861, new_n13863);
and_8  g13487(n11423, n10928, new_n13864);
and_8  g13488(n12591, n3627, new_n13865);
xor_4  g13489(new_n13865, new_n13864, new_n13866);
xor_4  g13490(new_n13866, new_n13863, new_n13867);
xor_4  g13491(new_n13867, new_n13860, new_n13868);
and_8  g13492(n11876, n4817, new_n13869);
nand_5 g13493(new_n6687_1, new_n6684, new_n13870);
and_8  g13494(new_n13870, new_n6688, new_n13871);
and_8  g13495(n10327, n4189, new_n13872);
and_8  g13496(n9920, n7456, new_n13873);
xor_4  g13497(new_n13873, new_n13872, new_n13874);
xor_4  g13498(new_n13874, new_n13871, new_n13875);
xor_4  g13499(new_n13875, new_n13869, new_n13876);
or_8   g13500(new_n13876, new_n13868, new_n13877);
not_8  g13501(new_n13867, new_n13878);
xor_4  g13502(new_n13878, new_n13860, new_n13879);
not_8  g13503(new_n13876, new_n13880);
or_8   g13504(new_n13880, new_n13879, new_n13881);
and_8  g13505(new_n13881, new_n13877, new_n13882);
and_8  g13506(new_n13882, new_n13856, new_n13883);
and_8  g13507(new_n13880, new_n13879, new_n13884);
and_8  g13508(new_n13876, new_n13868, new_n13885);
or_8   g13509(new_n13885, new_n13884, new_n13886);
and_8  g13510(new_n13886, new_n13855, new_n13887);
or_8   g13511(new_n13887, new_n13883, new_n13888);
or_8   g13512(new_n13888, new_n13854, new_n13889);
or_8   g13513(new_n13852, new_n13851, new_n13890);
or_8   g13514(new_n13849, new_n13840, new_n13891);
and_8  g13515(new_n13891, new_n13890, new_n13892);
or_8   g13516(new_n13886, new_n13855, new_n13893);
or_8   g13517(new_n13882, new_n13856, new_n13894);
and_8  g13518(new_n13894, new_n13893, new_n13895);
or_8   g13519(new_n13895, new_n13892, new_n13896);
and_8  g13520(new_n13896, new_n13889, new_n13897);
nor_6  g13521(new_n13897, new_n13785, new_n13898);
and_8  g13522(new_n13897, new_n13785, new_n13899);
or_8   g13523(new_n13899, new_n13898, new_n13900);
or_8   g13524(new_n13900, new_n13782, new_n13901);
and_8  g13525(new_n13780, new_n13771, new_n13902);
and_8  g13526(new_n13776, new_n13772, new_n13903);
or_8   g13527(new_n13903, new_n13902, new_n13904);
xor_4  g13528(new_n13897, new_n13785, new_n13905);
or_8   g13529(new_n13905, new_n13904, new_n13906);
and_8  g13530(new_n13906, new_n13901, new_n13907);
not_8  g13531(new_n6494, new_n13908);
or_8   g13532(new_n6496, new_n13908, new_n13909);
or_8   g13533(new_n6498, new_n6491, new_n13910);
and_8  g13534(new_n13910, new_n13909, new_n13911);
and_8  g13535(new_n6660, new_n6694, new_n13912);
nor_6  g13536(new_n6697, new_n13912, new_n13913);
xor_4  g13537(new_n13913, new_n13911, new_n13914);
not_8  g13538(new_n13914, new_n13915);
and_8  g13539(new_n6758, new_n6774, new_n13916);
and_8  g13540(new_n6796, new_n6776_1, new_n13917);
or_8   g13541(new_n13917, new_n13916, new_n13918);
and_8  g13542(n11023, n1094, new_n13919);
xnor_4 g13543(new_n13919, new_n13918, new_n13920);
and_8  g13544(new_n6782, new_n6777, new_n13921);
or_8   g13545(new_n6793, new_n13921, new_n13922);
not_8  g13546(new_n13922, new_n13923);
and_8  g13547(new_n6682, new_n6681, new_n13924);
and_8  g13548(new_n6690, new_n6683, new_n13925);
or_8   g13549(new_n13925, new_n13924, new_n13926);
or_8   g13550(new_n6780, new_n6779, new_n13927);
not_8  g13551(new_n6778, new_n13928);
or_8   g13552(new_n6781, new_n13928, new_n13929);
and_8  g13553(new_n13929, new_n13927, new_n13930);
or_8   g13554(new_n6789, new_n6788, new_n13931);
or_8   g13555(new_n6790, new_n6787, new_n13932);
and_8  g13556(new_n13932, new_n13931, new_n13933);
xor_4  g13557(new_n13933, new_n13930, new_n13934);
and_8  g13558(n12069, n10685, new_n13935);
and_8  g13559(n6578, n5645, new_n13936);
xor_4  g13560(new_n13936, new_n13935, new_n13937);
not_8  g13561(new_n13937, new_n13938);
nand_5 g13562(n5767, n2749, new_n13939);
and_8  g13563(n996, n159, new_n13940);
and_8  g13564(n5314, n1510, new_n13941);
xor_4  g13565(new_n13941, new_n13940, new_n13942);
xor_4  g13566(new_n13942, new_n13939, new_n13943);
xor_4  g13567(new_n13943, new_n13938, new_n13944);
xor_4  g13568(new_n13944, new_n13934, new_n13945);
nand_5 g13569(new_n6785, new_n6784, new_n13946);
or_8   g13570(new_n6791, new_n6786, new_n13947);
and_8  g13571(new_n13947, new_n13946, new_n13948);
or_8   g13572(new_n6628, new_n6663, new_n13949);
and_8  g13573(n9583, n2564, new_n13950);
and_8  g13574(n9640, n7320, new_n13951);
xor_4  g13575(new_n13951, new_n13950, new_n13952);
xor_4  g13576(new_n13952, new_n13949, new_n13953);
and_8  g13577(n1199, n1067, new_n13954);
and_8  g13578(n12247, n11153, new_n13955);
xor_4  g13579(new_n13955, new_n13954, new_n13956);
xor_4  g13580(new_n13956, new_n13953, new_n13957);
xor_4  g13581(new_n13957, new_n13948, new_n13958);
or_8   g13582(new_n13958, new_n13945, new_n13959);
xor_4  g13583(new_n13943, new_n13937, new_n13960);
xor_4  g13584(new_n13960, new_n13934, new_n13961);
not_8  g13585(new_n13956, new_n13962);
xor_4  g13586(new_n13962, new_n13953, new_n13963);
xor_4  g13587(new_n13963, new_n13948, new_n13964);
or_8   g13588(new_n13964, new_n13961, new_n13965);
and_8  g13589(new_n13965, new_n13959, new_n13966);
and_8  g13590(new_n13966, new_n13926, new_n13967);
not_8  g13591(new_n13926, new_n13968);
and_8  g13592(new_n13964, new_n13961, new_n13969);
and_8  g13593(new_n13958, new_n13945, new_n13970);
or_8   g13594(new_n13970, new_n13969, new_n13971);
and_8  g13595(new_n13971, new_n13968, new_n13972);
or_8   g13596(new_n13972, new_n13967, new_n13973);
not_8  g13597(new_n6679, new_n13974);
or_8   g13598(new_n13974, new_n6674, new_n13975);
or_8   g13599(new_n6691, new_n6680, new_n13976);
and_8  g13600(new_n13976, new_n13975, new_n13977);
or_8   g13601(new_n6677, new_n6676, new_n13978);
or_8   g13602(new_n6678, new_n6675, new_n13979);
and_8  g13603(new_n13979, new_n13978, new_n13980);
and_8  g13604(n6687, n753, new_n13981);
and_8  g13605(n2087, n1798, new_n13982);
xnor_4 g13606(new_n13982, new_n13981, new_n13983);
xor_4  g13607(new_n13983, new_n13980, new_n13984);
xor_4  g13608(new_n13984, new_n13977, new_n13985);
and_8  g13609(new_n13985, new_n13973, new_n13986);
nor_6  g13610(new_n13985, new_n13973, new_n13987);
or_8   g13611(new_n13987, new_n13986, new_n13988);
and_8  g13612(new_n13988, new_n13923, new_n13989);
xor_4  g13613(new_n13985, new_n13973, new_n13990);
and_8  g13614(new_n13990, new_n13922, new_n13991);
or_8   g13615(new_n13991, new_n13989, new_n13992);
or_8   g13616(new_n13992, new_n13920, new_n13993);
xor_4  g13617(new_n13919, new_n13918, new_n13994);
or_8   g13618(new_n13990, new_n13922, new_n13995);
or_8   g13619(new_n13988, new_n13923, new_n13996);
and_8  g13620(new_n13996, new_n13995, new_n13997);
or_8   g13621(new_n13997, new_n13994, new_n13998);
and_8  g13622(new_n13998, new_n13993, new_n13999);
and_8  g13623(new_n13999, new_n13915, new_n14000);
and_8  g13624(new_n13997, new_n13994, new_n14001);
and_8  g13625(new_n13992, new_n13920, new_n14002);
or_8   g13626(new_n14002, new_n14001, new_n14003);
and_8  g13627(new_n14003, new_n13914, new_n14004);
or_8   g13628(new_n14004, new_n14000, new_n14005);
or_8   g13629(new_n6814, new_n6816, new_n14006);
and_8  g13630(new_n6596, new_n6570, new_n14007);
and_8  g13631(new_n6617, new_n6602, new_n14008);
or_8   g13632(new_n14008, new_n14007, new_n14009);
xor_4  g13633(new_n14009, new_n14006, new_n14010);
or_8   g13634(new_n14010, new_n14005, new_n14011);
or_8   g13635(new_n14003, new_n13914, new_n14012);
or_8   g13636(new_n13999, new_n13915, new_n14013);
and_8  g13637(new_n14013, new_n14012, new_n14014);
nor_6  g13638(new_n6814, new_n6816, new_n14015);
xor_4  g13639(new_n14009, new_n14015, new_n14016);
or_8   g13640(new_n14016, new_n14014, new_n14017);
and_8  g13641(new_n14017, new_n14011, new_n14018);
or_8   g13642(new_n14018, new_n13907, new_n14019);
and_8  g13643(new_n13905, new_n13904, new_n14020);
and_8  g13644(new_n13900, new_n13782, new_n14021);
or_8   g13645(new_n14021, new_n14020, new_n14022);
and_8  g13646(new_n14016, new_n14014, new_n14023);
and_8  g13647(new_n14010, new_n14005, new_n14024);
or_8   g13648(new_n14024, new_n14023, new_n14025);
or_8   g13649(new_n14025, new_n14022, new_n14026);
and_8  g13650(new_n14026, new_n14019, new_n14027);
and_8  g13651(n11922, n4828, new_n14028);
not_8  g13652(new_n14028, new_n14029);
nor_6  g13653(new_n6857, new_n6835, new_n14030);
or_8   g13654(new_n14030, new_n6898, new_n14031);
or_8   g13655(new_n14031, new_n6862, new_n14032);
and_8  g13656(new_n6864, new_n14032, new_n14033);
or_8   g13657(new_n14033, new_n14029, new_n14034);
and_8  g13658(new_n6859, new_n6825, new_n14035);
and_8  g13659(new_n6860_1, new_n6719, new_n14036);
or_8   g13660(new_n14036, new_n14035, new_n14037);
or_8   g13661(new_n14037, new_n14028, new_n14038);
and_8  g13662(new_n14038, new_n14034, new_n14039);
nor_6  g13663(new_n14039, new_n14027, new_n14040);
and_8  g13664(new_n14039, new_n14027, new_n14041);
or_8   g13665(new_n14041, new_n14040, new_n14042);
and_8  g13666(new_n14042, new_n13770, new_n14043);
xor_4  g13667(new_n6865, new_n6618, new_n14044);
and_8  g13668(new_n6902, new_n14044, new_n14045);
or_8   g13669(new_n14045, new_n6866, new_n14046);
xor_4  g13670(new_n14039, new_n14027, new_n14047);
and_8  g13671(new_n14047, new_n14046, new_n14048);
or_8   g13672(new_n14048, new_n14043, new_n14049);
or_8   g13673(new_n14049, new_n13767, new_n14050);
not_8  g13674(new_n13767, new_n14051);
or_8   g13675(new_n14047, new_n14046, new_n14052);
or_8   g13676(new_n14042, new_n13770, new_n14053);
and_8  g13677(new_n14053, new_n14052, new_n14054);
or_8   g13678(new_n14054, new_n14051, new_n14055);
and_8  g13679(new_n14055, new_n14050, new_n14056);
xor_4  g13680(new_n14056, new_n13762, n9767);
xnor_4 g13681(new_n2094, new_n2093, n9820);
xor_4  g13682(new_n10040, new_n10037, new_n14059);
xor_4  g13683(new_n14059, new_n10036, n9938);
xor_4  g13684(new_n885, new_n884, n10476);
xnor_4 g13685(new_n882, new_n874, n10589);
xor_4  g13686(new_n1158, new_n1157, n10695);
xor_4  g13687(new_n3753, new_n3376, new_n14064);
xor_4  g13688(new_n14064, new_n3800, n10789);
xor_4  g13689(new_n3028, new_n3015, n10851);
xnor_4 g13690(new_n5174, new_n5165, n10913);
xor_4  g13691(new_n7412, new_n7622, n10949);
xnor_4 g13692(new_n11980, new_n11932, n11216);
xor_4  g13693(new_n5166, new_n5157, n11326);
and_8  g13694(new_n5792, new_n5496, new_n14071);
or_8   g13695(new_n5920, new_n14071, new_n14072);
or_8   g13696(new_n5842, new_n5840, new_n14073);
not_8  g13697(new_n5918, new_n14074);
or_8   g13698(new_n14074, new_n5845, new_n14075);
and_8  g13699(new_n14075, new_n14073, new_n14076);
and_8  g13700(new_n5835, new_n5806, new_n14077);
not_8  g13701(new_n5804, new_n14078);
or_8   g13702(new_n5674, new_n14078, new_n14079);
and_8  g13703(new_n5839, new_n14079, new_n14080);
or_8   g13704(new_n14080, new_n14077, new_n14081);
not_8  g13705(new_n5831, new_n14082);
or_8   g13706(new_n5834, new_n5828, new_n14083);
and_8  g13707(new_n14083, new_n14082, new_n14084);
and_8  g13708(n9763, n45, new_n14085);
and_8  g13709(n8759, n7823, new_n14086);
xor_4  g13710(new_n14086, new_n14085, new_n14087);
xor_4  g13711(new_n14087, new_n14084, new_n14088);
or_8   g13712(new_n5462, new_n5461, new_n14089);
or_8   g13713(new_n5463, new_n5460, new_n14090);
and_8  g13714(new_n14090, new_n14089, new_n14091);
nand_5 g13715(n9241, n9189, new_n14092);
xor_4  g13716(new_n14092, new_n14091, new_n14093);
and_8  g13717(n12705, n4634, new_n14094);
and_8  g13718(n12145, n7436, new_n14095);
xor_4  g13719(new_n14095, new_n14094, new_n14096);
and_8  g13720(n9195, n4312, new_n14097);
and_8  g13721(n10217, n6776, new_n14098);
xor_4  g13722(new_n14098, new_n14097, new_n14099);
xor_4  g13723(new_n14099, new_n14096, new_n14100);
xor_4  g13724(new_n14100, new_n14093, new_n14101);
nand_5 g13725(new_n5817, new_n5816, new_n14102);
or_8   g13726(new_n5823, new_n5818, new_n14103);
and_8  g13727(new_n14103, new_n14102, new_n14104);
or_8   g13728(new_n5812, new_n5811, new_n14105);
or_8   g13729(new_n5813, new_n5810, new_n14106);
and_8  g13730(new_n14106, new_n14105, new_n14107);
xor_4  g13731(new_n14107, new_n14104, new_n14108);
xor_4  g13732(new_n14108, new_n14101, new_n14109);
and_8  g13733(new_n5821, new_n5820, new_n14110);
or_8   g13734(new_n5821, new_n5820, new_n14111);
and_8  g13735(new_n14111, new_n5819, new_n14112);
or_8   g13736(new_n14112, new_n14110, new_n14113);
not_8  g13737(new_n14113, new_n14114);
xor_4  g13738(new_n14114, new_n14109, new_n14115);
and_8  g13739(n3986, n3342, new_n14116);
and_8  g13740(n8276, n2522, new_n14117);
and_8  g13741(n12299, n12221, new_n14118);
xor_4  g13742(new_n14118, new_n14117, new_n14119);
xor_4  g13743(new_n14119, new_n14116, new_n14120);
and_8  g13744(new_n14120, new_n14115, new_n14121);
xor_4  g13745(new_n14113, new_n14109, new_n14122);
not_8  g13746(new_n14120, new_n14123);
and_8  g13747(new_n14123, new_n14122, new_n14124);
nor_6  g13748(new_n14124, new_n14121, new_n14125);
and_8  g13749(new_n5814_1, new_n5809, new_n14126);
or_8   g13750(new_n5825, new_n14126, new_n14127);
and_8  g13751(new_n5746, new_n5897, new_n14128);
and_8  g13752(new_n5899, new_n5895, new_n14129);
or_8   g13753(new_n14129, new_n14128, new_n14130);
xor_4  g13754(new_n14130, new_n14127, new_n14131);
xor_4  g13755(new_n14131, new_n14125, new_n14132);
or_8   g13756(new_n14132, new_n14088, new_n14133);
not_8  g13757(new_n14087, new_n14134);
xor_4  g13758(new_n14134, new_n14084, new_n14135);
or_8   g13759(new_n14124, new_n14121, new_n14136);
xor_4  g13760(new_n14131, new_n14136, new_n14137);
or_8   g13761(new_n14137, new_n14135, new_n14138);
and_8  g13762(new_n14138, new_n14133, new_n14139);
and_8  g13763(new_n14139, new_n14081, new_n14140);
and_8  g13764(new_n5837, new_n5554, new_n14141);
or_8   g13765(new_n14077, new_n14141, new_n14142);
or_8   g13766(new_n14142, new_n5805, new_n14143);
and_8  g13767(new_n14143, new_n5838, new_n14144);
and_8  g13768(new_n14137, new_n14135, new_n14145);
and_8  g13769(new_n14132, new_n14088, new_n14146);
or_8   g13770(new_n14146, new_n14145, new_n14147);
and_8  g13771(new_n14147, new_n14144, new_n14148);
or_8   g13772(new_n14148, new_n14140, new_n14149);
and_8  g13773(n12025, n10223, new_n14150);
nand_5 g13774(new_n5458, new_n5457, new_n14151);
or_8   g13775(new_n5464, new_n5459, new_n14152);
and_8  g13776(new_n14152, new_n14151, new_n14153);
xor_4  g13777(new_n14153, new_n14150, new_n14154);
or_8   g13778(new_n14154, new_n14149, new_n14155);
or_8   g13779(new_n14147, new_n14144, new_n14156);
or_8   g13780(new_n14139, new_n14081, new_n14157);
and_8  g13781(new_n14157, new_n14156, new_n14158);
not_8  g13782(new_n14154, new_n14159);
or_8   g13783(new_n14159, new_n14158, new_n14160);
and_8  g13784(new_n14160, new_n14155, new_n14161);
nand_5 g13785(new_n5884, new_n5879, new_n14162);
not_8  g13786(new_n5885, new_n14163);
or_8   g13787(new_n5894, new_n14163, new_n14164);
and_8  g13788(new_n14164, new_n14162, new_n14165);
and_8  g13789(n7690, n5579, new_n14166);
and_8  g13790(n7388, n2507, new_n14167);
xor_4  g13791(new_n14167, new_n14166, new_n14168);
and_8  g13792(n7270, n2393, new_n14169);
and_8  g13793(n5331, n1576, new_n14170);
xor_4  g13794(new_n14170, new_n14169, new_n14171);
xor_4  g13795(new_n14171, new_n14168, new_n14172);
and_8  g13796(n3616, n2498, new_n14173);
and_8  g13797(n12648, n6016, new_n14174);
xor_4  g13798(new_n14174, new_n14173, new_n14175);
xor_4  g13799(new_n14175, new_n14172, new_n14176);
and_8  g13800(n5798, n2530, new_n14177);
and_8  g13801(n10644, n7946, new_n14178);
xor_4  g13802(new_n14178, new_n14177, new_n14179);
or_8   g13803(new_n5882, new_n5881, new_n14180);
or_8   g13804(new_n5883, new_n5880, new_n14181);
and_8  g13805(new_n14181, new_n14180, new_n14182);
or_8   g13806(new_n5453, new_n5452, new_n14183);
or_8   g13807(new_n5454, new_n5451, new_n14184);
and_8  g13808(new_n14184, new_n14183, new_n14185);
xor_4  g13809(new_n14185, new_n14182, new_n14186);
xor_4  g13810(new_n14186, new_n14179, new_n14187);
xor_4  g13811(new_n14187, new_n14176, new_n14188);
xor_4  g13812(new_n14188, new_n14165, new_n14189);
and_8  g13813(new_n5709, new_n5869, new_n14190);
and_8  g13814(new_n5871, new_n5867, new_n14191);
nor_6  g13815(new_n14191, new_n14190, new_n14192);
or_8   g13816(new_n5891, new_n5890, new_n14193);
or_8   g13817(new_n5892, new_n5889, new_n14194);
and_8  g13818(new_n14194, new_n14193, new_n14195);
and_8  g13819(new_n5887, new_n5886, new_n14196);
nor_6  g13820(new_n5893, new_n5888, new_n14197);
or_8   g13821(new_n14197, new_n14196, new_n14198);
and_8  g13822(n7965, n6431, new_n14199);
and_8  g13823(n9111, n5857, new_n14200);
xor_4  g13824(new_n14200, new_n14199, new_n14201);
and_8  g13825(n11892, n5153, new_n14202);
and_8  g13826(n5860, n806, new_n14203);
xor_4  g13827(new_n14203, new_n14202, new_n14204);
and_8  g13828(n10545, n521, new_n14205);
and_8  g13829(n10547, n7265, new_n14206);
xor_4  g13830(new_n14206, new_n14205, new_n14207);
xnor_4 g13831(new_n14207, new_n14204, new_n14208);
xor_4  g13832(new_n14208, new_n14201, new_n14209);
xor_4  g13833(new_n14209, new_n14198, new_n14210);
xor_4  g13834(new_n14210, new_n14195, new_n14211);
xor_4  g13835(new_n14211, new_n14192, new_n14212);
and_8  g13836(new_n5455, new_n5450, new_n14213);
and_8  g13837(new_n5465, new_n5456, new_n14214);
or_8   g13838(new_n14214, new_n14213, new_n14215);
nand_5 g13839(new_n5856, new_n5855, new_n14216);
or_8   g13840(new_n5862, new_n5857_1, new_n14217);
nand_5 g13841(new_n14217, new_n14216, new_n14218);
xor_4  g13842(new_n14218, new_n14215, new_n14219);
xor_4  g13843(new_n14219, new_n14212, new_n14220);
xor_4  g13844(new_n14220, new_n14189, new_n14221);
not_8  g13845(new_n5846, new_n14222);
and_8  g13846(new_n5872, new_n14222, new_n14223);
nor_6  g13847(new_n5908, new_n14223, new_n14224);
and_8  g13848(new_n5471, new_n5470, new_n14225);
or_8   g13849(new_n5474, new_n14225, new_n14226);
not_8  g13850(new_n5851, new_n14227);
or_8   g13851(new_n5853, new_n14227, new_n14228);
and_8  g13852(new_n5864, new_n14228, new_n14229);
not_8  g13853(new_n14229, new_n14230);
or_8   g13854(new_n5860_1, new_n5859, new_n14231);
or_8   g13855(new_n5861, new_n5858, new_n14232);
and_8  g13856(new_n14232, new_n14231, new_n14233);
and_8  g13857(n4499, n2558, new_n14234);
and_8  g13858(n5305, n2512, new_n14235);
xor_4  g13859(new_n14235, new_n14234, new_n14236);
xor_4  g13860(new_n14236, new_n14233, new_n14237);
or_8   g13861(new_n5850, new_n5847, new_n14238);
and_8  g13862(new_n14238, new_n5848, new_n14239);
and_8  g13863(n8476, n2347, new_n14240);
and_8  g13864(new_n14240, new_n14239, new_n14241);
and_8  g13865(new_n14240, new_n5716, new_n14242);
nor_6  g13866(new_n14242, new_n14239, new_n14243);
or_8   g13867(new_n14243, new_n14241, new_n14244);
and_8  g13868(n2253, n1097, new_n14245);
and_8  g13869(n5964, n3865, new_n14246);
xor_4  g13870(new_n14246, new_n14245, new_n14247);
xor_4  g13871(new_n14247, new_n14244, new_n14248);
xor_4  g13872(new_n14248, new_n14237, new_n14249);
xor_4  g13873(new_n14249, new_n14230, new_n14250);
and_8  g13874(n10510, n2024, new_n14251);
and_8  g13875(n11257, n2879, new_n14252);
xor_4  g13876(new_n14252, new_n14251, new_n14253);
not_8  g13877(new_n14253, new_n14254);
xor_4  g13878(new_n14254, new_n14250, new_n14255);
xor_4  g13879(new_n14255, new_n14226, new_n14256);
xor_4  g13880(new_n14256, new_n14224, new_n14257);
and_8  g13881(new_n14257, new_n14221, new_n14258);
not_8  g13882(new_n14189, new_n14259);
xor_4  g13883(new_n14220, new_n14259, new_n14260);
or_8   g13884(new_n5908, new_n14223, new_n14261);
xor_4  g13885(new_n14256, new_n14261, new_n14262);
and_8  g13886(new_n14262, new_n14260, new_n14263);
or_8   g13887(new_n14263, new_n14258, new_n14264);
or_8   g13888(new_n14264, new_n14161, new_n14265);
and_8  g13889(new_n14159, new_n14158, new_n14266);
and_8  g13890(new_n14154, new_n14149, new_n14267);
or_8   g13891(new_n14267, new_n14266, new_n14268);
or_8   g13892(new_n14262, new_n14260, new_n14269);
or_8   g13893(new_n14257, new_n14221, new_n14270);
and_8  g13894(new_n14270, new_n14269, new_n14271);
or_8   g13895(new_n14271, new_n14268, new_n14272);
and_8  g13896(new_n14272, new_n14265, new_n14273);
or_8   g13897(new_n5905, new_n5877, new_n14274);
or_8   g13898(new_n5915, new_n5914, new_n14275);
and_8  g13899(new_n14275, new_n14274, new_n14276);
or_8   g13900(new_n5478, new_n5446, new_n14277);
or_8   g13901(new_n5476, new_n5447, new_n14278);
and_8  g13902(new_n14278, new_n14277, new_n14279);
and_8  g13903(new_n5499, new_n5497, new_n14280);
or_8   g13904(new_n14280, new_n5490, new_n14281);
and_8  g13905(new_n14281, new_n14279, new_n14282);
or_8   g13906(new_n14282, new_n5479, new_n14283);
and_8  g13907(new_n5900, new_n5754, new_n14284);
or_8   g13908(new_n5911, new_n14284, new_n14285);
or_8   g13909(new_n14285, new_n14283, new_n14286);
or_8   g13910(new_n5494, new_n5480, new_n14287);
and_8  g13911(new_n14287, new_n14278, new_n14288);
not_8  g13912(new_n14285, new_n14289);
or_8   g13913(new_n14289, new_n14288, new_n14290);
and_8  g13914(new_n14290, new_n14286, new_n14291);
xor_4  g13915(new_n14291, new_n14276, new_n14292);
and_8  g13916(new_n14292, new_n14273, new_n14293);
and_8  g13917(new_n14271, new_n14268, new_n14294);
and_8  g13918(new_n14264, new_n14161, new_n14295);
or_8   g13919(new_n14295, new_n14294, new_n14296);
and_8  g13920(new_n14291, new_n14276, new_n14297);
nor_6  g13921(new_n14291, new_n14276, new_n14298);
or_8   g13922(new_n14298, new_n14297, new_n14299);
and_8  g13923(new_n14299, new_n14296, new_n14300);
or_8   g13924(new_n14300, new_n14293, new_n14301);
or_8   g13925(new_n14301, new_n14076, new_n14302);
nor_6  g13926(new_n14074, new_n5845, new_n14303);
or_8   g13927(new_n14303, new_n5844, new_n14304);
or_8   g13928(new_n14299, new_n14296, new_n14305);
or_8   g13929(new_n14292, new_n14273, new_n14306);
and_8  g13930(new_n14306, new_n14305, new_n14307);
or_8   g13931(new_n14307, new_n14304, new_n14308);
and_8  g13932(new_n14308, new_n14302, new_n14309);
xor_4  g13933(new_n14309, new_n14072, n11707);
xnor_4 g13934(new_n6399, new_n6398, n11755);
xor_4  g13935(new_n3793, new_n3792, n11780);
xor_4  g13936(new_n10451_1, new_n10438, n11919);
xor_4  g13937(new_n10453, new_n10446, n12005);
xnor_4 g13938(new_n10926, new_n10923, n12014);
xor_4  g13939(new_n9122, new_n9084, n12020);
xnor_4 g13940(new_n11973, new_n11944, n12076);
xor_4  g13941(new_n12558, new_n12557, n12111);
nor_6  g13942(new_n10928_1, new_n10911, new_n14319);
or_8   g13943(new_n14319, new_n10929, n12444);
xor_4  g13944(new_n5798_1, new_n5781, n12807);
endmodule


