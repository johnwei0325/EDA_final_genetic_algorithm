// Benchmark "top_809568696_809776567_809698999_863110837_1234615" written by ABC on Thu Jun 27 01:36:09 2024

module top_809568696_809776567_809698999_863110837_1234615 ( 
    n74, n203, n271, n394, n411, n427, n462, n498, n650, n656, n666, n674,
    n702, n730, n737, n760, n844, n977, n1027, n1093, n1222, n1265, n1268,
    n1347, n1568, n1637, n1702, n1763, n1776, n2048, n2061, n2164, n2166,
    n2201, n2334, n2454, n2573, n2615, n2674, n2699, n2895, n3130, n3166,
    n3263, n3367, n3388, n3506, n3532, n3652, n3655, n3673, n3775, n3799,
    n3804, n3833, n3893, n3910, n3972, n4000, n4022, n4039, n4117, n4131,
    n4147, n4154, n4172, n4175, n4225, n4282, n4292, n4615, n4659, n4755,
    n4774, n4785, n4895, n4907, n5009, n5014, n5023, n5033, n5046, n5077,
    n5184, n5185, n5225, n5430, n5449, n5467, n5502, n5601, n5725, n5786,
    n5943, n5950, n5960, n6007, n6054, n6114, n6147, n6251, n6258, n6270,
    n6362, n6436, n6460, n6480, n6517, n6555, n6586, n6680, n6693, n6703,
    n6758, n6791, n6810, n6873, n6946, n6999, n7104, n7272, n7282, n7354,
    n7450, n7652, n7667, n7748, n7832, n7941, n7972, n7988, n8002, n8044,
    n8073, n8204, n8262, n8302, n8315, n8397, n8439, n8463, n8486, n8550,
    n8552, n8598, n8635, n8649, n8737, n8746, n8780, n8799, n8800, n8873,
    n8892, n8926, n8997, n9026, n9110, n9154, n9186, n9252, n9314, n9543,
    n9544, n9555, n9589, n9830, n9893, n9921, n9936, n9977, n10050, n10051,
    n10061, n10080, n10112, n10147, n10255, n10278, n10283, n10378, n10407,
    n10426, n10446, n10466, n10470, n10573, n10615, n10630, n10736, n10750,
    n10765, n10862, n10912, n10945, n11143, n11158, n11269, n11345, n11404,
    n11529, n11590, n11605, n11666, n11756, n11776, n11842, n11854, n11875,
    n11902, n11930, n11933, n11961, n12009, n12012, n12025, n12142, n12218,
    n12270, n12321, n12336, n12573, n12614, n12782, n12829, n12885, n12927,
    n12976, n13000, n13093, n13102, n13109, n13186, n13224, n13231, n13295,
    n13363, n13364, n13509, n13511, n13561, n13625, n13636, n13814, n13882,
    n13890, n13944, n13992, n14072, n14163, n14293, n14303, n14408, n14464,
    n14475, n14483,
    n8, n46, n91, n126, n278, n389, n451, n490, n543, n682, n884, n948,
    n1094, n1122, n1124, n1329, n1545, n1739, n1827, n1900, n1927, n1951,
    n2027, n2126, n2175, n2223, n2311, n2407, n2556, n2559, n2572, n2672,
    n2734, n3090, n3242, n3340, n3603, n3854, n3901, n4125, n4279, n4305,
    n4345, n4437, n4541, n4604, n4672, n4858, n4971, n5479, n5550, n5586,
    n5806, n5851, n5987, n6012, n6198, n6275, n6314, n6682, n6696, n6786,
    n6853, n6952, n6979, n7071, n7073, n7132, n7152, n7246, n7265, n7382,
    n7655, n7771, n7825, n8068, n8085, n8124, n8144, n8215, n8306, n8471,
    n8604, n8909, n9096, n9342, n9437, n9447, n9570, n9665, n9717, n10515,
    n10591, n10791, n10802, n10915, n11122, n11393, n11463, n11534, n11627,
    n11664, n11822, n11847, n12032, n12166, n12232, n12355, n12535, n12989,
    n13010, n13045, n13114, n13141, n13316, n13577, n13639, n13658, n13693,
    n13760, n13853, n13870, n13953, n13959, n14289, n14307, n14330, n14399,
    n14463  );
  input  n74, n203, n271, n394, n411, n427, n462, n498, n650, n656, n666,
    n674, n702, n730, n737, n760, n844, n977, n1027, n1093, n1222, n1265,
    n1268, n1347, n1568, n1637, n1702, n1763, n1776, n2048, n2061, n2164,
    n2166, n2201, n2334, n2454, n2573, n2615, n2674, n2699, n2895, n3130,
    n3166, n3263, n3367, n3388, n3506, n3532, n3652, n3655, n3673, n3775,
    n3799, n3804, n3833, n3893, n3910, n3972, n4000, n4022, n4039, n4117,
    n4131, n4147, n4154, n4172, n4175, n4225, n4282, n4292, n4615, n4659,
    n4755, n4774, n4785, n4895, n4907, n5009, n5014, n5023, n5033, n5046,
    n5077, n5184, n5185, n5225, n5430, n5449, n5467, n5502, n5601, n5725,
    n5786, n5943, n5950, n5960, n6007, n6054, n6114, n6147, n6251, n6258,
    n6270, n6362, n6436, n6460, n6480, n6517, n6555, n6586, n6680, n6693,
    n6703, n6758, n6791, n6810, n6873, n6946, n6999, n7104, n7272, n7282,
    n7354, n7450, n7652, n7667, n7748, n7832, n7941, n7972, n7988, n8002,
    n8044, n8073, n8204, n8262, n8302, n8315, n8397, n8439, n8463, n8486,
    n8550, n8552, n8598, n8635, n8649, n8737, n8746, n8780, n8799, n8800,
    n8873, n8892, n8926, n8997, n9026, n9110, n9154, n9186, n9252, n9314,
    n9543, n9544, n9555, n9589, n9830, n9893, n9921, n9936, n9977, n10050,
    n10051, n10061, n10080, n10112, n10147, n10255, n10278, n10283, n10378,
    n10407, n10426, n10446, n10466, n10470, n10573, n10615, n10630, n10736,
    n10750, n10765, n10862, n10912, n10945, n11143, n11158, n11269, n11345,
    n11404, n11529, n11590, n11605, n11666, n11756, n11776, n11842, n11854,
    n11875, n11902, n11930, n11933, n11961, n12009, n12012, n12025, n12142,
    n12218, n12270, n12321, n12336, n12573, n12614, n12782, n12829, n12885,
    n12927, n12976, n13000, n13093, n13102, n13109, n13186, n13224, n13231,
    n13295, n13363, n13364, n13509, n13511, n13561, n13625, n13636, n13814,
    n13882, n13890, n13944, n13992, n14072, n14163, n14293, n14303, n14408,
    n14464, n14475, n14483;
  output n8, n46, n91, n126, n278, n389, n451, n490, n543, n682, n884, n948,
    n1094, n1122, n1124, n1329, n1545, n1739, n1827, n1900, n1927, n1951,
    n2027, n2126, n2175, n2223, n2311, n2407, n2556, n2559, n2572, n2672,
    n2734, n3090, n3242, n3340, n3603, n3854, n3901, n4125, n4279, n4305,
    n4345, n4437, n4541, n4604, n4672, n4858, n4971, n5479, n5550, n5586,
    n5806, n5851, n5987, n6012, n6198, n6275, n6314, n6682, n6696, n6786,
    n6853, n6952, n6979, n7071, n7073, n7132, n7152, n7246, n7265, n7382,
    n7655, n7771, n7825, n8068, n8085, n8124, n8144, n8215, n8306, n8471,
    n8604, n8909, n9096, n9342, n9437, n9447, n9570, n9665, n9717, n10515,
    n10591, n10791, n10802, n10915, n11122, n11393, n11463, n11534, n11627,
    n11664, n11822, n11847, n12032, n12166, n12232, n12355, n12535, n12989,
    n13010, n13045, n13114, n13141, n13316, n13577, n13639, n13658, n13693,
    n13760, n13853, n13870, n13953, n13959, n14289, n14307, n14330, n14399,
    n14463;
  wire new_n386, new_n387, new_n388, new_n389_1, new_n390, new_n391,
    new_n392, new_n393, new_n394_1, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411_1, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427_1, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451_1, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462_1, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490_1, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543_1, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650_1,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656_1, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666_1, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674_1, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682_1, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702_1, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730_1, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737_1, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760_1, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884_1, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948_1, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977_1, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027_1, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093_1, new_n1094_1, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122_1, new_n1123, new_n1124_1, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222_1, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265_1, new_n1266,
    new_n1267, new_n1268_1, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329_1, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347_1, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545_1, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568_1,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637_1, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702_1, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739_1, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763_1, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776_1, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827_1, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900_1, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927_1, new_n1928, new_n1929,
    new_n1931, new_n1932, new_n1933, new_n1934, new_n1935, new_n1936,
    new_n1937, new_n1938, new_n1939, new_n1940, new_n1941, new_n1942,
    new_n1943, new_n1944, new_n1945, new_n1946, new_n1947, new_n1948,
    new_n1949, new_n1950, new_n1951_1, new_n1952, new_n1953, new_n1954,
    new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960,
    new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966,
    new_n1967, new_n1968, new_n1969, new_n1970, new_n1971, new_n1972,
    new_n1973, new_n1974, new_n1975, new_n1976, new_n1977, new_n1978,
    new_n1979, new_n1980, new_n1981, new_n1982, new_n1983, new_n1984,
    new_n1985, new_n1986, new_n1987, new_n1988, new_n1989, new_n1990,
    new_n1991, new_n1992, new_n1993, new_n1994, new_n1995, new_n1996,
    new_n1997, new_n1998, new_n1999, new_n2000, new_n2001, new_n2002,
    new_n2003, new_n2004, new_n2005, new_n2006, new_n2007, new_n2008,
    new_n2009, new_n2010, new_n2011, new_n2012, new_n2013, new_n2014,
    new_n2015, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027_1,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2043, new_n2044, new_n2045,
    new_n2046, new_n2047, new_n2048_1, new_n2049, new_n2050, new_n2051,
    new_n2052, new_n2053, new_n2054, new_n2055, new_n2056, new_n2057,
    new_n2058, new_n2059, new_n2060, new_n2061_1, new_n2062, new_n2063,
    new_n2064, new_n2065, new_n2066, new_n2067, new_n2068, new_n2069,
    new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075,
    new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081,
    new_n2082, new_n2083, new_n2084, new_n2085, new_n2086, new_n2087,
    new_n2088, new_n2089, new_n2090, new_n2091, new_n2092, new_n2093,
    new_n2094, new_n2095, new_n2096, new_n2097, new_n2098, new_n2099,
    new_n2100, new_n2101, new_n2102, new_n2103, new_n2104, new_n2105,
    new_n2106, new_n2107, new_n2108, new_n2109, new_n2110, new_n2111,
    new_n2112, new_n2113, new_n2114, new_n2115, new_n2116, new_n2117,
    new_n2118, new_n2119, new_n2120, new_n2121, new_n2122, new_n2123,
    new_n2124, new_n2125, new_n2126_1, new_n2127, new_n2128, new_n2129,
    new_n2130, new_n2131, new_n2132, new_n2133, new_n2134, new_n2135,
    new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2141,
    new_n2142, new_n2143, new_n2144, new_n2145, new_n2146, new_n2147,
    new_n2148, new_n2149, new_n2150, new_n2151, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164_1, new_n2165, new_n2166_1,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175_1, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201_1, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223_1, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311_1,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334_1, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407_1, new_n2408,
    new_n2409, new_n2410, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454_1, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2498, new_n2499, new_n2500,
    new_n2501, new_n2502, new_n2503, new_n2504, new_n2505, new_n2506,
    new_n2507, new_n2508, new_n2509, new_n2510, new_n2511, new_n2512,
    new_n2513, new_n2514, new_n2515, new_n2516, new_n2517, new_n2518,
    new_n2519, new_n2520, new_n2521, new_n2522, new_n2523, new_n2524,
    new_n2525, new_n2526, new_n2527, new_n2528, new_n2529, new_n2530,
    new_n2531, new_n2532, new_n2533, new_n2534, new_n2535, new_n2536,
    new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2553, new_n2554,
    new_n2555, new_n2556_1, new_n2557, new_n2558, new_n2559_1, new_n2560,
    new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572_1,
    new_n2573_1, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615_1,
    new_n2616, new_n2617, new_n2618, new_n2619, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659, new_n2660, new_n2661, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2671, new_n2672_1, new_n2673, new_n2674_1, new_n2675, new_n2676,
    new_n2677, new_n2678, new_n2679, new_n2680, new_n2681, new_n2682,
    new_n2683, new_n2684, new_n2685, new_n2686, new_n2687, new_n2688,
    new_n2689, new_n2690, new_n2691, new_n2692, new_n2693, new_n2694,
    new_n2695, new_n2696, new_n2697, new_n2698, new_n2699_1, new_n2700,
    new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706,
    new_n2707, new_n2708, new_n2709, new_n2710, new_n2711, new_n2712,
    new_n2713, new_n2714, new_n2715, new_n2716, new_n2717, new_n2718,
    new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730,
    new_n2731, new_n2732, new_n2733, new_n2734_1, new_n2735, new_n2736,
    new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742,
    new_n2743, new_n2744, new_n2745, new_n2746, new_n2747, new_n2748,
    new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2759, new_n2760, new_n2761,
    new_n2762, new_n2763, new_n2764, new_n2765, new_n2766, new_n2767,
    new_n2768, new_n2769, new_n2770, new_n2771, new_n2772, new_n2773,
    new_n2774, new_n2775, new_n2776, new_n2777, new_n2778, new_n2779,
    new_n2780, new_n2781, new_n2782, new_n2783, new_n2784, new_n2785,
    new_n2786, new_n2787, new_n2788, new_n2789, new_n2790, new_n2791,
    new_n2792, new_n2793, new_n2794, new_n2795, new_n2796, new_n2797,
    new_n2798, new_n2799, new_n2800, new_n2801, new_n2802, new_n2803,
    new_n2804, new_n2805, new_n2806, new_n2807, new_n2808, new_n2809,
    new_n2810, new_n2811, new_n2812, new_n2813, new_n2814, new_n2815,
    new_n2816, new_n2817, new_n2818, new_n2819, new_n2820, new_n2821,
    new_n2822, new_n2823, new_n2824, new_n2825, new_n2826, new_n2827,
    new_n2828, new_n2829, new_n2830, new_n2831, new_n2832, new_n2833,
    new_n2834, new_n2835, new_n2836, new_n2837, new_n2838, new_n2839,
    new_n2840, new_n2841, new_n2842, new_n2843, new_n2844, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895_1, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2932, new_n2933, new_n2934, new_n2935, new_n2936, new_n2937,
    new_n2938, new_n2939, new_n2940, new_n2941, new_n2942, new_n2943,
    new_n2944, new_n2945, new_n2946, new_n2947, new_n2948, new_n2949,
    new_n2950, new_n2951, new_n2952, new_n2953, new_n2954, new_n2955,
    new_n2956, new_n2957, new_n2958, new_n2959, new_n2960, new_n2961,
    new_n2962, new_n2963, new_n2964, new_n2965, new_n2966, new_n2967,
    new_n2968, new_n2969, new_n2970, new_n2971, new_n2972, new_n2973,
    new_n2974, new_n2975, new_n2976, new_n2977, new_n2978, new_n2979,
    new_n2980, new_n2981, new_n2982, new_n2983, new_n2984, new_n2985,
    new_n2986, new_n2987, new_n2988, new_n2989, new_n2990, new_n2991,
    new_n2992, new_n2993, new_n2994, new_n2995, new_n2996, new_n2997,
    new_n2998, new_n2999, new_n3000, new_n3001, new_n3002, new_n3003,
    new_n3004, new_n3005, new_n3006, new_n3007, new_n3008, new_n3009,
    new_n3010, new_n3011, new_n3012, new_n3013, new_n3014, new_n3015,
    new_n3016, new_n3017, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090_1, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3105, new_n3106, new_n3107,
    new_n3108, new_n3109, new_n3110, new_n3111, new_n3112, new_n3113,
    new_n3114, new_n3115, new_n3116, new_n3117, new_n3118, new_n3119,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130_1, new_n3131,
    new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137,
    new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155,
    new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166_1, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242_1, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260, new_n3261, new_n3262, new_n3263_1, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3367_1, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388_1, new_n3389, new_n3390, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3453,
    new_n3454, new_n3455, new_n3456, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506_1, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532_1, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3540, new_n3541, new_n3542, new_n3543, new_n3544,
    new_n3545, new_n3546, new_n3547, new_n3548, new_n3549, new_n3550,
    new_n3551, new_n3552, new_n3553, new_n3554, new_n3555, new_n3556,
    new_n3557, new_n3558, new_n3559, new_n3560, new_n3561, new_n3562,
    new_n3563, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568,
    new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603_1, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3626, new_n3627, new_n3628, new_n3629,
    new_n3630, new_n3631, new_n3632, new_n3633, new_n3634, new_n3635,
    new_n3636, new_n3637, new_n3638, new_n3639, new_n3640, new_n3641,
    new_n3642, new_n3643, new_n3644, new_n3645, new_n3646, new_n3647,
    new_n3648, new_n3649, new_n3650, new_n3651, new_n3652_1, new_n3653,
    new_n3654, new_n3655_1, new_n3656, new_n3657, new_n3658, new_n3659,
    new_n3660, new_n3661, new_n3662, new_n3663, new_n3664, new_n3665,
    new_n3666, new_n3667, new_n3668, new_n3669, new_n3670, new_n3671,
    new_n3672, new_n3673_1, new_n3674, new_n3675, new_n3676, new_n3677,
    new_n3678, new_n3679, new_n3680, new_n3681, new_n3682, new_n3683,
    new_n3684, new_n3685, new_n3686, new_n3687, new_n3688, new_n3689,
    new_n3690, new_n3691, new_n3692, new_n3693, new_n3694, new_n3695,
    new_n3696, new_n3697, new_n3698, new_n3699, new_n3700, new_n3701,
    new_n3702, new_n3703, new_n3704, new_n3705, new_n3706, new_n3707,
    new_n3708, new_n3709, new_n3710, new_n3711, new_n3713, new_n3714,
    new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720,
    new_n3721, new_n3722, new_n3723, new_n3724, new_n3725, new_n3726,
    new_n3727, new_n3728, new_n3729, new_n3730, new_n3731, new_n3732,
    new_n3733, new_n3734, new_n3735, new_n3736, new_n3737, new_n3738,
    new_n3739, new_n3740, new_n3741, new_n3742, new_n3743, new_n3744,
    new_n3745, new_n3746, new_n3747, new_n3748, new_n3749, new_n3750,
    new_n3751, new_n3752, new_n3753, new_n3754, new_n3755, new_n3756,
    new_n3757, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762,
    new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768,
    new_n3769, new_n3770, new_n3771, new_n3772, new_n3773, new_n3774,
    new_n3775_1, new_n3776, new_n3777, new_n3778, new_n3779, new_n3780,
    new_n3781, new_n3782, new_n3783, new_n3784, new_n3785, new_n3786,
    new_n3787, new_n3788, new_n3789, new_n3790, new_n3791, new_n3792,
    new_n3793, new_n3794, new_n3795, new_n3796, new_n3797, new_n3798,
    new_n3800, new_n3801, new_n3802, new_n3803, new_n3804_1, new_n3805,
    new_n3806, new_n3807, new_n3808, new_n3809, new_n3810, new_n3811,
    new_n3812, new_n3813, new_n3814, new_n3815, new_n3816, new_n3817,
    new_n3818, new_n3819, new_n3820, new_n3821, new_n3822, new_n3823,
    new_n3824, new_n3825, new_n3826, new_n3827, new_n3828, new_n3829,
    new_n3830, new_n3831, new_n3832, new_n3833_1, new_n3834, new_n3835,
    new_n3836, new_n3837, new_n3838, new_n3839, new_n3840, new_n3841,
    new_n3842, new_n3843, new_n3844, new_n3845, new_n3846, new_n3847,
    new_n3848, new_n3849, new_n3850, new_n3851, new_n3852, new_n3853,
    new_n3854_1, new_n3855, new_n3856, new_n3857, new_n3858, new_n3859,
    new_n3860, new_n3861, new_n3862, new_n3863, new_n3864, new_n3865,
    new_n3866, new_n3867, new_n3868, new_n3869, new_n3870, new_n3871,
    new_n3872, new_n3873, new_n3874, new_n3875, new_n3876, new_n3877,
    new_n3878, new_n3879, new_n3880, new_n3881, new_n3882, new_n3883,
    new_n3884, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891, new_n3892, new_n3893_1, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901_1, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909, new_n3910_1, new_n3911, new_n3912, new_n3913, new_n3914,
    new_n3915, new_n3916, new_n3917, new_n3918, new_n3919, new_n3920,
    new_n3921, new_n3922, new_n3923, new_n3924, new_n3925, new_n3926,
    new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932,
    new_n3933, new_n3934, new_n3935, new_n3936, new_n3937, new_n3938,
    new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944,
    new_n3945, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950,
    new_n3951, new_n3952, new_n3953, new_n3954, new_n3955, new_n3956,
    new_n3957, new_n3958, new_n3959, new_n3960, new_n3961, new_n3962,
    new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968,
    new_n3969, new_n3970, new_n3971, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000_1, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022_1, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039_1, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117_1, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125_1, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131_1, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4146, new_n4147_1, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154_1, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172_1, new_n4173, new_n4174, new_n4175_1,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187,
    new_n4188, new_n4189, new_n4190, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4211,
    new_n4212, new_n4213, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225_1, new_n4226, new_n4227, new_n4228, new_n4229,
    new_n4230, new_n4231, new_n4232, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279_1, new_n4280, new_n4281, new_n4282_1, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292_1, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305_1, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325, new_n4326, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345_1,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374, new_n4375,
    new_n4376, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401, new_n4402, new_n4403, new_n4404, new_n4406,
    new_n4407, new_n4408, new_n4409, new_n4410, new_n4411, new_n4412,
    new_n4413, new_n4414, new_n4415, new_n4416, new_n4417, new_n4418,
    new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424,
    new_n4425, new_n4426, new_n4427, new_n4428, new_n4429, new_n4430,
    new_n4431, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437_1, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4494, new_n4495, new_n4496, new_n4497,
    new_n4498, new_n4499, new_n4500, new_n4501, new_n4502, new_n4503,
    new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509,
    new_n4510, new_n4511, new_n4512, new_n4513, new_n4514, new_n4515,
    new_n4516, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521,
    new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527,
    new_n4528, new_n4529, new_n4530, new_n4531, new_n4532, new_n4533,
    new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539,
    new_n4540, new_n4541_1, new_n4542, new_n4543, new_n4544, new_n4545,
    new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551,
    new_n4552, new_n4553, new_n4554, new_n4555, new_n4557, new_n4558,
    new_n4559, new_n4560, new_n4561, new_n4562, new_n4563, new_n4564,
    new_n4565, new_n4566, new_n4567, new_n4568, new_n4569, new_n4570,
    new_n4571, new_n4572, new_n4573, new_n4574, new_n4575, new_n4576,
    new_n4577, new_n4578, new_n4579, new_n4580, new_n4581, new_n4582,
    new_n4583, new_n4584, new_n4585, new_n4586, new_n4587, new_n4588,
    new_n4589, new_n4590, new_n4591, new_n4592, new_n4593, new_n4594,
    new_n4595, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604_1, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615_1, new_n4616, new_n4617, new_n4618,
    new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624,
    new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630,
    new_n4631, new_n4632, new_n4633, new_n4634, new_n4635, new_n4636,
    new_n4637, new_n4638, new_n4639, new_n4640, new_n4641, new_n4642,
    new_n4643, new_n4645, new_n4646, new_n4647, new_n4648, new_n4649,
    new_n4650, new_n4651, new_n4652, new_n4653, new_n4654, new_n4655,
    new_n4656, new_n4657, new_n4658, new_n4659_1, new_n4660, new_n4661,
    new_n4662, new_n4663, new_n4664, new_n4665, new_n4666, new_n4667,
    new_n4668, new_n4669, new_n4670, new_n4671, new_n4672_1, new_n4673,
    new_n4674, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686, new_n4687, new_n4688, new_n4689, new_n4690, new_n4691,
    new_n4692, new_n4693, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703,
    new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709,
    new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715,
    new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721,
    new_n4722, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727,
    new_n4728, new_n4729, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755_1, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774_1, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785_1, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4817, new_n4818, new_n4819,
    new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825,
    new_n4826, new_n4827, new_n4828, new_n4829, new_n4830, new_n4831,
    new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837,
    new_n4838, new_n4839, new_n4840, new_n4841, new_n4842, new_n4843,
    new_n4844, new_n4845, new_n4846, new_n4847, new_n4848, new_n4849,
    new_n4850, new_n4851, new_n4852, new_n4853, new_n4854, new_n4855,
    new_n4856, new_n4857, new_n4858_1, new_n4859, new_n4860, new_n4861,
    new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867,
    new_n4868, new_n4869, new_n4870, new_n4871, new_n4872, new_n4873,
    new_n4874, new_n4875, new_n4876, new_n4877, new_n4878, new_n4879,
    new_n4880, new_n4881, new_n4882, new_n4883, new_n4884, new_n4885,
    new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891,
    new_n4892, new_n4893, new_n4894, new_n4895_1, new_n4896, new_n4897,
    new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903,
    new_n4905, new_n4906, new_n4907_1, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938, new_n4939, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971_1, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009_1, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014_1, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023_1, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031,
    new_n5032, new_n5033_1, new_n5034, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046_1, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184_1, new_n5185_1, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211, new_n5212, new_n5213,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5218, new_n5219,
    new_n5220, new_n5221, new_n5222, new_n5223, new_n5224, new_n5225_1,
    new_n5226, new_n5227, new_n5228, new_n5229, new_n5230, new_n5231,
    new_n5232, new_n5233, new_n5234, new_n5235, new_n5236, new_n5237,
    new_n5238, new_n5239, new_n5240, new_n5241, new_n5242, new_n5243,
    new_n5244, new_n5245, new_n5246, new_n5247, new_n5248, new_n5249,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255, new_n5256,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273, new_n5274,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300, new_n5301, new_n5302, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337, new_n5339, new_n5340, new_n5341,
    new_n5342, new_n5343, new_n5344, new_n5345, new_n5346, new_n5347,
    new_n5348, new_n5349, new_n5350, new_n5351, new_n5352, new_n5353,
    new_n5354, new_n5355, new_n5356, new_n5357, new_n5358, new_n5359,
    new_n5360, new_n5361, new_n5362, new_n5363, new_n5364, new_n5365,
    new_n5366, new_n5367, new_n5368, new_n5369, new_n5370, new_n5371,
    new_n5372, new_n5373, new_n5374, new_n5375, new_n5376, new_n5377,
    new_n5378, new_n5379, new_n5380, new_n5381, new_n5382, new_n5383,
    new_n5384, new_n5385, new_n5386, new_n5387, new_n5388, new_n5389,
    new_n5390, new_n5391, new_n5392, new_n5393, new_n5394, new_n5395,
    new_n5396, new_n5397, new_n5398, new_n5399, new_n5400, new_n5401,
    new_n5402, new_n5403, new_n5404, new_n5405, new_n5406, new_n5407,
    new_n5408, new_n5409, new_n5410, new_n5411, new_n5412, new_n5413,
    new_n5414, new_n5415, new_n5416, new_n5417, new_n5418, new_n5419,
    new_n5420, new_n5421, new_n5422, new_n5423, new_n5424, new_n5426,
    new_n5427, new_n5428, new_n5429, new_n5430_1, new_n5431, new_n5432,
    new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438,
    new_n5439, new_n5440, new_n5441, new_n5442, new_n5443, new_n5444,
    new_n5445, new_n5446, new_n5447, new_n5448, new_n5449_1, new_n5450,
    new_n5451, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467_1, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479_1, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502_1, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5514, new_n5515, new_n5516, new_n5517,
    new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523,
    new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529,
    new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535,
    new_n5536, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541,
    new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547,
    new_n5548, new_n5549, new_n5550_1, new_n5551, new_n5552, new_n5553,
    new_n5554, new_n5555, new_n5556, new_n5557, new_n5558, new_n5559,
    new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565,
    new_n5566, new_n5567, new_n5568, new_n5569, new_n5570, new_n5571,
    new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577,
    new_n5578, new_n5579, new_n5580, new_n5581, new_n5582, new_n5583,
    new_n5584, new_n5585, new_n5586_1, new_n5587, new_n5588, new_n5589,
    new_n5590, new_n5591, new_n5592, new_n5593, new_n5594, new_n5595,
    new_n5596, new_n5597, new_n5598, new_n5599, new_n5600, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644,
    new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5688, new_n5689, new_n5690, new_n5691, new_n5692, new_n5693,
    new_n5694, new_n5695, new_n5696, new_n5697, new_n5698, new_n5699,
    new_n5700, new_n5701, new_n5702, new_n5703, new_n5704, new_n5705,
    new_n5706, new_n5707, new_n5708, new_n5709, new_n5710, new_n5711,
    new_n5712, new_n5713, new_n5714, new_n5715, new_n5716, new_n5717,
    new_n5718, new_n5719, new_n5720, new_n5721, new_n5722, new_n5723,
    new_n5724, new_n5725_1, new_n5726, new_n5727, new_n5728, new_n5729,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759,
    new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786_1, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806_1, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851_1, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5861, new_n5862, new_n5863,
    new_n5864, new_n5865, new_n5866, new_n5867, new_n5868, new_n5869,
    new_n5870, new_n5871, new_n5872, new_n5873, new_n5874, new_n5875,
    new_n5876, new_n5877, new_n5878, new_n5879, new_n5880, new_n5881,
    new_n5882, new_n5883, new_n5884, new_n5885, new_n5886, new_n5887,
    new_n5888, new_n5889, new_n5890, new_n5891, new_n5892, new_n5893,
    new_n5894, new_n5895, new_n5896, new_n5897, new_n5898, new_n5899,
    new_n5900, new_n5901, new_n5902, new_n5903, new_n5904, new_n5905,
    new_n5906, new_n5907, new_n5908, new_n5909, new_n5910, new_n5911,
    new_n5912, new_n5913, new_n5914, new_n5915, new_n5916, new_n5917,
    new_n5918, new_n5919, new_n5920, new_n5921, new_n5922, new_n5923,
    new_n5924, new_n5925, new_n5926, new_n5927, new_n5928, new_n5929,
    new_n5930, new_n5931, new_n5932, new_n5933, new_n5934, new_n5935,
    new_n5936, new_n5937, new_n5938, new_n5939, new_n5940, new_n5941,
    new_n5942, new_n5943_1, new_n5944, new_n5945, new_n5946, new_n5948,
    new_n5949, new_n5950_1, new_n5951, new_n5952, new_n5953, new_n5954,
    new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960_1,
    new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966,
    new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972,
    new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978,
    new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984,
    new_n5985, new_n5986, new_n5987_1, new_n5988, new_n5989, new_n5990,
    new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996,
    new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002,
    new_n6003, new_n6004, new_n6005, new_n6006, new_n6007_1, new_n6008,
    new_n6009, new_n6010, new_n6011, new_n6012_1, new_n6013, new_n6014,
    new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020,
    new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026,
    new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032,
    new_n6034, new_n6035, new_n6036, new_n6037, new_n6038, new_n6039,
    new_n6040, new_n6041, new_n6042, new_n6043, new_n6044, new_n6045,
    new_n6046, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051,
    new_n6052, new_n6053, new_n6054_1, new_n6055, new_n6056, new_n6057,
    new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063,
    new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069,
    new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075,
    new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081,
    new_n6082, new_n6083, new_n6084, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104, new_n6105,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114_1, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6121, new_n6122, new_n6123, new_n6124,
    new_n6125, new_n6126, new_n6127, new_n6128, new_n6129, new_n6130,
    new_n6131, new_n6132, new_n6133, new_n6134, new_n6135, new_n6136,
    new_n6137, new_n6138, new_n6139, new_n6140, new_n6141, new_n6142,
    new_n6143, new_n6144, new_n6145, new_n6146, new_n6147_1, new_n6148,
    new_n6149, new_n6150, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160,
    new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166,
    new_n6167, new_n6168, new_n6169, new_n6170, new_n6171, new_n6172,
    new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178,
    new_n6179, new_n6180, new_n6181, new_n6182, new_n6183, new_n6184,
    new_n6185, new_n6186, new_n6187, new_n6188, new_n6189, new_n6190,
    new_n6191, new_n6192, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198_1, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204, new_n6205, new_n6206, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251_1,
    new_n6252, new_n6253, new_n6254, new_n6255, new_n6256, new_n6257,
    new_n6258_1, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270_1, new_n6271, new_n6272, new_n6273, new_n6274, new_n6275_1,
    new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6288, new_n6289, new_n6290, new_n6291, new_n6292, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314_1, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362_1, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436_1, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460_1, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6466, new_n6467, new_n6468, new_n6469, new_n6470,
    new_n6471, new_n6472, new_n6473, new_n6474, new_n6475, new_n6476,
    new_n6477, new_n6478, new_n6479, new_n6480_1, new_n6481, new_n6482,
    new_n6483, new_n6484, new_n6485, new_n6486, new_n6487, new_n6488,
    new_n6489, new_n6490, new_n6491, new_n6492, new_n6493, new_n6494,
    new_n6495, new_n6496, new_n6497, new_n6498, new_n6499, new_n6500,
    new_n6501, new_n6502, new_n6503, new_n6504, new_n6505, new_n6506,
    new_n6507, new_n6508, new_n6509, new_n6510, new_n6511, new_n6512,
    new_n6513, new_n6514, new_n6515, new_n6516, new_n6517_1, new_n6518,
    new_n6519, new_n6520, new_n6521, new_n6522, new_n6523, new_n6524,
    new_n6525, new_n6526, new_n6527, new_n6528, new_n6529, new_n6530,
    new_n6531, new_n6532, new_n6533, new_n6534, new_n6535, new_n6536,
    new_n6537, new_n6538, new_n6539, new_n6540, new_n6541, new_n6542,
    new_n6543, new_n6544, new_n6545, new_n6546, new_n6547, new_n6548,
    new_n6549, new_n6550, new_n6551, new_n6552, new_n6554, new_n6555_1,
    new_n6556, new_n6557, new_n6558, new_n6559, new_n6560, new_n6561,
    new_n6562, new_n6563, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586_1, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6640,
    new_n6641, new_n6642, new_n6643, new_n6644, new_n6645, new_n6646,
    new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652,
    new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658,
    new_n6659, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664,
    new_n6665, new_n6666, new_n6667, new_n6668, new_n6669, new_n6670,
    new_n6671, new_n6672, new_n6673, new_n6674, new_n6675, new_n6676,
    new_n6677, new_n6678, new_n6679, new_n6680_1, new_n6681, new_n6682_1,
    new_n6683, new_n6684, new_n6685, new_n6686, new_n6687, new_n6688,
    new_n6689, new_n6690, new_n6691, new_n6692, new_n6693_1, new_n6694,
    new_n6695, new_n6696_1, new_n6697, new_n6698, new_n6699, new_n6700,
    new_n6701, new_n6702, new_n6703_1, new_n6704, new_n6705, new_n6706,
    new_n6707, new_n6708, new_n6709, new_n6710, new_n6711, new_n6712,
    new_n6713, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718,
    new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758_1, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786_1, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791_1,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810_1, new_n6812, new_n6813, new_n6814, new_n6815, new_n6816,
    new_n6817, new_n6818, new_n6819, new_n6820, new_n6821, new_n6822,
    new_n6823, new_n6824, new_n6825, new_n6826, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853_1, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860, new_n6861, new_n6862, new_n6863, new_n6864,
    new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873_1, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6898, new_n6899, new_n6900, new_n6901,
    new_n6902, new_n6903, new_n6904, new_n6905, new_n6906, new_n6907,
    new_n6908, new_n6909, new_n6910, new_n6911, new_n6912, new_n6913,
    new_n6914, new_n6915, new_n6916, new_n6917, new_n6918, new_n6919,
    new_n6920, new_n6921, new_n6922, new_n6923, new_n6924, new_n6925,
    new_n6926, new_n6927, new_n6928, new_n6929, new_n6930, new_n6931,
    new_n6932, new_n6933, new_n6934, new_n6935, new_n6936, new_n6937,
    new_n6938, new_n6939, new_n6940, new_n6941, new_n6942, new_n6943,
    new_n6944, new_n6945, new_n6946_1, new_n6947, new_n6948, new_n6949,
    new_n6950, new_n6951, new_n6952_1, new_n6953, new_n6954, new_n6955,
    new_n6956, new_n6957, new_n6958, new_n6959, new_n6960, new_n6961,
    new_n6962, new_n6963, new_n6964, new_n6965, new_n6966, new_n6967,
    new_n6968, new_n6969, new_n6970, new_n6971, new_n6972, new_n6973,
    new_n6974, new_n6975, new_n6976, new_n6977, new_n6978, new_n6979_1,
    new_n6980, new_n6981, new_n6982, new_n6984, new_n6985, new_n6986,
    new_n6987, new_n6988, new_n6989, new_n6990, new_n6991, new_n6992,
    new_n6993, new_n6994, new_n6995, new_n6996, new_n6997, new_n6998,
    new_n6999_1, new_n7000, new_n7001, new_n7002, new_n7003, new_n7004,
    new_n7005, new_n7006, new_n7007, new_n7008, new_n7009, new_n7010,
    new_n7011, new_n7012, new_n7013, new_n7014, new_n7015, new_n7016,
    new_n7017, new_n7018, new_n7019, new_n7020, new_n7021, new_n7022,
    new_n7023, new_n7024, new_n7025, new_n7026, new_n7027, new_n7028,
    new_n7029, new_n7030, new_n7031, new_n7032, new_n7033, new_n7034,
    new_n7035, new_n7036, new_n7037, new_n7038, new_n7039, new_n7040,
    new_n7041, new_n7042, new_n7043, new_n7044, new_n7045, new_n7046,
    new_n7047, new_n7048, new_n7049, new_n7050, new_n7051, new_n7052,
    new_n7053, new_n7054, new_n7055, new_n7056, new_n7057, new_n7058,
    new_n7059, new_n7060, new_n7061, new_n7062, new_n7063, new_n7064,
    new_n7065, new_n7066, new_n7067, new_n7068, new_n7070, new_n7071_1,
    new_n7072, new_n7073_1, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104_1, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132_1, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152_1, new_n7153, new_n7154, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190, new_n7191, new_n7192,
    new_n7193, new_n7194, new_n7195, new_n7196, new_n7197, new_n7198,
    new_n7199, new_n7200, new_n7201, new_n7202, new_n7203, new_n7204,
    new_n7205, new_n7206, new_n7207, new_n7208, new_n7209, new_n7210,
    new_n7211, new_n7212, new_n7213, new_n7214, new_n7215, new_n7216,
    new_n7217, new_n7218, new_n7219, new_n7220, new_n7221, new_n7222,
    new_n7223, new_n7224, new_n7225, new_n7226, new_n7227, new_n7228,
    new_n7229, new_n7230, new_n7231, new_n7232, new_n7233, new_n7234,
    new_n7235, new_n7236, new_n7237, new_n7238, new_n7239, new_n7240,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246_1, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265_1,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270, new_n7271,
    new_n7272_1, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282_1, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382_1, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7417,
    new_n7418, new_n7419, new_n7420, new_n7421, new_n7422, new_n7423,
    new_n7424, new_n7425, new_n7426, new_n7427, new_n7428, new_n7429,
    new_n7430, new_n7431, new_n7432, new_n7433, new_n7434, new_n7435,
    new_n7436, new_n7437, new_n7438, new_n7439, new_n7440, new_n7441,
    new_n7442, new_n7443, new_n7444, new_n7445, new_n7446, new_n7447,
    new_n7448, new_n7449, new_n7450_1, new_n7451, new_n7452, new_n7453,
    new_n7454, new_n7455, new_n7456, new_n7457, new_n7458, new_n7459,
    new_n7460, new_n7461, new_n7462, new_n7463, new_n7464, new_n7465,
    new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471,
    new_n7472, new_n7473, new_n7474, new_n7475, new_n7476, new_n7477,
    new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483,
    new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489,
    new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495,
    new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501,
    new_n7503, new_n7504, new_n7505, new_n7506, new_n7507, new_n7508,
    new_n7509, new_n7510, new_n7511, new_n7512, new_n7513, new_n7514,
    new_n7515, new_n7516, new_n7517, new_n7518, new_n7519, new_n7520,
    new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526,
    new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532,
    new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538,
    new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544,
    new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550,
    new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556,
    new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562,
    new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568,
    new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574,
    new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580,
    new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586,
    new_n7587, new_n7588, new_n7589, new_n7591, new_n7592, new_n7593,
    new_n7594, new_n7595, new_n7596, new_n7597, new_n7598, new_n7599,
    new_n7600, new_n7601, new_n7602, new_n7603, new_n7604, new_n7605,
    new_n7606, new_n7607, new_n7608, new_n7609, new_n7610, new_n7611,
    new_n7612, new_n7613, new_n7614, new_n7615, new_n7616, new_n7617,
    new_n7618, new_n7619, new_n7620, new_n7621, new_n7622, new_n7623,
    new_n7624, new_n7625, new_n7626, new_n7627, new_n7628, new_n7629,
    new_n7630, new_n7631, new_n7632, new_n7633, new_n7634, new_n7635,
    new_n7636, new_n7637, new_n7638, new_n7639, new_n7640, new_n7641,
    new_n7642, new_n7643, new_n7644, new_n7645, new_n7646, new_n7647,
    new_n7648, new_n7649, new_n7650, new_n7651, new_n7652_1, new_n7653,
    new_n7654, new_n7655_1, new_n7656, new_n7657, new_n7658, new_n7659,
    new_n7660, new_n7661, new_n7662, new_n7663, new_n7664, new_n7665,
    new_n7666, new_n7667_1, new_n7668, new_n7669, new_n7670, new_n7671,
    new_n7672, new_n7673, new_n7674, new_n7675, new_n7677, new_n7678,
    new_n7679, new_n7680, new_n7681, new_n7682, new_n7683, new_n7684,
    new_n7685, new_n7686, new_n7687, new_n7688, new_n7689, new_n7690,
    new_n7691, new_n7692, new_n7693, new_n7694, new_n7695, new_n7696,
    new_n7697, new_n7698, new_n7699, new_n7700, new_n7701, new_n7702,
    new_n7703, new_n7704, new_n7705, new_n7706, new_n7707, new_n7708,
    new_n7709, new_n7710, new_n7711, new_n7712, new_n7713, new_n7714,
    new_n7715, new_n7716, new_n7717, new_n7718, new_n7719, new_n7720,
    new_n7721, new_n7722, new_n7723, new_n7724, new_n7725, new_n7726,
    new_n7727, new_n7728, new_n7729, new_n7730, new_n7731, new_n7732,
    new_n7733, new_n7734, new_n7735, new_n7736, new_n7737, new_n7738,
    new_n7739, new_n7740, new_n7741, new_n7742, new_n7743, new_n7744,
    new_n7745, new_n7746, new_n7747, new_n7748_1, new_n7749, new_n7750,
    new_n7751, new_n7752, new_n7753, new_n7754, new_n7755, new_n7756,
    new_n7757, new_n7758, new_n7759, new_n7760, new_n7761, new_n7762,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771_1, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823,
    new_n7824, new_n7825_1, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832_1, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7936, new_n7937, new_n7938, new_n7939,
    new_n7940, new_n7941_1, new_n7942, new_n7943, new_n7944, new_n7945,
    new_n7946, new_n7947, new_n7948, new_n7949, new_n7950, new_n7951,
    new_n7952, new_n7953, new_n7954, new_n7955, new_n7956, new_n7957,
    new_n7958, new_n7959, new_n7960, new_n7961, new_n7962, new_n7963,
    new_n7964, new_n7965, new_n7966, new_n7967, new_n7968, new_n7969,
    new_n7970, new_n7971, new_n7972_1, new_n7973, new_n7974, new_n7975,
    new_n7976, new_n7977, new_n7978, new_n7979, new_n7980, new_n7981,
    new_n7982, new_n7983, new_n7984, new_n7985, new_n7986, new_n7987,
    new_n7988_1, new_n7989, new_n7990, new_n7991, new_n7992, new_n7993,
    new_n7994, new_n7995, new_n7996, new_n7997, new_n7998, new_n7999,
    new_n8000, new_n8001, new_n8002_1, new_n8003, new_n8004, new_n8005,
    new_n8006, new_n8007, new_n8008, new_n8009, new_n8010, new_n8011,
    new_n8012, new_n8013, new_n8014, new_n8015, new_n8016, new_n8017,
    new_n8018, new_n8019, new_n8020, new_n8021, new_n8022, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044_1, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068_1, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073_1, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085_1, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8110, new_n8111, new_n8112, new_n8113, new_n8114, new_n8115,
    new_n8116, new_n8117, new_n8118, new_n8119, new_n8120, new_n8121,
    new_n8122, new_n8123, new_n8124_1, new_n8125, new_n8126, new_n8127,
    new_n8128, new_n8129, new_n8130, new_n8131, new_n8132, new_n8133,
    new_n8134, new_n8135, new_n8136, new_n8137, new_n8138, new_n8139,
    new_n8140, new_n8141, new_n8142, new_n8143, new_n8144_1, new_n8145,
    new_n8146, new_n8147, new_n8148, new_n8149, new_n8150, new_n8151,
    new_n8152, new_n8153, new_n8154, new_n8155, new_n8156, new_n8157,
    new_n8158, new_n8159, new_n8160, new_n8161, new_n8162, new_n8163,
    new_n8164, new_n8165, new_n8166, new_n8167, new_n8168, new_n8169,
    new_n8170, new_n8171, new_n8172, new_n8173, new_n8174, new_n8175,
    new_n8176, new_n8177, new_n8178, new_n8179, new_n8180, new_n8181,
    new_n8182, new_n8183, new_n8184, new_n8185, new_n8186, new_n8187,
    new_n8188, new_n8189, new_n8190, new_n8191, new_n8192, new_n8193,
    new_n8194, new_n8196, new_n8197, new_n8198, new_n8199, new_n8200,
    new_n8201, new_n8202, new_n8203, new_n8204_1, new_n8205, new_n8206,
    new_n8207, new_n8208, new_n8209, new_n8210, new_n8211, new_n8212,
    new_n8213, new_n8214, new_n8215_1, new_n8216, new_n8217, new_n8218,
    new_n8219, new_n8220, new_n8221, new_n8222, new_n8223, new_n8224,
    new_n8225, new_n8226, new_n8227, new_n8228, new_n8229, new_n8230,
    new_n8231, new_n8232, new_n8233, new_n8234, new_n8235, new_n8236,
    new_n8237, new_n8238, new_n8239, new_n8240, new_n8241, new_n8242,
    new_n8243, new_n8244, new_n8245, new_n8246, new_n8247, new_n8248,
    new_n8249, new_n8250, new_n8251, new_n8252, new_n8253, new_n8254,
    new_n8255, new_n8256, new_n8257, new_n8258, new_n8259, new_n8260,
    new_n8261, new_n8262_1, new_n8263, new_n8264, new_n8265, new_n8266,
    new_n8267, new_n8268, new_n8269, new_n8270, new_n8271, new_n8272,
    new_n8273, new_n8274, new_n8275, new_n8276, new_n8277, new_n8278,
    new_n8279, new_n8280, new_n8281, new_n8283, new_n8284, new_n8285,
    new_n8286, new_n8287, new_n8288, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302_1, new_n8303,
    new_n8304, new_n8305, new_n8306_1, new_n8307, new_n8308, new_n8309,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315_1,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321,
    new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397_1, new_n8398, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8431, new_n8432, new_n8433, new_n8434, new_n8435, new_n8436,
    new_n8437, new_n8438, new_n8439_1, new_n8440, new_n8441, new_n8442,
    new_n8443, new_n8444, new_n8445, new_n8446, new_n8447, new_n8448,
    new_n8449, new_n8450, new_n8451, new_n8452, new_n8453, new_n8454,
    new_n8455, new_n8456, new_n8458, new_n8459, new_n8460, new_n8461,
    new_n8462, new_n8463_1, new_n8464, new_n8465, new_n8466, new_n8467,
    new_n8468, new_n8469, new_n8470, new_n8471_1, new_n8472, new_n8473,
    new_n8474, new_n8475, new_n8476, new_n8477, new_n8478, new_n8479,
    new_n8480, new_n8481, new_n8482, new_n8483, new_n8484, new_n8485,
    new_n8486_1, new_n8487, new_n8488, new_n8489, new_n8490, new_n8491,
    new_n8492, new_n8493, new_n8494, new_n8495, new_n8496, new_n8497,
    new_n8498, new_n8499, new_n8500, new_n8501, new_n8502, new_n8503,
    new_n8504, new_n8505, new_n8506, new_n8507, new_n8508, new_n8509,
    new_n8510, new_n8511, new_n8512, new_n8513, new_n8514, new_n8515,
    new_n8516, new_n8517, new_n8518, new_n8519, new_n8520, new_n8521,
    new_n8522, new_n8523, new_n8524, new_n8525, new_n8526, new_n8527,
    new_n8528, new_n8529, new_n8530, new_n8531, new_n8532, new_n8533,
    new_n8534, new_n8535, new_n8536, new_n8537, new_n8538, new_n8539,
    new_n8540, new_n8541, new_n8542, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550_1, new_n8551, new_n8552_1,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598_1, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604_1, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635_1, new_n8636, new_n8637,
    new_n8638, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8644, new_n8645, new_n8646, new_n8647, new_n8648, new_n8649_1,
    new_n8650, new_n8651, new_n8652, new_n8653, new_n8654, new_n8655,
    new_n8656, new_n8657, new_n8658, new_n8659, new_n8660, new_n8661,
    new_n8662, new_n8663, new_n8664, new_n8665, new_n8666, new_n8667,
    new_n8668, new_n8669, new_n8670, new_n8671, new_n8672, new_n8673,
    new_n8674, new_n8675, new_n8676, new_n8677, new_n8678, new_n8679,
    new_n8680, new_n8681, new_n8682, new_n8683, new_n8684, new_n8685,
    new_n8686, new_n8687, new_n8688, new_n8689, new_n8690, new_n8691,
    new_n8692, new_n8693, new_n8694, new_n8695, new_n8696, new_n8697,
    new_n8698, new_n8699, new_n8700, new_n8701, new_n8702, new_n8703,
    new_n8704, new_n8705, new_n8706, new_n8707, new_n8708, new_n8709,
    new_n8710, new_n8711, new_n8712, new_n8713, new_n8714, new_n8716,
    new_n8717, new_n8718, new_n8719, new_n8720, new_n8721, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737_1, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744, new_n8745, new_n8746_1,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780_1, new_n8781, new_n8782,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799_1, new_n8800_1,
    new_n8801, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873_1,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8890, new_n8891, new_n8892_1,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909_1, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926_1, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8977,
    new_n8978, new_n8979, new_n8980, new_n8981, new_n8982, new_n8983,
    new_n8984, new_n8985, new_n8986, new_n8987, new_n8988, new_n8989,
    new_n8990, new_n8991, new_n8992, new_n8993, new_n8994, new_n8995,
    new_n8996, new_n8997_1, new_n8998, new_n8999, new_n9000, new_n9001,
    new_n9002, new_n9003, new_n9004, new_n9005, new_n9006, new_n9007,
    new_n9008, new_n9009, new_n9010, new_n9011, new_n9012, new_n9013,
    new_n9014, new_n9015, new_n9016, new_n9017, new_n9018, new_n9019,
    new_n9020, new_n9021, new_n9022, new_n9023, new_n9024, new_n9025,
    new_n9026_1, new_n9027, new_n9028, new_n9029, new_n9030, new_n9031,
    new_n9032, new_n9033, new_n9034, new_n9035, new_n9036, new_n9037,
    new_n9038, new_n9039, new_n9040, new_n9041, new_n9042, new_n9043,
    new_n9044, new_n9045, new_n9046, new_n9047, new_n9048, new_n9049,
    new_n9050, new_n9051, new_n9052, new_n9053, new_n9054, new_n9055,
    new_n9056, new_n9057, new_n9058, new_n9059, new_n9060, new_n9061,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096_1, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110_1,
    new_n9111, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9150, new_n9151, new_n9152, new_n9153,
    new_n9154_1, new_n9155, new_n9156, new_n9157, new_n9158, new_n9159,
    new_n9160, new_n9161, new_n9162, new_n9163, new_n9164, new_n9165,
    new_n9166, new_n9167, new_n9168, new_n9169, new_n9170, new_n9171,
    new_n9172, new_n9173, new_n9174, new_n9175, new_n9176, new_n9177,
    new_n9178, new_n9179, new_n9180, new_n9181, new_n9182, new_n9183,
    new_n9184, new_n9185, new_n9186_1, new_n9187, new_n9188, new_n9189,
    new_n9190, new_n9191, new_n9192, new_n9193, new_n9194, new_n9195,
    new_n9196, new_n9197, new_n9198, new_n9199, new_n9200, new_n9201,
    new_n9202, new_n9203, new_n9204, new_n9205, new_n9206, new_n9207,
    new_n9208, new_n9209, new_n9210, new_n9211, new_n9212, new_n9213,
    new_n9214, new_n9215, new_n9216, new_n9217, new_n9218, new_n9219,
    new_n9220, new_n9221, new_n9222, new_n9223, new_n9224, new_n9225,
    new_n9226, new_n9227, new_n9228, new_n9229, new_n9230, new_n9231,
    new_n9232, new_n9233, new_n9234, new_n9236, new_n9237, new_n9238,
    new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244,
    new_n9245, new_n9246, new_n9247, new_n9248, new_n9249, new_n9250,
    new_n9251, new_n9252_1, new_n9253, new_n9254, new_n9255, new_n9256,
    new_n9257, new_n9258, new_n9259, new_n9260, new_n9261, new_n9262,
    new_n9263, new_n9264, new_n9265, new_n9266, new_n9267, new_n9268,
    new_n9269, new_n9270, new_n9271, new_n9272, new_n9273, new_n9274,
    new_n9275, new_n9276, new_n9277, new_n9278, new_n9279, new_n9280,
    new_n9281, new_n9282, new_n9283, new_n9284, new_n9285, new_n9286,
    new_n9287, new_n9288, new_n9289, new_n9290, new_n9291, new_n9292,
    new_n9293, new_n9294, new_n9295, new_n9296, new_n9297, new_n9298,
    new_n9299, new_n9300, new_n9301, new_n9302, new_n9303, new_n9304,
    new_n9305, new_n9306, new_n9307, new_n9308, new_n9309, new_n9310,
    new_n9311, new_n9312, new_n9313, new_n9314_1, new_n9315, new_n9316,
    new_n9317, new_n9318, new_n9319, new_n9320, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342_1, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437_1, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447_1, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9494, new_n9495, new_n9496, new_n9497, new_n9498, new_n9499,
    new_n9500, new_n9501, new_n9502, new_n9503, new_n9504, new_n9505,
    new_n9506, new_n9507, new_n9508, new_n9509, new_n9510, new_n9511,
    new_n9512, new_n9513, new_n9514, new_n9515, new_n9516, new_n9517,
    new_n9518, new_n9519, new_n9520, new_n9521, new_n9522, new_n9523,
    new_n9524, new_n9525, new_n9526, new_n9527, new_n9528, new_n9529,
    new_n9530, new_n9531, new_n9532, new_n9533, new_n9534, new_n9535,
    new_n9536, new_n9537, new_n9538, new_n9539, new_n9540, new_n9541,
    new_n9542, new_n9543_1, new_n9544_1, new_n9545, new_n9546, new_n9547,
    new_n9548, new_n9549, new_n9550, new_n9551, new_n9552, new_n9553,
    new_n9554, new_n9555_1, new_n9556, new_n9557, new_n9558, new_n9559,
    new_n9560, new_n9561, new_n9562, new_n9563, new_n9564, new_n9565,
    new_n9566, new_n9567, new_n9568, new_n9569, new_n9570_1, new_n9571,
    new_n9572, new_n9573, new_n9574, new_n9575, new_n9576, new_n9577,
    new_n9578, new_n9580, new_n9581, new_n9582, new_n9583, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589_1, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633, new_n9634, new_n9635, new_n9636, new_n9637, new_n9638,
    new_n9639, new_n9640, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9666, new_n9667, new_n9668, new_n9669,
    new_n9670, new_n9671, new_n9672, new_n9673, new_n9674, new_n9675,
    new_n9676, new_n9677, new_n9678, new_n9679, new_n9680, new_n9681,
    new_n9682, new_n9683, new_n9684, new_n9685, new_n9686, new_n9687,
    new_n9688, new_n9689, new_n9690, new_n9691, new_n9692, new_n9693,
    new_n9694, new_n9695, new_n9696, new_n9697, new_n9698, new_n9699,
    new_n9700, new_n9701, new_n9702, new_n9703, new_n9704, new_n9705,
    new_n9706, new_n9707, new_n9708, new_n9709, new_n9710, new_n9711,
    new_n9712, new_n9713, new_n9714, new_n9715, new_n9716, new_n9717_1,
    new_n9718, new_n9719, new_n9720, new_n9721, new_n9722, new_n9723,
    new_n9724, new_n9725, new_n9726, new_n9727, new_n9728, new_n9729,
    new_n9730, new_n9731, new_n9732, new_n9733, new_n9734, new_n9735,
    new_n9736, new_n9737, new_n9738, new_n9739, new_n9740, new_n9741,
    new_n9742, new_n9743, new_n9744, new_n9745, new_n9746, new_n9747,
    new_n9748, new_n9749, new_n9750, new_n9751, new_n9753, new_n9754,
    new_n9755, new_n9756, new_n9757, new_n9758, new_n9759, new_n9760,
    new_n9761, new_n9762, new_n9763, new_n9764, new_n9765, new_n9766,
    new_n9767, new_n9768, new_n9769, new_n9770, new_n9771, new_n9772,
    new_n9773, new_n9774, new_n9775, new_n9776, new_n9777, new_n9778,
    new_n9779, new_n9780, new_n9781, new_n9782, new_n9783, new_n9784,
    new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790,
    new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796,
    new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802,
    new_n9803, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808,
    new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814,
    new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820,
    new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826,
    new_n9827, new_n9828, new_n9829, new_n9830_1, new_n9831, new_n9832,
    new_n9833, new_n9834, new_n9835, new_n9836, new_n9837, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893_1,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920, new_n9921_1, new_n9922, new_n9923,
    new_n9925, new_n9926, new_n9927, new_n9928, new_n9929, new_n9930,
    new_n9931, new_n9932, new_n9933, new_n9934, new_n9935, new_n9936_1,
    new_n9937, new_n9938, new_n9939, new_n9940, new_n9941, new_n9942,
    new_n9943, new_n9944, new_n9945, new_n9946, new_n9947, new_n9948,
    new_n9949, new_n9950, new_n9951, new_n9952, new_n9953, new_n9954,
    new_n9955, new_n9956, new_n9957, new_n9958, new_n9959, new_n9960,
    new_n9961, new_n9962, new_n9963, new_n9964, new_n9965, new_n9966,
    new_n9967, new_n9968, new_n9969, new_n9970, new_n9971, new_n9972,
    new_n9973, new_n9974, new_n9975, new_n9976, new_n9977_1, new_n9978,
    new_n9979, new_n9980, new_n9981, new_n9982, new_n9983, new_n9984,
    new_n9985, new_n9986, new_n9987, new_n9988, new_n9989, new_n9990,
    new_n9991, new_n9992, new_n9993, new_n9994, new_n9995, new_n9996,
    new_n9997, new_n9998, new_n9999, new_n10000, new_n10001, new_n10002,
    new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015,
    new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050_1,
    new_n10051_1, new_n10052, new_n10053, new_n10054, new_n10055,
    new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061_1, new_n10062, new_n10063, new_n10064, new_n10065,
    new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071,
    new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077,
    new_n10078, new_n10079, new_n10080_1, new_n10081, new_n10082,
    new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088,
    new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094,
    new_n10095, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111, new_n10112_1,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117, new_n10118,
    new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125, new_n10126, new_n10127, new_n10128, new_n10129, new_n10130,
    new_n10131, new_n10132, new_n10133, new_n10134, new_n10135, new_n10136,
    new_n10137, new_n10138, new_n10139, new_n10140, new_n10141, new_n10142,
    new_n10143, new_n10144, new_n10145, new_n10146, new_n10147_1,
    new_n10148, new_n10149, new_n10150, new_n10151, new_n10152, new_n10153,
    new_n10154, new_n10155, new_n10156, new_n10157, new_n10158, new_n10159,
    new_n10160, new_n10161, new_n10162, new_n10163, new_n10164, new_n10165,
    new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177,
    new_n10178, new_n10179, new_n10180, new_n10181, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217, new_n10218, new_n10219, new_n10220,
    new_n10221, new_n10222, new_n10223, new_n10224, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255_1,
    new_n10256, new_n10257, new_n10258, new_n10259, new_n10260, new_n10261,
    new_n10262, new_n10263, new_n10264, new_n10265, new_n10266, new_n10267,
    new_n10268, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278_1, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283_1, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10357,
    new_n10358, new_n10359, new_n10360, new_n10361, new_n10362, new_n10363,
    new_n10364, new_n10365, new_n10366, new_n10367, new_n10368, new_n10369,
    new_n10370, new_n10371, new_n10372, new_n10373, new_n10374, new_n10375,
    new_n10376, new_n10377, new_n10378_1, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407_1, new_n10408, new_n10409,
    new_n10410, new_n10411, new_n10412, new_n10413, new_n10414, new_n10415,
    new_n10416, new_n10417, new_n10418, new_n10419, new_n10420, new_n10421,
    new_n10422, new_n10423, new_n10424, new_n10425, new_n10426_1,
    new_n10427, new_n10428, new_n10429, new_n10430, new_n10431, new_n10432,
    new_n10433, new_n10434, new_n10435, new_n10436, new_n10437, new_n10438,
    new_n10439, new_n10440, new_n10441, new_n10442, new_n10444, new_n10445,
    new_n10446_1, new_n10447, new_n10448, new_n10449, new_n10450,
    new_n10451, new_n10452, new_n10453, new_n10454, new_n10455, new_n10456,
    new_n10457, new_n10458, new_n10459, new_n10460, new_n10461, new_n10462,
    new_n10463, new_n10464, new_n10465, new_n10466_1, new_n10467,
    new_n10468, new_n10469, new_n10470_1, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484,
    new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490,
    new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496,
    new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502,
    new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508,
    new_n10509, new_n10510, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515_1, new_n10516, new_n10517, new_n10518, new_n10519,
    new_n10520, new_n10521, new_n10522, new_n10523, new_n10524, new_n10525,
    new_n10526, new_n10527, new_n10528, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561, new_n10562,
    new_n10563, new_n10564, new_n10565, new_n10566, new_n10567, new_n10568,
    new_n10569, new_n10570, new_n10571, new_n10572, new_n10573_1,
    new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579,
    new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585,
    new_n10586, new_n10587, new_n10588, new_n10589, new_n10590,
    new_n10591_1, new_n10592, new_n10593, new_n10594, new_n10595,
    new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601,
    new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607,
    new_n10608, new_n10609, new_n10610, new_n10611, new_n10612, new_n10613,
    new_n10614, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630_1, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649,
    new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655,
    new_n10656, new_n10657, new_n10658, new_n10659, new_n10660, new_n10661,
    new_n10662, new_n10663, new_n10664, new_n10665, new_n10666, new_n10667,
    new_n10668, new_n10669, new_n10670, new_n10671, new_n10672, new_n10673,
    new_n10674, new_n10675, new_n10676, new_n10677, new_n10678, new_n10679,
    new_n10680, new_n10681, new_n10682, new_n10683, new_n10684, new_n10685,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10702, new_n10703, new_n10704,
    new_n10705, new_n10706, new_n10707, new_n10708, new_n10709, new_n10710,
    new_n10711, new_n10712, new_n10713, new_n10714, new_n10715, new_n10716,
    new_n10717, new_n10718, new_n10719, new_n10720, new_n10721, new_n10722,
    new_n10723, new_n10724, new_n10725, new_n10726, new_n10727, new_n10728,
    new_n10729, new_n10730, new_n10731, new_n10732, new_n10733, new_n10734,
    new_n10735, new_n10736_1, new_n10737, new_n10738, new_n10739,
    new_n10740, new_n10741, new_n10742, new_n10743, new_n10744, new_n10745,
    new_n10746, new_n10747, new_n10748, new_n10749, new_n10750_1,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765_1, new_n10766, new_n10767,
    new_n10768, new_n10769, new_n10770, new_n10771, new_n10772, new_n10773,
    new_n10774, new_n10775, new_n10776, new_n10777, new_n10778, new_n10779,
    new_n10780, new_n10781, new_n10782, new_n10783, new_n10784, new_n10785,
    new_n10786, new_n10788, new_n10789, new_n10790, new_n10791_1,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802_1,
    new_n10803, new_n10804, new_n10805, new_n10806, new_n10807, new_n10808,
    new_n10809, new_n10810, new_n10811, new_n10812, new_n10813, new_n10814,
    new_n10815, new_n10816, new_n10817, new_n10818, new_n10819, new_n10820,
    new_n10821, new_n10822, new_n10823, new_n10824, new_n10825, new_n10826,
    new_n10827, new_n10828, new_n10829, new_n10830, new_n10831, new_n10832,
    new_n10833, new_n10834, new_n10835, new_n10836, new_n10837, new_n10838,
    new_n10839, new_n10840, new_n10841, new_n10842, new_n10843, new_n10844,
    new_n10845, new_n10846, new_n10847, new_n10848, new_n10849, new_n10850,
    new_n10851, new_n10852, new_n10853, new_n10854, new_n10855, new_n10856,
    new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862_1, new_n10863, new_n10864, new_n10865, new_n10866,
    new_n10867, new_n10868, new_n10869, new_n10870, new_n10871, new_n10872,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903,
    new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909,
    new_n10910, new_n10911, new_n10912_1, new_n10913, new_n10914,
    new_n10915_1, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10928, new_n10929, new_n10930, new_n10931,
    new_n10932, new_n10933, new_n10934, new_n10935, new_n10936, new_n10937,
    new_n10938, new_n10939, new_n10940, new_n10941, new_n10942, new_n10943,
    new_n10944, new_n10945_1, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10961,
    new_n10962, new_n10963, new_n10964, new_n10965, new_n10966, new_n10967,
    new_n10968, new_n10969, new_n10970, new_n10971, new_n10972, new_n10973,
    new_n10974, new_n10975, new_n10976, new_n10977, new_n10978, new_n10979,
    new_n10980, new_n10981, new_n10982, new_n10983, new_n10984, new_n10985,
    new_n10986, new_n10987, new_n10988, new_n10989, new_n10990, new_n10991,
    new_n10992, new_n10993, new_n10994, new_n10995, new_n10996, new_n10997,
    new_n10998, new_n10999, new_n11000, new_n11001, new_n11002, new_n11003,
    new_n11004, new_n11005, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011, new_n11012, new_n11013, new_n11014, new_n11015,
    new_n11016, new_n11017, new_n11018, new_n11019, new_n11020, new_n11021,
    new_n11022, new_n11023, new_n11024, new_n11025, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045,
    new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052,
    new_n11053, new_n11054, new_n11055, new_n11056, new_n11057, new_n11058,
    new_n11059, new_n11060, new_n11061, new_n11062, new_n11063, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078, new_n11079, new_n11080, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093, new_n11094,
    new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101, new_n11102, new_n11103, new_n11104, new_n11105, new_n11106,
    new_n11107, new_n11108, new_n11109, new_n11110, new_n11111, new_n11112,
    new_n11113, new_n11114, new_n11115, new_n11116, new_n11117, new_n11118,
    new_n11119, new_n11120, new_n11121, new_n11122_1, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129,
    new_n11130, new_n11131, new_n11133, new_n11134, new_n11135, new_n11136,
    new_n11137, new_n11138, new_n11139, new_n11140, new_n11141, new_n11142,
    new_n11143_1, new_n11144, new_n11145, new_n11146, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11153,
    new_n11154, new_n11155, new_n11156, new_n11157, new_n11158_1,
    new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164,
    new_n11165, new_n11166, new_n11167, new_n11168, new_n11169, new_n11170,
    new_n11171, new_n11172, new_n11173, new_n11174, new_n11175, new_n11176,
    new_n11177, new_n11178, new_n11179, new_n11180, new_n11181, new_n11182,
    new_n11183, new_n11184, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192, new_n11193, new_n11194,
    new_n11195, new_n11196, new_n11197, new_n11198, new_n11199, new_n11200,
    new_n11201, new_n11202, new_n11203, new_n11204, new_n11205, new_n11206,
    new_n11207, new_n11208, new_n11209, new_n11210, new_n11211, new_n11212,
    new_n11213, new_n11214, new_n11215, new_n11216, new_n11217, new_n11219,
    new_n11220, new_n11221, new_n11222, new_n11223, new_n11224, new_n11225,
    new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231,
    new_n11232, new_n11233, new_n11234, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245, new_n11246, new_n11247, new_n11248, new_n11249,
    new_n11250, new_n11251, new_n11252, new_n11253, new_n11254, new_n11255,
    new_n11256, new_n11257, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269_1, new_n11270, new_n11271, new_n11272,
    new_n11273, new_n11274, new_n11275, new_n11276, new_n11277, new_n11278,
    new_n11279, new_n11280, new_n11281, new_n11282, new_n11283, new_n11284,
    new_n11285, new_n11286, new_n11287, new_n11288, new_n11289, new_n11290,
    new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11305, new_n11306, new_n11307, new_n11308, new_n11309,
    new_n11310, new_n11311, new_n11312, new_n11313, new_n11314, new_n11315,
    new_n11316, new_n11317, new_n11318, new_n11319, new_n11320, new_n11321,
    new_n11322, new_n11323, new_n11324, new_n11325, new_n11326, new_n11327,
    new_n11328, new_n11329, new_n11330, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344,
    new_n11345_1, new_n11346, new_n11347, new_n11348, new_n11349,
    new_n11350, new_n11351, new_n11352, new_n11353, new_n11354, new_n11355,
    new_n11356, new_n11357, new_n11358, new_n11359, new_n11360, new_n11361,
    new_n11362, new_n11363, new_n11364, new_n11365, new_n11366, new_n11367,
    new_n11368, new_n11369, new_n11370, new_n11371, new_n11372, new_n11373,
    new_n11374, new_n11375, new_n11376, new_n11377, new_n11378, new_n11379,
    new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385,
    new_n11386, new_n11387, new_n11388, new_n11389, new_n11391, new_n11392,
    new_n11393_1, new_n11394, new_n11395, new_n11396, new_n11397,
    new_n11398, new_n11399, new_n11400, new_n11401, new_n11402, new_n11403,
    new_n11404_1, new_n11405, new_n11406, new_n11407, new_n11408,
    new_n11409, new_n11410, new_n11411, new_n11412, new_n11413, new_n11414,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419, new_n11420,
    new_n11421, new_n11422, new_n11423, new_n11424, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444,
    new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450,
    new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462,
    new_n11463_1, new_n11464, new_n11465, new_n11466, new_n11467,
    new_n11468, new_n11469, new_n11470, new_n11471, new_n11472, new_n11473,
    new_n11474, new_n11475, new_n11476, new_n11478, new_n11479, new_n11480,
    new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496, new_n11497, new_n11498,
    new_n11499, new_n11500, new_n11501, new_n11502, new_n11503, new_n11504,
    new_n11505, new_n11506, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515, new_n11516,
    new_n11517, new_n11518, new_n11519, new_n11520, new_n11521, new_n11522,
    new_n11523, new_n11524, new_n11525, new_n11526, new_n11527, new_n11528,
    new_n11529_1, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534_1, new_n11535, new_n11536, new_n11537, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11564, new_n11565, new_n11566, new_n11567, new_n11568, new_n11569,
    new_n11570, new_n11571, new_n11572, new_n11573, new_n11574, new_n11575,
    new_n11576, new_n11577, new_n11578, new_n11579, new_n11580, new_n11581,
    new_n11582, new_n11583, new_n11584, new_n11585, new_n11586, new_n11587,
    new_n11588, new_n11589, new_n11590_1, new_n11591, new_n11592,
    new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605_1, new_n11606, new_n11607, new_n11608, new_n11609,
    new_n11610, new_n11611, new_n11612, new_n11613, new_n11614, new_n11615,
    new_n11616, new_n11617, new_n11618, new_n11619, new_n11620, new_n11621,
    new_n11622, new_n11623, new_n11624, new_n11625, new_n11626,
    new_n11627_1, new_n11628, new_n11629, new_n11630, new_n11631,
    new_n11632, new_n11633, new_n11634, new_n11635, new_n11636, new_n11637,
    new_n11638, new_n11639, new_n11640, new_n11641, new_n11642, new_n11643,
    new_n11644, new_n11645, new_n11646, new_n11647, new_n11648, new_n11650,
    new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656,
    new_n11657, new_n11658, new_n11659, new_n11660, new_n11661, new_n11662,
    new_n11663, new_n11664_1, new_n11665, new_n11666_1, new_n11667,
    new_n11668, new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674, new_n11675, new_n11676, new_n11677, new_n11678, new_n11679,
    new_n11680, new_n11681, new_n11682, new_n11683, new_n11684, new_n11685,
    new_n11686, new_n11687, new_n11688, new_n11689, new_n11690, new_n11691,
    new_n11692, new_n11693, new_n11694, new_n11695, new_n11696, new_n11697,
    new_n11698, new_n11699, new_n11700, new_n11701, new_n11702, new_n11703,
    new_n11704, new_n11705, new_n11706, new_n11707, new_n11708, new_n11709,
    new_n11710, new_n11711, new_n11712, new_n11713, new_n11714, new_n11715,
    new_n11716, new_n11717, new_n11718, new_n11719, new_n11720, new_n11721,
    new_n11722, new_n11723, new_n11724, new_n11725, new_n11726, new_n11727,
    new_n11728, new_n11729, new_n11730, new_n11731, new_n11732, new_n11733,
    new_n11734, new_n11735, new_n11736, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755, new_n11756_1, new_n11757,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776_1, new_n11777, new_n11778, new_n11779, new_n11780,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791, new_n11792,
    new_n11793, new_n11794, new_n11795, new_n11796, new_n11797, new_n11798,
    new_n11799, new_n11800, new_n11801, new_n11802, new_n11803, new_n11804,
    new_n11805, new_n11806, new_n11807, new_n11808, new_n11809, new_n11810,
    new_n11811, new_n11812, new_n11813, new_n11814, new_n11815, new_n11816,
    new_n11817, new_n11818, new_n11819, new_n11820, new_n11821,
    new_n11822_1, new_n11823, new_n11825, new_n11826, new_n11827,
    new_n11828, new_n11829, new_n11830, new_n11831, new_n11832, new_n11833,
    new_n11834, new_n11835, new_n11836, new_n11837, new_n11838, new_n11839,
    new_n11840, new_n11841, new_n11842_1, new_n11843, new_n11844,
    new_n11845, new_n11846, new_n11847_1, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854_1,
    new_n11855, new_n11856, new_n11857, new_n11858, new_n11859, new_n11860,
    new_n11861, new_n11862, new_n11863, new_n11864, new_n11865, new_n11866,
    new_n11867, new_n11868, new_n11869, new_n11870, new_n11871, new_n11872,
    new_n11873, new_n11874, new_n11875_1, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902_1, new_n11903, new_n11904, new_n11905, new_n11906,
    new_n11907, new_n11908, new_n11909, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926, new_n11927, new_n11928, new_n11929, new_n11930_1,
    new_n11931, new_n11932, new_n11933_1, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961_1, new_n11962, new_n11963, new_n11964,
    new_n11965, new_n11966, new_n11967, new_n11968, new_n11969, new_n11970,
    new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976,
    new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11999, new_n12000, new_n12001,
    new_n12002, new_n12003, new_n12004, new_n12005, new_n12006, new_n12007,
    new_n12008, new_n12009_1, new_n12010, new_n12011, new_n12012_1,
    new_n12013, new_n12014, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020, new_n12021, new_n12022, new_n12023, new_n12024,
    new_n12025_1, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032_1, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044, new_n12045, new_n12046,
    new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052,
    new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058,
    new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064,
    new_n12065, new_n12066, new_n12067, new_n12068, new_n12069, new_n12070,
    new_n12071, new_n12072, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12085, new_n12086, new_n12087, new_n12088, new_n12089,
    new_n12090, new_n12091, new_n12092, new_n12093, new_n12094, new_n12095,
    new_n12096, new_n12097, new_n12098, new_n12099, new_n12100, new_n12101,
    new_n12102, new_n12103, new_n12104, new_n12105, new_n12106, new_n12107,
    new_n12108, new_n12109, new_n12110, new_n12111, new_n12112, new_n12113,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121, new_n12122, new_n12123, new_n12124, new_n12125,
    new_n12126, new_n12127, new_n12128, new_n12129, new_n12130, new_n12131,
    new_n12132, new_n12133, new_n12134, new_n12135, new_n12136, new_n12137,
    new_n12138, new_n12139, new_n12140, new_n12141, new_n12142_1,
    new_n12143, new_n12144, new_n12145, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166_1, new_n12167, new_n12168, new_n12169, new_n12171,
    new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177,
    new_n12178, new_n12179, new_n12180, new_n12181, new_n12182, new_n12183,
    new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189,
    new_n12190, new_n12191, new_n12192, new_n12193, new_n12194, new_n12195,
    new_n12196, new_n12197, new_n12198, new_n12199, new_n12200, new_n12201,
    new_n12202, new_n12203, new_n12204, new_n12205, new_n12206, new_n12207,
    new_n12208, new_n12209, new_n12210, new_n12211, new_n12212, new_n12213,
    new_n12214, new_n12215, new_n12216, new_n12217, new_n12218_1,
    new_n12219, new_n12220, new_n12221, new_n12222, new_n12223, new_n12224,
    new_n12225, new_n12226, new_n12227, new_n12228, new_n12229, new_n12230,
    new_n12231, new_n12232_1, new_n12233, new_n12234, new_n12235,
    new_n12236, new_n12237, new_n12238, new_n12239, new_n12240, new_n12241,
    new_n12242, new_n12243, new_n12244, new_n12245, new_n12246, new_n12247,
    new_n12248, new_n12249, new_n12250, new_n12251, new_n12252, new_n12253,
    new_n12254, new_n12255, new_n12256, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270_1, new_n12271,
    new_n12272, new_n12273, new_n12274, new_n12275, new_n12276, new_n12277,
    new_n12278, new_n12279, new_n12280, new_n12281, new_n12282, new_n12283,
    new_n12284, new_n12285, new_n12286, new_n12287, new_n12288, new_n12289,
    new_n12290, new_n12291, new_n12292, new_n12293, new_n12294, new_n12295,
    new_n12296, new_n12297, new_n12298, new_n12299, new_n12300, new_n12301,
    new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315, new_n12316, new_n12317, new_n12318, new_n12319,
    new_n12320, new_n12321_1, new_n12322, new_n12323, new_n12324,
    new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335,
    new_n12336_1, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341, new_n12342, new_n12344, new_n12345, new_n12346, new_n12347,
    new_n12348, new_n12349, new_n12350, new_n12351, new_n12352, new_n12353,
    new_n12354, new_n12355_1, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370,
    new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382,
    new_n12383, new_n12384, new_n12385, new_n12386, new_n12387, new_n12388,
    new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394,
    new_n12395, new_n12396, new_n12397, new_n12398, new_n12399, new_n12400,
    new_n12401, new_n12402, new_n12403, new_n12404, new_n12405, new_n12406,
    new_n12407, new_n12408, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444, new_n12445, new_n12446, new_n12447, new_n12448, new_n12449,
    new_n12450, new_n12451, new_n12452, new_n12453, new_n12454, new_n12455,
    new_n12456, new_n12457, new_n12458, new_n12459, new_n12460, new_n12461,
    new_n12462, new_n12463, new_n12464, new_n12465, new_n12466, new_n12467,
    new_n12468, new_n12469, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495, new_n12496, new_n12497,
    new_n12498, new_n12499, new_n12500, new_n12501, new_n12502, new_n12503,
    new_n12504, new_n12505, new_n12506, new_n12507, new_n12508, new_n12509,
    new_n12510, new_n12511, new_n12512, new_n12513, new_n12514, new_n12516,
    new_n12517, new_n12518, new_n12519, new_n12520, new_n12521, new_n12522,
    new_n12523, new_n12524, new_n12525, new_n12526, new_n12527, new_n12528,
    new_n12529, new_n12530, new_n12531, new_n12532, new_n12533, new_n12534,
    new_n12535_1, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545,
    new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573_1, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591, new_n12592,
    new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598,
    new_n12599, new_n12600, new_n12601;
not_4  g00000(n2674, new_n386);
nor_5  g00001(n10426, new_n386, new_n387);
not_4  g00002(n4895, new_n388);
nor_5  g00003(n8598, new_n388, new_n389_1);
nor_5  g00004(n12270, n8780, new_n390);
not_4  g00005(new_n390, new_n391);
nor_5  g00006(new_n391, new_n389_1, new_n392);
not_4  g00007(n1268, new_n393);
nor_5  g00008(new_n393, n1265, new_n394_1);
nor_5  g00009(n8892, n1265, new_n395);
nor_5  g00010(new_n395, new_n394_1, new_n396);
nor_5  g00011(new_n396, n8598, new_n397);
not_4  g00012(n5046, new_n398);
nor_5  g00013(n6362, new_n398, new_n399);
nor_5  g00014(n1268, n394, new_n400);
not_4  g00015(new_n400, new_n401);
nor_5  g00016(new_n401, new_n399, new_n402);
not_4  g00017(n8649, new_n403);
nor_5  g00018(new_n403, n5950, new_n404);
nor_5  g00019(n12927, n10050, new_n405);
not_4  g00020(new_n405, new_n406);
nor_5  g00021(new_n406, new_n404, new_n407);
not_4  g00022(n8439, new_n408);
nor_5  g00023(new_n408, n702, new_n409);
nor_5  g00024(n3910, n844, new_n410);
not_4  g00025(new_n410, new_n411_1);
nor_5  g00026(new_n411_1, new_n409, new_n412);
not_4  g00027(n2061, new_n413);
nor_5  g00028(n9026, new_n413, new_n414);
nor_5  g00029(n12336, n9186, new_n415);
not_4  g00030(new_n415, new_n416);
nor_5  g00031(new_n416, new_n414, new_n417);
not_4  g00032(n10147, new_n418);
nor_5  g00033(new_n418, n8397, new_n419);
nor_5  g00034(n14464, n12976, new_n420);
not_4  g00035(new_n420, new_n421);
nor_5  g00036(new_n421, new_n419, new_n422);
not_4  g00037(n7667, new_n423);
nor_5  g00038(n11930, new_n423, new_n424);
nor_5  g00039(n13636, n11930, new_n425);
nor_5  g00040(new_n425, new_n424, new_n426);
nor_5  g00041(new_n426, n8397, new_n427_1);
not_4  g00042(n14408, new_n428);
nor_5  g00043(n14483, new_n428, new_n429);
nor_5  g00044(n14303, n7667, new_n430);
not_4  g00045(new_n430, new_n431);
nor_5  g00046(new_n431, new_n429, new_n432);
not_4  g00047(n12025, new_n433);
nor_5  g00048(new_n433, n6460, new_n434);
nor_5  g00049(n5023, n3673, new_n435);
not_4  g00050(new_n435, new_n436);
nor_5  g00051(new_n436, new_n434, new_n437);
not_4  g00052(n3130, new_n438);
nor_5  g00053(n13000, new_n438, new_n439);
nor_5  g00054(n13000, n10446, new_n440);
nor_5  g00055(new_n440, new_n439, new_n441);
nor_5  g00056(new_n441, n6460, new_n442);
not_4  g00057(n5786, new_n443);
nor_5  g00058(n8486, new_n443, new_n444);
nor_5  g00059(n9589, n8552, new_n445);
not_4  g00060(new_n445, new_n446);
nor_5  g00061(new_n446, new_n444, new_n447);
nor_5  g00062(n8997, n3532, new_n448);
not_4  g00063(n3532, new_n449);
nand_5 g00064(n11345, new_n449, new_n450);
not_4  g00065(new_n450, new_n451_1);
nor_5  g00066(new_n451_1, new_n448, new_n452);
nor_5  g00067(new_n452, n8486, new_n453);
not_4  g00068(n6480, new_n454);
nor_5  g00069(n6791, new_n454, new_n455);
nor_5  g00070(n11345, n3263, new_n456);
not_4  g00071(new_n456, new_n457);
nor_5  g00072(new_n457, new_n455, new_n458);
not_4  g00073(n4615, new_n459);
nor_5  g00074(n4785, new_n459, new_n460);
nor_5  g00075(n9921, n730, new_n461);
not_4  g00076(new_n461, new_n462_1);
nor_5  g00077(new_n462_1, new_n460, new_n463);
not_4  g00078(n427, new_n464);
nor_5  g00079(n9893, new_n464, new_n465);
nor_5  g00080(n6999, n6517, new_n466);
not_4  g00081(new_n466, new_n467);
nor_5  g00082(new_n467, new_n465, new_n468);
not_4  g00083(n12321, new_n469);
nor_5  g00084(new_n469, n5502, new_n470);
nor_5  g00085(n14072, n9544, new_n471);
not_4  g00086(new_n471, new_n472);
nor_5  g00087(new_n472, new_n470, new_n473);
not_4  g00088(n6555, new_n474);
nor_5  g00089(n9555, new_n474, new_n475);
nor_5  g00090(n10736, n7972, new_n476);
not_4  g00091(new_n476, new_n477);
nor_5  g00092(new_n477, new_n475, new_n478);
not_4  g00093(n4659, new_n479);
nor_5  g00094(new_n479, n4131, new_n480);
nor_5  g00095(n12573, n10470, new_n481);
not_4  g00096(new_n481, new_n482);
nor_5  g00097(new_n482, new_n480, new_n483);
not_4  g00098(n11590, new_n484);
nor_5  g00099(new_n484, n5014, new_n485);
nor_5  g00100(n11158, n10407, new_n486);
not_4  g00101(new_n486, new_n487);
nor_5  g00102(new_n487, new_n485, new_n488);
not_4  g00103(n9154, new_n489);
nor_5  g00104(n11933, new_n489, new_n490_1);
nor_5  g00105(n6436, n3833, new_n491);
not_4  g00106(new_n491, new_n492);
nor_5  g00107(new_n492, new_n490_1, new_n493);
not_4  g00108(n11875, new_n494);
nor_5  g00109(new_n494, n8262, new_n495);
nor_5  g00110(n10061, n4117, new_n496);
not_4  g00111(new_n496, new_n497);
nor_5  g00112(new_n497, new_n495, new_n498_1);
not_4  g00113(n4022, new_n499);
not_4  g00114(n1568, new_n500);
nand_5 g00115(n8635, new_n500, new_n501);
nand_5 g00116(new_n501, new_n499, new_n502);
nor_5  g00117(new_n502, n13814, new_n503);
not_4  g00118(n8800, new_n504);
nor_5  g00119(new_n504, n8463, new_n505);
nor_5  g00120(n5184, n203, new_n506);
not_4  g00121(new_n506, new_n507);
nor_5  g00122(new_n507, new_n505, new_n508);
not_4  g00123(n4154, new_n509);
nor_5  g00124(new_n509, n4000, new_n510);
nor_5  g00125(n6703, n3506, new_n511);
not_4  g00126(new_n511, new_n512);
nor_5  g00127(new_n512, new_n510, new_n513);
not_4  g00128(n7652, new_n514);
nor_5  g00129(n8073, new_n514, new_n515);
nor_5  g00130(n13093, n650, new_n516);
not_4  g00131(new_n516, new_n517);
nor_5  g00132(new_n517, new_n515, new_n518);
not_4  g00133(n3804, new_n519);
nor_5  g00134(n10112, new_n519, new_n520);
nor_5  g00135(n10466, n10112, new_n521);
nor_5  g00136(new_n521, new_n520, new_n522);
nor_5  g00137(new_n522, n8073, new_n523);
not_4  g00138(n13882, new_n524);
nor_5  g00139(new_n524, n5943, new_n525);
nor_5  g00140(n6680, n3804, new_n526);
not_4  g00141(new_n526, new_n527);
nor_5  g00142(new_n527, new_n525, new_n528);
not_4  g00143(n8746, new_n529);
nor_5  g00144(new_n529, n5430, new_n530);
nor_5  g00145(n8550, n5725, new_n531);
not_4  g00146(new_n531, new_n532);
nor_5  g00147(new_n532, new_n530, new_n533);
nor_5  g00148(n5430, n760, new_n534);
not_4  g00149(new_n534, new_n535);
not_4  g00150(n13295, new_n536);
nor_5  g00151(new_n536, n3799, new_n537);
nor_5  g00152(new_n537, new_n535, new_n538);
not_4  g00153(n3367, new_n539);
nor_5  g00154(n9543, new_n539, new_n540);
nor_5  g00155(n11776, n6873, new_n541);
not_4  g00156(new_n541, new_n542);
nor_5  g00157(new_n542, new_n540, new_n543_1);
not_4  g00158(n271, new_n544);
nor_5  g00159(n6007, new_n544, new_n545);
nor_5  g00160(n6007, n5960, new_n546);
nor_5  g00161(new_n546, new_n545, new_n547);
nor_5  g00162(new_n547, n9543, new_n548);
not_4  g00163(n13224, new_n549);
nor_5  g00164(new_n549, n11605, new_n550);
nor_5  g00165(n9977, n5225, new_n551);
not_4  g00166(new_n551, new_n552);
nor_5  g00167(new_n552, new_n550, new_n553);
not_4  g00168(n74, new_n554);
nor_5  g00169(n9314, new_n554, new_n555);
nor_5  g00170(n13109, n9110, new_n556);
not_4  g00171(new_n556, new_n557);
nor_5  g00172(new_n557, new_n555, new_n558);
not_4  g00173(n1763, new_n559);
nor_5  g00174(n12009, new_n559, new_n560);
nor_5  g00175(n5033, n4172, new_n561);
not_4  g00176(new_n561, new_n562);
nor_5  g00177(new_n562, new_n560, new_n563);
not_4  g00178(n1222, new_n564);
nor_5  g00179(n11961, new_n564, new_n565);
nor_5  g00180(n7832, n1776, new_n566);
not_4  g00181(new_n566, new_n567);
nor_5  g00182(new_n567, new_n565, new_n568);
not_4  g00183(n1027, new_n569);
nand_5 g00184(n11842, new_n569, new_n570);
not_4  g00185(new_n570, new_n571);
nor_5  g00186(n2048, n1027, new_n572);
nor_5  g00187(new_n572, new_n571, new_n573);
nor_5  g00188(new_n573, n11961, new_n574);
nor_5  g00189(n8002, n2166, new_n575);
not_4  g00190(new_n575, new_n576);
not_4  g00191(n6147, new_n577);
not_4  g00192(n2166, new_n578);
nand_5 g00193(n2201, new_n578, new_n579);
nand_5 g00194(new_n579, new_n577, new_n580);
nor_5  g00195(new_n580, n11842, new_n581);
nand_5 g00196(new_n581, new_n576, new_n582);
nand_5 g00197(new_n582, new_n574, new_n583);
nand_5 g00198(new_n583, new_n568, new_n584);
not_4  g00199(n1776, new_n585);
nor_5  g00200(n14475, new_n585, new_n586);
nor_5  g00201(n14475, n13625, new_n587);
nor_5  g00202(new_n587, new_n586, new_n588);
nor_5  g00203(new_n588, n10573, new_n589);
nand_5 g00204(new_n589, new_n584, new_n590);
not_4  g00205(n13102, new_n591);
nor_5  g00206(new_n591, n10573, new_n592);
nor_5  g00207(n13363, n7354, new_n593);
not_4  g00208(new_n593, new_n594);
nor_5  g00209(new_n594, new_n592, new_n595);
nand_5 g00210(new_n595, new_n590, new_n596);
not_4  g00211(n13363, new_n597);
nor_5  g00212(new_n597, n6054, new_n598);
nor_5  g00213(n6054, n2573, new_n599);
nor_5  g00214(new_n599, new_n598, new_n600);
nor_5  g00215(new_n600, n12009, new_n601);
nand_5 g00216(new_n601, new_n596, new_n602);
nand_5 g00217(new_n602, new_n563, new_n603);
not_4  g00218(n4172, new_n604);
nor_5  g00219(n4774, new_n604, new_n605);
nor_5  g00220(n4774, n4755, new_n606);
nor_5  g00221(new_n606, new_n605, new_n607);
nor_5  g00222(new_n607, n9314, new_n608);
nand_5 g00223(new_n608, new_n603, new_n609);
nand_5 g00224(new_n609, new_n558, new_n610);
not_4  g00225(n9110, new_n611);
nor_5  g00226(new_n611, n7104, new_n612);
nor_5  g00227(n13231, n7104, new_n613);
nor_5  g00228(new_n613, new_n612, new_n614);
nor_5  g00229(new_n614, n11605, new_n615);
nand_5 g00230(new_n615, new_n610, new_n616);
nand_5 g00231(new_n616, new_n553, new_n617);
not_4  g00232(n9977, new_n618);
nor_5  g00233(new_n618, n1347, new_n619);
nor_5  g00234(n8315, n1347, new_n620);
nor_5  g00235(new_n620, new_n619, new_n621);
nor_5  g00236(new_n621, n6258, new_n622);
nand_5 g00237(new_n622, new_n617, new_n623);
not_4  g00238(n13890, new_n624);
nor_5  g00239(new_n624, n6258, new_n625);
nor_5  g00240(n2334, n271, new_n626);
not_4  g00241(new_n626, new_n627);
nor_5  g00242(new_n627, new_n625, new_n628);
nand_5 g00243(new_n628, new_n623, new_n629);
nand_5 g00244(new_n629, new_n548, new_n630);
nand_5 g00245(new_n630, new_n543_1, new_n631);
not_4  g00246(n6873, new_n632);
nor_5  g00247(n7988, new_n632, new_n633);
nor_5  g00248(n10912, n7988, new_n634);
nor_5  g00249(new_n634, new_n633, new_n635);
nor_5  g00250(new_n635, n10630, new_n636);
nand_5 g00251(new_n636, new_n631, new_n637);
not_4  g00252(n5185, new_n638);
nor_5  g00253(n10630, new_n638, new_n639);
nor_5  g00254(n3799, n3652, new_n640);
not_4  g00255(new_n640, new_n641);
nor_5  g00256(new_n641, new_n639, new_n642);
nand_5 g00257(new_n642, new_n637, new_n643);
nand_5 g00258(new_n643, new_n538, new_n644);
nand_5 g00259(new_n644, new_n533, new_n645);
not_4  g00260(n5725, new_n646);
nor_5  g00261(new_n646, n2164, new_n647);
nor_5  g00262(n14163, n2164, new_n648);
nor_5  g00263(new_n648, new_n647, new_n649);
nor_5  g00264(new_n649, n5943, new_n650_1);
nand_5 g00265(new_n650_1, new_n645, new_n651);
nand_5 g00266(new_n651, new_n528, new_n652);
nand_5 g00267(new_n652, new_n523, new_n653);
nand_5 g00268(new_n653, new_n518, new_n654);
not_4  g00269(n650, new_n655);
nor_5  g00270(n9252, new_n655, new_n656_1);
nor_5  g00271(n11902, n9252, new_n657);
nor_5  g00272(new_n657, new_n656_1, new_n658);
nor_5  g00273(new_n658, n411, new_n659);
nand_5 g00274(new_n659, new_n654, new_n660);
not_4  g00275(n8799, new_n661);
nor_5  g00276(new_n661, n411, new_n662);
nor_5  g00277(n12614, n10765, new_n663);
not_4  g00278(new_n663, new_n664);
nor_5  g00279(new_n664, new_n662, new_n665);
nand_5 g00280(new_n665, new_n660, new_n666_1);
nor_5  g00281(n4000, n3388, new_n667);
not_4  g00282(new_n667, new_n668);
not_4  g00283(n10765, new_n669);
nand_5 g00284(n12142, new_n669, new_n670);
not_4  g00285(new_n670, new_n671);
nor_5  g00286(new_n671, new_n668, new_n672);
nand_5 g00287(new_n672, new_n666_1, new_n673);
nand_5 g00288(new_n673, new_n513, new_n674_1);
not_4  g00289(n6703, new_n675);
nor_5  g00290(n11269, new_n675, new_n676);
nor_5  g00291(n11269, n462, new_n677);
nor_5  g00292(new_n677, new_n676, new_n678);
nor_5  g00293(new_n678, n8926, new_n679);
nand_5 g00294(new_n679, new_n674_1, new_n680);
not_4  g00295(n3893, new_n681);
nor_5  g00296(n8926, new_n681, new_n682_1);
nor_5  g00297(n8044, n2454, new_n683);
not_4  g00298(new_n683, new_n684);
nor_5  g00299(new_n684, new_n682_1, new_n685);
nand_5 g00300(new_n685, new_n680, new_n686);
not_4  g00301(n8044, new_n687);
nor_5  g00302(n8204, new_n687, new_n688);
nor_5  g00303(n14293, n8204, new_n689);
nor_5  g00304(new_n689, new_n688, new_n690);
nor_5  g00305(new_n690, n8463, new_n691);
nand_5 g00306(new_n691, new_n686, new_n692);
nand_5 g00307(new_n692, new_n508, new_n693);
not_4  g00308(n5184, new_n694);
nor_5  g00309(new_n694, n2895, new_n695);
nor_5  g00310(n2895, n737, new_n696);
nor_5  g00311(new_n696, new_n695, new_n697);
nor_5  g00312(new_n697, n1568, new_n698);
nand_5 g00313(new_n698, new_n693, new_n699);
nand_5 g00314(new_n699, new_n503, new_n700);
nor_5  g00315(n10255, new_n499, new_n701);
nor_5  g00316(n10255, n5449, new_n702_1);
nor_5  g00317(new_n702_1, new_n701, new_n703);
nor_5  g00318(new_n703, n8262, new_n704);
nand_5 g00319(new_n704, new_n700, new_n705);
nand_5 g00320(new_n705, new_n498_1, new_n706);
not_4  g00321(n10061, new_n707);
nor_5  g00322(n12885, new_n707, new_n708);
nor_5  g00323(n12885, n11666, new_n709);
nor_5  g00324(new_n709, new_n708, new_n710);
nor_5  g00325(new_n710, n11933, new_n711);
nand_5 g00326(new_n711, new_n706, new_n712);
nand_5 g00327(new_n712, new_n493, new_n713);
nor_5  g00328(n11143, n5014, new_n714);
not_4  g00329(new_n714, new_n715);
not_4  g00330(n2699, new_n716);
nor_5  g00331(n6436, new_n716, new_n717);
nor_5  g00332(new_n717, new_n715, new_n718);
nand_5 g00333(new_n718, new_n713, new_n719);
nand_5 g00334(new_n719, new_n488, new_n720);
nor_5  g00335(n10051, n4131, new_n721);
not_4  g00336(new_n721, new_n722);
not_4  g00337(n13992, new_n723);
nor_5  g00338(new_n723, n10407, new_n724);
nor_5  g00339(new_n724, new_n722, new_n725);
nand_5 g00340(new_n725, new_n720, new_n726);
nand_5 g00341(new_n726, new_n483, new_n727);
not_4  g00342(n10470, new_n728);
nor_5  g00343(new_n728, n6693, new_n729);
nor_5  g00344(n12829, n6693, new_n730_1);
nor_5  g00345(new_n730_1, new_n729, new_n731);
nor_5  g00346(new_n731, n9555, new_n732);
nand_5 g00347(new_n732, new_n727, new_n733);
nand_5 g00348(new_n733, new_n478, new_n734);
not_4  g00349(n7972, new_n735);
nor_5  g00350(new_n735, n3972, new_n736);
nor_5  g00351(n10945, n3972, new_n737_1);
nor_5  g00352(new_n737_1, new_n736, new_n738);
nor_5  g00353(new_n738, n7450, new_n739);
nand_5 g00354(new_n739, new_n734, new_n740);
not_4  g00355(n10615, new_n741);
nor_5  g00356(new_n741, n7450, new_n742);
nor_5  g00357(n9830, n8302, new_n743);
not_4  g00358(new_n743, new_n744);
nor_5  g00359(new_n744, new_n742, new_n745);
nand_5 g00360(new_n745, new_n740, new_n746);
not_4  g00361(n8302, new_n747);
nor_5  g00362(new_n747, n3166, new_n748);
nor_5  g00363(n6270, n3166, new_n749);
nor_5  g00364(new_n749, new_n748, new_n750);
nor_5  g00365(new_n750, n5502, new_n751);
nand_5 g00366(new_n751, new_n746, new_n752);
nand_5 g00367(new_n752, new_n473, new_n753);
not_4  g00368(n14072, new_n754);
nor_5  g00369(new_n754, n6251, new_n755);
nor_5  g00370(n6251, n1702, new_n756);
nor_5  g00371(new_n756, new_n755, new_n757);
nor_5  g00372(new_n757, n6758, new_n758);
nand_5 g00373(new_n758, new_n753, new_n759);
not_4  g00374(n4147, new_n760_1);
nor_5  g00375(n6758, new_n760_1, new_n761);
nor_5  g00376(n10378, n10080, new_n762);
not_4  g00377(new_n762, new_n763);
nor_5  g00378(new_n763, new_n761, new_n764);
nand_5 g00379(new_n764, new_n759, new_n765);
not_4  g00380(n10080, new_n766);
nor_5  g00381(new_n766, n977, new_n767);
nor_5  g00382(n4282, n977, new_n768);
nor_5  g00383(new_n768, new_n767, new_n769);
nor_5  g00384(new_n769, n9893, new_n770);
nand_5 g00385(new_n770, new_n765, new_n771);
nand_5 g00386(new_n771, new_n468, new_n772);
not_4  g00387(n6999, new_n773);
nor_5  g00388(n10862, new_n773, new_n774);
nor_5  g00389(n12218, n10862, new_n775);
nor_5  g00390(new_n775, new_n774, new_n776);
nor_5  g00391(new_n776, n9936, new_n777);
nand_5 g00392(new_n777, new_n772, new_n778);
not_4  g00393(n1093, new_n779);
nor_5  g00394(n9936, new_n779, new_n780);
nor_5  g00395(n8737, n2615, new_n781);
not_4  g00396(new_n781, new_n782);
nor_5  g00397(new_n782, new_n780, new_n783);
nand_5 g00398(new_n783, new_n778, new_n784);
not_4  g00399(n8737, new_n785);
nor_5  g00400(n13561, new_n785, new_n786);
nor_5  g00401(n13561, n656, new_n787);
nor_5  g00402(new_n787, new_n786, new_n788);
nor_5  g00403(new_n788, n4785, new_n789);
nand_5 g00404(new_n789, new_n784, new_n790);
nand_5 g00405(new_n790, new_n463, new_n791);
not_4  g00406(n9921, new_n792);
nor_5  g00407(n10283, new_n792, new_n793);
nor_5  g00408(n10283, n3775, new_n794);
nor_5  g00409(new_n794, new_n793, new_n795);
nor_5  g00410(new_n795, n6791, new_n796);
nand_5 g00411(new_n796, new_n791, new_n797);
nand_5 g00412(new_n797, new_n458, new_n798);
nand_5 g00413(new_n798, new_n453, new_n799);
nand_5 g00414(new_n799, new_n447, new_n800);
not_4  g00415(n9589, new_n801);
nor_5  g00416(n10750, new_n801, new_n802);
nor_5  g00417(n10750, n1637, new_n803);
nor_5  g00418(new_n803, new_n802, new_n804);
nor_5  g00419(new_n804, n498, new_n805);
nand_5 g00420(new_n805, new_n800, new_n806);
not_4  g00421(n11404, new_n807);
nor_5  g00422(new_n807, n498, new_n808);
nor_5  g00423(n4175, n3130, new_n809);
not_4  g00424(new_n809, new_n810);
nor_5  g00425(new_n810, new_n808, new_n811);
nand_5 g00426(new_n811, new_n806, new_n812);
nand_5 g00427(new_n812, new_n442, new_n813);
nand_5 g00428(new_n813, new_n437, new_n814);
not_4  g00429(n5023, new_n815);
nor_5  g00430(new_n815, n4225, new_n816);
nor_5  g00431(n6586, n4225, new_n817);
nor_5  g00432(new_n817, new_n816, new_n818);
nor_5  g00433(new_n818, n14483, new_n819);
nand_5 g00434(new_n819, new_n814, new_n820);
nand_5 g00435(new_n820, new_n432, new_n821);
nand_5 g00436(new_n821, new_n427_1, new_n822);
nand_5 g00437(new_n822, new_n422, new_n823);
not_4  g00438(n12976, new_n824);
nor_5  g00439(new_n824, n6810, new_n825);
nor_5  g00440(n12012, n6810, new_n826);
nor_5  g00441(new_n826, new_n825, new_n827);
nor_5  g00442(new_n827, n11756, new_n828);
nand_5 g00443(new_n828, new_n823, new_n829);
not_4  g00444(n666, new_n830);
nor_5  g00445(n11756, new_n830, new_n831);
nor_5  g00446(n13511, n13364, new_n832);
not_4  g00447(new_n832, new_n833);
nor_5  g00448(new_n833, new_n831, new_n834);
nand_5 g00449(new_n834, new_n829, new_n835);
nor_5  g00450(n9026, n3655, new_n836);
not_4  g00451(new_n836, new_n837);
not_4  g00452(n4907, new_n838);
nor_5  g00453(n13364, new_n838, new_n839);
nor_5  g00454(new_n839, new_n837, new_n840);
nand_5 g00455(new_n840, new_n835, new_n841);
nand_5 g00456(new_n841, new_n417, new_n842);
not_4  g00457(n12336, new_n843);
nor_5  g00458(new_n843, n4292, new_n844_1);
nor_5  g00459(n6114, n4292, new_n845);
nor_5  g00460(new_n845, new_n844_1, new_n846);
nor_5  g00461(new_n846, n7272, new_n847);
nand_5 g00462(new_n847, new_n842, new_n848);
not_4  g00463(n7748, new_n849);
not_4  g00464(n7272, new_n850);
nand_5 g00465(n12782, new_n850, new_n851);
nand_5 g00466(new_n851, new_n849, new_n852);
nor_5  g00467(new_n852, n13186, new_n853);
nand_5 g00468(new_n853, new_n848, new_n854);
not_4  g00469(n11854, new_n855);
not_4  g00470(n13186, new_n856);
nand_5 g00471(new_n856, n10278, new_n857);
nand_5 g00472(new_n857, new_n855, new_n858);
nor_5  g00473(new_n858, n702, new_n859);
nand_5 g00474(new_n859, new_n854, new_n860);
nand_5 g00475(new_n860, new_n412, new_n861);
nor_5  g00476(n5077, n674, new_n862);
not_4  g00477(new_n862, new_n863);
not_4  g00478(n8873, new_n864);
nor_5  g00479(new_n864, n3910, new_n865);
nor_5  g00480(new_n865, new_n863, new_n866);
nand_5 g00481(new_n866, new_n861, new_n867);
not_4  g00482(n5467, new_n868);
nor_5  g00483(new_n868, n5077, new_n869);
nor_5  g00484(n13944, n7282, new_n870);
not_4  g00485(new_n870, new_n871);
nor_5  g00486(new_n871, new_n869, new_n872);
nand_5 g00487(new_n872, new_n867, new_n873);
not_4  g00488(n13944, new_n874);
nor_5  g00489(new_n874, n7941, new_n875);
nor_5  g00490(n7941, n6946, new_n876);
nor_5  g00491(new_n876, new_n875, new_n877);
nor_5  g00492(new_n877, n5950, new_n878);
nand_5 g00493(new_n878, new_n873, new_n879);
nand_5 g00494(new_n879, new_n407, new_n880);
not_4  g00495(n10050, new_n881);
nor_5  g00496(new_n881, n4039, new_n882);
nor_5  g00497(n11529, n4039, new_n883);
nor_5  g00498(new_n883, new_n882, new_n884_1);
nor_5  g00499(new_n884_1, n6362, new_n885);
nand_5 g00500(new_n885, new_n880, new_n886);
nand_5 g00501(new_n886, new_n402, new_n887);
nand_5 g00502(new_n887, new_n397, new_n888);
nand_5 g00503(new_n888, new_n392, new_n889);
not_4  g00504(n12270, new_n890);
nor_5  g00505(new_n890, n5601, new_n891);
nor_5  g00506(n5601, n5009, new_n892);
nor_5  g00507(new_n892, new_n891, new_n893);
nor_5  g00508(new_n893, n10426, new_n894);
nand_5 g00509(new_n894, new_n889, new_n895);
nand_5 g00510(new_n895, n13509, new_n896);
nor_5  g00511(new_n896, new_n387, n8);
not_4  g00512(n10378, new_n898);
nor_5  g00513(new_n898, n4282, new_n899);
not_4  g00514(n6758, new_n900);
nand_5 g00515(n6251, new_n760_1, new_n901);
nand_5 g00516(new_n901, new_n900, new_n902);
nor_5  g00517(new_n902, n4282, new_n903);
not_4  g00518(n1702, new_n904);
nand_5 g00519(n9544, new_n904, new_n905);
nand_5 g00520(new_n905, new_n760_1, new_n906);
nor_5  g00521(new_n906, n14072, new_n907);
nor_5  g00522(n5502, n1702, new_n908);
not_4  g00523(new_n908, new_n909);
nand_5 g00524(new_n469, n3166, new_n910);
not_4  g00525(new_n910, new_n911);
nor_5  g00526(new_n911, new_n909, new_n912);
not_4  g00527(n9830, new_n913);
nor_5  g00528(new_n913, n6270, new_n914);
nor_5  g00529(n12321, n8302, new_n915);
not_4  g00530(new_n915, new_n916);
nor_5  g00531(new_n916, new_n914, new_n917);
nor_5  g00532(n7450, n6270, new_n918);
not_4  g00533(new_n918, new_n919);
nand_5 g00534(new_n741, n3972, new_n920);
not_4  g00535(new_n920, new_n921);
nor_5  g00536(new_n921, new_n919, new_n922);
not_4  g00537(n10736, new_n923);
nor_5  g00538(n10945, new_n923, new_n924);
nor_5  g00539(n10615, n7972, new_n925);
not_4  g00540(new_n925, new_n926);
nor_5  g00541(new_n926, new_n924, new_n927);
not_4  g00542(n9555, new_n928);
nand_5 g00543(n6693, new_n474, new_n929);
nand_5 g00544(new_n929, new_n928, new_n930);
nor_5  g00545(new_n930, n10945, new_n931);
not_4  g00546(n12573, new_n932);
nor_5  g00547(n12829, new_n932, new_n933);
nor_5  g00548(n10470, n6555, new_n934);
not_4  g00549(new_n934, new_n935);
nor_5  g00550(new_n935, new_n933, new_n936);
nor_5  g00551(new_n721, new_n480, new_n937);
nor_5  g00552(new_n937, n12829, new_n938);
nand_5 g00553(new_n723, n11158, new_n939);
nand_5 g00554(new_n939, new_n479, new_n940);
nor_5  g00555(new_n940, n10407, new_n941);
nor_5  g00556(new_n714, new_n485, new_n942);
nor_5  g00557(new_n942, n13992, new_n943);
not_4  g00558(n3833, new_n944);
nor_5  g00559(new_n944, n2699, new_n945);
nor_5  g00560(n11590, n6436, new_n946);
not_4  g00561(new_n946, new_n947);
nor_5  g00562(new_n947, new_n945, new_n948_1);
not_4  g00563(n11933, new_n949);
nand_5 g00564(n12885, new_n489, new_n950);
nand_5 g00565(new_n950, new_n949, new_n951);
nor_5  g00566(new_n951, n2699, new_n952);
not_4  g00567(n4117, new_n953);
nor_5  g00568(n11666, new_n953, new_n954);
nor_5  g00569(n10061, n9154, new_n955);
not_4  g00570(new_n955, new_n956);
nor_5  g00571(new_n956, new_n954, new_n957);
not_4  g00572(n8262, new_n958);
nand_5 g00573(new_n494, n10255, new_n959);
nand_5 g00574(new_n959, new_n958, new_n960);
nor_5  g00575(new_n960, n11666, new_n961);
not_4  g00576(n13814, new_n962);
nor_5  g00577(new_n962, n5449, new_n963);
nor_5  g00578(n11875, n4022, new_n964);
not_4  g00579(new_n964, new_n965);
nor_5  g00580(new_n965, new_n963, new_n966);
nor_5  g00581(n5449, n1568, new_n967);
not_4  g00582(new_n967, new_n968);
not_4  g00583(n2895, new_n969);
nor_5  g00584(n8635, new_n969, new_n970);
nor_5  g00585(new_n970, new_n968, new_n971);
not_4  g00586(n203, new_n972);
nor_5  g00587(n737, new_n972, new_n973);
nor_5  g00588(n8635, n5184, new_n974);
not_4  g00589(new_n974, new_n975);
nor_5  g00590(new_n975, new_n973, new_n976);
not_4  g00591(n2454, new_n977_1);
nor_5  g00592(n14293, new_n977_1, new_n978);
nor_5  g00593(n8800, n8044, new_n979);
not_4  g00594(new_n979, new_n980);
nor_5  g00595(new_n980, new_n978, new_n981);
not_4  g00596(n8926, new_n982);
nand_5 g00597(n11269, new_n681, new_n983);
nand_5 g00598(new_n983, new_n982, new_n984);
nor_5  g00599(new_n984, n14293, new_n985);
not_4  g00600(n3506, new_n986);
nor_5  g00601(new_n986, n462, new_n987);
nor_5  g00602(n6703, n3893, new_n988);
not_4  g00603(new_n988, new_n989);
nor_5  g00604(new_n989, new_n987, new_n990);
nor_5  g00605(n4000, n462, new_n991);
not_4  g00606(new_n991, new_n992);
not_4  g00607(n3388, new_n993);
nor_5  g00608(n4154, new_n993, new_n994);
nor_5  g00609(new_n994, new_n992, new_n995);
not_4  g00610(n12614, new_n996);
nor_5  g00611(new_n996, n12142, new_n997);
nor_5  g00612(n10765, n4154, new_n998);
not_4  g00613(new_n998, new_n999);
nor_5  g00614(new_n999, new_n997, new_n1000);
not_4  g00615(n411, new_n1001);
nand_5 g00616(n9252, new_n661, new_n1002);
nand_5 g00617(new_n1002, new_n1001, new_n1003);
nor_5  g00618(new_n1003, n12142, new_n1004);
not_4  g00619(n13093, new_n1005);
nor_5  g00620(new_n1005, n11902, new_n1006);
nor_5  g00621(n8799, n650, new_n1007);
not_4  g00622(new_n1007, new_n1008);
nor_5  g00623(new_n1008, new_n1006, new_n1009);
nor_5  g00624(n10112, n8073, new_n1010);
nor_5  g00625(new_n1010, new_n515, new_n1011);
nor_5  g00626(new_n1011, n11902, new_n1012);
not_4  g00627(n6680, new_n1013);
nor_5  g00628(n10466, new_n1013, new_n1014);
nor_5  g00629(n7652, n3804, new_n1015);
not_4  g00630(new_n1015, new_n1016);
nor_5  g00631(new_n1016, new_n1014, new_n1017);
not_4  g00632(n5943, new_n1018);
nand_5 g00633(new_n524, n2164, new_n1019);
nand_5 g00634(new_n1019, new_n1018, new_n1020);
nor_5  g00635(new_n1020, n10466, new_n1021);
not_4  g00636(n8550, new_n1022);
nor_5  g00637(n14163, new_n1022, new_n1023);
nor_5  g00638(n13882, n5725, new_n1024);
not_4  g00639(new_n1024, new_n1025);
nor_5  g00640(new_n1025, new_n1023, new_n1026);
nor_5  g00641(new_n534, new_n530, new_n1027_1);
nor_5  g00642(new_n1027_1, n14163, new_n1028);
not_4  g00643(n3652, new_n1029);
nor_5  g00644(n13295, new_n1029, new_n1030);
nor_5  g00645(n8746, n3799, new_n1031);
not_4  g00646(new_n1031, new_n1032);
nor_5  g00647(new_n1032, new_n1030, new_n1033);
nor_5  g00648(n10630, n7988, new_n1034);
nor_5  g00649(new_n1034, new_n639, new_n1035);
nor_5  g00650(new_n1035, n13295, new_n1036);
not_4  g00651(n10912, new_n1037);
nand_5 g00652(n11776, new_n1037, new_n1038);
nand_5 g00653(new_n1038, new_n638, new_n1039);
nor_5  g00654(new_n1039, n6873, new_n1040);
nor_5  g00655(n10912, n9543, new_n1041);
not_4  g00656(new_n1041, new_n1042);
nand_5 g00657(n6007, new_n539, new_n1043);
not_4  g00658(new_n1043, new_n1044);
nor_5  g00659(new_n1044, new_n1042, new_n1045);
not_4  g00660(n2334, new_n1046);
nor_5  g00661(n5960, new_n1046, new_n1047);
nor_5  g00662(n3367, n271, new_n1048);
not_4  g00663(new_n1048, new_n1049);
nor_5  g00664(new_n1049, new_n1047, new_n1050);
nor_5  g00665(n6258, n1347, new_n1051);
nor_5  g00666(new_n1051, new_n625, new_n1052);
nor_5  g00667(new_n1052, n5960, new_n1053);
not_4  g00668(n8315, new_n1054);
nand_5 g00669(new_n1054, n5225, new_n1055);
nand_5 g00670(new_n1055, new_n618, new_n1056);
nor_5  g00671(new_n1056, n13890, new_n1057);
not_4  g00672(n13109, new_n1058);
nor_5  g00673(n13231, new_n1058, new_n1059);
nor_5  g00674(n13224, n9110, new_n1060);
not_4  g00675(new_n1060, new_n1061);
nor_5  g00676(new_n1061, new_n1059, new_n1062);
nor_5  g00677(n9314, n4774, new_n1063);
nor_5  g00678(new_n1063, new_n555, new_n1064);
nor_5  g00679(new_n1064, n13231, new_n1065);
not_4  g00680(n7354, new_n1066);
nor_5  g00681(new_n1066, n2573, new_n1067);
nor_5  g00682(n13363, n1763, new_n1068);
not_4  g00683(new_n1068, new_n1069);
nor_5  g00684(new_n1069, new_n1067, new_n1070);
nor_5  g00685(n10573, n2573, new_n1071);
not_4  g00686(new_n1071, new_n1072);
nand_5 g00687(n14475, new_n591, new_n1073);
not_4  g00688(new_n1073, new_n1074);
nor_5  g00689(new_n1074, new_n1072, new_n1075);
not_4  g00690(n7832, new_n1076);
nor_5  g00691(n13625, new_n1076, new_n1077);
nor_5  g00692(n13102, n1776, new_n1078);
not_4  g00693(new_n1078, new_n1079);
nor_5  g00694(new_n1079, new_n1077, new_n1080);
nor_5  g00695(new_n577, n2048, new_n1081);
nor_5  g00696(n11842, n1222, new_n1082);
not_4  g00697(new_n1082, new_n1083);
nor_5  g00698(new_n1083, new_n1081, new_n1084);
nor_5  g00699(n13509, n2201, new_n1085);
not_4  g00700(new_n1085, new_n1086);
nor_5  g00701(new_n1086, new_n387, new_n1087);
nor_5  g00702(n9893, n977, new_n1088);
nor_5  g00703(new_n1088, new_n465, new_n1089);
nand_5 g00704(new_n1089, new_n466, new_n1090);
nand_5 g00705(new_n1090, new_n777, new_n1091);
nand_5 g00706(new_n1091, new_n783, new_n1092);
nand_5 g00707(new_n1092, new_n789, new_n1093_1);
nand_5 g00708(new_n1093_1, new_n463, new_n1094_1);
nand_5 g00709(new_n1094_1, new_n796, new_n1095);
nand_5 g00710(new_n1095, new_n458, new_n1096);
nand_5 g00711(new_n1096, new_n453, new_n1097);
nand_5 g00712(new_n1097, new_n447, new_n1098);
nand_5 g00713(new_n1098, new_n805, new_n1099);
nand_5 g00714(new_n1099, new_n811, new_n1100);
nand_5 g00715(new_n1100, new_n442, new_n1101);
nand_5 g00716(new_n1101, new_n437, new_n1102);
nand_5 g00717(new_n1102, new_n819, new_n1103);
nand_5 g00718(new_n1103, new_n432, new_n1104);
nand_5 g00719(new_n1104, new_n427_1, new_n1105);
nand_5 g00720(new_n1105, new_n422, new_n1106);
nand_5 g00721(new_n1106, new_n828, new_n1107);
nand_5 g00722(new_n1107, new_n834, new_n1108);
nand_5 g00723(new_n1108, new_n840, new_n1109);
nand_5 g00724(new_n1109, new_n417, new_n1110);
nand_5 g00725(new_n1110, new_n847, new_n1111);
nand_5 g00726(new_n1111, new_n853, new_n1112);
nand_5 g00727(new_n1112, new_n859, new_n1113);
nand_5 g00728(new_n1113, new_n412, new_n1114);
nand_5 g00729(new_n1114, new_n866, new_n1115);
nand_5 g00730(new_n1115, new_n872, new_n1116);
nand_5 g00731(new_n1116, new_n878, new_n1117);
nand_5 g00732(new_n1117, new_n407, new_n1118);
nand_5 g00733(new_n1118, new_n885, new_n1119);
nand_5 g00734(new_n1119, new_n402, new_n1120);
nand_5 g00735(new_n1120, new_n397, new_n1121);
nand_5 g00736(new_n1121, new_n392, new_n1122_1);
nand_5 g00737(new_n1122_1, new_n894, new_n1123);
nand_5 g00738(new_n1123, new_n1087, new_n1124_1);
nor_5  g00739(n2166, n2048, new_n1125);
not_4  g00740(new_n1125, new_n1126);
not_4  g00741(n8002, new_n1127);
nor_5  g00742(new_n1127, n2201, new_n1128);
nor_5  g00743(new_n1128, new_n1126, new_n1129);
nand_5 g00744(new_n1129, new_n1124_1, new_n1130);
nand_5 g00745(new_n1130, new_n1084, new_n1131);
nor_5  g00746(n11961, n1027, new_n1132);
nor_5  g00747(new_n1132, new_n565, new_n1133);
nor_5  g00748(new_n1133, n13625, new_n1134);
nand_5 g00749(new_n1134, new_n1131, new_n1135);
nand_5 g00750(new_n1135, new_n1080, new_n1136);
nand_5 g00751(new_n1136, new_n1075, new_n1137);
nand_5 g00752(new_n1137, new_n1070, new_n1138);
nor_5  g00753(n12009, n4755, new_n1139);
not_4  g00754(new_n1139, new_n1140);
nand_5 g00755(n6054, new_n559, new_n1141);
not_4  g00756(new_n1141, new_n1142);
nor_5  g00757(new_n1142, new_n1140, new_n1143);
nand_5 g00758(new_n1143, new_n1138, new_n1144);
not_4  g00759(n4755, new_n1145);
nand_5 g00760(n5033, new_n1145, new_n1146);
nand_5 g00761(new_n1146, new_n554, new_n1147);
nor_5  g00762(new_n1147, n4172, new_n1148);
nand_5 g00763(new_n1148, new_n1144, new_n1149);
nand_5 g00764(new_n1149, new_n1065, new_n1150);
nand_5 g00765(new_n1150, new_n1062, new_n1151);
nor_5  g00766(n11605, n8315, new_n1152);
not_4  g00767(new_n1152, new_n1153);
nand_5 g00768(new_n549, n7104, new_n1154);
not_4  g00769(new_n1154, new_n1155);
nor_5  g00770(new_n1155, new_n1153, new_n1156);
nand_5 g00771(new_n1156, new_n1151, new_n1157);
nand_5 g00772(new_n1157, new_n1057, new_n1158);
nand_5 g00773(new_n1158, new_n1053, new_n1159);
nand_5 g00774(new_n1159, new_n1050, new_n1160);
nand_5 g00775(new_n1160, new_n1045, new_n1161);
nand_5 g00776(new_n1161, new_n1040, new_n1162);
nand_5 g00777(new_n1162, new_n1036, new_n1163);
nand_5 g00778(new_n1163, new_n1033, new_n1164);
nand_5 g00779(new_n1164, new_n1028, new_n1165);
nand_5 g00780(new_n1165, new_n1026, new_n1166);
nand_5 g00781(new_n1166, new_n1021, new_n1167);
nand_5 g00782(new_n1167, new_n1017, new_n1168);
nand_5 g00783(new_n1168, new_n1012, new_n1169);
nand_5 g00784(new_n1169, new_n1009, new_n1170);
nand_5 g00785(new_n1170, new_n1004, new_n1171);
nand_5 g00786(new_n1171, new_n1000, new_n1172);
nand_5 g00787(new_n1172, new_n995, new_n1173);
nand_5 g00788(new_n1173, new_n990, new_n1174);
nand_5 g00789(new_n1174, new_n985, new_n1175);
nand_5 g00790(new_n1175, new_n981, new_n1176);
nor_5  g00791(n8463, n8204, new_n1177);
nor_5  g00792(new_n1177, new_n505, new_n1178);
nor_5  g00793(new_n1178, n737, new_n1179);
nand_5 g00794(new_n1179, new_n1176, new_n1180);
nand_5 g00795(new_n1180, new_n976, new_n1181);
nand_5 g00796(new_n1181, new_n971, new_n1182);
nand_5 g00797(new_n1182, new_n966, new_n1183);
nand_5 g00798(new_n1183, new_n961, new_n1184);
nand_5 g00799(new_n1184, new_n957, new_n1185);
nand_5 g00800(new_n1185, new_n952, new_n1186);
nand_5 g00801(new_n1186, new_n948_1, new_n1187);
nand_5 g00802(new_n1187, new_n943, new_n1188);
nand_5 g00803(new_n1188, new_n941, new_n1189);
nand_5 g00804(new_n1189, new_n938, new_n1190);
nand_5 g00805(new_n1190, new_n936, new_n1191);
nand_5 g00806(new_n1191, new_n931, new_n1192);
nand_5 g00807(new_n1192, new_n927, new_n1193);
nand_5 g00808(new_n1193, new_n922, new_n1194);
nand_5 g00809(new_n1194, new_n917, new_n1195);
nand_5 g00810(new_n1195, new_n912, new_n1196);
nand_5 g00811(new_n1196, new_n907, new_n1197);
nand_5 g00812(new_n1197, new_n903, new_n1198);
nand_5 g00813(new_n1198, n10080, new_n1199);
nor_5  g00814(new_n1199, new_n899, n46);
nor_5  g00815(n13509, n2674, new_n1201);
not_4  g00816(new_n1201, new_n1202);
nor_5  g00817(new_n1202, new_n891, new_n1203);
nor_5  g00818(n5046, n394, new_n1204);
not_4  g00819(new_n1204, new_n1205);
nor_5  g00820(new_n1205, new_n882, new_n1206);
not_4  g00821(new_n883, new_n1207);
not_4  g00822(n5950, new_n1208);
nor_5  g00823(n12927, new_n1208, new_n1209);
nor_5  g00824(new_n1209, new_n1207, new_n1210);
nor_5  g00825(n12927, n8649, new_n1211);
not_4  g00826(new_n1211, new_n1212);
nor_5  g00827(new_n1212, new_n875, new_n1213);
not_4  g00828(n7282, new_n1214);
nor_5  g00829(new_n1214, n6946, new_n1215);
nor_5  g00830(n6946, n5077, new_n1216);
nor_5  g00831(new_n1216, new_n1215, new_n1217);
nor_5  g00832(new_n1217, n7941, new_n1218);
not_4  g00833(n3910, new_n1219);
nor_5  g00834(new_n1219, n674, new_n1220);
nor_5  g00835(n7282, n5467, new_n1221);
not_4  g00836(new_n1221, new_n1222_1);
nor_5  g00837(new_n1222_1, new_n1220, new_n1223);
nor_5  g00838(new_n856, n11854, new_n1224);
nor_5  g00839(n8439, n844, new_n1225);
not_4  g00840(new_n1225, new_n1226);
nor_5  g00841(new_n1226, new_n1224, new_n1227);
nor_5  g00842(n10278, new_n849, new_n1228);
nor_5  g00843(n10278, n7272, new_n1229);
nor_5  g00844(new_n1229, new_n1228, new_n1230);
nor_5  g00845(new_n1230, n11854, new_n1231);
nor_5  g00846(n12782, n7748, new_n1232);
not_4  g00847(new_n1232, new_n1233);
nor_5  g00848(new_n1233, new_n844_1, new_n1234);
not_4  g00849(n6114, new_n1235);
nand_5 g00850(n9186, new_n1235, new_n1236);
not_4  g00851(new_n1236, new_n1237);
nor_5  g00852(n9026, n6114, new_n1238);
nor_5  g00853(new_n1238, new_n1237, new_n1239);
nor_5  g00854(new_n1239, n4292, new_n1240);
not_4  g00855(n3655, new_n1241);
nand_5 g00856(n13364, new_n1241, new_n1242);
nand_5 g00857(new_n1242, new_n413, new_n1243);
nor_5  g00858(new_n1243, n9186, new_n1244);
nor_5  g00859(n4907, n3655, new_n1245);
not_4  g00860(new_n1245, new_n1246);
not_4  g00861(n11756, new_n1247);
nor_5  g00862(n13511, new_n1247, new_n1248);
nor_5  g00863(new_n1248, new_n1246, new_n1249);
nor_5  g00864(n13511, n666, new_n1250);
not_4  g00865(new_n1250, new_n1251);
nor_5  g00866(new_n1251, new_n825, new_n1252);
not_4  g00867(new_n826, new_n1253);
not_4  g00868(n8397, new_n1254);
nor_5  g00869(n14464, new_n1254, new_n1255);
nor_5  g00870(new_n1255, new_n1253, new_n1256);
nor_5  g00871(n14408, n14303, new_n1257);
not_4  g00872(new_n1257, new_n1258);
nor_5  g00873(new_n1258, new_n816, new_n1259);
not_4  g00874(n3673, new_n1260);
nor_5  g00875(n6586, new_n1260, new_n1261);
nor_5  g00876(n6586, n6460, new_n1262);
nor_5  g00877(new_n1262, new_n1261, new_n1263);
nor_5  g00878(new_n1263, n4225, new_n1264);
not_4  g00879(n10446, new_n1265_1);
not_4  g00880(n4175, new_n1266);
nand_5 g00881(new_n1266, n498, new_n1267);
nand_5 g00882(new_n1267, new_n1265_1, new_n1268_1);
nor_5  g00883(new_n1268_1, n13000, new_n1269);
nor_5  g00884(n11404, n4175, new_n1270);
not_4  g00885(new_n1270, new_n1271);
nor_5  g00886(new_n1271, new_n802, new_n1272);
not_4  g00887(n1637, new_n1273);
not_4  g00888(n8552, new_n1274);
nand_5 g00889(new_n1274, n8486, new_n1275);
nand_5 g00890(new_n1275, new_n1273, new_n1276);
nor_5  g00891(new_n1276, n10750, new_n1277);
nor_5  g00892(n6480, n3263, new_n1278);
not_4  g00893(new_n1278, new_n1279);
nor_5  g00894(new_n1279, new_n793, new_n1280);
nor_5  g00895(n4615, n730, new_n1281);
not_4  g00896(new_n1281, new_n1282);
nor_5  g00897(new_n1282, new_n786, new_n1283);
not_4  g00898(new_n787, new_n1284);
not_4  g00899(n2615, new_n1285);
nand_5 g00900(n9936, new_n1285, new_n1286);
not_4  g00901(new_n1286, new_n1287);
nor_5  g00902(new_n1287, new_n1284, new_n1288);
nor_5  g00903(n2615, n1093, new_n1289);
not_4  g00904(new_n1289, new_n1290);
nor_5  g00905(new_n1290, new_n774, new_n1291);
nor_5  g00906(n6517, n427, new_n1292);
not_4  g00907(new_n1292, new_n1293);
nor_5  g00908(new_n1293, new_n767, new_n1294);
nor_5  g00909(n6758, n4282, new_n1295);
nor_5  g00910(new_n1295, new_n899, new_n1296);
nor_5  g00911(new_n1296, n977, new_n1297);
nor_5  g00912(n10378, n4147, new_n1298);
not_4  g00913(new_n1298, new_n1299);
nor_5  g00914(new_n1299, new_n755, new_n1300);
not_4  g00915(new_n756, new_n1301);
not_4  g00916(n5502, new_n1302);
nor_5  g00917(n9544, new_n1302, new_n1303);
nor_5  g00918(new_n1303, new_n1301, new_n1304);
nor_5  g00919(n12321, n9544, new_n1305);
not_4  g00920(new_n1305, new_n1306);
nor_5  g00921(new_n1306, new_n748, new_n1307);
nor_5  g00922(new_n918, new_n914, new_n1308);
nor_5  g00923(new_n1308, n3166, new_n1309);
nor_5  g00924(n10615, n9830, new_n1310);
not_4  g00925(new_n1310, new_n1311);
nor_5  g00926(new_n1311, new_n736, new_n1312);
nor_5  g00927(n10945, n9555, new_n1313);
nor_5  g00928(new_n1313, new_n924, new_n1314);
nor_5  g00929(new_n1314, n3972, new_n1315);
nor_5  g00930(n10736, n6555, new_n1316);
not_4  g00931(new_n1316, new_n1317);
nor_5  g00932(new_n1317, new_n729, new_n1318);
nor_5  g00933(n12829, n4131, new_n1319);
nor_5  g00934(new_n1319, new_n933, new_n1320);
nor_5  g00935(new_n1320, n6693, new_n1321);
not_4  g00936(n10407, new_n1322);
nor_5  g00937(new_n1322, n10051, new_n1323);
nor_5  g00938(n12573, n4659, new_n1324);
not_4  g00939(new_n1324, new_n1325);
nor_5  g00940(new_n1325, new_n1323, new_n1326);
nor_5  g00941(n13992, n10051, new_n1327);
not_4  g00942(new_n1327, new_n1328);
not_4  g00943(n5014, new_n1329_1);
nor_5  g00944(n11158, new_n1329_1, new_n1330);
nor_5  g00945(new_n1330, new_n1328, new_n1331);
nor_5  g00946(n11143, n2699, new_n1332);
not_4  g00947(new_n1332, new_n1333);
not_4  g00948(n11158, new_n1334);
not_4  g00949(n11143, new_n1335);
nand_5 g00950(new_n1335, n6436, new_n1336);
nand_5 g00951(new_n1336, new_n1334, new_n1337);
nor_5  g00952(new_n1337, n11590, new_n1338);
nand_5 g00953(new_n1338, new_n1333, new_n1339);
nand_5 g00954(new_n1339, new_n1331, new_n1340);
nand_5 g00955(new_n1340, new_n1326, new_n1341);
nand_5 g00956(new_n1341, new_n1321, new_n1342);
nand_5 g00957(new_n1342, new_n1318, new_n1343);
nand_5 g00958(new_n1343, new_n1315, new_n1344);
nand_5 g00959(new_n1344, new_n1312, new_n1345);
nand_5 g00960(new_n1345, new_n1309, new_n1346);
nand_5 g00961(new_n1346, new_n1307, new_n1347_1);
nand_5 g00962(new_n1347_1, new_n1304, new_n1348);
nand_5 g00963(new_n1348, new_n1300, new_n1349);
nand_5 g00964(new_n1349, new_n1297, new_n1350);
nand_5 g00965(new_n1350, new_n1294, new_n1351);
not_4  g00966(new_n775, new_n1352);
not_4  g00967(n9893, new_n1353);
nor_5  g00968(new_n1353, n6517, new_n1354);
nor_5  g00969(new_n1354, new_n1352, new_n1355);
nand_5 g00970(new_n1355, new_n1351, new_n1356);
nand_5 g00971(new_n1356, new_n1291, new_n1357);
nand_5 g00972(new_n1357, new_n1288, new_n1358);
nand_5 g00973(new_n1358, new_n1283, new_n1359);
not_4  g00974(new_n794, new_n1360);
not_4  g00975(n4785, new_n1361);
nor_5  g00976(new_n1361, n730, new_n1362);
nor_5  g00977(new_n1362, new_n1360, new_n1363);
nand_5 g00978(new_n1363, new_n1359, new_n1364);
nand_5 g00979(new_n1364, new_n1280, new_n1365);
not_4  g00980(n3263, new_n1366);
nor_5  g00981(n8997, new_n1366, new_n1367);
nor_5  g00982(n8997, n6791, new_n1368);
nor_5  g00983(new_n1368, new_n1367, new_n1369);
nor_5  g00984(new_n1369, n3532, new_n1370);
nand_5 g00985(new_n1370, new_n1365, new_n1371);
nand_5 g00986(new_n450, new_n443, new_n1372);
nor_5  g00987(new_n1372, n8552, new_n1373);
nand_5 g00988(new_n1373, new_n1371, new_n1374);
nand_5 g00989(new_n1374, new_n1277, new_n1375);
nand_5 g00990(new_n1375, new_n1272, new_n1376);
nand_5 g00991(new_n1376, new_n1269, new_n1377);
nor_5  g00992(n12025, n3673, new_n1378);
not_4  g00993(new_n1378, new_n1379);
nor_5  g00994(new_n1379, new_n439, new_n1380);
nand_5 g00995(new_n1380, new_n1377, new_n1381);
nand_5 g00996(new_n1381, new_n1264, new_n1382);
nand_5 g00997(new_n1382, new_n1259, new_n1383);
not_4  g00998(n13636, new_n1384);
not_4  g00999(n14303, new_n1385);
nand_5 g01000(n14483, new_n1385, new_n1386);
nand_5 g01001(new_n1386, new_n1384, new_n1387);
nor_5  g01002(new_n1387, n11930, new_n1388);
nand_5 g01003(new_n1388, new_n1383, new_n1389);
nor_5  g01004(n14464, n10147, new_n1390);
not_4  g01005(new_n1390, new_n1391);
nor_5  g01006(new_n1391, new_n424, new_n1392);
nand_5 g01007(new_n1392, new_n1389, new_n1393);
nand_5 g01008(new_n1393, new_n1256, new_n1394);
nand_5 g01009(new_n1394, new_n1252, new_n1395);
nand_5 g01010(new_n1395, new_n1249, new_n1396);
nand_5 g01011(new_n1396, new_n1244, new_n1397);
nand_5 g01012(new_n1397, new_n1240, new_n1398);
nand_5 g01013(new_n1398, new_n1234, new_n1399);
nand_5 g01014(new_n1399, new_n1231, new_n1400);
nand_5 g01015(new_n1400, new_n1227, new_n1401);
nor_5  g01016(n8873, n674, new_n1402);
not_4  g01017(new_n1402, new_n1403);
not_4  g01018(n844, new_n1404);
nand_5 g01019(new_n1404, n702, new_n1405);
not_4  g01020(new_n1405, new_n1406);
nor_5  g01021(new_n1406, new_n1403, new_n1407);
nand_5 g01022(new_n1407, new_n1401, new_n1408);
nand_5 g01023(new_n1408, new_n1223, new_n1409);
nand_5 g01024(new_n1409, new_n1218, new_n1410);
nand_5 g01025(new_n1410, new_n1213, new_n1411);
nand_5 g01026(new_n1411, new_n1210, new_n1412);
nand_5 g01027(new_n1412, new_n1206, new_n1413);
not_4  g01028(n394, new_n1414);
nor_5  g01029(n8892, new_n1414, new_n1415);
nor_5  g01030(n8892, n6362, new_n1416);
nor_5  g01031(new_n1416, new_n1415, new_n1417);
nor_5  g01032(new_n1417, n1265, new_n1418);
nand_5 g01033(new_n1418, new_n1413, new_n1419);
nor_5  g01034(n8780, n4895, new_n1420);
not_4  g01035(new_n1420, new_n1421);
nor_5  g01036(new_n1421, new_n394_1, new_n1422);
nand_5 g01037(new_n1422, new_n1419, new_n1423);
not_4  g01038(n8780, new_n1424);
nor_5  g01039(new_n1424, n5009, new_n1425);
nor_5  g01040(n8598, n5009, new_n1426);
nor_5  g01041(new_n1426, new_n1425, new_n1427);
nor_5  g01042(new_n1427, n5601, new_n1428);
nand_5 g01043(new_n1428, new_n1423, new_n1429);
nand_5 g01044(new_n1429, new_n1203, new_n1430);
not_4  g01045(n10426, new_n1431);
nor_5  g01046(n13509, new_n1431, new_n1432);
nor_5  g01047(new_n1432, new_n576, new_n1433);
nand_5 g01048(new_n1433, new_n1430, new_n1434);
nand_5 g01049(new_n1434, new_n581, new_n1435);
nand_5 g01050(new_n1435, new_n574, new_n1436);
nand_5 g01051(new_n1436, new_n568, new_n1437);
nand_5 g01052(new_n1437, new_n589, new_n1438);
nand_5 g01053(new_n1438, new_n595, new_n1439);
nand_5 g01054(new_n1439, new_n601, new_n1440);
nand_5 g01055(new_n1440, new_n563, new_n1441);
nand_5 g01056(new_n1441, new_n608, new_n1442);
nand_5 g01057(new_n1442, new_n558, new_n1443);
nand_5 g01058(new_n1443, new_n615, new_n1444);
nand_5 g01059(new_n1444, new_n553, new_n1445);
nand_5 g01060(new_n1445, new_n622, new_n1446);
nand_5 g01061(new_n1446, new_n628, new_n1447);
nand_5 g01062(new_n1447, new_n548, new_n1448);
nand_5 g01063(new_n1448, new_n543_1, new_n1449);
nand_5 g01064(new_n1449, new_n636, new_n1450);
nand_5 g01065(new_n1450, new_n642, new_n1451);
nand_5 g01066(new_n1451, new_n538, new_n1452);
nand_5 g01067(new_n1452, new_n533, new_n1453);
nand_5 g01068(new_n1453, new_n650_1, new_n1454);
nand_5 g01069(new_n1454, new_n528, new_n1455);
nand_5 g01070(new_n1455, new_n523, new_n1456);
nand_5 g01071(new_n1456, new_n518, new_n1457);
nand_5 g01072(new_n1457, new_n659, new_n1458);
nand_5 g01073(new_n1458, new_n665, new_n1459);
nand_5 g01074(new_n1459, new_n672, new_n1460);
nand_5 g01075(new_n1460, new_n513, new_n1461);
nand_5 g01076(new_n1461, new_n679, new_n1462);
nand_5 g01077(new_n1462, new_n685, new_n1463);
nand_5 g01078(new_n1463, new_n691, new_n1464);
nand_5 g01079(new_n1464, new_n508, new_n1465);
nand_5 g01080(new_n1465, new_n698, new_n1466);
nand_5 g01081(new_n1466, new_n503, new_n1467);
nand_5 g01082(new_n1467, new_n704, new_n1468);
nand_5 g01083(new_n1468, new_n498_1, new_n1469);
nand_5 g01084(new_n1469, new_n711, new_n1470);
nand_5 g01085(new_n1470, n3833, new_n1471);
nor_5  g01086(new_n1471, new_n490_1, n91);
nand_5 g01087(new_n960, new_n496, new_n1473);
nand_5 g01088(new_n1473, new_n711, new_n1474);
nand_5 g01089(new_n1474, new_n493, new_n1475);
nand_5 g01090(new_n1475, new_n718, new_n1476);
nand_5 g01091(new_n1476, new_n488, new_n1477);
nand_5 g01092(new_n1477, new_n725, new_n1478);
nand_5 g01093(new_n1478, new_n483, new_n1479);
nand_5 g01094(new_n1479, new_n732, new_n1480);
nand_5 g01095(new_n1480, new_n478, new_n1481);
nand_5 g01096(new_n1481, new_n739, new_n1482);
nand_5 g01097(new_n1482, new_n745, new_n1483);
nand_5 g01098(new_n1483, new_n751, new_n1484);
nand_5 g01099(new_n1484, new_n473, new_n1485);
nand_5 g01100(new_n1485, new_n758, new_n1486);
nand_5 g01101(new_n1486, new_n764, new_n1487);
nand_5 g01102(new_n1487, new_n770, new_n1488);
nand_5 g01103(new_n1488, new_n468, new_n1489);
nand_5 g01104(new_n1489, new_n777, new_n1490);
nand_5 g01105(new_n1490, new_n783, new_n1491);
nand_5 g01106(new_n1491, new_n789, new_n1492);
nand_5 g01107(new_n1492, new_n463, new_n1493);
nand_5 g01108(new_n1493, new_n796, new_n1494);
nand_5 g01109(new_n1494, new_n458, new_n1495);
nand_5 g01110(new_n1495, new_n453, new_n1496);
nand_5 g01111(new_n1496, new_n447, new_n1497);
nand_5 g01112(new_n1497, new_n805, new_n1498);
nand_5 g01113(new_n1498, new_n811, new_n1499);
nand_5 g01114(new_n1499, new_n442, new_n1500);
nand_5 g01115(new_n1500, new_n437, new_n1501);
nand_5 g01116(new_n1501, new_n819, new_n1502);
nand_5 g01117(new_n1502, new_n432, new_n1503);
nand_5 g01118(new_n1503, new_n427_1, new_n1504);
nand_5 g01119(new_n1504, new_n422, new_n1505);
nand_5 g01120(new_n1505, new_n828, new_n1506);
nand_5 g01121(new_n1506, new_n834, new_n1507);
nand_5 g01122(new_n1507, new_n840, new_n1508);
nand_5 g01123(new_n1508, new_n417, new_n1509);
nand_5 g01124(new_n1509, new_n847, new_n1510);
nand_5 g01125(new_n1510, new_n853, new_n1511);
nand_5 g01126(new_n1511, new_n859, new_n1512);
nand_5 g01127(new_n1512, new_n412, new_n1513);
nand_5 g01128(new_n1513, new_n866, new_n1514);
nand_5 g01129(new_n1514, new_n872, new_n1515);
nand_5 g01130(new_n1515, new_n878, new_n1516);
nand_5 g01131(new_n1516, new_n407, new_n1517);
nand_5 g01132(new_n1517, new_n885, new_n1518);
nand_5 g01133(new_n1518, new_n402, new_n1519);
nand_5 g01134(new_n1519, new_n397, new_n1520);
nand_5 g01135(new_n1520, new_n392, new_n1521);
nand_5 g01136(new_n1521, new_n894, new_n1522);
nand_5 g01137(new_n1522, new_n1087, new_n1523);
nand_5 g01138(new_n1523, new_n1129, new_n1524);
nand_5 g01139(new_n1524, new_n1084, new_n1525);
nand_5 g01140(new_n1525, new_n1134, new_n1526);
nand_5 g01141(new_n1526, new_n1080, new_n1527);
nand_5 g01142(new_n1527, new_n1075, new_n1528);
nand_5 g01143(new_n1528, new_n1070, new_n1529);
nand_5 g01144(new_n1529, new_n1143, new_n1530);
nand_5 g01145(new_n1530, new_n1148, new_n1531);
nand_5 g01146(new_n1531, new_n1065, new_n1532);
nand_5 g01147(new_n1532, new_n1062, new_n1533);
nand_5 g01148(new_n1533, new_n1156, new_n1534);
nand_5 g01149(new_n1534, new_n1057, new_n1535);
nand_5 g01150(new_n1535, new_n1053, new_n1536);
nand_5 g01151(new_n1536, new_n1050, new_n1537);
nand_5 g01152(new_n1537, new_n1045, new_n1538);
nand_5 g01153(new_n1538, new_n1040, new_n1539);
nand_5 g01154(new_n1539, new_n1036, new_n1540);
nand_5 g01155(new_n1540, new_n1033, new_n1541);
nand_5 g01156(new_n1541, new_n1028, new_n1542);
nand_5 g01157(new_n1542, new_n1026, new_n1543);
nand_5 g01158(new_n1543, new_n1021, new_n1544);
nand_5 g01159(new_n1544, new_n1017, new_n1545_1);
nand_5 g01160(new_n1545_1, new_n1012, new_n1546);
nand_5 g01161(new_n1546, new_n1009, new_n1547);
nand_5 g01162(new_n1547, new_n1004, new_n1548);
nand_5 g01163(new_n1548, new_n1000, new_n1549);
nand_5 g01164(new_n1549, new_n995, new_n1550);
nand_5 g01165(new_n1550, new_n990, new_n1551);
nand_5 g01166(new_n1551, new_n985, new_n1552);
nand_5 g01167(new_n1552, new_n981, new_n1553);
nand_5 g01168(new_n1553, new_n1179, new_n1554);
nand_5 g01169(new_n1554, new_n976, new_n1555);
nand_5 g01170(new_n1555, new_n971, new_n1556);
nand_5 g01171(new_n1556, n4022, new_n1557);
nor_5  g01172(new_n1557, new_n963, n126);
nor_5  g01173(n11933, n2699, new_n1559);
nor_5  g01174(new_n1559, new_n945, new_n1560);
nor_5  g01175(new_n1560, n11143, new_n1561);
nor_5  g01176(n9154, n3833, new_n1562);
not_4  g01177(new_n1562, new_n1563);
nor_5  g01178(new_n1563, new_n708, new_n1564);
nor_5  g01179(n11666, n8262, new_n1565);
nor_5  g01180(new_n1565, new_n954, new_n1566);
nor_5  g01181(new_n1566, n12885, new_n1567);
nor_5  g01182(n11875, n4117, new_n1568_1);
not_4  g01183(new_n1568_1, new_n1569);
nor_5  g01184(new_n1569, new_n701, new_n1570);
not_4  g01185(new_n702_1, new_n1571);
nor_5  g01186(n13814, new_n500, new_n1572);
nor_5  g01187(new_n1572, new_n1571, new_n1573);
nor_5  g01188(n13814, n8635, new_n1574);
not_4  g01189(new_n1574, new_n1575);
nor_5  g01190(new_n1575, new_n695, new_n1576);
not_4  g01191(n737, new_n1577);
nand_5 g01192(n8463, new_n972, new_n1578);
nand_5 g01193(new_n1578, new_n1577, new_n1579);
nor_5  g01194(new_n1579, n2895, new_n1580);
nor_5  g01195(n8800, n203, new_n1581);
not_4  g01196(new_n1581, new_n1582);
nor_5  g01197(new_n1582, new_n688, new_n1583);
nor_5  g01198(n14293, n8926, new_n1584);
nor_5  g01199(new_n1584, new_n978, new_n1585);
nor_5  g01200(new_n1585, n8204, new_n1586);
nor_5  g01201(n3893, n2454, new_n1587);
not_4  g01202(new_n1587, new_n1588);
nor_5  g01203(new_n1588, new_n676, new_n1589);
nor_5  g01204(new_n669, n3388, new_n1590);
nor_5  g01205(n4154, n3506, new_n1591);
not_4  g01206(new_n1591, new_n1592);
nor_5  g01207(new_n1592, new_n1590, new_n1593);
nor_5  g01208(n12142, n411, new_n1594);
nor_5  g01209(new_n1594, new_n997, new_n1595);
nor_5  g01210(new_n1595, n3388, new_n1596);
nor_5  g01211(n12614, n8799, new_n1597);
not_4  g01212(new_n1597, new_n1598);
nor_5  g01213(new_n1598, new_n656_1, new_n1599);
nor_5  g01214(n11902, n8073, new_n1600);
nor_5  g01215(new_n1600, new_n1006, new_n1601);
nor_5  g01216(new_n1601, n9252, new_n1602);
nor_5  g01217(n13882, n6680, new_n1603);
not_4  g01218(new_n1603, new_n1604);
nor_5  g01219(new_n1604, new_n647, new_n1605);
nor_5  g01220(n14163, n5430, new_n1606);
nor_5  g01221(new_n1606, new_n1023, new_n1607);
nor_5  g01222(new_n1607, n2164, new_n1608);
nor_5  g01223(n13295, n10630, new_n1609);
nor_5  g01224(new_n1609, new_n1030, new_n1610);
nor_5  g01225(new_n1610, n760, new_n1611);
nor_5  g01226(n5185, n3652, new_n1612);
not_4  g01227(new_n1612, new_n1613);
nor_5  g01228(new_n1613, new_n633, new_n1614);
not_4  g01229(n5960, new_n1615);
nand_5 g01230(n6258, new_n1046, new_n1616);
nand_5 g01231(new_n1616, new_n1615, new_n1617);
nor_5  g01232(new_n1617, n6007, new_n1618);
nor_5  g01233(n13890, n2334, new_n1619);
not_4  g01234(new_n1619, new_n1620);
nor_5  g01235(new_n1620, new_n619, new_n1621);
not_4  g01236(new_n620, new_n1622);
not_4  g01237(n11605, new_n1623);
nor_5  g01238(new_n1623, n5225, new_n1624);
nor_5  g01239(new_n1624, new_n1622, new_n1625);
nor_5  g01240(n13224, n5225, new_n1626);
not_4  g01241(new_n1626, new_n1627);
nor_5  g01242(new_n1627, new_n612, new_n1628);
not_4  g01243(new_n613, new_n1629);
nand_5 g01244(new_n1058, n9314, new_n1630);
not_4  g01245(new_n1630, new_n1631);
nor_5  g01246(new_n1631, new_n1629, new_n1632);
nor_5  g01247(n13109, n74, new_n1633);
not_4  g01248(new_n1633, new_n1634);
nor_5  g01249(new_n1634, new_n605, new_n1635);
not_4  g01250(new_n1146, new_n1636);
nor_5  g01251(new_n1636, new_n1139, new_n1637_1);
nor_5  g01252(new_n1637_1, n4774, new_n1638);
nor_5  g01253(n5033, n1763, new_n1639);
not_4  g01254(new_n1639, new_n1640);
nor_5  g01255(new_n1640, new_n598, new_n1641);
nor_5  g01256(new_n1071, new_n1067, new_n1642);
nor_5  g01257(new_n1642, n6054, new_n1643);
nor_5  g01258(n13102, n7354, new_n1644);
not_4  g01259(new_n1644, new_n1645);
nor_5  g01260(new_n1645, new_n586, new_n1646);
nor_5  g01261(n13625, n11961, new_n1647);
nor_5  g01262(new_n1647, new_n1077, new_n1648);
nor_5  g01263(new_n1648, n14475, new_n1649);
nand_5 g01264(new_n570, new_n564, new_n1650);
nor_5  g01265(new_n1650, n7832, new_n1651);
nor_5  g01266(new_n1125, new_n1081, new_n1652);
nor_5  g01267(new_n1652, n1027, new_n1653);
not_4  g01268(n13509, new_n1654);
nor_5  g01269(new_n1654, n8002, new_n1655);
nor_5  g01270(n6147, n2201, new_n1656);
not_4  g01271(new_n1656, new_n1657);
nor_5  g01272(new_n1657, new_n1655, new_n1658);
nor_5  g01273(n10426, n8002, new_n1659);
not_4  g01274(new_n1659, new_n1660);
nand_5 g01275(n5601, new_n386, new_n1661);
not_4  g01276(new_n1661, new_n1662);
nor_5  g01277(new_n1662, new_n1660, new_n1663);
nor_5  g01278(n12270, n2674, new_n1664);
not_4  g01279(new_n1664, new_n1665);
nor_5  g01280(new_n1665, new_n1425, new_n1666);
nor_5  g01281(n8598, n1265, new_n1667);
nor_5  g01282(new_n1667, new_n389_1, new_n1668);
nor_5  g01283(new_n1668, n5009, new_n1669);
nor_5  g01284(n4895, n1268, new_n1670);
not_4  g01285(new_n1670, new_n1671);
nor_5  g01286(new_n1671, new_n1415, new_n1672);
not_4  g01287(new_n1416, new_n1673);
nand_5 g01288(new_n398, n4039, new_n1674);
not_4  g01289(new_n1674, new_n1675);
nor_5  g01290(new_n1675, new_n1673, new_n1676);
not_4  g01291(n11529, new_n1677);
nand_5 g01292(n12927, new_n1677, new_n1678);
nand_5 g01293(new_n1678, new_n398, new_n1679);
nor_5  g01294(new_n1679, n10050, new_n1680);
nor_5  g01295(n11529, n5950, new_n1681);
not_4  g01296(new_n1681, new_n1682);
nand_5 g01297(new_n403, n7941, new_n1683);
not_4  g01298(new_n1683, new_n1684);
nor_5  g01299(new_n1684, new_n1682, new_n1685);
nor_5  g01300(n13944, n8649, new_n1686);
not_4  g01301(new_n1686, new_n1687);
nor_5  g01302(new_n1687, new_n1215, new_n1688);
nor_5  g01303(n8873, new_n1404, new_n1689);
nor_5  g01304(n5467, n3910, new_n1690);
not_4  g01305(new_n1690, new_n1691);
nor_5  g01306(new_n1691, new_n1689, new_n1692);
nor_5  g01307(n11854, n702, new_n1693);
nor_5  g01308(new_n1693, new_n409, new_n1694);
nor_5  g01309(new_n1694, n8873, new_n1695);
nor_5  g01310(n13186, n8439, new_n1696);
not_4  g01311(new_n1696, new_n1697);
nor_5  g01312(new_n1697, new_n1228, new_n1698);
not_4  g01313(new_n851, new_n1699);
nor_5  g01314(n7272, n4292, new_n1700);
nor_5  g01315(new_n1700, new_n1699, new_n1701);
nor_5  g01316(new_n1701, n10278, new_n1702_1);
nand_5 g01317(new_n1236, new_n843, new_n1703);
nor_5  g01318(new_n1703, n12782, new_n1704);
not_4  g01319(n13511, new_n1705);
nor_5  g01320(new_n1705, n4907, new_n1706);
nor_5  g01321(n13364, n2061, new_n1707);
not_4  g01322(new_n1707, new_n1708);
nor_5  g01323(new_n1708, new_n1706, new_n1709);
not_4  g01324(n12012, new_n1710);
nand_5 g01325(n14464, new_n1710, new_n1711);
nand_5 g01326(new_n1711, new_n830, new_n1712);
nor_5  g01327(new_n1712, n12976, new_n1713);
nor_5  g01328(n12012, n8397, new_n1714);
not_4  g01329(new_n1714, new_n1715);
nand_5 g01330(n11930, new_n418, new_n1716);
not_4  g01331(new_n1716, new_n1717);
nor_5  g01332(new_n1717, new_n1715, new_n1718);
nor_5  g01333(new_n1385, n13636, new_n1719);
nor_5  g01334(n10147, n7667, new_n1720);
not_4  g01335(new_n1720, new_n1721);
nor_5  g01336(new_n1721, new_n1719, new_n1722);
not_4  g01337(n14483, new_n1723);
nand_5 g01338(new_n428, n4225, new_n1724);
nand_5 g01339(new_n1724, new_n1723, new_n1725);
nor_5  g01340(new_n1725, n13636, new_n1726);
nor_5  g01341(n14408, n5023, new_n1727);
nand_5 g01342(new_n1727, new_n1263, new_n1728);
nand_5 g01343(new_n1728, new_n1726, new_n1729);
nand_5 g01344(new_n1729, new_n1722, new_n1730);
nand_5 g01345(new_n1730, new_n1718, new_n1731);
nand_5 g01346(new_n1731, new_n1713, new_n1732);
nor_5  g01347(n11756, n4907, new_n1733);
not_4  g01348(new_n1733, new_n1734);
nand_5 g01349(n6810, new_n830, new_n1735);
not_4  g01350(new_n1735, new_n1736);
nor_5  g01351(new_n1736, new_n1734, new_n1737);
nand_5 g01352(new_n1737, new_n1732, new_n1738);
nand_5 g01353(new_n1738, new_n1709, new_n1739_1);
not_4  g01354(new_n1238, new_n1740);
nor_5  g01355(new_n1241, n2061, new_n1741);
nor_5  g01356(new_n1741, new_n1740, new_n1742);
nand_5 g01357(new_n1742, new_n1739_1, new_n1743);
nand_5 g01358(new_n1743, new_n1704, new_n1744);
nand_5 g01359(new_n1744, new_n1702_1, new_n1745);
nand_5 g01360(new_n1745, new_n1698, new_n1746);
nand_5 g01361(new_n1746, new_n1695, new_n1747);
nand_5 g01362(new_n1747, new_n1692, new_n1748);
not_4  g01363(new_n1216, new_n1749);
not_4  g01364(n674, new_n1750);
nor_5  g01365(n5467, new_n1750, new_n1751);
nor_5  g01366(new_n1751, new_n1749, new_n1752);
nand_5 g01367(new_n1752, new_n1748, new_n1753);
nand_5 g01368(new_n1753, new_n1688, new_n1754);
nand_5 g01369(new_n1754, new_n1685, new_n1755);
nand_5 g01370(new_n1755, new_n1680, new_n1756);
nand_5 g01371(new_n1756, new_n1676, new_n1757);
nand_5 g01372(new_n1757, new_n1672, new_n1758);
nand_5 g01373(new_n1758, new_n1669, new_n1759);
nand_5 g01374(new_n1759, new_n1666, new_n1760);
nand_5 g01375(new_n1760, new_n1663, new_n1761);
nand_5 g01376(new_n1761, new_n1658, new_n1762);
nand_5 g01377(new_n1762, new_n1653, new_n1763_1);
nand_5 g01378(new_n1763_1, new_n1651, new_n1764);
nand_5 g01379(new_n1764, new_n1649, new_n1765);
nand_5 g01380(new_n1765, new_n1646, new_n1766);
nand_5 g01381(new_n1766, new_n1643, new_n1767);
nand_5 g01382(new_n1767, new_n1641, new_n1768);
nand_5 g01383(new_n1768, new_n1638, new_n1769);
nand_5 g01384(new_n1769, new_n1635, new_n1770);
nand_5 g01385(new_n1770, new_n1632, new_n1771);
nand_5 g01386(new_n1771, new_n1628, new_n1772);
nand_5 g01387(new_n1772, new_n1625, new_n1773);
nand_5 g01388(new_n1773, new_n1621, new_n1774);
nand_5 g01389(new_n1774, new_n1618, new_n1775);
nor_5  g01390(n11776, n3367, new_n1776_1);
not_4  g01391(new_n1776_1, new_n1777);
nor_5  g01392(new_n1777, new_n545, new_n1778);
nand_5 g01393(new_n1778, new_n1775, new_n1779);
not_4  g01394(new_n1038, new_n1780);
nor_5  g01395(new_n1041, new_n1780, new_n1781);
nor_5  g01396(new_n1781, n7988, new_n1782);
nand_5 g01397(new_n1782, new_n1779, new_n1783);
nand_5 g01398(new_n1783, new_n1614, new_n1784);
nand_5 g01399(new_n1784, new_n1611, new_n1785);
not_4  g01400(n760, new_n1786);
nand_5 g01401(n3799, new_n1786, new_n1787);
nand_5 g01402(new_n1787, new_n1022, new_n1788);
nor_5  g01403(new_n1788, n8746, new_n1789);
nand_5 g01404(new_n1789, new_n1785, new_n1790);
nand_5 g01405(new_n1790, new_n1608, new_n1791);
nand_5 g01406(new_n1791, new_n1605, new_n1792);
nor_5  g01407(n10466, n5943, new_n1793);
nor_5  g01408(new_n1793, new_n1014, new_n1794);
nor_5  g01409(new_n1794, n10112, new_n1795);
nand_5 g01410(new_n1795, new_n1792, new_n1796);
nor_5  g01411(n13093, n7652, new_n1797);
not_4  g01412(new_n1797, new_n1798);
nor_5  g01413(new_n1798, new_n520, new_n1799);
nand_5 g01414(new_n1799, new_n1796, new_n1800);
nand_5 g01415(new_n1800, new_n1602, new_n1801);
nand_5 g01416(new_n1801, new_n1599, new_n1802);
nand_5 g01417(new_n1802, new_n1596, new_n1803);
nand_5 g01418(new_n1803, new_n1593, new_n1804);
nor_5  g01419(new_n991, new_n987, new_n1805);
nor_5  g01420(new_n1805, n11269, new_n1806);
nand_5 g01421(new_n1806, new_n1804, new_n1807);
nand_5 g01422(new_n1807, new_n1589, new_n1808);
nand_5 g01423(new_n1808, new_n1586, new_n1809);
nand_5 g01424(new_n1809, new_n1583, new_n1810);
nand_5 g01425(new_n1810, new_n1580, new_n1811);
nand_5 g01426(new_n1811, new_n1576, new_n1812);
nand_5 g01427(new_n1812, new_n1573, new_n1813);
nand_5 g01428(new_n1813, new_n1570, new_n1814);
nand_5 g01429(new_n1814, new_n1567, new_n1815);
nand_5 g01430(new_n1815, new_n1564, new_n1816);
nand_5 g01431(new_n1816, new_n1561, new_n1817);
nand_5 g01432(new_n1817, new_n1338, new_n1818);
nand_5 g01433(new_n1818, new_n1331, new_n1819);
nand_5 g01434(new_n1819, new_n1326, new_n1820);
nand_5 g01435(new_n1820, new_n1321, new_n1821);
nand_5 g01436(new_n1821, new_n1318, new_n1822);
nand_5 g01437(new_n1822, new_n1315, new_n1823);
nand_5 g01438(new_n1823, new_n1312, new_n1824);
nand_5 g01439(new_n1824, new_n1309, new_n1825);
nand_5 g01440(new_n1825, new_n1307, new_n1826);
nand_5 g01441(new_n1826, new_n1304, new_n1827_1);
nand_5 g01442(new_n1827_1, new_n1300, new_n1828);
nand_5 g01443(new_n1828, new_n1297, new_n1829);
nand_5 g01444(new_n1829, new_n1294, new_n1830);
nand_5 g01445(new_n1830, new_n1355, new_n1831);
nand_5 g01446(new_n1831, new_n1291, new_n1832);
nand_5 g01447(new_n1832, new_n1288, new_n1833);
nand_5 g01448(new_n1833, new_n1283, new_n1834);
nand_5 g01449(new_n1834, new_n1363, new_n1835);
nand_5 g01450(new_n1835, new_n1280, new_n1836);
nand_5 g01451(new_n1836, new_n1370, new_n1837);
nand_5 g01452(new_n1837, new_n1373, new_n1838);
nand_5 g01453(new_n1838, new_n1277, new_n1839);
nand_5 g01454(new_n1839, new_n1272, new_n1840);
nand_5 g01455(new_n1840, new_n1269, new_n1841);
nand_5 g01456(new_n1841, n12025, new_n1842);
nor_5  g01457(new_n1842, new_n439, n278);
not_4  g01458(new_n1242, new_n1844);
nand_5 g01459(new_n1704, new_n1740, new_n1845);
nand_5 g01460(new_n1845, new_n1702_1, new_n1846);
nand_5 g01461(new_n1846, new_n1698, new_n1847);
nand_5 g01462(new_n1847, new_n1695, new_n1848);
nand_5 g01463(new_n1848, new_n1692, new_n1849);
nand_5 g01464(new_n1849, new_n1752, new_n1850);
nand_5 g01465(new_n1850, new_n1688, new_n1851);
nand_5 g01466(new_n1851, new_n1685, new_n1852);
nand_5 g01467(new_n1852, new_n1680, new_n1853);
nand_5 g01468(new_n1853, new_n1676, new_n1854);
nand_5 g01469(new_n1854, new_n1672, new_n1855);
nand_5 g01470(new_n1855, new_n1669, new_n1856);
nand_5 g01471(new_n1856, new_n1666, new_n1857);
nand_5 g01472(new_n1857, new_n1663, new_n1858);
nand_5 g01473(new_n1858, new_n1658, new_n1859);
nand_5 g01474(new_n1859, new_n1653, new_n1860);
nand_5 g01475(new_n1860, new_n1651, new_n1861);
nand_5 g01476(new_n1861, new_n1649, new_n1862);
nand_5 g01477(new_n1862, new_n1646, new_n1863);
nand_5 g01478(new_n1863, new_n1643, new_n1864);
nand_5 g01479(new_n1864, new_n1641, new_n1865);
nand_5 g01480(new_n1865, new_n1638, new_n1866);
nand_5 g01481(new_n1866, new_n1635, new_n1867);
nand_5 g01482(new_n1867, new_n1632, new_n1868);
nand_5 g01483(new_n1868, new_n1628, new_n1869);
nand_5 g01484(new_n1869, new_n1625, new_n1870);
nand_5 g01485(new_n1870, new_n1621, new_n1871);
nand_5 g01486(new_n1871, new_n1618, new_n1872);
nand_5 g01487(new_n1872, new_n1778, new_n1873);
nand_5 g01488(new_n1873, new_n1782, new_n1874);
nand_5 g01489(new_n1874, new_n1614, new_n1875);
nand_5 g01490(new_n1875, new_n1611, new_n1876);
nand_5 g01491(new_n1876, new_n1789, new_n1877);
nand_5 g01492(new_n1877, new_n1608, new_n1878);
nand_5 g01493(new_n1878, new_n1605, new_n1879);
nand_5 g01494(new_n1879, new_n1795, new_n1880);
nand_5 g01495(new_n1880, new_n1799, new_n1881);
nand_5 g01496(new_n1881, new_n1602, new_n1882);
nand_5 g01497(new_n1882, new_n1599, new_n1883);
nand_5 g01498(new_n1883, new_n1596, new_n1884);
nand_5 g01499(new_n1884, new_n1593, new_n1885);
nand_5 g01500(new_n1885, new_n1806, new_n1886);
nand_5 g01501(new_n1886, new_n1589, new_n1887);
nand_5 g01502(new_n1887, new_n1586, new_n1888);
nand_5 g01503(new_n1888, new_n1583, new_n1889);
nand_5 g01504(new_n1889, new_n1580, new_n1890);
nand_5 g01505(new_n1890, new_n1576, new_n1891);
nand_5 g01506(new_n1891, new_n1573, new_n1892);
nand_5 g01507(new_n1892, new_n1570, new_n1893);
nand_5 g01508(new_n1893, new_n1567, new_n1894);
nand_5 g01509(new_n1894, new_n1564, new_n1895);
nand_5 g01510(new_n1895, new_n1561, new_n1896);
nand_5 g01511(new_n1896, new_n1338, new_n1897);
nand_5 g01512(new_n1897, new_n1331, new_n1898);
nand_5 g01513(new_n1898, new_n1326, new_n1899);
nand_5 g01514(new_n1899, new_n1321, new_n1900_1);
nand_5 g01515(new_n1900_1, new_n1318, new_n1901);
nand_5 g01516(new_n1901, new_n1315, new_n1902);
nand_5 g01517(new_n1902, new_n1312, new_n1903);
nand_5 g01518(new_n1903, new_n1309, new_n1904);
nand_5 g01519(new_n1904, new_n1307, new_n1905);
nand_5 g01520(new_n1905, new_n1304, new_n1906);
nand_5 g01521(new_n1906, new_n1300, new_n1907);
nand_5 g01522(new_n1907, new_n1297, new_n1908);
nand_5 g01523(new_n1908, new_n1294, new_n1909);
nand_5 g01524(new_n1909, new_n1355, new_n1910);
nand_5 g01525(new_n1910, new_n1291, new_n1911);
nand_5 g01526(new_n1911, new_n1288, new_n1912);
nand_5 g01527(new_n1912, new_n1283, new_n1913);
nand_5 g01528(new_n1913, new_n1363, new_n1914);
nand_5 g01529(new_n1914, new_n1280, new_n1915);
nand_5 g01530(new_n1915, new_n1370, new_n1916);
nand_5 g01531(new_n1916, new_n1373, new_n1917);
nand_5 g01532(new_n1917, new_n1277, new_n1918);
nand_5 g01533(new_n1918, new_n1272, new_n1919);
nand_5 g01534(new_n1919, new_n1269, new_n1920);
nand_5 g01535(new_n1920, new_n1380, new_n1921);
nand_5 g01536(new_n1921, new_n1264, new_n1922);
nand_5 g01537(new_n1922, new_n1259, new_n1923);
nand_5 g01538(new_n1923, new_n1388, new_n1924);
nand_5 g01539(new_n1924, new_n1392, new_n1925);
nand_5 g01540(new_n1925, new_n1256, new_n1926);
nand_5 g01541(new_n1926, new_n1252, new_n1927_1);
nand_5 g01542(new_n1927_1, new_n1249, new_n1928);
nand_5 g01543(new_n1928, n2061, new_n1929);
nor_5  g01544(new_n1929, new_n1844, n389);
nand_5 g01545(new_n1133, new_n566, new_n1931);
nand_5 g01546(new_n1931, new_n589, new_n1932);
nand_5 g01547(new_n1932, new_n595, new_n1933);
nand_5 g01548(new_n1933, new_n601, new_n1934);
nand_5 g01549(new_n1934, new_n563, new_n1935);
nand_5 g01550(new_n1935, new_n608, new_n1936);
nand_5 g01551(new_n1936, new_n558, new_n1937);
nand_5 g01552(new_n1937, new_n615, new_n1938);
nand_5 g01553(new_n1938, new_n553, new_n1939);
nand_5 g01554(new_n1939, new_n622, new_n1940);
nand_5 g01555(new_n1940, new_n628, new_n1941);
nand_5 g01556(new_n1941, new_n548, new_n1942);
nand_5 g01557(new_n1942, new_n543_1, new_n1943);
nand_5 g01558(new_n1943, new_n636, new_n1944);
nand_5 g01559(new_n1944, new_n642, new_n1945);
nand_5 g01560(new_n1945, new_n538, new_n1946);
nand_5 g01561(new_n1946, new_n533, new_n1947);
nand_5 g01562(new_n1947, new_n650_1, new_n1948);
nand_5 g01563(new_n1948, new_n528, new_n1949);
nand_5 g01564(new_n1949, new_n523, new_n1950);
nand_5 g01565(new_n1950, new_n518, new_n1951_1);
nand_5 g01566(new_n1951_1, new_n659, new_n1952);
nand_5 g01567(new_n1952, new_n665, new_n1953);
nand_5 g01568(new_n1953, new_n672, new_n1954);
nand_5 g01569(new_n1954, new_n513, new_n1955);
nand_5 g01570(new_n1955, new_n679, new_n1956);
nand_5 g01571(new_n1956, new_n685, new_n1957);
nand_5 g01572(new_n1957, new_n691, new_n1958);
nand_5 g01573(new_n1958, new_n508, new_n1959);
nand_5 g01574(new_n1959, new_n698, new_n1960);
nand_5 g01575(new_n1960, new_n503, new_n1961);
nand_5 g01576(new_n1961, new_n704, new_n1962);
nand_5 g01577(new_n1962, new_n498_1, new_n1963);
nand_5 g01578(new_n1963, new_n711, new_n1964);
nand_5 g01579(new_n1964, new_n493, new_n1965);
nand_5 g01580(new_n1965, new_n718, new_n1966);
nand_5 g01581(new_n1966, new_n488, new_n1967);
nand_5 g01582(new_n1967, new_n725, new_n1968);
nand_5 g01583(new_n1968, new_n483, new_n1969);
nand_5 g01584(new_n1969, new_n732, new_n1970);
nand_5 g01585(new_n1970, new_n478, new_n1971);
nand_5 g01586(new_n1971, new_n739, new_n1972);
nand_5 g01587(new_n1972, new_n745, new_n1973);
nand_5 g01588(new_n1973, new_n751, new_n1974);
nand_5 g01589(new_n1974, new_n473, new_n1975);
nand_5 g01590(new_n1975, new_n758, new_n1976);
nand_5 g01591(new_n1976, new_n764, new_n1977);
nand_5 g01592(new_n1977, new_n770, new_n1978);
nand_5 g01593(new_n1978, new_n468, new_n1979);
nand_5 g01594(new_n1979, new_n777, new_n1980);
nand_5 g01595(new_n1980, new_n783, new_n1981);
nand_5 g01596(new_n1981, new_n789, new_n1982);
nand_5 g01597(new_n1982, new_n463, new_n1983);
nand_5 g01598(new_n1983, new_n796, new_n1984);
nand_5 g01599(new_n1984, new_n458, new_n1985);
nand_5 g01600(new_n1985, new_n453, new_n1986);
nand_5 g01601(new_n1986, new_n447, new_n1987);
nand_5 g01602(new_n1987, new_n805, new_n1988);
nand_5 g01603(new_n1988, new_n811, new_n1989);
nand_5 g01604(new_n1989, new_n442, new_n1990);
nand_5 g01605(new_n1990, new_n437, new_n1991);
nand_5 g01606(new_n1991, new_n819, new_n1992);
nand_5 g01607(new_n1992, new_n432, new_n1993);
nand_5 g01608(new_n1993, new_n427_1, new_n1994);
nand_5 g01609(new_n1994, new_n422, new_n1995);
nand_5 g01610(new_n1995, new_n828, new_n1996);
nand_5 g01611(new_n1996, new_n834, new_n1997);
nand_5 g01612(new_n1997, new_n840, new_n1998);
nand_5 g01613(new_n1998, new_n417, new_n1999);
nand_5 g01614(new_n1999, new_n847, new_n2000);
nand_5 g01615(new_n2000, new_n853, new_n2001);
nand_5 g01616(new_n2001, new_n859, new_n2002);
nand_5 g01617(new_n2002, new_n412, new_n2003);
nand_5 g01618(new_n2003, new_n866, new_n2004);
nand_5 g01619(new_n2004, new_n872, new_n2005);
nand_5 g01620(new_n2005, new_n878, new_n2006);
nand_5 g01621(new_n2006, new_n407, new_n2007);
nand_5 g01622(new_n2007, new_n885, new_n2008);
nand_5 g01623(new_n2008, new_n402, new_n2009);
nand_5 g01624(new_n2009, new_n397, new_n2010);
nand_5 g01625(new_n2010, new_n392, new_n2011);
nand_5 g01626(new_n2011, new_n894, new_n2012);
nand_5 g01627(new_n2012, new_n1087, new_n2013);
nand_5 g01628(new_n2013, new_n1129, new_n2014);
nand_5 g01629(new_n2014, n11842, new_n2015);
nor_5  g01630(new_n2015, new_n1081, n451);
not_4  g01631(new_n1727, new_n2017);
nor_5  g01632(new_n2017, new_n1261, new_n2018);
not_4  g01633(new_n1262, new_n2019);
nand_5 g01634(n13000, new_n433, new_n2020);
not_4  g01635(new_n2020, new_n2021);
nor_5  g01636(new_n2021, new_n2019, new_n2022);
nor_5  g01637(n10446, new_n1266, new_n2023);
nor_5  g01638(n12025, n3130, new_n2024);
not_4  g01639(new_n2024, new_n2025);
nor_5  g01640(new_n2025, new_n2023, new_n2026);
nor_5  g01641(n10750, n498, new_n2027_1);
nor_5  g01642(new_n2027_1, new_n808, new_n2028);
nor_5  g01643(new_n2028, n10446, new_n2029);
nor_5  g01644(new_n1274, n1637, new_n2030);
nor_5  g01645(n11404, n9589, new_n2031);
not_4  g01646(new_n2031, new_n2032);
nor_5  g01647(new_n2032, new_n2030, new_n2033);
nor_5  g01648(n8486, n3532, new_n2034);
nor_5  g01649(new_n2034, new_n444, new_n2035);
nor_5  g01650(new_n2035, n1637, new_n2036);
nor_5  g01651(n11345, n5786, new_n2037);
not_4  g01652(new_n2037, new_n2038);
nor_5  g01653(new_n2038, new_n1367, new_n2039);
nor_5  g01654(n10283, n6791, new_n2040);
nor_5  g01655(new_n2040, new_n455, new_n2041);
nor_5  g01656(new_n2041, n8997, new_n2042);
not_4  g01657(n3775, new_n2043);
nand_5 g01658(new_n2043, n730, new_n2044);
nand_5 g01659(new_n2044, new_n454, new_n2045);
nor_5  g01660(new_n2045, n9921, new_n2046);
nor_5  g01661(n4785, n3775, new_n2047);
not_4  g01662(new_n2047, new_n2048_1);
nand_5 g01663(n13561, new_n459, new_n2049);
not_4  g01664(new_n2049, new_n2050);
nor_5  g01665(new_n2050, new_n2048_1, new_n2051);
nor_5  g01666(new_n1285, n656, new_n2052);
nor_5  g01667(n8737, n4615, new_n2053);
not_4  g01668(new_n2053, new_n2054);
nor_5  g01669(new_n2054, new_n2052, new_n2055);
nor_5  g01670(n10862, n9936, new_n2056);
nor_5  g01671(new_n2056, new_n780, new_n2057);
nor_5  g01672(new_n2057, n656, new_n2058);
not_4  g01673(n12218, new_n2059);
nand_5 g01674(new_n2059, n6517, new_n2060);
nand_5 g01675(new_n2060, new_n779, new_n2061_1);
nor_5  g01676(new_n2061_1, n6999, new_n2062);
nor_5  g01677(new_n1089, n12218, new_n2063);
nor_5  g01678(n10080, n427, new_n2064);
not_4  g01679(new_n2064, new_n2065);
nor_5  g01680(new_n2065, new_n899, new_n2066);
nand_5 g01681(new_n919, new_n917, new_n2067);
nand_5 g01682(new_n2067, new_n912, new_n2068);
nand_5 g01683(new_n2068, new_n907, new_n2069);
nand_5 g01684(new_n2069, new_n903, new_n2070);
nand_5 g01685(new_n2070, new_n2066, new_n2071);
nand_5 g01686(new_n2071, new_n2063, new_n2072);
nand_5 g01687(new_n2072, new_n2062, new_n2073);
nand_5 g01688(new_n2073, new_n2058, new_n2074);
nand_5 g01689(new_n2074, new_n2055, new_n2075);
nand_5 g01690(new_n2075, new_n2051, new_n2076);
nand_5 g01691(new_n2076, new_n2046, new_n2077);
nand_5 g01692(new_n2077, new_n2042, new_n2078);
nand_5 g01693(new_n2078, new_n2039, new_n2079);
nand_5 g01694(new_n2079, new_n2036, new_n2080);
nand_5 g01695(new_n2080, new_n2033, new_n2081);
nand_5 g01696(new_n2081, new_n2029, new_n2082);
nand_5 g01697(new_n2082, new_n2026, new_n2083);
nand_5 g01698(new_n2083, new_n2022, new_n2084);
nand_5 g01699(new_n2084, new_n2018, new_n2085);
nand_5 g01700(new_n2085, new_n1726, new_n2086);
nand_5 g01701(new_n2086, new_n1722, new_n2087);
nand_5 g01702(new_n2087, new_n1718, new_n2088);
nand_5 g01703(new_n2088, new_n1713, new_n2089);
nand_5 g01704(new_n2089, new_n1737, new_n2090);
nand_5 g01705(new_n2090, new_n1709, new_n2091);
nand_5 g01706(new_n2091, new_n1742, new_n2092);
nand_5 g01707(new_n2092, new_n1704, new_n2093);
nand_5 g01708(new_n2093, new_n1702_1, new_n2094);
nand_5 g01709(new_n2094, new_n1698, new_n2095);
nand_5 g01710(new_n2095, new_n1695, new_n2096);
nand_5 g01711(new_n2096, new_n1692, new_n2097);
nand_5 g01712(new_n2097, new_n1752, new_n2098);
nand_5 g01713(new_n2098, new_n1688, new_n2099);
nand_5 g01714(new_n2099, new_n1685, new_n2100);
nand_5 g01715(new_n2100, new_n1680, new_n2101);
nand_5 g01716(new_n2101, new_n1676, new_n2102);
nand_5 g01717(new_n2102, new_n1672, new_n2103);
nand_5 g01718(new_n2103, new_n1669, new_n2104);
nand_5 g01719(new_n2104, new_n1666, new_n2105);
nand_5 g01720(new_n2105, new_n1663, new_n2106);
nand_5 g01721(new_n2106, new_n1658, new_n2107);
nand_5 g01722(new_n2107, new_n1653, new_n2108);
nand_5 g01723(new_n2108, new_n1651, new_n2109);
nand_5 g01724(new_n2109, new_n1649, new_n2110);
nand_5 g01725(new_n2110, new_n1646, new_n2111);
nand_5 g01726(new_n2111, new_n1643, new_n2112);
nand_5 g01727(new_n2112, new_n1641, new_n2113);
nand_5 g01728(new_n2113, new_n1638, new_n2114);
nand_5 g01729(new_n2114, new_n1635, new_n2115);
nand_5 g01730(new_n2115, new_n1632, new_n2116);
nand_5 g01731(new_n2116, new_n1628, new_n2117);
nand_5 g01732(new_n2117, new_n1625, new_n2118);
nand_5 g01733(new_n2118, new_n1621, new_n2119);
nand_5 g01734(new_n2119, new_n1618, new_n2120);
nand_5 g01735(new_n2120, new_n1778, new_n2121);
nand_5 g01736(new_n2121, new_n1782, new_n2122);
nand_5 g01737(new_n2122, new_n1614, new_n2123);
nand_5 g01738(new_n2123, new_n1611, new_n2124);
nand_5 g01739(new_n2124, new_n1789, new_n2125);
nand_5 g01740(new_n2125, new_n1608, new_n2126_1);
nand_5 g01741(new_n2126_1, new_n1605, new_n2127);
nand_5 g01742(new_n2127, new_n1795, new_n2128);
nand_5 g01743(new_n2128, new_n1799, new_n2129);
nand_5 g01744(new_n2129, new_n1602, new_n2130);
nand_5 g01745(new_n2130, new_n1599, new_n2131);
nand_5 g01746(new_n2131, new_n1596, new_n2132);
nand_5 g01747(new_n2132, new_n1593, new_n2133);
nand_5 g01748(new_n2133, new_n1806, new_n2134);
nand_5 g01749(new_n2134, new_n1589, new_n2135);
nand_5 g01750(new_n2135, new_n1586, new_n2136);
nand_5 g01751(new_n2136, new_n1583, new_n2137);
nand_5 g01752(new_n2137, new_n1580, new_n2138);
nand_5 g01753(new_n2138, new_n1576, new_n2139);
nand_5 g01754(new_n2139, new_n1573, new_n2140);
nand_5 g01755(new_n2140, new_n1570, new_n2141);
nand_5 g01756(new_n2141, new_n1567, new_n2142);
nand_5 g01757(new_n2142, new_n1564, new_n2143);
nand_5 g01758(new_n2143, new_n1561, new_n2144);
nand_5 g01759(new_n2144, new_n1338, new_n2145);
nand_5 g01760(new_n2145, new_n1331, new_n2146);
nand_5 g01761(new_n2146, new_n1326, new_n2147);
nand_5 g01762(new_n2147, new_n1321, new_n2148);
nand_5 g01763(new_n2148, new_n1318, new_n2149);
nand_5 g01764(new_n2149, new_n1315, new_n2150);
nand_5 g01765(new_n2150, n10615, new_n2151);
nor_5  g01766(new_n2151, new_n736, n490);
not_4  g01767(new_n1609, new_n2153);
nand_5 g01768(new_n2153, new_n1033, new_n2154);
nand_5 g01769(new_n2154, new_n1028, new_n2155);
nand_5 g01770(new_n2155, new_n1026, new_n2156);
nand_5 g01771(new_n2156, new_n1021, new_n2157);
nand_5 g01772(new_n2157, new_n1017, new_n2158);
nand_5 g01773(new_n2158, new_n1012, new_n2159);
nand_5 g01774(new_n2159, new_n1009, new_n2160);
nand_5 g01775(new_n2160, new_n1004, new_n2161);
nand_5 g01776(new_n2161, new_n1000, new_n2162);
nand_5 g01777(new_n2162, new_n995, new_n2163);
nand_5 g01778(new_n2163, new_n990, new_n2164_1);
nand_5 g01779(new_n2164_1, new_n985, new_n2165);
nand_5 g01780(new_n2165, new_n981, new_n2166_1);
nand_5 g01781(new_n2166_1, new_n1179, new_n2167);
nand_5 g01782(new_n2167, new_n976, new_n2168);
nand_5 g01783(new_n2168, new_n971, new_n2169);
nand_5 g01784(new_n2169, new_n966, new_n2170);
nand_5 g01785(new_n2170, new_n961, new_n2171);
nand_5 g01786(new_n2171, new_n957, new_n2172);
nand_5 g01787(new_n2172, new_n952, new_n2173);
nand_5 g01788(new_n2173, new_n948_1, new_n2174);
nand_5 g01789(new_n2174, new_n943, new_n2175_1);
nand_5 g01790(new_n2175_1, new_n941, new_n2176);
nand_5 g01791(new_n2176, new_n938, new_n2177);
nand_5 g01792(new_n2177, new_n936, new_n2178);
nand_5 g01793(new_n2178, new_n931, new_n2179);
nand_5 g01794(new_n2179, new_n927, new_n2180);
nand_5 g01795(new_n2180, new_n922, new_n2181);
nand_5 g01796(new_n2181, new_n917, new_n2182);
nand_5 g01797(new_n2182, new_n912, new_n2183);
nand_5 g01798(new_n2183, new_n907, new_n2184);
nand_5 g01799(new_n2184, new_n903, new_n2185);
nand_5 g01800(new_n2185, new_n2066, new_n2186);
nand_5 g01801(new_n2186, new_n2063, new_n2187);
nand_5 g01802(new_n2187, new_n2062, new_n2188);
nand_5 g01803(new_n2188, new_n2058, new_n2189);
nand_5 g01804(new_n2189, new_n2055, new_n2190);
nand_5 g01805(new_n2190, new_n2051, new_n2191);
nand_5 g01806(new_n2191, new_n2046, new_n2192);
nand_5 g01807(new_n2192, new_n2042, new_n2193);
nand_5 g01808(new_n2193, new_n2039, new_n2194);
nand_5 g01809(new_n2194, new_n2036, new_n2195);
nand_5 g01810(new_n2195, new_n2033, new_n2196);
nand_5 g01811(new_n2196, new_n2029, new_n2197);
nand_5 g01812(new_n2197, new_n2026, new_n2198);
nand_5 g01813(new_n2198, new_n2022, new_n2199);
nand_5 g01814(new_n2199, new_n2018, new_n2200);
nand_5 g01815(new_n2200, new_n1726, new_n2201_1);
nand_5 g01816(new_n2201_1, new_n1722, new_n2202);
nand_5 g01817(new_n2202, new_n1718, new_n2203);
nand_5 g01818(new_n2203, new_n1713, new_n2204);
nand_5 g01819(new_n2204, new_n1737, new_n2205);
nand_5 g01820(new_n2205, new_n1709, new_n2206);
nand_5 g01821(new_n2206, new_n1742, new_n2207);
nand_5 g01822(new_n2207, new_n1704, new_n2208);
nand_5 g01823(new_n2208, new_n1702_1, new_n2209);
nand_5 g01824(new_n2209, new_n1698, new_n2210);
nand_5 g01825(new_n2210, new_n1695, new_n2211);
nand_5 g01826(new_n2211, new_n1692, new_n2212);
nand_5 g01827(new_n2212, new_n1752, new_n2213);
nand_5 g01828(new_n2213, new_n1688, new_n2214);
nand_5 g01829(new_n2214, new_n1685, new_n2215);
nand_5 g01830(new_n2215, new_n1680, new_n2216);
nand_5 g01831(new_n2216, new_n1676, new_n2217);
nand_5 g01832(new_n2217, new_n1672, new_n2218);
nand_5 g01833(new_n2218, new_n1669, new_n2219);
nand_5 g01834(new_n2219, new_n1666, new_n2220);
nand_5 g01835(new_n2220, new_n1663, new_n2221);
nand_5 g01836(new_n2221, new_n1658, new_n2222);
nand_5 g01837(new_n2222, new_n1653, new_n2223_1);
nand_5 g01838(new_n2223_1, new_n1651, new_n2224);
nand_5 g01839(new_n2224, new_n1649, new_n2225);
nand_5 g01840(new_n2225, new_n1646, new_n2226);
nand_5 g01841(new_n2226, new_n1643, new_n2227);
nand_5 g01842(new_n2227, new_n1641, new_n2228);
nand_5 g01843(new_n2228, new_n1638, new_n2229);
nand_5 g01844(new_n2229, new_n1635, new_n2230);
nand_5 g01845(new_n2230, new_n1632, new_n2231);
nand_5 g01846(new_n2231, new_n1628, new_n2232);
nand_5 g01847(new_n2232, new_n1625, new_n2233);
nand_5 g01848(new_n2233, new_n1621, new_n2234);
nand_5 g01849(new_n2234, new_n1618, new_n2235);
nand_5 g01850(new_n2235, new_n1778, new_n2236);
nand_5 g01851(new_n2236, new_n1782, new_n2237);
nand_5 g01852(new_n2237, n5185, new_n2238);
nor_5  g01853(new_n2238, new_n633, n543);
nand_5 g01854(new_n1633, new_n607, new_n2240);
nand_5 g01855(new_n2240, new_n1632, new_n2241);
nand_5 g01856(new_n2241, new_n1628, new_n2242);
nand_5 g01857(new_n2242, new_n1625, new_n2243);
nand_5 g01858(new_n2243, new_n1621, new_n2244);
nand_5 g01859(new_n2244, new_n1618, new_n2245);
nand_5 g01860(new_n2245, new_n1778, new_n2246);
nand_5 g01861(new_n2246, new_n1782, new_n2247);
nand_5 g01862(new_n2247, new_n1614, new_n2248);
nand_5 g01863(new_n2248, new_n1611, new_n2249);
nand_5 g01864(new_n2249, new_n1789, new_n2250);
nand_5 g01865(new_n2250, new_n1608, new_n2251);
nand_5 g01866(new_n2251, new_n1605, new_n2252);
nand_5 g01867(new_n2252, new_n1795, new_n2253);
nand_5 g01868(new_n2253, new_n1799, new_n2254);
nand_5 g01869(new_n2254, new_n1602, new_n2255);
nand_5 g01870(new_n2255, new_n1599, new_n2256);
nand_5 g01871(new_n2256, new_n1596, new_n2257);
nand_5 g01872(new_n2257, new_n1593, new_n2258);
nand_5 g01873(new_n2258, new_n1806, new_n2259);
nand_5 g01874(new_n2259, new_n1589, new_n2260);
nand_5 g01875(new_n2260, new_n1586, new_n2261);
nand_5 g01876(new_n2261, new_n1583, new_n2262);
nand_5 g01877(new_n2262, new_n1580, new_n2263);
nand_5 g01878(new_n2263, new_n1576, new_n2264);
nand_5 g01879(new_n2264, new_n1573, new_n2265);
nand_5 g01880(new_n2265, new_n1570, new_n2266);
nand_5 g01881(new_n2266, new_n1567, new_n2267);
nand_5 g01882(new_n2267, new_n1564, new_n2268);
nand_5 g01883(new_n2268, new_n1561, new_n2269);
nand_5 g01884(new_n2269, new_n1338, new_n2270);
nand_5 g01885(new_n2270, new_n1331, new_n2271);
nand_5 g01886(new_n2271, new_n1326, new_n2272);
nand_5 g01887(new_n2272, new_n1321, new_n2273);
nand_5 g01888(new_n2273, new_n1318, new_n2274);
nand_5 g01889(new_n2274, new_n1315, new_n2275);
nand_5 g01890(new_n2275, new_n1312, new_n2276);
nand_5 g01891(new_n2276, new_n1309, new_n2277);
nand_5 g01892(new_n2277, new_n1307, new_n2278);
nand_5 g01893(new_n2278, new_n1304, new_n2279);
nand_5 g01894(new_n2279, new_n1300, new_n2280);
nand_5 g01895(new_n2280, new_n1297, new_n2281);
nand_5 g01896(new_n2281, new_n1294, new_n2282);
nand_5 g01897(new_n2282, new_n1355, new_n2283);
nand_5 g01898(new_n2283, new_n1291, new_n2284);
nand_5 g01899(new_n2284, new_n1288, new_n2285);
nand_5 g01900(new_n2285, new_n1283, new_n2286);
nand_5 g01901(new_n2286, new_n1363, new_n2287);
nand_5 g01902(new_n2287, new_n1280, new_n2288);
nand_5 g01903(new_n2288, new_n1370, new_n2289);
nand_5 g01904(new_n2289, new_n1373, new_n2290);
nand_5 g01905(new_n2290, new_n1277, new_n2291);
nand_5 g01906(new_n2291, new_n1272, new_n2292);
nand_5 g01907(new_n2292, new_n1269, new_n2293);
nand_5 g01908(new_n2293, new_n1380, new_n2294);
nand_5 g01909(new_n2294, new_n1264, new_n2295);
nand_5 g01910(new_n2295, new_n1259, new_n2296);
nand_5 g01911(new_n2296, new_n1388, new_n2297);
nand_5 g01912(new_n2297, new_n1392, new_n2298);
nand_5 g01913(new_n2298, new_n1256, new_n2299);
nand_5 g01914(new_n2299, new_n1252, new_n2300);
nand_5 g01915(new_n2300, new_n1249, new_n2301);
nand_5 g01916(new_n2301, new_n1244, new_n2302);
nand_5 g01917(new_n2302, new_n1240, new_n2303);
nand_5 g01918(new_n2303, new_n1234, new_n2304);
nand_5 g01919(new_n2304, new_n1231, new_n2305);
nand_5 g01920(new_n2305, new_n1227, new_n2306);
nand_5 g01921(new_n2306, new_n1407, new_n2307);
nand_5 g01922(new_n2307, new_n1223, new_n2308);
nand_5 g01923(new_n2308, new_n1218, new_n2309);
nand_5 g01924(new_n2309, new_n1213, new_n2310);
nand_5 g01925(new_n2310, new_n1210, new_n2311_1);
nand_5 g01926(new_n2311_1, new_n1206, new_n2312);
nand_5 g01927(new_n2312, new_n1418, new_n2313);
nand_5 g01928(new_n2313, new_n1422, new_n2314);
nand_5 g01929(new_n2314, new_n1428, new_n2315);
nand_5 g01930(new_n2315, new_n1203, new_n2316);
nand_5 g01931(new_n2316, new_n1433, new_n2317);
nand_5 g01932(new_n2317, new_n581, new_n2318);
nand_5 g01933(new_n2318, new_n574, new_n2319);
nand_5 g01934(new_n2319, new_n568, new_n2320);
nand_5 g01935(new_n2320, new_n589, new_n2321);
nand_5 g01936(new_n2321, new_n595, new_n2322);
nand_5 g01937(new_n2322, new_n601, new_n2323);
nand_5 g01938(new_n2323, n5033, new_n2324);
nor_5  g01939(new_n2324, new_n560, n682);
nand_5 g01940(new_n1153, new_n1057, new_n2326);
nand_5 g01941(new_n2326, new_n1053, new_n2327);
nand_5 g01942(new_n2327, new_n1050, new_n2328);
nand_5 g01943(new_n2328, new_n1045, new_n2329);
nand_5 g01944(new_n2329, new_n1040, new_n2330);
nand_5 g01945(new_n2330, new_n1036, new_n2331);
nand_5 g01946(new_n2331, new_n1033, new_n2332);
nand_5 g01947(new_n2332, new_n1028, new_n2333);
nand_5 g01948(new_n2333, new_n1026, new_n2334_1);
nand_5 g01949(new_n2334_1, new_n1021, new_n2335);
nand_5 g01950(new_n2335, new_n1017, new_n2336);
nand_5 g01951(new_n2336, new_n1012, new_n2337);
nand_5 g01952(new_n2337, new_n1009, new_n2338);
nand_5 g01953(new_n2338, new_n1004, new_n2339);
nand_5 g01954(new_n2339, new_n1000, new_n2340);
nand_5 g01955(new_n2340, new_n995, new_n2341);
nand_5 g01956(new_n2341, new_n990, new_n2342);
nand_5 g01957(new_n2342, new_n985, new_n2343);
nand_5 g01958(new_n2343, new_n981, new_n2344);
nand_5 g01959(new_n2344, new_n1179, new_n2345);
nand_5 g01960(new_n2345, new_n976, new_n2346);
nand_5 g01961(new_n2346, new_n971, new_n2347);
nand_5 g01962(new_n2347, new_n966, new_n2348);
nand_5 g01963(new_n2348, new_n961, new_n2349);
nand_5 g01964(new_n2349, new_n957, new_n2350);
nand_5 g01965(new_n2350, new_n952, new_n2351);
nand_5 g01966(new_n2351, new_n948_1, new_n2352);
nand_5 g01967(new_n2352, new_n943, new_n2353);
nand_5 g01968(new_n2353, new_n941, new_n2354);
nand_5 g01969(new_n2354, new_n938, new_n2355);
nand_5 g01970(new_n2355, new_n936, new_n2356);
nand_5 g01971(new_n2356, new_n931, new_n2357);
nand_5 g01972(new_n2357, new_n927, new_n2358);
nand_5 g01973(new_n2358, new_n922, new_n2359);
nand_5 g01974(new_n2359, new_n917, new_n2360);
nand_5 g01975(new_n2360, new_n912, new_n2361);
nand_5 g01976(new_n2361, new_n907, new_n2362);
nand_5 g01977(new_n2362, new_n903, new_n2363);
nand_5 g01978(new_n2363, new_n2066, new_n2364);
nand_5 g01979(new_n2364, new_n2063, new_n2365);
nand_5 g01980(new_n2365, new_n2062, new_n2366);
nand_5 g01981(new_n2366, new_n2058, new_n2367);
nand_5 g01982(new_n2367, new_n2055, new_n2368);
nand_5 g01983(new_n2368, new_n2051, new_n2369);
nand_5 g01984(new_n2369, new_n2046, new_n2370);
nand_5 g01985(new_n2370, new_n2042, new_n2371);
nand_5 g01986(new_n2371, new_n2039, new_n2372);
nand_5 g01987(new_n2372, new_n2036, new_n2373);
nand_5 g01988(new_n2373, new_n2033, new_n2374);
nand_5 g01989(new_n2374, new_n2029, new_n2375);
nand_5 g01990(new_n2375, new_n2026, new_n2376);
nand_5 g01991(new_n2376, new_n2022, new_n2377);
nand_5 g01992(new_n2377, new_n2018, new_n2378);
nand_5 g01993(new_n2378, new_n1726, new_n2379);
nand_5 g01994(new_n2379, new_n1722, new_n2380);
nand_5 g01995(new_n2380, new_n1718, new_n2381);
nand_5 g01996(new_n2381, new_n1713, new_n2382);
nand_5 g01997(new_n2382, new_n1737, new_n2383);
nand_5 g01998(new_n2383, new_n1709, new_n2384);
nand_5 g01999(new_n2384, new_n1742, new_n2385);
nand_5 g02000(new_n2385, new_n1704, new_n2386);
nand_5 g02001(new_n2386, new_n1702_1, new_n2387);
nand_5 g02002(new_n2387, new_n1698, new_n2388);
nand_5 g02003(new_n2388, new_n1695, new_n2389);
nand_5 g02004(new_n2389, new_n1692, new_n2390);
nand_5 g02005(new_n2390, new_n1752, new_n2391);
nand_5 g02006(new_n2391, new_n1688, new_n2392);
nand_5 g02007(new_n2392, new_n1685, new_n2393);
nand_5 g02008(new_n2393, new_n1680, new_n2394);
nand_5 g02009(new_n2394, new_n1676, new_n2395);
nand_5 g02010(new_n2395, new_n1672, new_n2396);
nand_5 g02011(new_n2396, new_n1669, new_n2397);
nand_5 g02012(new_n2397, new_n1666, new_n2398);
nand_5 g02013(new_n2398, new_n1663, new_n2399);
nand_5 g02014(new_n2399, new_n1658, new_n2400);
nand_5 g02015(new_n2400, new_n1653, new_n2401);
nand_5 g02016(new_n2401, new_n1651, new_n2402);
nand_5 g02017(new_n2402, new_n1649, new_n2403);
nand_5 g02018(new_n2403, new_n1646, new_n2404);
nand_5 g02019(new_n2404, new_n1643, new_n2405);
nand_5 g02020(new_n2405, new_n1641, new_n2406);
nand_5 g02021(new_n2406, new_n1638, new_n2407_1);
nand_5 g02022(new_n2407_1, new_n1635, new_n2408);
nand_5 g02023(new_n2408, new_n1632, new_n2409);
nand_5 g02024(new_n2409, n13224, new_n2410);
nor_5  g02025(new_n2410, new_n612, n884);
nand_5 g02026(new_n1660, new_n1658, new_n2412);
nand_5 g02027(new_n2412, new_n1653, new_n2413);
nand_5 g02028(new_n2413, new_n1651, new_n2414);
nand_5 g02029(new_n2414, new_n1649, new_n2415);
nand_5 g02030(new_n2415, new_n1646, new_n2416);
nand_5 g02031(new_n2416, new_n1643, new_n2417);
nand_5 g02032(new_n2417, new_n1641, new_n2418);
nand_5 g02033(new_n2418, new_n1638, new_n2419);
nand_5 g02034(new_n2419, new_n1635, new_n2420);
nand_5 g02035(new_n2420, new_n1632, new_n2421);
nand_5 g02036(new_n2421, new_n1628, new_n2422);
nand_5 g02037(new_n2422, new_n1625, new_n2423);
nand_5 g02038(new_n2423, new_n1621, new_n2424);
nand_5 g02039(new_n2424, new_n1618, new_n2425);
nand_5 g02040(new_n2425, new_n1778, new_n2426);
nand_5 g02041(new_n2426, new_n1782, new_n2427);
nand_5 g02042(new_n2427, new_n1614, new_n2428);
nand_5 g02043(new_n2428, new_n1611, new_n2429);
nand_5 g02044(new_n2429, new_n1789, new_n2430);
nand_5 g02045(new_n2430, new_n1608, new_n2431);
nand_5 g02046(new_n2431, new_n1605, new_n2432);
nand_5 g02047(new_n2432, new_n1795, new_n2433);
nand_5 g02048(new_n2433, new_n1799, new_n2434);
nand_5 g02049(new_n2434, new_n1602, new_n2435);
nand_5 g02050(new_n2435, new_n1599, new_n2436);
nand_5 g02051(new_n2436, new_n1596, new_n2437);
nand_5 g02052(new_n2437, new_n1593, new_n2438);
nand_5 g02053(new_n2438, new_n1806, new_n2439);
nand_5 g02054(new_n2439, new_n1589, new_n2440);
nand_5 g02055(new_n2440, new_n1586, new_n2441);
nand_5 g02056(new_n2441, new_n1583, new_n2442);
nand_5 g02057(new_n2442, new_n1580, new_n2443);
nand_5 g02058(new_n2443, new_n1576, new_n2444);
nand_5 g02059(new_n2444, new_n1573, new_n2445);
nand_5 g02060(new_n2445, new_n1570, new_n2446);
nand_5 g02061(new_n2446, new_n1567, new_n2447);
nand_5 g02062(new_n2447, new_n1564, new_n2448);
nand_5 g02063(new_n2448, new_n1561, new_n2449);
nand_5 g02064(new_n2449, new_n1338, new_n2450);
nand_5 g02065(new_n2450, new_n1331, new_n2451);
nand_5 g02066(new_n2451, new_n1326, new_n2452);
nand_5 g02067(new_n2452, new_n1321, new_n2453);
nand_5 g02068(new_n2453, new_n1318, new_n2454_1);
nand_5 g02069(new_n2454_1, new_n1315, new_n2455);
nand_5 g02070(new_n2455, new_n1312, new_n2456);
nand_5 g02071(new_n2456, new_n1309, new_n2457);
nand_5 g02072(new_n2457, new_n1307, new_n2458);
nand_5 g02073(new_n2458, new_n1304, new_n2459);
nand_5 g02074(new_n2459, new_n1300, new_n2460);
nand_5 g02075(new_n2460, new_n1297, new_n2461);
nand_5 g02076(new_n2461, new_n1294, new_n2462);
nand_5 g02077(new_n2462, new_n1355, new_n2463);
nand_5 g02078(new_n2463, new_n1291, new_n2464);
nand_5 g02079(new_n2464, new_n1288, new_n2465);
nand_5 g02080(new_n2465, new_n1283, new_n2466);
nand_5 g02081(new_n2466, new_n1363, new_n2467);
nand_5 g02082(new_n2467, new_n1280, new_n2468);
nand_5 g02083(new_n2468, new_n1370, new_n2469);
nand_5 g02084(new_n2469, new_n1373, new_n2470);
nand_5 g02085(new_n2470, new_n1277, new_n2471);
nand_5 g02086(new_n2471, new_n1272, new_n2472);
nand_5 g02087(new_n2472, new_n1269, new_n2473);
nand_5 g02088(new_n2473, new_n1380, new_n2474);
nand_5 g02089(new_n2474, new_n1264, new_n2475);
nand_5 g02090(new_n2475, new_n1259, new_n2476);
nand_5 g02091(new_n2476, new_n1388, new_n2477);
nand_5 g02092(new_n2477, new_n1392, new_n2478);
nand_5 g02093(new_n2478, new_n1256, new_n2479);
nand_5 g02094(new_n2479, new_n1252, new_n2480);
nand_5 g02095(new_n2480, new_n1249, new_n2481);
nand_5 g02096(new_n2481, new_n1244, new_n2482);
nand_5 g02097(new_n2482, new_n1240, new_n2483);
nand_5 g02098(new_n2483, new_n1234, new_n2484);
nand_5 g02099(new_n2484, new_n1231, new_n2485);
nand_5 g02100(new_n2485, new_n1227, new_n2486);
nand_5 g02101(new_n2486, new_n1407, new_n2487);
nand_5 g02102(new_n2487, new_n1223, new_n2488);
nand_5 g02103(new_n2488, new_n1218, new_n2489);
nand_5 g02104(new_n2489, new_n1213, new_n2490);
nand_5 g02105(new_n2490, new_n1210, new_n2491);
nand_5 g02106(new_n2491, new_n1206, new_n2492);
nand_5 g02107(new_n2492, new_n1418, new_n2493);
nand_5 g02108(new_n2493, new_n1422, new_n2494);
nand_5 g02109(new_n2494, new_n1428, new_n2495);
nand_5 g02110(new_n2495, n2674, new_n2496);
nor_5  g02111(new_n2496, new_n891, n948);
nand_5 g02112(new_n1314, new_n925, new_n2498);
nand_5 g02113(new_n2498, new_n922, new_n2499);
nand_5 g02114(new_n2499, new_n917, new_n2500);
nand_5 g02115(new_n2500, new_n912, new_n2501);
nand_5 g02116(new_n2501, new_n907, new_n2502);
nand_5 g02117(new_n2502, new_n903, new_n2503);
nand_5 g02118(new_n2503, new_n2066, new_n2504);
nand_5 g02119(new_n2504, new_n2063, new_n2505);
nand_5 g02120(new_n2505, new_n2062, new_n2506);
nand_5 g02121(new_n2506, new_n2058, new_n2507);
nand_5 g02122(new_n2507, new_n2055, new_n2508);
nand_5 g02123(new_n2508, new_n2051, new_n2509);
nand_5 g02124(new_n2509, new_n2046, new_n2510);
nand_5 g02125(new_n2510, new_n2042, new_n2511);
nand_5 g02126(new_n2511, new_n2039, new_n2512);
nand_5 g02127(new_n2512, new_n2036, new_n2513);
nand_5 g02128(new_n2513, new_n2033, new_n2514);
nand_5 g02129(new_n2514, new_n2029, new_n2515);
nand_5 g02130(new_n2515, new_n2026, new_n2516);
nand_5 g02131(new_n2516, new_n2022, new_n2517);
nand_5 g02132(new_n2517, new_n2018, new_n2518);
nand_5 g02133(new_n2518, new_n1726, new_n2519);
nand_5 g02134(new_n2519, new_n1722, new_n2520);
nand_5 g02135(new_n2520, new_n1718, new_n2521);
nand_5 g02136(new_n2521, new_n1713, new_n2522);
nand_5 g02137(new_n2522, new_n1737, new_n2523);
nand_5 g02138(new_n2523, new_n1709, new_n2524);
nand_5 g02139(new_n2524, new_n1742, new_n2525);
nand_5 g02140(new_n2525, new_n1704, new_n2526);
nand_5 g02141(new_n2526, new_n1702_1, new_n2527);
nand_5 g02142(new_n2527, new_n1698, new_n2528);
nand_5 g02143(new_n2528, new_n1695, new_n2529);
nand_5 g02144(new_n2529, new_n1692, new_n2530);
nand_5 g02145(new_n2530, new_n1752, new_n2531);
nand_5 g02146(new_n2531, new_n1688, new_n2532);
nand_5 g02147(new_n2532, new_n1685, new_n2533);
nand_5 g02148(new_n2533, new_n1680, new_n2534);
nand_5 g02149(new_n2534, new_n1676, new_n2535);
nand_5 g02150(new_n2535, new_n1672, new_n2536);
nand_5 g02151(new_n2536, new_n1669, new_n2537);
nand_5 g02152(new_n2537, new_n1666, new_n2538);
nand_5 g02153(new_n2538, new_n1663, new_n2539);
nand_5 g02154(new_n2539, new_n1658, new_n2540);
nand_5 g02155(new_n2540, new_n1653, new_n2541);
nand_5 g02156(new_n2541, new_n1651, new_n2542);
nand_5 g02157(new_n2542, new_n1649, new_n2543);
nand_5 g02158(new_n2543, new_n1646, new_n2544);
nand_5 g02159(new_n2544, new_n1643, new_n2545);
nand_5 g02160(new_n2545, new_n1641, new_n2546);
nand_5 g02161(new_n2546, new_n1638, new_n2547);
nand_5 g02162(new_n2547, new_n1635, new_n2548);
nand_5 g02163(new_n2548, new_n1632, new_n2549);
nand_5 g02164(new_n2549, new_n1628, new_n2550);
nand_5 g02165(new_n2550, new_n1625, new_n2551);
nand_5 g02166(new_n2551, new_n1621, new_n2552);
nand_5 g02167(new_n2552, new_n1618, new_n2553);
nand_5 g02168(new_n2553, new_n1778, new_n2554);
nand_5 g02169(new_n2554, new_n1782, new_n2555);
nand_5 g02170(new_n2555, new_n1614, new_n2556_1);
nand_5 g02171(new_n2556_1, new_n1611, new_n2557);
nand_5 g02172(new_n2557, new_n1789, new_n2558);
nand_5 g02173(new_n2558, new_n1608, new_n2559_1);
nand_5 g02174(new_n2559_1, new_n1605, new_n2560);
nand_5 g02175(new_n2560, new_n1795, new_n2561);
nand_5 g02176(new_n2561, new_n1799, new_n2562);
nand_5 g02177(new_n2562, new_n1602, new_n2563);
nand_5 g02178(new_n2563, new_n1599, new_n2564);
nand_5 g02179(new_n2564, new_n1596, new_n2565);
nand_5 g02180(new_n2565, new_n1593, new_n2566);
nand_5 g02181(new_n2566, new_n1806, new_n2567);
nand_5 g02182(new_n2567, new_n1589, new_n2568);
nand_5 g02183(new_n2568, new_n1586, new_n2569);
nand_5 g02184(new_n2569, new_n1583, new_n2570);
nand_5 g02185(new_n2570, new_n1580, new_n2571);
nand_5 g02186(new_n2571, new_n1576, new_n2572_1);
nand_5 g02187(new_n2572_1, new_n1573, new_n2573_1);
nand_5 g02188(new_n2573_1, new_n1570, new_n2574);
nand_5 g02189(new_n2574, new_n1567, new_n2575);
nand_5 g02190(new_n2575, new_n1564, new_n2576);
nand_5 g02191(new_n2576, new_n1561, new_n2577);
nand_5 g02192(new_n2577, new_n1338, new_n2578);
nand_5 g02193(new_n2578, new_n1331, new_n2579);
nand_5 g02194(new_n2579, new_n1326, new_n2580);
nand_5 g02195(new_n2580, new_n1321, new_n2581);
nand_5 g02196(new_n2581, n6555, new_n2582);
nor_5  g02197(new_n2582, new_n729, n1094);
nand_5 g02198(new_n1661, new_n1431, new_n2584);
nand_5 g02199(new_n2584, new_n1085, new_n2585);
nand_5 g02200(new_n2585, new_n1129, new_n2586);
nand_5 g02201(new_n2586, new_n1084, new_n2587);
nand_5 g02202(new_n2587, new_n1134, new_n2588);
nand_5 g02203(new_n2588, new_n1080, new_n2589);
nand_5 g02204(new_n2589, new_n1075, new_n2590);
nand_5 g02205(new_n2590, new_n1070, new_n2591);
nand_5 g02206(new_n2591, new_n1143, new_n2592);
nand_5 g02207(new_n2592, new_n1148, new_n2593);
nand_5 g02208(new_n2593, new_n1065, new_n2594);
nand_5 g02209(new_n2594, new_n1062, new_n2595);
nand_5 g02210(new_n2595, new_n1156, new_n2596);
nand_5 g02211(new_n2596, new_n1057, new_n2597);
nand_5 g02212(new_n2597, new_n1053, new_n2598);
nand_5 g02213(new_n2598, new_n1050, new_n2599);
nand_5 g02214(new_n2599, new_n1045, new_n2600);
nand_5 g02215(new_n2600, new_n1040, new_n2601);
nand_5 g02216(new_n2601, new_n1036, new_n2602);
nand_5 g02217(new_n2602, new_n1033, new_n2603);
nand_5 g02218(new_n2603, new_n1028, new_n2604);
nand_5 g02219(new_n2604, new_n1026, new_n2605);
nand_5 g02220(new_n2605, new_n1021, new_n2606);
nand_5 g02221(new_n2606, new_n1017, new_n2607);
nand_5 g02222(new_n2607, new_n1012, new_n2608);
nand_5 g02223(new_n2608, new_n1009, new_n2609);
nand_5 g02224(new_n2609, new_n1004, new_n2610);
nand_5 g02225(new_n2610, new_n1000, new_n2611);
nand_5 g02226(new_n2611, new_n995, new_n2612);
nand_5 g02227(new_n2612, new_n990, new_n2613);
nand_5 g02228(new_n2613, new_n985, new_n2614);
nand_5 g02229(new_n2614, new_n981, new_n2615_1);
nand_5 g02230(new_n2615_1, new_n1179, new_n2616);
nand_5 g02231(new_n2616, new_n976, new_n2617);
nand_5 g02232(new_n2617, new_n971, new_n2618);
nand_5 g02233(new_n2618, new_n966, new_n2619);
nand_5 g02234(new_n2619, new_n961, new_n2620);
nand_5 g02235(new_n2620, new_n957, new_n2621);
nand_5 g02236(new_n2621, new_n952, new_n2622);
nand_5 g02237(new_n2622, new_n948_1, new_n2623);
nand_5 g02238(new_n2623, new_n943, new_n2624);
nand_5 g02239(new_n2624, new_n941, new_n2625);
nand_5 g02240(new_n2625, new_n938, new_n2626);
nand_5 g02241(new_n2626, new_n936, new_n2627);
nand_5 g02242(new_n2627, new_n931, new_n2628);
nand_5 g02243(new_n2628, new_n927, new_n2629);
nand_5 g02244(new_n2629, new_n922, new_n2630);
nand_5 g02245(new_n2630, new_n917, new_n2631);
nand_5 g02246(new_n2631, new_n912, new_n2632);
nand_5 g02247(new_n2632, new_n907, new_n2633);
nand_5 g02248(new_n2633, new_n903, new_n2634);
nand_5 g02249(new_n2634, new_n2066, new_n2635);
nand_5 g02250(new_n2635, new_n2063, new_n2636);
nand_5 g02251(new_n2636, new_n2062, new_n2637);
nand_5 g02252(new_n2637, new_n2058, new_n2638);
nand_5 g02253(new_n2638, new_n2055, new_n2639);
nand_5 g02254(new_n2639, new_n2051, new_n2640);
nand_5 g02255(new_n2640, new_n2046, new_n2641);
nand_5 g02256(new_n2641, new_n2042, new_n2642);
nand_5 g02257(new_n2642, new_n2039, new_n2643);
nand_5 g02258(new_n2643, new_n2036, new_n2644);
nand_5 g02259(new_n2644, new_n2033, new_n2645);
nand_5 g02260(new_n2645, new_n2029, new_n2646);
nand_5 g02261(new_n2646, new_n2026, new_n2647);
nand_5 g02262(new_n2647, new_n2022, new_n2648);
nand_5 g02263(new_n2648, new_n2018, new_n2649);
nand_5 g02264(new_n2649, new_n1726, new_n2650);
nand_5 g02265(new_n2650, new_n1722, new_n2651);
nand_5 g02266(new_n2651, new_n1718, new_n2652);
nand_5 g02267(new_n2652, new_n1713, new_n2653);
nand_5 g02268(new_n2653, new_n1737, new_n2654);
nand_5 g02269(new_n2654, new_n1709, new_n2655);
nand_5 g02270(new_n2655, new_n1742, new_n2656);
nand_5 g02271(new_n2656, new_n1704, new_n2657);
nand_5 g02272(new_n2657, new_n1702_1, new_n2658);
nand_5 g02273(new_n2658, new_n1698, new_n2659);
nand_5 g02274(new_n2659, new_n1695, new_n2660);
nand_5 g02275(new_n2660, new_n1692, new_n2661);
nand_5 g02276(new_n2661, new_n1752, new_n2662);
nand_5 g02277(new_n2662, new_n1688, new_n2663);
nand_5 g02278(new_n2663, new_n1685, new_n2664);
nand_5 g02279(new_n2664, new_n1680, new_n2665);
nand_5 g02280(new_n2665, new_n1676, new_n2666);
nand_5 g02281(new_n2666, new_n1672, new_n2667);
nand_5 g02282(new_n2667, new_n1669, new_n2668);
nand_5 g02283(new_n2668, n12270, new_n2669);
nor_5  g02284(new_n2669, new_n1425, n1122);
not_4  g02285(n9543, new_n2671);
nand_5 g02286(new_n1043, new_n2671, new_n2672_1);
nand_5 g02287(new_n2672_1, new_n541, new_n2673);
nand_5 g02288(new_n2673, new_n636, new_n2674_1);
nand_5 g02289(new_n2674_1, new_n642, new_n2675);
nand_5 g02290(new_n2675, new_n538, new_n2676);
nand_5 g02291(new_n2676, new_n533, new_n2677);
nand_5 g02292(new_n2677, new_n650_1, new_n2678);
nand_5 g02293(new_n2678, new_n528, new_n2679);
nand_5 g02294(new_n2679, new_n523, new_n2680);
nand_5 g02295(new_n2680, new_n518, new_n2681);
nand_5 g02296(new_n2681, new_n659, new_n2682);
nand_5 g02297(new_n2682, new_n665, new_n2683);
nand_5 g02298(new_n2683, new_n672, new_n2684);
nand_5 g02299(new_n2684, new_n513, new_n2685);
nand_5 g02300(new_n2685, new_n679, new_n2686);
nand_5 g02301(new_n2686, new_n685, new_n2687);
nand_5 g02302(new_n2687, new_n691, new_n2688);
nand_5 g02303(new_n2688, new_n508, new_n2689);
nand_5 g02304(new_n2689, new_n698, new_n2690);
nand_5 g02305(new_n2690, new_n503, new_n2691);
nand_5 g02306(new_n2691, new_n704, new_n2692);
nand_5 g02307(new_n2692, new_n498_1, new_n2693);
nand_5 g02308(new_n2693, new_n711, new_n2694);
nand_5 g02309(new_n2694, new_n493, new_n2695);
nand_5 g02310(new_n2695, new_n718, new_n2696);
nand_5 g02311(new_n2696, new_n488, new_n2697);
nand_5 g02312(new_n2697, new_n725, new_n2698);
nand_5 g02313(new_n2698, new_n483, new_n2699_1);
nand_5 g02314(new_n2699_1, new_n732, new_n2700);
nand_5 g02315(new_n2700, new_n478, new_n2701);
nand_5 g02316(new_n2701, new_n739, new_n2702);
nand_5 g02317(new_n2702, new_n745, new_n2703);
nand_5 g02318(new_n2703, new_n751, new_n2704);
nand_5 g02319(new_n2704, new_n473, new_n2705);
nand_5 g02320(new_n2705, new_n758, new_n2706);
nand_5 g02321(new_n2706, new_n764, new_n2707);
nand_5 g02322(new_n2707, new_n770, new_n2708);
nand_5 g02323(new_n2708, new_n468, new_n2709);
nand_5 g02324(new_n2709, new_n777, new_n2710);
nand_5 g02325(new_n2710, new_n783, new_n2711);
nand_5 g02326(new_n2711, new_n789, new_n2712);
nand_5 g02327(new_n2712, new_n463, new_n2713);
nand_5 g02328(new_n2713, new_n796, new_n2714);
nand_5 g02329(new_n2714, new_n458, new_n2715);
nand_5 g02330(new_n2715, new_n453, new_n2716);
nand_5 g02331(new_n2716, new_n447, new_n2717);
nand_5 g02332(new_n2717, new_n805, new_n2718);
nand_5 g02333(new_n2718, new_n811, new_n2719);
nand_5 g02334(new_n2719, new_n442, new_n2720);
nand_5 g02335(new_n2720, new_n437, new_n2721);
nand_5 g02336(new_n2721, new_n819, new_n2722);
nand_5 g02337(new_n2722, new_n432, new_n2723);
nand_5 g02338(new_n2723, new_n427_1, new_n2724);
nand_5 g02339(new_n2724, new_n422, new_n2725);
nand_5 g02340(new_n2725, new_n828, new_n2726);
nand_5 g02341(new_n2726, new_n834, new_n2727);
nand_5 g02342(new_n2727, new_n840, new_n2728);
nand_5 g02343(new_n2728, new_n417, new_n2729);
nand_5 g02344(new_n2729, new_n847, new_n2730);
nand_5 g02345(new_n2730, new_n853, new_n2731);
nand_5 g02346(new_n2731, new_n859, new_n2732);
nand_5 g02347(new_n2732, new_n412, new_n2733);
nand_5 g02348(new_n2733, new_n866, new_n2734_1);
nand_5 g02349(new_n2734_1, new_n872, new_n2735);
nand_5 g02350(new_n2735, new_n878, new_n2736);
nand_5 g02351(new_n2736, new_n407, new_n2737);
nand_5 g02352(new_n2737, new_n885, new_n2738);
nand_5 g02353(new_n2738, new_n402, new_n2739);
nand_5 g02354(new_n2739, new_n397, new_n2740);
nand_5 g02355(new_n2740, new_n392, new_n2741);
nand_5 g02356(new_n2741, new_n894, new_n2742);
nand_5 g02357(new_n2742, new_n1087, new_n2743);
nand_5 g02358(new_n2743, new_n1129, new_n2744);
nand_5 g02359(new_n2744, new_n1084, new_n2745);
nand_5 g02360(new_n2745, new_n1134, new_n2746);
nand_5 g02361(new_n2746, new_n1080, new_n2747);
nand_5 g02362(new_n2747, new_n1075, new_n2748);
nand_5 g02363(new_n2748, new_n1070, new_n2749);
nand_5 g02364(new_n2749, new_n1143, new_n2750);
nand_5 g02365(new_n2750, new_n1148, new_n2751);
nand_5 g02366(new_n2751, new_n1065, new_n2752);
nand_5 g02367(new_n2752, new_n1062, new_n2753);
nand_5 g02368(new_n2753, new_n1156, new_n2754);
nand_5 g02369(new_n2754, new_n1057, new_n2755);
nand_5 g02370(new_n2755, new_n1053, new_n2756);
nand_5 g02371(new_n2756, n271, new_n2757);
nor_5  g02372(new_n2757, new_n1047, n1124);
not_4  g02373(new_n1667, new_n2759);
nand_5 g02374(new_n2759, new_n392, new_n2760);
nand_5 g02375(new_n2760, new_n894, new_n2761);
nand_5 g02376(new_n2761, new_n1087, new_n2762);
nand_5 g02377(new_n2762, new_n1129, new_n2763);
nand_5 g02378(new_n2763, new_n1084, new_n2764);
nand_5 g02379(new_n2764, new_n1134, new_n2765);
nand_5 g02380(new_n2765, new_n1080, new_n2766);
nand_5 g02381(new_n2766, new_n1075, new_n2767);
nand_5 g02382(new_n2767, new_n1070, new_n2768);
nand_5 g02383(new_n2768, new_n1143, new_n2769);
nand_5 g02384(new_n2769, new_n1148, new_n2770);
nand_5 g02385(new_n2770, new_n1065, new_n2771);
nand_5 g02386(new_n2771, new_n1062, new_n2772);
nand_5 g02387(new_n2772, new_n1156, new_n2773);
nand_5 g02388(new_n2773, new_n1057, new_n2774);
nand_5 g02389(new_n2774, new_n1053, new_n2775);
nand_5 g02390(new_n2775, new_n1050, new_n2776);
nand_5 g02391(new_n2776, new_n1045, new_n2777);
nand_5 g02392(new_n2777, new_n1040, new_n2778);
nand_5 g02393(new_n2778, new_n1036, new_n2779);
nand_5 g02394(new_n2779, new_n1033, new_n2780);
nand_5 g02395(new_n2780, new_n1028, new_n2781);
nand_5 g02396(new_n2781, new_n1026, new_n2782);
nand_5 g02397(new_n2782, new_n1021, new_n2783);
nand_5 g02398(new_n2783, new_n1017, new_n2784);
nand_5 g02399(new_n2784, new_n1012, new_n2785);
nand_5 g02400(new_n2785, new_n1009, new_n2786);
nand_5 g02401(new_n2786, new_n1004, new_n2787);
nand_5 g02402(new_n2787, new_n1000, new_n2788);
nand_5 g02403(new_n2788, new_n995, new_n2789);
nand_5 g02404(new_n2789, new_n990, new_n2790);
nand_5 g02405(new_n2790, new_n985, new_n2791);
nand_5 g02406(new_n2791, new_n981, new_n2792);
nand_5 g02407(new_n2792, new_n1179, new_n2793);
nand_5 g02408(new_n2793, new_n976, new_n2794);
nand_5 g02409(new_n2794, new_n971, new_n2795);
nand_5 g02410(new_n2795, new_n966, new_n2796);
nand_5 g02411(new_n2796, new_n961, new_n2797);
nand_5 g02412(new_n2797, new_n957, new_n2798);
nand_5 g02413(new_n2798, new_n952, new_n2799);
nand_5 g02414(new_n2799, new_n948_1, new_n2800);
nand_5 g02415(new_n2800, new_n943, new_n2801);
nand_5 g02416(new_n2801, new_n941, new_n2802);
nand_5 g02417(new_n2802, new_n938, new_n2803);
nand_5 g02418(new_n2803, new_n936, new_n2804);
nand_5 g02419(new_n2804, new_n931, new_n2805);
nand_5 g02420(new_n2805, new_n927, new_n2806);
nand_5 g02421(new_n2806, new_n922, new_n2807);
nand_5 g02422(new_n2807, new_n917, new_n2808);
nand_5 g02423(new_n2808, new_n912, new_n2809);
nand_5 g02424(new_n2809, new_n907, new_n2810);
nand_5 g02425(new_n2810, new_n903, new_n2811);
nand_5 g02426(new_n2811, new_n2066, new_n2812);
nand_5 g02427(new_n2812, new_n2063, new_n2813);
nand_5 g02428(new_n2813, new_n2062, new_n2814);
nand_5 g02429(new_n2814, new_n2058, new_n2815);
nand_5 g02430(new_n2815, new_n2055, new_n2816);
nand_5 g02431(new_n2816, new_n2051, new_n2817);
nand_5 g02432(new_n2817, new_n2046, new_n2818);
nand_5 g02433(new_n2818, new_n2042, new_n2819);
nand_5 g02434(new_n2819, new_n2039, new_n2820);
nand_5 g02435(new_n2820, new_n2036, new_n2821);
nand_5 g02436(new_n2821, new_n2033, new_n2822);
nand_5 g02437(new_n2822, new_n2029, new_n2823);
nand_5 g02438(new_n2823, new_n2026, new_n2824);
nand_5 g02439(new_n2824, new_n2022, new_n2825);
nand_5 g02440(new_n2825, new_n2018, new_n2826);
nand_5 g02441(new_n2826, new_n1726, new_n2827);
nand_5 g02442(new_n2827, new_n1722, new_n2828);
nand_5 g02443(new_n2828, new_n1718, new_n2829);
nand_5 g02444(new_n2829, new_n1713, new_n2830);
nand_5 g02445(new_n2830, new_n1737, new_n2831);
nand_5 g02446(new_n2831, new_n1709, new_n2832);
nand_5 g02447(new_n2832, new_n1742, new_n2833);
nand_5 g02448(new_n2833, new_n1704, new_n2834);
nand_5 g02449(new_n2834, new_n1702_1, new_n2835);
nand_5 g02450(new_n2835, new_n1698, new_n2836);
nand_5 g02451(new_n2836, new_n1695, new_n2837);
nand_5 g02452(new_n2837, new_n1692, new_n2838);
nand_5 g02453(new_n2838, new_n1752, new_n2839);
nand_5 g02454(new_n2839, new_n1688, new_n2840);
nand_5 g02455(new_n2840, new_n1685, new_n2841);
nand_5 g02456(new_n2841, new_n1680, new_n2842);
nand_5 g02457(new_n2842, new_n1676, new_n2843);
nand_5 g02458(new_n2843, n1268, new_n2844);
nor_5  g02459(new_n2844, new_n1415, n1329);
nand_5 g02460(new_n1562, new_n710, new_n2846);
nand_5 g02461(new_n2846, new_n1561, new_n2847);
nand_5 g02462(new_n2847, new_n1338, new_n2848);
nand_5 g02463(new_n2848, new_n1331, new_n2849);
nand_5 g02464(new_n2849, new_n1326, new_n2850);
nand_5 g02465(new_n2850, new_n1321, new_n2851);
nand_5 g02466(new_n2851, new_n1318, new_n2852);
nand_5 g02467(new_n2852, new_n1315, new_n2853);
nand_5 g02468(new_n2853, new_n1312, new_n2854);
nand_5 g02469(new_n2854, new_n1309, new_n2855);
nand_5 g02470(new_n2855, new_n1307, new_n2856);
nand_5 g02471(new_n2856, new_n1304, new_n2857);
nand_5 g02472(new_n2857, new_n1300, new_n2858);
nand_5 g02473(new_n2858, new_n1297, new_n2859);
nand_5 g02474(new_n2859, new_n1294, new_n2860);
nand_5 g02475(new_n2860, new_n1355, new_n2861);
nand_5 g02476(new_n2861, new_n1291, new_n2862);
nand_5 g02477(new_n2862, new_n1288, new_n2863);
nand_5 g02478(new_n2863, new_n1283, new_n2864);
nand_5 g02479(new_n2864, new_n1363, new_n2865);
nand_5 g02480(new_n2865, new_n1280, new_n2866);
nand_5 g02481(new_n2866, new_n1370, new_n2867);
nand_5 g02482(new_n2867, new_n1373, new_n2868);
nand_5 g02483(new_n2868, new_n1277, new_n2869);
nand_5 g02484(new_n2869, new_n1272, new_n2870);
nand_5 g02485(new_n2870, new_n1269, new_n2871);
nand_5 g02486(new_n2871, new_n1380, new_n2872);
nand_5 g02487(new_n2872, new_n1264, new_n2873);
nand_5 g02488(new_n2873, new_n1259, new_n2874);
nand_5 g02489(new_n2874, new_n1388, new_n2875);
nand_5 g02490(new_n2875, new_n1392, new_n2876);
nand_5 g02491(new_n2876, new_n1256, new_n2877);
nand_5 g02492(new_n2877, new_n1252, new_n2878);
nand_5 g02493(new_n2878, new_n1249, new_n2879);
nand_5 g02494(new_n2879, new_n1244, new_n2880);
nand_5 g02495(new_n2880, new_n1240, new_n2881);
nand_5 g02496(new_n2881, new_n1234, new_n2882);
nand_5 g02497(new_n2882, new_n1231, new_n2883);
nand_5 g02498(new_n2883, new_n1227, new_n2884);
nand_5 g02499(new_n2884, new_n1407, new_n2885);
nand_5 g02500(new_n2885, new_n1223, new_n2886);
nand_5 g02501(new_n2886, new_n1218, new_n2887);
nand_5 g02502(new_n2887, new_n1213, new_n2888);
nand_5 g02503(new_n2888, new_n1210, new_n2889);
nand_5 g02504(new_n2889, new_n1206, new_n2890);
nand_5 g02505(new_n2890, new_n1418, new_n2891);
nand_5 g02506(new_n2891, new_n1422, new_n2892);
nand_5 g02507(new_n2892, new_n1428, new_n2893);
nand_5 g02508(new_n2893, new_n1203, new_n2894);
nand_5 g02509(new_n2894, new_n1433, new_n2895_1);
nand_5 g02510(new_n2895_1, new_n581, new_n2896);
nand_5 g02511(new_n2896, new_n574, new_n2897);
nand_5 g02512(new_n2897, new_n568, new_n2898);
nand_5 g02513(new_n2898, new_n589, new_n2899);
nand_5 g02514(new_n2899, new_n595, new_n2900);
nand_5 g02515(new_n2900, new_n601, new_n2901);
nand_5 g02516(new_n2901, new_n563, new_n2902);
nand_5 g02517(new_n2902, new_n608, new_n2903);
nand_5 g02518(new_n2903, new_n558, new_n2904);
nand_5 g02519(new_n2904, new_n615, new_n2905);
nand_5 g02520(new_n2905, new_n553, new_n2906);
nand_5 g02521(new_n2906, new_n622, new_n2907);
nand_5 g02522(new_n2907, new_n628, new_n2908);
nand_5 g02523(new_n2908, new_n548, new_n2909);
nand_5 g02524(new_n2909, new_n543_1, new_n2910);
nand_5 g02525(new_n2910, new_n636, new_n2911);
nand_5 g02526(new_n2911, new_n642, new_n2912);
nand_5 g02527(new_n2912, new_n538, new_n2913);
nand_5 g02528(new_n2913, new_n533, new_n2914);
nand_5 g02529(new_n2914, new_n650_1, new_n2915);
nand_5 g02530(new_n2915, new_n528, new_n2916);
nand_5 g02531(new_n2916, new_n523, new_n2917);
nand_5 g02532(new_n2917, new_n518, new_n2918);
nand_5 g02533(new_n2918, new_n659, new_n2919);
nand_5 g02534(new_n2919, new_n665, new_n2920);
nand_5 g02535(new_n2920, new_n672, new_n2921);
nand_5 g02536(new_n2921, new_n513, new_n2922);
nand_5 g02537(new_n2922, new_n679, new_n2923);
nand_5 g02538(new_n2923, new_n685, new_n2924);
nand_5 g02539(new_n2924, new_n691, new_n2925);
nand_5 g02540(new_n2925, new_n508, new_n2926);
nand_5 g02541(new_n2926, new_n698, new_n2927);
nand_5 g02542(new_n2927, new_n503, new_n2928);
nand_5 g02543(new_n2928, new_n704, new_n2929);
nand_5 g02544(new_n2929, n4117, new_n2930);
nor_5  g02545(new_n2930, new_n495, n1545);
not_4  g02546(new_n1700, new_n2932);
nand_5 g02547(new_n2932, new_n853, new_n2933);
nand_5 g02548(new_n2933, new_n859, new_n2934);
nand_5 g02549(new_n2934, new_n412, new_n2935);
nand_5 g02550(new_n2935, new_n866, new_n2936);
nand_5 g02551(new_n2936, new_n872, new_n2937);
nand_5 g02552(new_n2937, new_n878, new_n2938);
nand_5 g02553(new_n2938, new_n407, new_n2939);
nand_5 g02554(new_n2939, new_n885, new_n2940);
nand_5 g02555(new_n2940, new_n402, new_n2941);
nand_5 g02556(new_n2941, new_n397, new_n2942);
nand_5 g02557(new_n2942, new_n392, new_n2943);
nand_5 g02558(new_n2943, new_n894, new_n2944);
nand_5 g02559(new_n2944, new_n1087, new_n2945);
nand_5 g02560(new_n2945, new_n1129, new_n2946);
nand_5 g02561(new_n2946, new_n1084, new_n2947);
nand_5 g02562(new_n2947, new_n1134, new_n2948);
nand_5 g02563(new_n2948, new_n1080, new_n2949);
nand_5 g02564(new_n2949, new_n1075, new_n2950);
nand_5 g02565(new_n2950, new_n1070, new_n2951);
nand_5 g02566(new_n2951, new_n1143, new_n2952);
nand_5 g02567(new_n2952, new_n1148, new_n2953);
nand_5 g02568(new_n2953, new_n1065, new_n2954);
nand_5 g02569(new_n2954, new_n1062, new_n2955);
nand_5 g02570(new_n2955, new_n1156, new_n2956);
nand_5 g02571(new_n2956, new_n1057, new_n2957);
nand_5 g02572(new_n2957, new_n1053, new_n2958);
nand_5 g02573(new_n2958, new_n1050, new_n2959);
nand_5 g02574(new_n2959, new_n1045, new_n2960);
nand_5 g02575(new_n2960, new_n1040, new_n2961);
nand_5 g02576(new_n2961, new_n1036, new_n2962);
nand_5 g02577(new_n2962, new_n1033, new_n2963);
nand_5 g02578(new_n2963, new_n1028, new_n2964);
nand_5 g02579(new_n2964, new_n1026, new_n2965);
nand_5 g02580(new_n2965, new_n1021, new_n2966);
nand_5 g02581(new_n2966, new_n1017, new_n2967);
nand_5 g02582(new_n2967, new_n1012, new_n2968);
nand_5 g02583(new_n2968, new_n1009, new_n2969);
nand_5 g02584(new_n2969, new_n1004, new_n2970);
nand_5 g02585(new_n2970, new_n1000, new_n2971);
nand_5 g02586(new_n2971, new_n995, new_n2972);
nand_5 g02587(new_n2972, new_n990, new_n2973);
nand_5 g02588(new_n2973, new_n985, new_n2974);
nand_5 g02589(new_n2974, new_n981, new_n2975);
nand_5 g02590(new_n2975, new_n1179, new_n2976);
nand_5 g02591(new_n2976, new_n976, new_n2977);
nand_5 g02592(new_n2977, new_n971, new_n2978);
nand_5 g02593(new_n2978, new_n966, new_n2979);
nand_5 g02594(new_n2979, new_n961, new_n2980);
nand_5 g02595(new_n2980, new_n957, new_n2981);
nand_5 g02596(new_n2981, new_n952, new_n2982);
nand_5 g02597(new_n2982, new_n948_1, new_n2983);
nand_5 g02598(new_n2983, new_n943, new_n2984);
nand_5 g02599(new_n2984, new_n941, new_n2985);
nand_5 g02600(new_n2985, new_n938, new_n2986);
nand_5 g02601(new_n2986, new_n936, new_n2987);
nand_5 g02602(new_n2987, new_n931, new_n2988);
nand_5 g02603(new_n2988, new_n927, new_n2989);
nand_5 g02604(new_n2989, new_n922, new_n2990);
nand_5 g02605(new_n2990, new_n917, new_n2991);
nand_5 g02606(new_n2991, new_n912, new_n2992);
nand_5 g02607(new_n2992, new_n907, new_n2993);
nand_5 g02608(new_n2993, new_n903, new_n2994);
nand_5 g02609(new_n2994, new_n2066, new_n2995);
nand_5 g02610(new_n2995, new_n2063, new_n2996);
nand_5 g02611(new_n2996, new_n2062, new_n2997);
nand_5 g02612(new_n2997, new_n2058, new_n2998);
nand_5 g02613(new_n2998, new_n2055, new_n2999);
nand_5 g02614(new_n2999, new_n2051, new_n3000);
nand_5 g02615(new_n3000, new_n2046, new_n3001);
nand_5 g02616(new_n3001, new_n2042, new_n3002);
nand_5 g02617(new_n3002, new_n2039, new_n3003);
nand_5 g02618(new_n3003, new_n2036, new_n3004);
nand_5 g02619(new_n3004, new_n2033, new_n3005);
nand_5 g02620(new_n3005, new_n2029, new_n3006);
nand_5 g02621(new_n3006, new_n2026, new_n3007);
nand_5 g02622(new_n3007, new_n2022, new_n3008);
nand_5 g02623(new_n3008, new_n2018, new_n3009);
nand_5 g02624(new_n3009, new_n1726, new_n3010);
nand_5 g02625(new_n3010, new_n1722, new_n3011);
nand_5 g02626(new_n3011, new_n1718, new_n3012);
nand_5 g02627(new_n3012, new_n1713, new_n3013);
nand_5 g02628(new_n3013, new_n1737, new_n3014);
nand_5 g02629(new_n3014, new_n1709, new_n3015);
nand_5 g02630(new_n3015, new_n1742, new_n3016);
nand_5 g02631(new_n3016, n12336, new_n3017);
nor_5  g02632(new_n3017, new_n1237, n1739);
nand_5 g02633(new_n1420, new_n396, new_n3019);
nand_5 g02634(new_n3019, new_n1428, new_n3020);
nand_5 g02635(new_n3020, new_n1203, new_n3021);
nand_5 g02636(new_n3021, new_n1433, new_n3022);
nand_5 g02637(new_n3022, new_n581, new_n3023);
nand_5 g02638(new_n3023, new_n574, new_n3024);
nand_5 g02639(new_n3024, new_n568, new_n3025);
nand_5 g02640(new_n3025, new_n589, new_n3026);
nand_5 g02641(new_n3026, new_n595, new_n3027);
nand_5 g02642(new_n3027, new_n601, new_n3028);
nand_5 g02643(new_n3028, new_n563, new_n3029);
nand_5 g02644(new_n3029, new_n608, new_n3030);
nand_5 g02645(new_n3030, new_n558, new_n3031);
nand_5 g02646(new_n3031, new_n615, new_n3032);
nand_5 g02647(new_n3032, new_n553, new_n3033);
nand_5 g02648(new_n3033, new_n622, new_n3034);
nand_5 g02649(new_n3034, new_n628, new_n3035);
nand_5 g02650(new_n3035, new_n548, new_n3036);
nand_5 g02651(new_n3036, new_n543_1, new_n3037);
nand_5 g02652(new_n3037, new_n636, new_n3038);
nand_5 g02653(new_n3038, new_n642, new_n3039);
nand_5 g02654(new_n3039, new_n538, new_n3040);
nand_5 g02655(new_n3040, new_n533, new_n3041);
nand_5 g02656(new_n3041, new_n650_1, new_n3042);
nand_5 g02657(new_n3042, new_n528, new_n3043);
nand_5 g02658(new_n3043, new_n523, new_n3044);
nand_5 g02659(new_n3044, new_n518, new_n3045);
nand_5 g02660(new_n3045, new_n659, new_n3046);
nand_5 g02661(new_n3046, new_n665, new_n3047);
nand_5 g02662(new_n3047, new_n672, new_n3048);
nand_5 g02663(new_n3048, new_n513, new_n3049);
nand_5 g02664(new_n3049, new_n679, new_n3050);
nand_5 g02665(new_n3050, new_n685, new_n3051);
nand_5 g02666(new_n3051, new_n691, new_n3052);
nand_5 g02667(new_n3052, new_n508, new_n3053);
nand_5 g02668(new_n3053, new_n698, new_n3054);
nand_5 g02669(new_n3054, new_n503, new_n3055);
nand_5 g02670(new_n3055, new_n704, new_n3056);
nand_5 g02671(new_n3056, new_n498_1, new_n3057);
nand_5 g02672(new_n3057, new_n711, new_n3058);
nand_5 g02673(new_n3058, new_n493, new_n3059);
nand_5 g02674(new_n3059, new_n718, new_n3060);
nand_5 g02675(new_n3060, new_n488, new_n3061);
nand_5 g02676(new_n3061, new_n725, new_n3062);
nand_5 g02677(new_n3062, new_n483, new_n3063);
nand_5 g02678(new_n3063, new_n732, new_n3064);
nand_5 g02679(new_n3064, new_n478, new_n3065);
nand_5 g02680(new_n3065, new_n739, new_n3066);
nand_5 g02681(new_n3066, new_n745, new_n3067);
nand_5 g02682(new_n3067, new_n751, new_n3068);
nand_5 g02683(new_n3068, new_n473, new_n3069);
nand_5 g02684(new_n3069, new_n758, new_n3070);
nand_5 g02685(new_n3070, new_n764, new_n3071);
nand_5 g02686(new_n3071, new_n770, new_n3072);
nand_5 g02687(new_n3072, new_n468, new_n3073);
nand_5 g02688(new_n3073, new_n777, new_n3074);
nand_5 g02689(new_n3074, new_n783, new_n3075);
nand_5 g02690(new_n3075, new_n789, new_n3076);
nand_5 g02691(new_n3076, new_n463, new_n3077);
nand_5 g02692(new_n3077, new_n796, new_n3078);
nand_5 g02693(new_n3078, new_n458, new_n3079);
nand_5 g02694(new_n3079, new_n453, new_n3080);
nand_5 g02695(new_n3080, new_n447, new_n3081);
nand_5 g02696(new_n3081, new_n805, new_n3082);
nand_5 g02697(new_n3082, new_n811, new_n3083);
nand_5 g02698(new_n3083, new_n442, new_n3084);
nand_5 g02699(new_n3084, new_n437, new_n3085);
nand_5 g02700(new_n3085, new_n819, new_n3086);
nand_5 g02701(new_n3086, new_n432, new_n3087);
nand_5 g02702(new_n3087, new_n427_1, new_n3088);
nand_5 g02703(new_n3088, new_n422, new_n3089);
nand_5 g02704(new_n3089, new_n828, new_n3090_1);
nand_5 g02705(new_n3090_1, new_n834, new_n3091);
nand_5 g02706(new_n3091, new_n840, new_n3092);
nand_5 g02707(new_n3092, new_n417, new_n3093);
nand_5 g02708(new_n3093, new_n847, new_n3094);
nand_5 g02709(new_n3094, new_n853, new_n3095);
nand_5 g02710(new_n3095, new_n859, new_n3096);
nand_5 g02711(new_n3096, new_n412, new_n3097);
nand_5 g02712(new_n3097, new_n866, new_n3098);
nand_5 g02713(new_n3098, new_n872, new_n3099);
nand_5 g02714(new_n3099, new_n878, new_n3100);
nand_5 g02715(new_n3100, new_n407, new_n3101);
nand_5 g02716(new_n3101, new_n885, new_n3102);
nand_5 g02717(new_n3102, n394, new_n3103);
nor_5  g02718(new_n3103, new_n399, n1827);
nand_5 g02719(new_n1278, new_n795, new_n3105);
nand_5 g02720(new_n3105, new_n1370, new_n3106);
nand_5 g02721(new_n3106, new_n1373, new_n3107);
nand_5 g02722(new_n3107, new_n1277, new_n3108);
nand_5 g02723(new_n3108, new_n1272, new_n3109);
nand_5 g02724(new_n3109, new_n1269, new_n3110);
nand_5 g02725(new_n3110, new_n1380, new_n3111);
nand_5 g02726(new_n3111, new_n1264, new_n3112);
nand_5 g02727(new_n3112, new_n1259, new_n3113);
nand_5 g02728(new_n3113, new_n1388, new_n3114);
nand_5 g02729(new_n3114, new_n1392, new_n3115);
nand_5 g02730(new_n3115, new_n1256, new_n3116);
nand_5 g02731(new_n3116, new_n1252, new_n3117);
nand_5 g02732(new_n3117, new_n1249, new_n3118);
nand_5 g02733(new_n3118, new_n1244, new_n3119);
nand_5 g02734(new_n3119, new_n1240, new_n3120);
nand_5 g02735(new_n3120, new_n1234, new_n3121);
nand_5 g02736(new_n3121, new_n1231, new_n3122);
nand_5 g02737(new_n3122, new_n1227, new_n3123);
nand_5 g02738(new_n3123, new_n1407, new_n3124);
nand_5 g02739(new_n3124, new_n1223, new_n3125);
nand_5 g02740(new_n3125, new_n1218, new_n3126);
nand_5 g02741(new_n3126, new_n1213, new_n3127);
nand_5 g02742(new_n3127, new_n1210, new_n3128);
nand_5 g02743(new_n3128, new_n1206, new_n3129);
nand_5 g02744(new_n3129, new_n1418, new_n3130_1);
nand_5 g02745(new_n3130_1, new_n1422, new_n3131);
nand_5 g02746(new_n3131, new_n1428, new_n3132);
nand_5 g02747(new_n3132, new_n1203, new_n3133);
nand_5 g02748(new_n3133, new_n1433, new_n3134);
nand_5 g02749(new_n3134, new_n581, new_n3135);
nand_5 g02750(new_n3135, new_n574, new_n3136);
nand_5 g02751(new_n3136, new_n568, new_n3137);
nand_5 g02752(new_n3137, new_n589, new_n3138);
nand_5 g02753(new_n3138, new_n595, new_n3139);
nand_5 g02754(new_n3139, new_n601, new_n3140);
nand_5 g02755(new_n3140, new_n563, new_n3141);
nand_5 g02756(new_n3141, new_n608, new_n3142);
nand_5 g02757(new_n3142, new_n558, new_n3143);
nand_5 g02758(new_n3143, new_n615, new_n3144);
nand_5 g02759(new_n3144, new_n553, new_n3145);
nand_5 g02760(new_n3145, new_n622, new_n3146);
nand_5 g02761(new_n3146, new_n628, new_n3147);
nand_5 g02762(new_n3147, new_n548, new_n3148);
nand_5 g02763(new_n3148, new_n543_1, new_n3149);
nand_5 g02764(new_n3149, new_n636, new_n3150);
nand_5 g02765(new_n3150, new_n642, new_n3151);
nand_5 g02766(new_n3151, new_n538, new_n3152);
nand_5 g02767(new_n3152, new_n533, new_n3153);
nand_5 g02768(new_n3153, new_n650_1, new_n3154);
nand_5 g02769(new_n3154, new_n528, new_n3155);
nand_5 g02770(new_n3155, new_n523, new_n3156);
nand_5 g02771(new_n3156, new_n518, new_n3157);
nand_5 g02772(new_n3157, new_n659, new_n3158);
nand_5 g02773(new_n3158, new_n665, new_n3159);
nand_5 g02774(new_n3159, new_n672, new_n3160);
nand_5 g02775(new_n3160, new_n513, new_n3161);
nand_5 g02776(new_n3161, new_n679, new_n3162);
nand_5 g02777(new_n3162, new_n685, new_n3163);
nand_5 g02778(new_n3163, new_n691, new_n3164);
nand_5 g02779(new_n3164, new_n508, new_n3165);
nand_5 g02780(new_n3165, new_n698, new_n3166_1);
nand_5 g02781(new_n3166_1, new_n503, new_n3167);
nand_5 g02782(new_n3167, new_n704, new_n3168);
nand_5 g02783(new_n3168, new_n498_1, new_n3169);
nand_5 g02784(new_n3169, new_n711, new_n3170);
nand_5 g02785(new_n3170, new_n493, new_n3171);
nand_5 g02786(new_n3171, new_n718, new_n3172);
nand_5 g02787(new_n3172, new_n488, new_n3173);
nand_5 g02788(new_n3173, new_n725, new_n3174);
nand_5 g02789(new_n3174, new_n483, new_n3175);
nand_5 g02790(new_n3175, new_n732, new_n3176);
nand_5 g02791(new_n3176, new_n478, new_n3177);
nand_5 g02792(new_n3177, new_n739, new_n3178);
nand_5 g02793(new_n3178, new_n745, new_n3179);
nand_5 g02794(new_n3179, new_n751, new_n3180);
nand_5 g02795(new_n3180, new_n473, new_n3181);
nand_5 g02796(new_n3181, new_n758, new_n3182);
nand_5 g02797(new_n3182, new_n764, new_n3183);
nand_5 g02798(new_n3183, new_n770, new_n3184);
nand_5 g02799(new_n3184, new_n468, new_n3185);
nand_5 g02800(new_n3185, new_n777, new_n3186);
nand_5 g02801(new_n3186, new_n783, new_n3187);
nand_5 g02802(new_n3187, new_n789, new_n3188);
nand_5 g02803(new_n3188, n730, new_n3189);
nor_5  g02804(new_n3189, new_n460, n1900);
nand_5 g02805(new_n2049, new_n1361, new_n3191);
nand_5 g02806(new_n3191, new_n461, new_n3192);
nand_5 g02807(new_n3192, new_n796, new_n3193);
nand_5 g02808(new_n3193, new_n458, new_n3194);
nand_5 g02809(new_n3194, new_n453, new_n3195);
nand_5 g02810(new_n3195, new_n447, new_n3196);
nand_5 g02811(new_n3196, new_n805, new_n3197);
nand_5 g02812(new_n3197, new_n811, new_n3198);
nand_5 g02813(new_n3198, new_n442, new_n3199);
nand_5 g02814(new_n3199, new_n437, new_n3200);
nand_5 g02815(new_n3200, new_n819, new_n3201);
nand_5 g02816(new_n3201, new_n432, new_n3202);
nand_5 g02817(new_n3202, new_n427_1, new_n3203);
nand_5 g02818(new_n3203, new_n422, new_n3204);
nand_5 g02819(new_n3204, new_n828, new_n3205);
nand_5 g02820(new_n3205, new_n834, new_n3206);
nand_5 g02821(new_n3206, new_n840, new_n3207);
nand_5 g02822(new_n3207, new_n417, new_n3208);
nand_5 g02823(new_n3208, new_n847, new_n3209);
nand_5 g02824(new_n3209, new_n853, new_n3210);
nand_5 g02825(new_n3210, new_n859, new_n3211);
nand_5 g02826(new_n3211, new_n412, new_n3212);
nand_5 g02827(new_n3212, new_n866, new_n3213);
nand_5 g02828(new_n3213, new_n872, new_n3214);
nand_5 g02829(new_n3214, new_n878, new_n3215);
nand_5 g02830(new_n3215, new_n407, new_n3216);
nand_5 g02831(new_n3216, new_n885, new_n3217);
nand_5 g02832(new_n3217, new_n402, new_n3218);
nand_5 g02833(new_n3218, new_n397, new_n3219);
nand_5 g02834(new_n3219, new_n392, new_n3220);
nand_5 g02835(new_n3220, new_n894, new_n3221);
nand_5 g02836(new_n3221, new_n1087, new_n3222);
nand_5 g02837(new_n3222, new_n1129, new_n3223);
nand_5 g02838(new_n3223, new_n1084, new_n3224);
nand_5 g02839(new_n3224, new_n1134, new_n3225);
nand_5 g02840(new_n3225, new_n1080, new_n3226);
nand_5 g02841(new_n3226, new_n1075, new_n3227);
nand_5 g02842(new_n3227, new_n1070, new_n3228);
nand_5 g02843(new_n3228, new_n1143, new_n3229);
nand_5 g02844(new_n3229, new_n1148, new_n3230);
nand_5 g02845(new_n3230, new_n1065, new_n3231);
nand_5 g02846(new_n3231, new_n1062, new_n3232);
nand_5 g02847(new_n3232, new_n1156, new_n3233);
nand_5 g02848(new_n3233, new_n1057, new_n3234);
nand_5 g02849(new_n3234, new_n1053, new_n3235);
nand_5 g02850(new_n3235, new_n1050, new_n3236);
nand_5 g02851(new_n3236, new_n1045, new_n3237);
nand_5 g02852(new_n3237, new_n1040, new_n3238);
nand_5 g02853(new_n3238, new_n1036, new_n3239);
nand_5 g02854(new_n3239, new_n1033, new_n3240);
nand_5 g02855(new_n3240, new_n1028, new_n3241);
nand_5 g02856(new_n3241, new_n1026, new_n3242_1);
nand_5 g02857(new_n3242_1, new_n1021, new_n3243);
nand_5 g02858(new_n3243, new_n1017, new_n3244);
nand_5 g02859(new_n3244, new_n1012, new_n3245);
nand_5 g02860(new_n3245, new_n1009, new_n3246);
nand_5 g02861(new_n3246, new_n1004, new_n3247);
nand_5 g02862(new_n3247, new_n1000, new_n3248);
nand_5 g02863(new_n3248, new_n995, new_n3249);
nand_5 g02864(new_n3249, new_n990, new_n3250);
nand_5 g02865(new_n3250, new_n985, new_n3251);
nand_5 g02866(new_n3251, new_n981, new_n3252);
nand_5 g02867(new_n3252, new_n1179, new_n3253);
nand_5 g02868(new_n3253, new_n976, new_n3254);
nand_5 g02869(new_n3254, new_n971, new_n3255);
nand_5 g02870(new_n3255, new_n966, new_n3256);
nand_5 g02871(new_n3256, new_n961, new_n3257);
nand_5 g02872(new_n3257, new_n957, new_n3258);
nand_5 g02873(new_n3258, new_n952, new_n3259);
nand_5 g02874(new_n3259, new_n948_1, new_n3260);
nand_5 g02875(new_n3260, new_n943, new_n3261);
nand_5 g02876(new_n3261, new_n941, new_n3262);
nand_5 g02877(new_n3262, new_n938, new_n3263_1);
nand_5 g02878(new_n3263_1, new_n936, new_n3264);
nand_5 g02879(new_n3264, new_n931, new_n3265);
nand_5 g02880(new_n3265, new_n927, new_n3266);
nand_5 g02881(new_n3266, new_n922, new_n3267);
nand_5 g02882(new_n3267, new_n917, new_n3268);
nand_5 g02883(new_n3268, new_n912, new_n3269);
nand_5 g02884(new_n3269, new_n907, new_n3270);
nand_5 g02885(new_n3270, new_n903, new_n3271);
nand_5 g02886(new_n3271, new_n2066, new_n3272);
nand_5 g02887(new_n3272, new_n2063, new_n3273);
nand_5 g02888(new_n3273, new_n2062, new_n3274);
nand_5 g02889(new_n3274, new_n2058, new_n3275);
nand_5 g02890(new_n3275, n8737, new_n3276);
nor_5  g02891(new_n3276, new_n2052, n1927);
not_4  g02892(new_n1678, new_n3278);
not_4  g02893(n6362, new_n3279);
nand_5 g02894(new_n1674, new_n3279, new_n3280);
nand_5 g02895(new_n3280, new_n400, new_n3281);
nand_5 g02896(new_n3281, new_n397, new_n3282);
nand_5 g02897(new_n3282, new_n392, new_n3283);
nand_5 g02898(new_n3283, new_n894, new_n3284);
nand_5 g02899(new_n3284, new_n1087, new_n3285);
nand_5 g02900(new_n3285, new_n1129, new_n3286);
nand_5 g02901(new_n3286, new_n1084, new_n3287);
nand_5 g02902(new_n3287, new_n1134, new_n3288);
nand_5 g02903(new_n3288, new_n1080, new_n3289);
nand_5 g02904(new_n3289, new_n1075, new_n3290);
nand_5 g02905(new_n3290, new_n1070, new_n3291);
nand_5 g02906(new_n3291, new_n1143, new_n3292);
nand_5 g02907(new_n3292, new_n1148, new_n3293);
nand_5 g02908(new_n3293, new_n1065, new_n3294);
nand_5 g02909(new_n3294, new_n1062, new_n3295);
nand_5 g02910(new_n3295, new_n1156, new_n3296);
nand_5 g02911(new_n3296, new_n1057, new_n3297);
nand_5 g02912(new_n3297, new_n1053, new_n3298);
nand_5 g02913(new_n3298, new_n1050, new_n3299);
nand_5 g02914(new_n3299, new_n1045, new_n3300);
nand_5 g02915(new_n3300, new_n1040, new_n3301);
nand_5 g02916(new_n3301, new_n1036, new_n3302);
nand_5 g02917(new_n3302, new_n1033, new_n3303);
nand_5 g02918(new_n3303, new_n1028, new_n3304);
nand_5 g02919(new_n3304, new_n1026, new_n3305);
nand_5 g02920(new_n3305, new_n1021, new_n3306);
nand_5 g02921(new_n3306, new_n1017, new_n3307);
nand_5 g02922(new_n3307, new_n1012, new_n3308);
nand_5 g02923(new_n3308, new_n1009, new_n3309);
nand_5 g02924(new_n3309, new_n1004, new_n3310);
nand_5 g02925(new_n3310, new_n1000, new_n3311);
nand_5 g02926(new_n3311, new_n995, new_n3312);
nand_5 g02927(new_n3312, new_n990, new_n3313);
nand_5 g02928(new_n3313, new_n985, new_n3314);
nand_5 g02929(new_n3314, new_n981, new_n3315);
nand_5 g02930(new_n3315, new_n1179, new_n3316);
nand_5 g02931(new_n3316, new_n976, new_n3317);
nand_5 g02932(new_n3317, new_n971, new_n3318);
nand_5 g02933(new_n3318, new_n966, new_n3319);
nand_5 g02934(new_n3319, new_n961, new_n3320);
nand_5 g02935(new_n3320, new_n957, new_n3321);
nand_5 g02936(new_n3321, new_n952, new_n3322);
nand_5 g02937(new_n3322, new_n948_1, new_n3323);
nand_5 g02938(new_n3323, new_n943, new_n3324);
nand_5 g02939(new_n3324, new_n941, new_n3325);
nand_5 g02940(new_n3325, new_n938, new_n3326);
nand_5 g02941(new_n3326, new_n936, new_n3327);
nand_5 g02942(new_n3327, new_n931, new_n3328);
nand_5 g02943(new_n3328, new_n927, new_n3329);
nand_5 g02944(new_n3329, new_n922, new_n3330);
nand_5 g02945(new_n3330, new_n917, new_n3331);
nand_5 g02946(new_n3331, new_n912, new_n3332);
nand_5 g02947(new_n3332, new_n907, new_n3333);
nand_5 g02948(new_n3333, new_n903, new_n3334);
nand_5 g02949(new_n3334, new_n2066, new_n3335);
nand_5 g02950(new_n3335, new_n2063, new_n3336);
nand_5 g02951(new_n3336, new_n2062, new_n3337);
nand_5 g02952(new_n3337, new_n2058, new_n3338);
nand_5 g02953(new_n3338, new_n2055, new_n3339);
nand_5 g02954(new_n3339, new_n2051, new_n3340_1);
nand_5 g02955(new_n3340_1, new_n2046, new_n3341);
nand_5 g02956(new_n3341, new_n2042, new_n3342);
nand_5 g02957(new_n3342, new_n2039, new_n3343);
nand_5 g02958(new_n3343, new_n2036, new_n3344);
nand_5 g02959(new_n3344, new_n2033, new_n3345);
nand_5 g02960(new_n3345, new_n2029, new_n3346);
nand_5 g02961(new_n3346, new_n2026, new_n3347);
nand_5 g02962(new_n3347, new_n2022, new_n3348);
nand_5 g02963(new_n3348, new_n2018, new_n3349);
nand_5 g02964(new_n3349, new_n1726, new_n3350);
nand_5 g02965(new_n3350, new_n1722, new_n3351);
nand_5 g02966(new_n3351, new_n1718, new_n3352);
nand_5 g02967(new_n3352, new_n1713, new_n3353);
nand_5 g02968(new_n3353, new_n1737, new_n3354);
nand_5 g02969(new_n3354, new_n1709, new_n3355);
nand_5 g02970(new_n3355, new_n1742, new_n3356);
nand_5 g02971(new_n3356, new_n1704, new_n3357);
nand_5 g02972(new_n3357, new_n1702_1, new_n3358);
nand_5 g02973(new_n3358, new_n1698, new_n3359);
nand_5 g02974(new_n3359, new_n1695, new_n3360);
nand_5 g02975(new_n3360, new_n1692, new_n3361);
nand_5 g02976(new_n3361, new_n1752, new_n3362);
nand_5 g02977(new_n3362, new_n1688, new_n3363);
nand_5 g02978(new_n3363, new_n1685, new_n3364);
nand_5 g02979(new_n3364, n10050, new_n3365);
nor_5  g02980(new_n3365, new_n3278, n1951);
nand_5 g02981(new_n2048_1, new_n2046, new_n3367_1);
nand_5 g02982(new_n3367_1, new_n2042, new_n3368);
nand_5 g02983(new_n3368, new_n2039, new_n3369);
nand_5 g02984(new_n3369, new_n2036, new_n3370);
nand_5 g02985(new_n3370, new_n2033, new_n3371);
nand_5 g02986(new_n3371, new_n2029, new_n3372);
nand_5 g02987(new_n3372, new_n2026, new_n3373);
nand_5 g02988(new_n3373, new_n2022, new_n3374);
nand_5 g02989(new_n3374, new_n2018, new_n3375);
nand_5 g02990(new_n3375, new_n1726, new_n3376);
nand_5 g02991(new_n3376, new_n1722, new_n3377);
nand_5 g02992(new_n3377, new_n1718, new_n3378);
nand_5 g02993(new_n3378, new_n1713, new_n3379);
nand_5 g02994(new_n3379, new_n1737, new_n3380);
nand_5 g02995(new_n3380, new_n1709, new_n3381);
nand_5 g02996(new_n3381, new_n1742, new_n3382);
nand_5 g02997(new_n3382, new_n1704, new_n3383);
nand_5 g02998(new_n3383, new_n1702_1, new_n3384);
nand_5 g02999(new_n3384, new_n1698, new_n3385);
nand_5 g03000(new_n3385, new_n1695, new_n3386);
nand_5 g03001(new_n3386, new_n1692, new_n3387);
nand_5 g03002(new_n3387, new_n1752, new_n3388_1);
nand_5 g03003(new_n3388_1, new_n1688, new_n3389);
nand_5 g03004(new_n3389, new_n1685, new_n3390);
nand_5 g03005(new_n3390, new_n1680, new_n3391);
nand_5 g03006(new_n3391, new_n1676, new_n3392);
nand_5 g03007(new_n3392, new_n1672, new_n3393);
nand_5 g03008(new_n3393, new_n1669, new_n3394);
nand_5 g03009(new_n3394, new_n1666, new_n3395);
nand_5 g03010(new_n3395, new_n1663, new_n3396);
nand_5 g03011(new_n3396, new_n1658, new_n3397);
nand_5 g03012(new_n3397, new_n1653, new_n3398);
nand_5 g03013(new_n3398, new_n1651, new_n3399);
nand_5 g03014(new_n3399, new_n1649, new_n3400);
nand_5 g03015(new_n3400, new_n1646, new_n3401);
nand_5 g03016(new_n3401, new_n1643, new_n3402);
nand_5 g03017(new_n3402, new_n1641, new_n3403);
nand_5 g03018(new_n3403, new_n1638, new_n3404);
nand_5 g03019(new_n3404, new_n1635, new_n3405);
nand_5 g03020(new_n3405, new_n1632, new_n3406);
nand_5 g03021(new_n3406, new_n1628, new_n3407);
nand_5 g03022(new_n3407, new_n1625, new_n3408);
nand_5 g03023(new_n3408, new_n1621, new_n3409);
nand_5 g03024(new_n3409, new_n1618, new_n3410);
nand_5 g03025(new_n3410, new_n1778, new_n3411);
nand_5 g03026(new_n3411, new_n1782, new_n3412);
nand_5 g03027(new_n3412, new_n1614, new_n3413);
nand_5 g03028(new_n3413, new_n1611, new_n3414);
nand_5 g03029(new_n3414, new_n1789, new_n3415);
nand_5 g03030(new_n3415, new_n1608, new_n3416);
nand_5 g03031(new_n3416, new_n1605, new_n3417);
nand_5 g03032(new_n3417, new_n1795, new_n3418);
nand_5 g03033(new_n3418, new_n1799, new_n3419);
nand_5 g03034(new_n3419, new_n1602, new_n3420);
nand_5 g03035(new_n3420, new_n1599, new_n3421);
nand_5 g03036(new_n3421, new_n1596, new_n3422);
nand_5 g03037(new_n3422, new_n1593, new_n3423);
nand_5 g03038(new_n3423, new_n1806, new_n3424);
nand_5 g03039(new_n3424, new_n1589, new_n3425);
nand_5 g03040(new_n3425, new_n1586, new_n3426);
nand_5 g03041(new_n3426, new_n1583, new_n3427);
nand_5 g03042(new_n3427, new_n1580, new_n3428);
nand_5 g03043(new_n3428, new_n1576, new_n3429);
nand_5 g03044(new_n3429, new_n1573, new_n3430);
nand_5 g03045(new_n3430, new_n1570, new_n3431);
nand_5 g03046(new_n3431, new_n1567, new_n3432);
nand_5 g03047(new_n3432, new_n1564, new_n3433);
nand_5 g03048(new_n3433, new_n1561, new_n3434);
nand_5 g03049(new_n3434, new_n1338, new_n3435);
nand_5 g03050(new_n3435, new_n1331, new_n3436);
nand_5 g03051(new_n3436, new_n1326, new_n3437);
nand_5 g03052(new_n3437, new_n1321, new_n3438);
nand_5 g03053(new_n3438, new_n1318, new_n3439);
nand_5 g03054(new_n3439, new_n1315, new_n3440);
nand_5 g03055(new_n3440, new_n1312, new_n3441);
nand_5 g03056(new_n3441, new_n1309, new_n3442);
nand_5 g03057(new_n3442, new_n1307, new_n3443);
nand_5 g03058(new_n3443, new_n1304, new_n3444);
nand_5 g03059(new_n3444, new_n1300, new_n3445);
nand_5 g03060(new_n3445, new_n1297, new_n3446);
nand_5 g03061(new_n3446, new_n1294, new_n3447);
nand_5 g03062(new_n3447, new_n1355, new_n3448);
nand_5 g03063(new_n3448, new_n1291, new_n3449);
nand_5 g03064(new_n3449, new_n1288, new_n3450);
nand_5 g03065(new_n3450, n4615, new_n3451);
nor_5  g03066(new_n3451, new_n786, n2027);
not_4  g03067(new_n1426, new_n3453);
nand_5 g03068(new_n1666, new_n3453, new_n3454);
nand_5 g03069(new_n3454, new_n1663, new_n3455);
nand_5 g03070(new_n3455, new_n1658, new_n3456);
nand_5 g03071(new_n3456, new_n1653, new_n3457);
nand_5 g03072(new_n3457, new_n1651, new_n3458);
nand_5 g03073(new_n3458, new_n1649, new_n3459);
nand_5 g03074(new_n3459, new_n1646, new_n3460);
nand_5 g03075(new_n3460, new_n1643, new_n3461);
nand_5 g03076(new_n3461, new_n1641, new_n3462);
nand_5 g03077(new_n3462, new_n1638, new_n3463);
nand_5 g03078(new_n3463, new_n1635, new_n3464);
nand_5 g03079(new_n3464, new_n1632, new_n3465);
nand_5 g03080(new_n3465, new_n1628, new_n3466);
nand_5 g03081(new_n3466, new_n1625, new_n3467);
nand_5 g03082(new_n3467, new_n1621, new_n3468);
nand_5 g03083(new_n3468, new_n1618, new_n3469);
nand_5 g03084(new_n3469, new_n1778, new_n3470);
nand_5 g03085(new_n3470, new_n1782, new_n3471);
nand_5 g03086(new_n3471, new_n1614, new_n3472);
nand_5 g03087(new_n3472, new_n1611, new_n3473);
nand_5 g03088(new_n3473, new_n1789, new_n3474);
nand_5 g03089(new_n3474, new_n1608, new_n3475);
nand_5 g03090(new_n3475, new_n1605, new_n3476);
nand_5 g03091(new_n3476, new_n1795, new_n3477);
nand_5 g03092(new_n3477, new_n1799, new_n3478);
nand_5 g03093(new_n3478, new_n1602, new_n3479);
nand_5 g03094(new_n3479, new_n1599, new_n3480);
nand_5 g03095(new_n3480, new_n1596, new_n3481);
nand_5 g03096(new_n3481, new_n1593, new_n3482);
nand_5 g03097(new_n3482, new_n1806, new_n3483);
nand_5 g03098(new_n3483, new_n1589, new_n3484);
nand_5 g03099(new_n3484, new_n1586, new_n3485);
nand_5 g03100(new_n3485, new_n1583, new_n3486);
nand_5 g03101(new_n3486, new_n1580, new_n3487);
nand_5 g03102(new_n3487, new_n1576, new_n3488);
nand_5 g03103(new_n3488, new_n1573, new_n3489);
nand_5 g03104(new_n3489, new_n1570, new_n3490);
nand_5 g03105(new_n3490, new_n1567, new_n3491);
nand_5 g03106(new_n3491, new_n1564, new_n3492);
nand_5 g03107(new_n3492, new_n1561, new_n3493);
nand_5 g03108(new_n3493, new_n1338, new_n3494);
nand_5 g03109(new_n3494, new_n1331, new_n3495);
nand_5 g03110(new_n3495, new_n1326, new_n3496);
nand_5 g03111(new_n3496, new_n1321, new_n3497);
nand_5 g03112(new_n3497, new_n1318, new_n3498);
nand_5 g03113(new_n3498, new_n1315, new_n3499);
nand_5 g03114(new_n3499, new_n1312, new_n3500);
nand_5 g03115(new_n3500, new_n1309, new_n3501);
nand_5 g03116(new_n3501, new_n1307, new_n3502);
nand_5 g03117(new_n3502, new_n1304, new_n3503);
nand_5 g03118(new_n3503, new_n1300, new_n3504);
nand_5 g03119(new_n3504, new_n1297, new_n3505);
nand_5 g03120(new_n3505, new_n1294, new_n3506_1);
nand_5 g03121(new_n3506_1, new_n1355, new_n3507);
nand_5 g03122(new_n3507, new_n1291, new_n3508);
nand_5 g03123(new_n3508, new_n1288, new_n3509);
nand_5 g03124(new_n3509, new_n1283, new_n3510);
nand_5 g03125(new_n3510, new_n1363, new_n3511);
nand_5 g03126(new_n3511, new_n1280, new_n3512);
nand_5 g03127(new_n3512, new_n1370, new_n3513);
nand_5 g03128(new_n3513, new_n1373, new_n3514);
nand_5 g03129(new_n3514, new_n1277, new_n3515);
nand_5 g03130(new_n3515, new_n1272, new_n3516);
nand_5 g03131(new_n3516, new_n1269, new_n3517);
nand_5 g03132(new_n3517, new_n1380, new_n3518);
nand_5 g03133(new_n3518, new_n1264, new_n3519);
nand_5 g03134(new_n3519, new_n1259, new_n3520);
nand_5 g03135(new_n3520, new_n1388, new_n3521);
nand_5 g03136(new_n3521, new_n1392, new_n3522);
nand_5 g03137(new_n3522, new_n1256, new_n3523);
nand_5 g03138(new_n3523, new_n1252, new_n3524);
nand_5 g03139(new_n3524, new_n1249, new_n3525);
nand_5 g03140(new_n3525, new_n1244, new_n3526);
nand_5 g03141(new_n3526, new_n1240, new_n3527);
nand_5 g03142(new_n3527, new_n1234, new_n3528);
nand_5 g03143(new_n3528, new_n1231, new_n3529);
nand_5 g03144(new_n3529, new_n1227, new_n3530);
nand_5 g03145(new_n3530, new_n1407, new_n3531);
nand_5 g03146(new_n3531, new_n1223, new_n3532_1);
nand_5 g03147(new_n3532_1, new_n1218, new_n3533);
nand_5 g03148(new_n3533, new_n1213, new_n3534);
nand_5 g03149(new_n3534, new_n1210, new_n3535);
nand_5 g03150(new_n3535, new_n1206, new_n3536);
nand_5 g03151(new_n3536, new_n1418, new_n3537);
nand_5 g03152(new_n3537, n4895, new_n3538);
nor_5  g03153(new_n3538, new_n394_1, n2126);
nand_5 g03154(new_n1617, new_n1048, new_n3540);
nand_5 g03155(new_n3540, new_n1045, new_n3541);
nand_5 g03156(new_n3541, new_n1040, new_n3542);
nand_5 g03157(new_n3542, new_n1036, new_n3543);
nand_5 g03158(new_n3543, new_n1033, new_n3544);
nand_5 g03159(new_n3544, new_n1028, new_n3545);
nand_5 g03160(new_n3545, new_n1026, new_n3546);
nand_5 g03161(new_n3546, new_n1021, new_n3547);
nand_5 g03162(new_n3547, new_n1017, new_n3548);
nand_5 g03163(new_n3548, new_n1012, new_n3549);
nand_5 g03164(new_n3549, new_n1009, new_n3550);
nand_5 g03165(new_n3550, new_n1004, new_n3551);
nand_5 g03166(new_n3551, new_n1000, new_n3552);
nand_5 g03167(new_n3552, new_n995, new_n3553);
nand_5 g03168(new_n3553, new_n990, new_n3554);
nand_5 g03169(new_n3554, new_n985, new_n3555);
nand_5 g03170(new_n3555, new_n981, new_n3556);
nand_5 g03171(new_n3556, new_n1179, new_n3557);
nand_5 g03172(new_n3557, new_n976, new_n3558);
nand_5 g03173(new_n3558, new_n971, new_n3559);
nand_5 g03174(new_n3559, new_n966, new_n3560);
nand_5 g03175(new_n3560, new_n961, new_n3561);
nand_5 g03176(new_n3561, new_n957, new_n3562);
nand_5 g03177(new_n3562, new_n952, new_n3563);
nand_5 g03178(new_n3563, new_n948_1, new_n3564);
nand_5 g03179(new_n3564, new_n943, new_n3565);
nand_5 g03180(new_n3565, new_n941, new_n3566);
nand_5 g03181(new_n3566, new_n938, new_n3567);
nand_5 g03182(new_n3567, new_n936, new_n3568);
nand_5 g03183(new_n3568, new_n931, new_n3569);
nand_5 g03184(new_n3569, new_n927, new_n3570);
nand_5 g03185(new_n3570, new_n922, new_n3571);
nand_5 g03186(new_n3571, new_n917, new_n3572);
nand_5 g03187(new_n3572, new_n912, new_n3573);
nand_5 g03188(new_n3573, new_n907, new_n3574);
nand_5 g03189(new_n3574, new_n903, new_n3575);
nand_5 g03190(new_n3575, new_n2066, new_n3576);
nand_5 g03191(new_n3576, new_n2063, new_n3577);
nand_5 g03192(new_n3577, new_n2062, new_n3578);
nand_5 g03193(new_n3578, new_n2058, new_n3579);
nand_5 g03194(new_n3579, new_n2055, new_n3580);
nand_5 g03195(new_n3580, new_n2051, new_n3581);
nand_5 g03196(new_n3581, new_n2046, new_n3582);
nand_5 g03197(new_n3582, new_n2042, new_n3583);
nand_5 g03198(new_n3583, new_n2039, new_n3584);
nand_5 g03199(new_n3584, new_n2036, new_n3585);
nand_5 g03200(new_n3585, new_n2033, new_n3586);
nand_5 g03201(new_n3586, new_n2029, new_n3587);
nand_5 g03202(new_n3587, new_n2026, new_n3588);
nand_5 g03203(new_n3588, new_n2022, new_n3589);
nand_5 g03204(new_n3589, new_n2018, new_n3590);
nand_5 g03205(new_n3590, new_n1726, new_n3591);
nand_5 g03206(new_n3591, new_n1722, new_n3592);
nand_5 g03207(new_n3592, new_n1718, new_n3593);
nand_5 g03208(new_n3593, new_n1713, new_n3594);
nand_5 g03209(new_n3594, new_n1737, new_n3595);
nand_5 g03210(new_n3595, new_n1709, new_n3596);
nand_5 g03211(new_n3596, new_n1742, new_n3597);
nand_5 g03212(new_n3597, new_n1704, new_n3598);
nand_5 g03213(new_n3598, new_n1702_1, new_n3599);
nand_5 g03214(new_n3599, new_n1698, new_n3600);
nand_5 g03215(new_n3600, new_n1695, new_n3601);
nand_5 g03216(new_n3601, new_n1692, new_n3602);
nand_5 g03217(new_n3602, new_n1752, new_n3603_1);
nand_5 g03218(new_n3603_1, new_n1688, new_n3604);
nand_5 g03219(new_n3604, new_n1685, new_n3605);
nand_5 g03220(new_n3605, new_n1680, new_n3606);
nand_5 g03221(new_n3606, new_n1676, new_n3607);
nand_5 g03222(new_n3607, new_n1672, new_n3608);
nand_5 g03223(new_n3608, new_n1669, new_n3609);
nand_5 g03224(new_n3609, new_n1666, new_n3610);
nand_5 g03225(new_n3610, new_n1663, new_n3611);
nand_5 g03226(new_n3611, new_n1658, new_n3612);
nand_5 g03227(new_n3612, new_n1653, new_n3613);
nand_5 g03228(new_n3613, new_n1651, new_n3614);
nand_5 g03229(new_n3614, new_n1649, new_n3615);
nand_5 g03230(new_n3615, new_n1646, new_n3616);
nand_5 g03231(new_n3616, new_n1643, new_n3617);
nand_5 g03232(new_n3617, new_n1641, new_n3618);
nand_5 g03233(new_n3618, new_n1638, new_n3619);
nand_5 g03234(new_n3619, new_n1635, new_n3620);
nand_5 g03235(new_n3620, new_n1632, new_n3621);
nand_5 g03236(new_n3621, new_n1628, new_n3622);
nand_5 g03237(new_n3622, new_n1625, new_n3623);
nand_5 g03238(new_n3623, n13890, new_n3624);
nor_5  g03239(new_n3624, new_n619, n2175);
not_4  g03240(new_n440, new_n3626);
nand_5 g03241(new_n1380, new_n3626, new_n3627);
nand_5 g03242(new_n3627, new_n1264, new_n3628);
nand_5 g03243(new_n3628, new_n1259, new_n3629);
nand_5 g03244(new_n3629, new_n1388, new_n3630);
nand_5 g03245(new_n3630, new_n1392, new_n3631);
nand_5 g03246(new_n3631, new_n1256, new_n3632);
nand_5 g03247(new_n3632, new_n1252, new_n3633);
nand_5 g03248(new_n3633, new_n1249, new_n3634);
nand_5 g03249(new_n3634, new_n1244, new_n3635);
nand_5 g03250(new_n3635, new_n1240, new_n3636);
nand_5 g03251(new_n3636, new_n1234, new_n3637);
nand_5 g03252(new_n3637, new_n1231, new_n3638);
nand_5 g03253(new_n3638, new_n1227, new_n3639);
nand_5 g03254(new_n3639, new_n1407, new_n3640);
nand_5 g03255(new_n3640, new_n1223, new_n3641);
nand_5 g03256(new_n3641, new_n1218, new_n3642);
nand_5 g03257(new_n3642, new_n1213, new_n3643);
nand_5 g03258(new_n3643, new_n1210, new_n3644);
nand_5 g03259(new_n3644, new_n1206, new_n3645);
nand_5 g03260(new_n3645, new_n1418, new_n3646);
nand_5 g03261(new_n3646, new_n1422, new_n3647);
nand_5 g03262(new_n3647, new_n1428, new_n3648);
nand_5 g03263(new_n3648, new_n1203, new_n3649);
nand_5 g03264(new_n3649, new_n1433, new_n3650);
nand_5 g03265(new_n3650, new_n581, new_n3651);
nand_5 g03266(new_n3651, new_n574, new_n3652_1);
nand_5 g03267(new_n3652_1, new_n568, new_n3653);
nand_5 g03268(new_n3653, new_n589, new_n3654);
nand_5 g03269(new_n3654, new_n595, new_n3655_1);
nand_5 g03270(new_n3655_1, new_n601, new_n3656);
nand_5 g03271(new_n3656, new_n563, new_n3657);
nand_5 g03272(new_n3657, new_n608, new_n3658);
nand_5 g03273(new_n3658, new_n558, new_n3659);
nand_5 g03274(new_n3659, new_n615, new_n3660);
nand_5 g03275(new_n3660, new_n553, new_n3661);
nand_5 g03276(new_n3661, new_n622, new_n3662);
nand_5 g03277(new_n3662, new_n628, new_n3663);
nand_5 g03278(new_n3663, new_n548, new_n3664);
nand_5 g03279(new_n3664, new_n543_1, new_n3665);
nand_5 g03280(new_n3665, new_n636, new_n3666);
nand_5 g03281(new_n3666, new_n642, new_n3667);
nand_5 g03282(new_n3667, new_n538, new_n3668);
nand_5 g03283(new_n3668, new_n533, new_n3669);
nand_5 g03284(new_n3669, new_n650_1, new_n3670);
nand_5 g03285(new_n3670, new_n528, new_n3671);
nand_5 g03286(new_n3671, new_n523, new_n3672);
nand_5 g03287(new_n3672, new_n518, new_n3673_1);
nand_5 g03288(new_n3673_1, new_n659, new_n3674);
nand_5 g03289(new_n3674, new_n665, new_n3675);
nand_5 g03290(new_n3675, new_n672, new_n3676);
nand_5 g03291(new_n3676, new_n513, new_n3677);
nand_5 g03292(new_n3677, new_n679, new_n3678);
nand_5 g03293(new_n3678, new_n685, new_n3679);
nand_5 g03294(new_n3679, new_n691, new_n3680);
nand_5 g03295(new_n3680, new_n508, new_n3681);
nand_5 g03296(new_n3681, new_n698, new_n3682);
nand_5 g03297(new_n3682, new_n503, new_n3683);
nand_5 g03298(new_n3683, new_n704, new_n3684);
nand_5 g03299(new_n3684, new_n498_1, new_n3685);
nand_5 g03300(new_n3685, new_n711, new_n3686);
nand_5 g03301(new_n3686, new_n493, new_n3687);
nand_5 g03302(new_n3687, new_n718, new_n3688);
nand_5 g03303(new_n3688, new_n488, new_n3689);
nand_5 g03304(new_n3689, new_n725, new_n3690);
nand_5 g03305(new_n3690, new_n483, new_n3691);
nand_5 g03306(new_n3691, new_n732, new_n3692);
nand_5 g03307(new_n3692, new_n478, new_n3693);
nand_5 g03308(new_n3693, new_n739, new_n3694);
nand_5 g03309(new_n3694, new_n745, new_n3695);
nand_5 g03310(new_n3695, new_n751, new_n3696);
nand_5 g03311(new_n3696, new_n473, new_n3697);
nand_5 g03312(new_n3697, new_n758, new_n3698);
nand_5 g03313(new_n3698, new_n764, new_n3699);
nand_5 g03314(new_n3699, new_n770, new_n3700);
nand_5 g03315(new_n3700, new_n468, new_n3701);
nand_5 g03316(new_n3701, new_n777, new_n3702);
nand_5 g03317(new_n3702, new_n783, new_n3703);
nand_5 g03318(new_n3703, new_n789, new_n3704);
nand_5 g03319(new_n3704, new_n463, new_n3705);
nand_5 g03320(new_n3705, new_n796, new_n3706);
nand_5 g03321(new_n3706, new_n458, new_n3707);
nand_5 g03322(new_n3707, new_n453, new_n3708);
nand_5 g03323(new_n3708, new_n447, new_n3709);
nand_5 g03324(new_n3709, new_n805, new_n3710);
nand_5 g03325(new_n3710, n4175, new_n3711);
nor_5  g03326(new_n3711, new_n808, n2223);
not_4  g03327(new_n1010, new_n3713);
nand_5 g03328(new_n3713, new_n518, new_n3714);
nand_5 g03329(new_n3714, new_n659, new_n3715);
nand_5 g03330(new_n3715, new_n665, new_n3716);
nand_5 g03331(new_n3716, new_n672, new_n3717);
nand_5 g03332(new_n3717, new_n513, new_n3718);
nand_5 g03333(new_n3718, new_n679, new_n3719);
nand_5 g03334(new_n3719, new_n685, new_n3720);
nand_5 g03335(new_n3720, new_n691, new_n3721);
nand_5 g03336(new_n3721, new_n508, new_n3722);
nand_5 g03337(new_n3722, new_n698, new_n3723);
nand_5 g03338(new_n3723, new_n503, new_n3724);
nand_5 g03339(new_n3724, new_n704, new_n3725);
nand_5 g03340(new_n3725, new_n498_1, new_n3726);
nand_5 g03341(new_n3726, new_n711, new_n3727);
nand_5 g03342(new_n3727, new_n493, new_n3728);
nand_5 g03343(new_n3728, new_n718, new_n3729);
nand_5 g03344(new_n3729, new_n488, new_n3730);
nand_5 g03345(new_n3730, new_n725, new_n3731);
nand_5 g03346(new_n3731, new_n483, new_n3732);
nand_5 g03347(new_n3732, new_n732, new_n3733);
nand_5 g03348(new_n3733, new_n478, new_n3734);
nand_5 g03349(new_n3734, new_n739, new_n3735);
nand_5 g03350(new_n3735, new_n745, new_n3736);
nand_5 g03351(new_n3736, new_n751, new_n3737);
nand_5 g03352(new_n3737, new_n473, new_n3738);
nand_5 g03353(new_n3738, new_n758, new_n3739);
nand_5 g03354(new_n3739, new_n764, new_n3740);
nand_5 g03355(new_n3740, new_n770, new_n3741);
nand_5 g03356(new_n3741, new_n468, new_n3742);
nand_5 g03357(new_n3742, new_n777, new_n3743);
nand_5 g03358(new_n3743, new_n783, new_n3744);
nand_5 g03359(new_n3744, new_n789, new_n3745);
nand_5 g03360(new_n3745, new_n463, new_n3746);
nand_5 g03361(new_n3746, new_n796, new_n3747);
nand_5 g03362(new_n3747, new_n458, new_n3748);
nand_5 g03363(new_n3748, new_n453, new_n3749);
nand_5 g03364(new_n3749, new_n447, new_n3750);
nand_5 g03365(new_n3750, new_n805, new_n3751);
nand_5 g03366(new_n3751, new_n811, new_n3752);
nand_5 g03367(new_n3752, new_n442, new_n3753);
nand_5 g03368(new_n3753, new_n437, new_n3754);
nand_5 g03369(new_n3754, new_n819, new_n3755);
nand_5 g03370(new_n3755, new_n432, new_n3756);
nand_5 g03371(new_n3756, new_n427_1, new_n3757);
nand_5 g03372(new_n3757, new_n422, new_n3758);
nand_5 g03373(new_n3758, new_n828, new_n3759);
nand_5 g03374(new_n3759, new_n834, new_n3760);
nand_5 g03375(new_n3760, new_n840, new_n3761);
nand_5 g03376(new_n3761, new_n417, new_n3762);
nand_5 g03377(new_n3762, new_n847, new_n3763);
nand_5 g03378(new_n3763, new_n853, new_n3764);
nand_5 g03379(new_n3764, new_n859, new_n3765);
nand_5 g03380(new_n3765, new_n412, new_n3766);
nand_5 g03381(new_n3766, new_n866, new_n3767);
nand_5 g03382(new_n3767, new_n872, new_n3768);
nand_5 g03383(new_n3768, new_n878, new_n3769);
nand_5 g03384(new_n3769, new_n407, new_n3770);
nand_5 g03385(new_n3770, new_n885, new_n3771);
nand_5 g03386(new_n3771, new_n402, new_n3772);
nand_5 g03387(new_n3772, new_n397, new_n3773);
nand_5 g03388(new_n3773, new_n392, new_n3774);
nand_5 g03389(new_n3774, new_n894, new_n3775_1);
nand_5 g03390(new_n3775_1, new_n1087, new_n3776);
nand_5 g03391(new_n3776, new_n1129, new_n3777);
nand_5 g03392(new_n3777, new_n1084, new_n3778);
nand_5 g03393(new_n3778, new_n1134, new_n3779);
nand_5 g03394(new_n3779, new_n1080, new_n3780);
nand_5 g03395(new_n3780, new_n1075, new_n3781);
nand_5 g03396(new_n3781, new_n1070, new_n3782);
nand_5 g03397(new_n3782, new_n1143, new_n3783);
nand_5 g03398(new_n3783, new_n1148, new_n3784);
nand_5 g03399(new_n3784, new_n1065, new_n3785);
nand_5 g03400(new_n3785, new_n1062, new_n3786);
nand_5 g03401(new_n3786, new_n1156, new_n3787);
nand_5 g03402(new_n3787, new_n1057, new_n3788);
nand_5 g03403(new_n3788, new_n1053, new_n3789);
nand_5 g03404(new_n3789, new_n1050, new_n3790);
nand_5 g03405(new_n3790, new_n1045, new_n3791);
nand_5 g03406(new_n3791, new_n1040, new_n3792);
nand_5 g03407(new_n3792, new_n1036, new_n3793);
nand_5 g03408(new_n3793, new_n1033, new_n3794);
nand_5 g03409(new_n3794, new_n1028, new_n3795);
nand_5 g03410(new_n3795, new_n1026, new_n3796);
nand_5 g03411(new_n3796, new_n1021, new_n3797);
nand_5 g03412(new_n3797, n3804, new_n3798);
nor_5  g03413(new_n3798, new_n1014, n2311);
nand_5 g03414(new_n1715, new_n1713, new_n3800);
nand_5 g03415(new_n3800, new_n1737, new_n3801);
nand_5 g03416(new_n3801, new_n1709, new_n3802);
nand_5 g03417(new_n3802, new_n1742, new_n3803);
nand_5 g03418(new_n3803, new_n1704, new_n3804_1);
nand_5 g03419(new_n3804_1, new_n1702_1, new_n3805);
nand_5 g03420(new_n3805, new_n1698, new_n3806);
nand_5 g03421(new_n3806, new_n1695, new_n3807);
nand_5 g03422(new_n3807, new_n1692, new_n3808);
nand_5 g03423(new_n3808, new_n1752, new_n3809);
nand_5 g03424(new_n3809, new_n1688, new_n3810);
nand_5 g03425(new_n3810, new_n1685, new_n3811);
nand_5 g03426(new_n3811, new_n1680, new_n3812);
nand_5 g03427(new_n3812, new_n1676, new_n3813);
nand_5 g03428(new_n3813, new_n1672, new_n3814);
nand_5 g03429(new_n3814, new_n1669, new_n3815);
nand_5 g03430(new_n3815, new_n1666, new_n3816);
nand_5 g03431(new_n3816, new_n1663, new_n3817);
nand_5 g03432(new_n3817, new_n1658, new_n3818);
nand_5 g03433(new_n3818, new_n1653, new_n3819);
nand_5 g03434(new_n3819, new_n1651, new_n3820);
nand_5 g03435(new_n3820, new_n1649, new_n3821);
nand_5 g03436(new_n3821, new_n1646, new_n3822);
nand_5 g03437(new_n3822, new_n1643, new_n3823);
nand_5 g03438(new_n3823, new_n1641, new_n3824);
nand_5 g03439(new_n3824, new_n1638, new_n3825);
nand_5 g03440(new_n3825, new_n1635, new_n3826);
nand_5 g03441(new_n3826, new_n1632, new_n3827);
nand_5 g03442(new_n3827, new_n1628, new_n3828);
nand_5 g03443(new_n3828, new_n1625, new_n3829);
nand_5 g03444(new_n3829, new_n1621, new_n3830);
nand_5 g03445(new_n3830, new_n1618, new_n3831);
nand_5 g03446(new_n3831, new_n1778, new_n3832);
nand_5 g03447(new_n3832, new_n1782, new_n3833_1);
nand_5 g03448(new_n3833_1, new_n1614, new_n3834);
nand_5 g03449(new_n3834, new_n1611, new_n3835);
nand_5 g03450(new_n3835, new_n1789, new_n3836);
nand_5 g03451(new_n3836, new_n1608, new_n3837);
nand_5 g03452(new_n3837, new_n1605, new_n3838);
nand_5 g03453(new_n3838, new_n1795, new_n3839);
nand_5 g03454(new_n3839, new_n1799, new_n3840);
nand_5 g03455(new_n3840, new_n1602, new_n3841);
nand_5 g03456(new_n3841, new_n1599, new_n3842);
nand_5 g03457(new_n3842, new_n1596, new_n3843);
nand_5 g03458(new_n3843, new_n1593, new_n3844);
nand_5 g03459(new_n3844, new_n1806, new_n3845);
nand_5 g03460(new_n3845, new_n1589, new_n3846);
nand_5 g03461(new_n3846, new_n1586, new_n3847);
nand_5 g03462(new_n3847, new_n1583, new_n3848);
nand_5 g03463(new_n3848, new_n1580, new_n3849);
nand_5 g03464(new_n3849, new_n1576, new_n3850);
nand_5 g03465(new_n3850, new_n1573, new_n3851);
nand_5 g03466(new_n3851, new_n1570, new_n3852);
nand_5 g03467(new_n3852, new_n1567, new_n3853);
nand_5 g03468(new_n3853, new_n1564, new_n3854_1);
nand_5 g03469(new_n3854_1, new_n1561, new_n3855);
nand_5 g03470(new_n3855, new_n1338, new_n3856);
nand_5 g03471(new_n3856, new_n1331, new_n3857);
nand_5 g03472(new_n3857, new_n1326, new_n3858);
nand_5 g03473(new_n3858, new_n1321, new_n3859);
nand_5 g03474(new_n3859, new_n1318, new_n3860);
nand_5 g03475(new_n3860, new_n1315, new_n3861);
nand_5 g03476(new_n3861, new_n1312, new_n3862);
nand_5 g03477(new_n3862, new_n1309, new_n3863);
nand_5 g03478(new_n3863, new_n1307, new_n3864);
nand_5 g03479(new_n3864, new_n1304, new_n3865);
nand_5 g03480(new_n3865, new_n1300, new_n3866);
nand_5 g03481(new_n3866, new_n1297, new_n3867);
nand_5 g03482(new_n3867, new_n1294, new_n3868);
nand_5 g03483(new_n3868, new_n1355, new_n3869);
nand_5 g03484(new_n3869, new_n1291, new_n3870);
nand_5 g03485(new_n3870, new_n1288, new_n3871);
nand_5 g03486(new_n3871, new_n1283, new_n3872);
nand_5 g03487(new_n3872, new_n1363, new_n3873);
nand_5 g03488(new_n3873, new_n1280, new_n3874);
nand_5 g03489(new_n3874, new_n1370, new_n3875);
nand_5 g03490(new_n3875, new_n1373, new_n3876);
nand_5 g03491(new_n3876, new_n1277, new_n3877);
nand_5 g03492(new_n3877, new_n1272, new_n3878);
nand_5 g03493(new_n3878, new_n1269, new_n3879);
nand_5 g03494(new_n3879, new_n1380, new_n3880);
nand_5 g03495(new_n3880, new_n1264, new_n3881);
nand_5 g03496(new_n3881, new_n1259, new_n3882);
nand_5 g03497(new_n3882, new_n1388, new_n3883);
nand_5 g03498(new_n3883, n10147, new_n3884);
nor_5  g03499(new_n3884, new_n424, n2407);
not_4  g03500(new_n1594, new_n3886);
nand_5 g03501(new_n3886, new_n1000, new_n3887);
nand_5 g03502(new_n3887, new_n995, new_n3888);
nand_5 g03503(new_n3888, new_n990, new_n3889);
nand_5 g03504(new_n3889, new_n985, new_n3890);
nand_5 g03505(new_n3890, new_n981, new_n3891);
nand_5 g03506(new_n3891, new_n1179, new_n3892);
nand_5 g03507(new_n3892, new_n976, new_n3893_1);
nand_5 g03508(new_n3893_1, new_n971, new_n3894);
nand_5 g03509(new_n3894, new_n966, new_n3895);
nand_5 g03510(new_n3895, new_n961, new_n3896);
nand_5 g03511(new_n3896, new_n957, new_n3897);
nand_5 g03512(new_n3897, new_n952, new_n3898);
nand_5 g03513(new_n3898, new_n948_1, new_n3899);
nand_5 g03514(new_n3899, new_n943, new_n3900);
nand_5 g03515(new_n3900, new_n941, new_n3901_1);
nand_5 g03516(new_n3901_1, new_n938, new_n3902);
nand_5 g03517(new_n3902, new_n936, new_n3903);
nand_5 g03518(new_n3903, new_n931, new_n3904);
nand_5 g03519(new_n3904, new_n927, new_n3905);
nand_5 g03520(new_n3905, new_n922, new_n3906);
nand_5 g03521(new_n3906, new_n917, new_n3907);
nand_5 g03522(new_n3907, new_n912, new_n3908);
nand_5 g03523(new_n3908, new_n907, new_n3909);
nand_5 g03524(new_n3909, new_n903, new_n3910_1);
nand_5 g03525(new_n3910_1, new_n2066, new_n3911);
nand_5 g03526(new_n3911, new_n2063, new_n3912);
nand_5 g03527(new_n3912, new_n2062, new_n3913);
nand_5 g03528(new_n3913, new_n2058, new_n3914);
nand_5 g03529(new_n3914, new_n2055, new_n3915);
nand_5 g03530(new_n3915, new_n2051, new_n3916);
nand_5 g03531(new_n3916, new_n2046, new_n3917);
nand_5 g03532(new_n3917, new_n2042, new_n3918);
nand_5 g03533(new_n3918, new_n2039, new_n3919);
nand_5 g03534(new_n3919, new_n2036, new_n3920);
nand_5 g03535(new_n3920, new_n2033, new_n3921);
nand_5 g03536(new_n3921, new_n2029, new_n3922);
nand_5 g03537(new_n3922, new_n2026, new_n3923);
nand_5 g03538(new_n3923, new_n2022, new_n3924);
nand_5 g03539(new_n3924, new_n2018, new_n3925);
nand_5 g03540(new_n3925, new_n1726, new_n3926);
nand_5 g03541(new_n3926, new_n1722, new_n3927);
nand_5 g03542(new_n3927, new_n1718, new_n3928);
nand_5 g03543(new_n3928, new_n1713, new_n3929);
nand_5 g03544(new_n3929, new_n1737, new_n3930);
nand_5 g03545(new_n3930, new_n1709, new_n3931);
nand_5 g03546(new_n3931, new_n1742, new_n3932);
nand_5 g03547(new_n3932, new_n1704, new_n3933);
nand_5 g03548(new_n3933, new_n1702_1, new_n3934);
nand_5 g03549(new_n3934, new_n1698, new_n3935);
nand_5 g03550(new_n3935, new_n1695, new_n3936);
nand_5 g03551(new_n3936, new_n1692, new_n3937);
nand_5 g03552(new_n3937, new_n1752, new_n3938);
nand_5 g03553(new_n3938, new_n1688, new_n3939);
nand_5 g03554(new_n3939, new_n1685, new_n3940);
nand_5 g03555(new_n3940, new_n1680, new_n3941);
nand_5 g03556(new_n3941, new_n1676, new_n3942);
nand_5 g03557(new_n3942, new_n1672, new_n3943);
nand_5 g03558(new_n3943, new_n1669, new_n3944);
nand_5 g03559(new_n3944, new_n1666, new_n3945);
nand_5 g03560(new_n3945, new_n1663, new_n3946);
nand_5 g03561(new_n3946, new_n1658, new_n3947);
nand_5 g03562(new_n3947, new_n1653, new_n3948);
nand_5 g03563(new_n3948, new_n1651, new_n3949);
nand_5 g03564(new_n3949, new_n1649, new_n3950);
nand_5 g03565(new_n3950, new_n1646, new_n3951);
nand_5 g03566(new_n3951, new_n1643, new_n3952);
nand_5 g03567(new_n3952, new_n1641, new_n3953);
nand_5 g03568(new_n3953, new_n1638, new_n3954);
nand_5 g03569(new_n3954, new_n1635, new_n3955);
nand_5 g03570(new_n3955, new_n1632, new_n3956);
nand_5 g03571(new_n3956, new_n1628, new_n3957);
nand_5 g03572(new_n3957, new_n1625, new_n3958);
nand_5 g03573(new_n3958, new_n1621, new_n3959);
nand_5 g03574(new_n3959, new_n1618, new_n3960);
nand_5 g03575(new_n3960, new_n1778, new_n3961);
nand_5 g03576(new_n3961, new_n1782, new_n3962);
nand_5 g03577(new_n3962, new_n1614, new_n3963);
nand_5 g03578(new_n3963, new_n1611, new_n3964);
nand_5 g03579(new_n3964, new_n1789, new_n3965);
nand_5 g03580(new_n3965, new_n1608, new_n3966);
nand_5 g03581(new_n3966, new_n1605, new_n3967);
nand_5 g03582(new_n3967, new_n1795, new_n3968);
nand_5 g03583(new_n3968, new_n1799, new_n3969);
nand_5 g03584(new_n3969, new_n1602, new_n3970);
nand_5 g03585(new_n3970, n8799, new_n3971);
nor_5  g03586(new_n3971, new_n656_1, n2556);
nand_5 g03587(new_n1644, new_n588, new_n3973);
nand_5 g03588(new_n3973, new_n1643, new_n3974);
nand_5 g03589(new_n3974, new_n1641, new_n3975);
nand_5 g03590(new_n3975, new_n1638, new_n3976);
nand_5 g03591(new_n3976, new_n1635, new_n3977);
nand_5 g03592(new_n3977, new_n1632, new_n3978);
nand_5 g03593(new_n3978, new_n1628, new_n3979);
nand_5 g03594(new_n3979, new_n1625, new_n3980);
nand_5 g03595(new_n3980, new_n1621, new_n3981);
nand_5 g03596(new_n3981, new_n1618, new_n3982);
nand_5 g03597(new_n3982, new_n1778, new_n3983);
nand_5 g03598(new_n3983, new_n1782, new_n3984);
nand_5 g03599(new_n3984, new_n1614, new_n3985);
nand_5 g03600(new_n3985, new_n1611, new_n3986);
nand_5 g03601(new_n3986, new_n1789, new_n3987);
nand_5 g03602(new_n3987, new_n1608, new_n3988);
nand_5 g03603(new_n3988, new_n1605, new_n3989);
nand_5 g03604(new_n3989, new_n1795, new_n3990);
nand_5 g03605(new_n3990, new_n1799, new_n3991);
nand_5 g03606(new_n3991, new_n1602, new_n3992);
nand_5 g03607(new_n3992, new_n1599, new_n3993);
nand_5 g03608(new_n3993, new_n1596, new_n3994);
nand_5 g03609(new_n3994, new_n1593, new_n3995);
nand_5 g03610(new_n3995, new_n1806, new_n3996);
nand_5 g03611(new_n3996, new_n1589, new_n3997);
nand_5 g03612(new_n3997, new_n1586, new_n3998);
nand_5 g03613(new_n3998, new_n1583, new_n3999);
nand_5 g03614(new_n3999, new_n1580, new_n4000_1);
nand_5 g03615(new_n4000_1, new_n1576, new_n4001);
nand_5 g03616(new_n4001, new_n1573, new_n4002);
nand_5 g03617(new_n4002, new_n1570, new_n4003);
nand_5 g03618(new_n4003, new_n1567, new_n4004);
nand_5 g03619(new_n4004, new_n1564, new_n4005);
nand_5 g03620(new_n4005, new_n1561, new_n4006);
nand_5 g03621(new_n4006, new_n1338, new_n4007);
nand_5 g03622(new_n4007, new_n1331, new_n4008);
nand_5 g03623(new_n4008, new_n1326, new_n4009);
nand_5 g03624(new_n4009, new_n1321, new_n4010);
nand_5 g03625(new_n4010, new_n1318, new_n4011);
nand_5 g03626(new_n4011, new_n1315, new_n4012);
nand_5 g03627(new_n4012, new_n1312, new_n4013);
nand_5 g03628(new_n4013, new_n1309, new_n4014);
nand_5 g03629(new_n4014, new_n1307, new_n4015);
nand_5 g03630(new_n4015, new_n1304, new_n4016);
nand_5 g03631(new_n4016, new_n1300, new_n4017);
nand_5 g03632(new_n4017, new_n1297, new_n4018);
nand_5 g03633(new_n4018, new_n1294, new_n4019);
nand_5 g03634(new_n4019, new_n1355, new_n4020);
nand_5 g03635(new_n4020, new_n1291, new_n4021);
nand_5 g03636(new_n4021, new_n1288, new_n4022_1);
nand_5 g03637(new_n4022_1, new_n1283, new_n4023);
nand_5 g03638(new_n4023, new_n1363, new_n4024);
nand_5 g03639(new_n4024, new_n1280, new_n4025);
nand_5 g03640(new_n4025, new_n1370, new_n4026);
nand_5 g03641(new_n4026, new_n1373, new_n4027);
nand_5 g03642(new_n4027, new_n1277, new_n4028);
nand_5 g03643(new_n4028, new_n1272, new_n4029);
nand_5 g03644(new_n4029, new_n1269, new_n4030);
nand_5 g03645(new_n4030, new_n1380, new_n4031);
nand_5 g03646(new_n4031, new_n1264, new_n4032);
nand_5 g03647(new_n4032, new_n1259, new_n4033);
nand_5 g03648(new_n4033, new_n1388, new_n4034);
nand_5 g03649(new_n4034, new_n1392, new_n4035);
nand_5 g03650(new_n4035, new_n1256, new_n4036);
nand_5 g03651(new_n4036, new_n1252, new_n4037);
nand_5 g03652(new_n4037, new_n1249, new_n4038);
nand_5 g03653(new_n4038, new_n1244, new_n4039_1);
nand_5 g03654(new_n4039_1, new_n1240, new_n4040);
nand_5 g03655(new_n4040, new_n1234, new_n4041);
nand_5 g03656(new_n4041, new_n1231, new_n4042);
nand_5 g03657(new_n4042, new_n1227, new_n4043);
nand_5 g03658(new_n4043, new_n1407, new_n4044);
nand_5 g03659(new_n4044, new_n1223, new_n4045);
nand_5 g03660(new_n4045, new_n1218, new_n4046);
nand_5 g03661(new_n4046, new_n1213, new_n4047);
nand_5 g03662(new_n4047, new_n1210, new_n4048);
nand_5 g03663(new_n4048, new_n1206, new_n4049);
nand_5 g03664(new_n4049, new_n1418, new_n4050);
nand_5 g03665(new_n4050, new_n1422, new_n4051);
nand_5 g03666(new_n4051, new_n1428, new_n4052);
nand_5 g03667(new_n4052, new_n1203, new_n4053);
nand_5 g03668(new_n4053, new_n1433, new_n4054);
nand_5 g03669(new_n4054, new_n581, new_n4055);
nand_5 g03670(new_n4055, new_n574, new_n4056);
nand_5 g03671(new_n4056, n7832, new_n4057);
nor_5  g03672(new_n4057, new_n565, n2559);
not_4  g03673(new_n448, new_n4059);
nand_5 g03674(new_n1373, new_n4059, new_n4060);
nand_5 g03675(new_n4060, new_n1277, new_n4061);
nand_5 g03676(new_n4061, new_n1272, new_n4062);
nand_5 g03677(new_n4062, new_n1269, new_n4063);
nand_5 g03678(new_n4063, new_n1380, new_n4064);
nand_5 g03679(new_n4064, new_n1264, new_n4065);
nand_5 g03680(new_n4065, new_n1259, new_n4066);
nand_5 g03681(new_n4066, new_n1388, new_n4067);
nand_5 g03682(new_n4067, new_n1392, new_n4068);
nand_5 g03683(new_n4068, new_n1256, new_n4069);
nand_5 g03684(new_n4069, new_n1252, new_n4070);
nand_5 g03685(new_n4070, new_n1249, new_n4071);
nand_5 g03686(new_n4071, new_n1244, new_n4072);
nand_5 g03687(new_n4072, new_n1240, new_n4073);
nand_5 g03688(new_n4073, new_n1234, new_n4074);
nand_5 g03689(new_n4074, new_n1231, new_n4075);
nand_5 g03690(new_n4075, new_n1227, new_n4076);
nand_5 g03691(new_n4076, new_n1407, new_n4077);
nand_5 g03692(new_n4077, new_n1223, new_n4078);
nand_5 g03693(new_n4078, new_n1218, new_n4079);
nand_5 g03694(new_n4079, new_n1213, new_n4080);
nand_5 g03695(new_n4080, new_n1210, new_n4081);
nand_5 g03696(new_n4081, new_n1206, new_n4082);
nand_5 g03697(new_n4082, new_n1418, new_n4083);
nand_5 g03698(new_n4083, new_n1422, new_n4084);
nand_5 g03699(new_n4084, new_n1428, new_n4085);
nand_5 g03700(new_n4085, new_n1203, new_n4086);
nand_5 g03701(new_n4086, new_n1433, new_n4087);
nand_5 g03702(new_n4087, new_n581, new_n4088);
nand_5 g03703(new_n4088, new_n574, new_n4089);
nand_5 g03704(new_n4089, new_n568, new_n4090);
nand_5 g03705(new_n4090, new_n589, new_n4091);
nand_5 g03706(new_n4091, new_n595, new_n4092);
nand_5 g03707(new_n4092, new_n601, new_n4093);
nand_5 g03708(new_n4093, new_n563, new_n4094);
nand_5 g03709(new_n4094, new_n608, new_n4095);
nand_5 g03710(new_n4095, new_n558, new_n4096);
nand_5 g03711(new_n4096, new_n615, new_n4097);
nand_5 g03712(new_n4097, new_n553, new_n4098);
nand_5 g03713(new_n4098, new_n622, new_n4099);
nand_5 g03714(new_n4099, new_n628, new_n4100);
nand_5 g03715(new_n4100, new_n548, new_n4101);
nand_5 g03716(new_n4101, new_n543_1, new_n4102);
nand_5 g03717(new_n4102, new_n636, new_n4103);
nand_5 g03718(new_n4103, new_n642, new_n4104);
nand_5 g03719(new_n4104, new_n538, new_n4105);
nand_5 g03720(new_n4105, new_n533, new_n4106);
nand_5 g03721(new_n4106, new_n650_1, new_n4107);
nand_5 g03722(new_n4107, new_n528, new_n4108);
nand_5 g03723(new_n4108, new_n523, new_n4109);
nand_5 g03724(new_n4109, new_n518, new_n4110);
nand_5 g03725(new_n4110, new_n659, new_n4111);
nand_5 g03726(new_n4111, new_n665, new_n4112);
nand_5 g03727(new_n4112, new_n672, new_n4113);
nand_5 g03728(new_n4113, new_n513, new_n4114);
nand_5 g03729(new_n4114, new_n679, new_n4115);
nand_5 g03730(new_n4115, new_n685, new_n4116);
nand_5 g03731(new_n4116, new_n691, new_n4117_1);
nand_5 g03732(new_n4117_1, new_n508, new_n4118);
nand_5 g03733(new_n4118, new_n698, new_n4119);
nand_5 g03734(new_n4119, new_n503, new_n4120);
nand_5 g03735(new_n4120, new_n704, new_n4121);
nand_5 g03736(new_n4121, new_n498_1, new_n4122);
nand_5 g03737(new_n4122, new_n711, new_n4123);
nand_5 g03738(new_n4123, new_n493, new_n4124);
nand_5 g03739(new_n4124, new_n718, new_n4125_1);
nand_5 g03740(new_n4125_1, new_n488, new_n4126);
nand_5 g03741(new_n4126, new_n725, new_n4127);
nand_5 g03742(new_n4127, new_n483, new_n4128);
nand_5 g03743(new_n4128, new_n732, new_n4129);
nand_5 g03744(new_n4129, new_n478, new_n4130);
nand_5 g03745(new_n4130, new_n739, new_n4131_1);
nand_5 g03746(new_n4131_1, new_n745, new_n4132);
nand_5 g03747(new_n4132, new_n751, new_n4133);
nand_5 g03748(new_n4133, new_n473, new_n4134);
nand_5 g03749(new_n4134, new_n758, new_n4135);
nand_5 g03750(new_n4135, new_n764, new_n4136);
nand_5 g03751(new_n4136, new_n770, new_n4137);
nand_5 g03752(new_n4137, new_n468, new_n4138);
nand_5 g03753(new_n4138, new_n777, new_n4139);
nand_5 g03754(new_n4139, new_n783, new_n4140);
nand_5 g03755(new_n4140, new_n789, new_n4141);
nand_5 g03756(new_n4141, new_n463, new_n4142);
nand_5 g03757(new_n4142, new_n796, new_n4143);
nand_5 g03758(new_n4143, n3263, new_n4144);
nor_5  g03759(new_n4144, new_n455, n2572);
not_4  g03760(new_n1055, new_n4146);
not_4  g03761(new_n1051, new_n4147_1);
nand_5 g03762(new_n4147_1, new_n628, new_n4148);
nand_5 g03763(new_n4148, new_n548, new_n4149);
nand_5 g03764(new_n4149, new_n543_1, new_n4150);
nand_5 g03765(new_n4150, new_n636, new_n4151);
nand_5 g03766(new_n4151, new_n642, new_n4152);
nand_5 g03767(new_n4152, new_n538, new_n4153);
nand_5 g03768(new_n4153, new_n533, new_n4154_1);
nand_5 g03769(new_n4154_1, new_n650_1, new_n4155);
nand_5 g03770(new_n4155, new_n528, new_n4156);
nand_5 g03771(new_n4156, new_n523, new_n4157);
nand_5 g03772(new_n4157, new_n518, new_n4158);
nand_5 g03773(new_n4158, new_n659, new_n4159);
nand_5 g03774(new_n4159, new_n665, new_n4160);
nand_5 g03775(new_n4160, new_n672, new_n4161);
nand_5 g03776(new_n4161, new_n513, new_n4162);
nand_5 g03777(new_n4162, new_n679, new_n4163);
nand_5 g03778(new_n4163, new_n685, new_n4164);
nand_5 g03779(new_n4164, new_n691, new_n4165);
nand_5 g03780(new_n4165, new_n508, new_n4166);
nand_5 g03781(new_n4166, new_n698, new_n4167);
nand_5 g03782(new_n4167, new_n503, new_n4168);
nand_5 g03783(new_n4168, new_n704, new_n4169);
nand_5 g03784(new_n4169, new_n498_1, new_n4170);
nand_5 g03785(new_n4170, new_n711, new_n4171);
nand_5 g03786(new_n4171, new_n493, new_n4172_1);
nand_5 g03787(new_n4172_1, new_n718, new_n4173);
nand_5 g03788(new_n4173, new_n488, new_n4174);
nand_5 g03789(new_n4174, new_n725, new_n4175_1);
nand_5 g03790(new_n4175_1, new_n483, new_n4176);
nand_5 g03791(new_n4176, new_n732, new_n4177);
nand_5 g03792(new_n4177, new_n478, new_n4178);
nand_5 g03793(new_n4178, new_n739, new_n4179);
nand_5 g03794(new_n4179, new_n745, new_n4180);
nand_5 g03795(new_n4180, new_n751, new_n4181);
nand_5 g03796(new_n4181, new_n473, new_n4182);
nand_5 g03797(new_n4182, new_n758, new_n4183);
nand_5 g03798(new_n4183, new_n764, new_n4184);
nand_5 g03799(new_n4184, new_n770, new_n4185);
nand_5 g03800(new_n4185, new_n468, new_n4186);
nand_5 g03801(new_n4186, new_n777, new_n4187);
nand_5 g03802(new_n4187, new_n783, new_n4188);
nand_5 g03803(new_n4188, new_n789, new_n4189);
nand_5 g03804(new_n4189, new_n463, new_n4190);
nand_5 g03805(new_n4190, new_n796, new_n4191);
nand_5 g03806(new_n4191, new_n458, new_n4192);
nand_5 g03807(new_n4192, new_n453, new_n4193);
nand_5 g03808(new_n4193, new_n447, new_n4194);
nand_5 g03809(new_n4194, new_n805, new_n4195);
nand_5 g03810(new_n4195, new_n811, new_n4196);
nand_5 g03811(new_n4196, new_n442, new_n4197);
nand_5 g03812(new_n4197, new_n437, new_n4198);
nand_5 g03813(new_n4198, new_n819, new_n4199);
nand_5 g03814(new_n4199, new_n432, new_n4200);
nand_5 g03815(new_n4200, new_n427_1, new_n4201);
nand_5 g03816(new_n4201, new_n422, new_n4202);
nand_5 g03817(new_n4202, new_n828, new_n4203);
nand_5 g03818(new_n4203, new_n834, new_n4204);
nand_5 g03819(new_n4204, new_n840, new_n4205);
nand_5 g03820(new_n4205, new_n417, new_n4206);
nand_5 g03821(new_n4206, new_n847, new_n4207);
nand_5 g03822(new_n4207, new_n853, new_n4208);
nand_5 g03823(new_n4208, new_n859, new_n4209);
nand_5 g03824(new_n4209, new_n412, new_n4210);
nand_5 g03825(new_n4210, new_n866, new_n4211);
nand_5 g03826(new_n4211, new_n872, new_n4212);
nand_5 g03827(new_n4212, new_n878, new_n4213);
nand_5 g03828(new_n4213, new_n407, new_n4214);
nand_5 g03829(new_n4214, new_n885, new_n4215);
nand_5 g03830(new_n4215, new_n402, new_n4216);
nand_5 g03831(new_n4216, new_n397, new_n4217);
nand_5 g03832(new_n4217, new_n392, new_n4218);
nand_5 g03833(new_n4218, new_n894, new_n4219);
nand_5 g03834(new_n4219, new_n1087, new_n4220);
nand_5 g03835(new_n4220, new_n1129, new_n4221);
nand_5 g03836(new_n4221, new_n1084, new_n4222);
nand_5 g03837(new_n4222, new_n1134, new_n4223);
nand_5 g03838(new_n4223, new_n1080, new_n4224);
nand_5 g03839(new_n4224, new_n1075, new_n4225_1);
nand_5 g03840(new_n4225_1, new_n1070, new_n4226);
nand_5 g03841(new_n4226, new_n1143, new_n4227);
nand_5 g03842(new_n4227, new_n1148, new_n4228);
nand_5 g03843(new_n4228, new_n1065, new_n4229);
nand_5 g03844(new_n4229, new_n1062, new_n4230);
nand_5 g03845(new_n4230, new_n1156, new_n4231);
nand_5 g03846(new_n4231, n9977, new_n4232);
nor_5  g03847(new_n4232, new_n4146, n2672);
nand_5 g03848(new_n984, new_n683, new_n4234);
nand_5 g03849(new_n4234, new_n691, new_n4235);
nand_5 g03850(new_n4235, new_n508, new_n4236);
nand_5 g03851(new_n4236, new_n698, new_n4237);
nand_5 g03852(new_n4237, new_n503, new_n4238);
nand_5 g03853(new_n4238, new_n704, new_n4239);
nand_5 g03854(new_n4239, new_n498_1, new_n4240);
nand_5 g03855(new_n4240, new_n711, new_n4241);
nand_5 g03856(new_n4241, new_n493, new_n4242);
nand_5 g03857(new_n4242, new_n718, new_n4243);
nand_5 g03858(new_n4243, new_n488, new_n4244);
nand_5 g03859(new_n4244, new_n725, new_n4245);
nand_5 g03860(new_n4245, new_n483, new_n4246);
nand_5 g03861(new_n4246, new_n732, new_n4247);
nand_5 g03862(new_n4247, new_n478, new_n4248);
nand_5 g03863(new_n4248, new_n739, new_n4249);
nand_5 g03864(new_n4249, new_n745, new_n4250);
nand_5 g03865(new_n4250, new_n751, new_n4251);
nand_5 g03866(new_n4251, new_n473, new_n4252);
nand_5 g03867(new_n4252, new_n758, new_n4253);
nand_5 g03868(new_n4253, new_n764, new_n4254);
nand_5 g03869(new_n4254, new_n770, new_n4255);
nand_5 g03870(new_n4255, new_n468, new_n4256);
nand_5 g03871(new_n4256, new_n777, new_n4257);
nand_5 g03872(new_n4257, new_n783, new_n4258);
nand_5 g03873(new_n4258, new_n789, new_n4259);
nand_5 g03874(new_n4259, new_n463, new_n4260);
nand_5 g03875(new_n4260, new_n796, new_n4261);
nand_5 g03876(new_n4261, new_n458, new_n4262);
nand_5 g03877(new_n4262, new_n453, new_n4263);
nand_5 g03878(new_n4263, new_n447, new_n4264);
nand_5 g03879(new_n4264, new_n805, new_n4265);
nand_5 g03880(new_n4265, new_n811, new_n4266);
nand_5 g03881(new_n4266, new_n442, new_n4267);
nand_5 g03882(new_n4267, new_n437, new_n4268);
nand_5 g03883(new_n4268, new_n819, new_n4269);
nand_5 g03884(new_n4269, new_n432, new_n4270);
nand_5 g03885(new_n4270, new_n427_1, new_n4271);
nand_5 g03886(new_n4271, new_n422, new_n4272);
nand_5 g03887(new_n4272, new_n828, new_n4273);
nand_5 g03888(new_n4273, new_n834, new_n4274);
nand_5 g03889(new_n4274, new_n840, new_n4275);
nand_5 g03890(new_n4275, new_n417, new_n4276);
nand_5 g03891(new_n4276, new_n847, new_n4277);
nand_5 g03892(new_n4277, new_n853, new_n4278);
nand_5 g03893(new_n4278, new_n859, new_n4279_1);
nand_5 g03894(new_n4279_1, new_n412, new_n4280);
nand_5 g03895(new_n4280, new_n866, new_n4281);
nand_5 g03896(new_n4281, new_n872, new_n4282_1);
nand_5 g03897(new_n4282_1, new_n878, new_n4283);
nand_5 g03898(new_n4283, new_n407, new_n4284);
nand_5 g03899(new_n4284, new_n885, new_n4285);
nand_5 g03900(new_n4285, new_n402, new_n4286);
nand_5 g03901(new_n4286, new_n397, new_n4287);
nand_5 g03902(new_n4287, new_n392, new_n4288);
nand_5 g03903(new_n4288, new_n894, new_n4289);
nand_5 g03904(new_n4289, new_n1087, new_n4290);
nand_5 g03905(new_n4290, new_n1129, new_n4291);
nand_5 g03906(new_n4291, new_n1084, new_n4292_1);
nand_5 g03907(new_n4292_1, new_n1134, new_n4293);
nand_5 g03908(new_n4293, new_n1080, new_n4294);
nand_5 g03909(new_n4294, new_n1075, new_n4295);
nand_5 g03910(new_n4295, new_n1070, new_n4296);
nand_5 g03911(new_n4296, new_n1143, new_n4297);
nand_5 g03912(new_n4297, new_n1148, new_n4298);
nand_5 g03913(new_n4298, new_n1065, new_n4299);
nand_5 g03914(new_n4299, new_n1062, new_n4300);
nand_5 g03915(new_n4300, new_n1156, new_n4301);
nand_5 g03916(new_n4301, new_n1057, new_n4302);
nand_5 g03917(new_n4302, new_n1053, new_n4303);
nand_5 g03918(new_n4303, new_n1050, new_n4304);
nand_5 g03919(new_n4304, new_n1045, new_n4305_1);
nand_5 g03920(new_n4305_1, new_n1040, new_n4306);
nand_5 g03921(new_n4306, new_n1036, new_n4307);
nand_5 g03922(new_n4307, new_n1033, new_n4308);
nand_5 g03923(new_n4308, new_n1028, new_n4309);
nand_5 g03924(new_n4309, new_n1026, new_n4310);
nand_5 g03925(new_n4310, new_n1021, new_n4311);
nand_5 g03926(new_n4311, new_n1017, new_n4312);
nand_5 g03927(new_n4312, new_n1012, new_n4313);
nand_5 g03928(new_n4313, new_n1009, new_n4314);
nand_5 g03929(new_n4314, new_n1004, new_n4315);
nand_5 g03930(new_n4315, new_n1000, new_n4316);
nand_5 g03931(new_n4316, new_n995, new_n4317);
nand_5 g03932(new_n4317, n6703, new_n4318);
nor_5  g03933(new_n4318, new_n987, n2734);
nand_5 g03934(new_n1003, new_n663, new_n4320);
nand_5 g03935(new_n4320, new_n672, new_n4321);
nand_5 g03936(new_n4321, new_n513, new_n4322);
nand_5 g03937(new_n4322, new_n679, new_n4323);
nand_5 g03938(new_n4323, new_n685, new_n4324);
nand_5 g03939(new_n4324, new_n691, new_n4325);
nand_5 g03940(new_n4325, new_n508, new_n4326);
nand_5 g03941(new_n4326, new_n698, new_n4327);
nand_5 g03942(new_n4327, new_n503, new_n4328);
nand_5 g03943(new_n4328, new_n704, new_n4329);
nand_5 g03944(new_n4329, new_n498_1, new_n4330);
nand_5 g03945(new_n4330, new_n711, new_n4331);
nand_5 g03946(new_n4331, new_n493, new_n4332);
nand_5 g03947(new_n4332, new_n718, new_n4333);
nand_5 g03948(new_n4333, new_n488, new_n4334);
nand_5 g03949(new_n4334, new_n725, new_n4335);
nand_5 g03950(new_n4335, new_n483, new_n4336);
nand_5 g03951(new_n4336, new_n732, new_n4337);
nand_5 g03952(new_n4337, new_n478, new_n4338);
nand_5 g03953(new_n4338, new_n739, new_n4339);
nand_5 g03954(new_n4339, new_n745, new_n4340);
nand_5 g03955(new_n4340, new_n751, new_n4341);
nand_5 g03956(new_n4341, new_n473, new_n4342);
nand_5 g03957(new_n4342, new_n758, new_n4343);
nand_5 g03958(new_n4343, new_n764, new_n4344);
nand_5 g03959(new_n4344, new_n770, new_n4345_1);
nand_5 g03960(new_n4345_1, new_n468, new_n4346);
nand_5 g03961(new_n4346, new_n777, new_n4347);
nand_5 g03962(new_n4347, new_n783, new_n4348);
nand_5 g03963(new_n4348, new_n789, new_n4349);
nand_5 g03964(new_n4349, new_n463, new_n4350);
nand_5 g03965(new_n4350, new_n796, new_n4351);
nand_5 g03966(new_n4351, new_n458, new_n4352);
nand_5 g03967(new_n4352, new_n453, new_n4353);
nand_5 g03968(new_n4353, new_n447, new_n4354);
nand_5 g03969(new_n4354, new_n805, new_n4355);
nand_5 g03970(new_n4355, new_n811, new_n4356);
nand_5 g03971(new_n4356, new_n442, new_n4357);
nand_5 g03972(new_n4357, new_n437, new_n4358);
nand_5 g03973(new_n4358, new_n819, new_n4359);
nand_5 g03974(new_n4359, new_n432, new_n4360);
nand_5 g03975(new_n4360, new_n427_1, new_n4361);
nand_5 g03976(new_n4361, new_n422, new_n4362);
nand_5 g03977(new_n4362, new_n828, new_n4363);
nand_5 g03978(new_n4363, new_n834, new_n4364);
nand_5 g03979(new_n4364, new_n840, new_n4365);
nand_5 g03980(new_n4365, new_n417, new_n4366);
nand_5 g03981(new_n4366, new_n847, new_n4367);
nand_5 g03982(new_n4367, new_n853, new_n4368);
nand_5 g03983(new_n4368, new_n859, new_n4369);
nand_5 g03984(new_n4369, new_n412, new_n4370);
nand_5 g03985(new_n4370, new_n866, new_n4371);
nand_5 g03986(new_n4371, new_n872, new_n4372);
nand_5 g03987(new_n4372, new_n878, new_n4373);
nand_5 g03988(new_n4373, new_n407, new_n4374);
nand_5 g03989(new_n4374, new_n885, new_n4375);
nand_5 g03990(new_n4375, new_n402, new_n4376);
nand_5 g03991(new_n4376, new_n397, new_n4377);
nand_5 g03992(new_n4377, new_n392, new_n4378);
nand_5 g03993(new_n4378, new_n894, new_n4379);
nand_5 g03994(new_n4379, new_n1087, new_n4380);
nand_5 g03995(new_n4380, new_n1129, new_n4381);
nand_5 g03996(new_n4381, new_n1084, new_n4382);
nand_5 g03997(new_n4382, new_n1134, new_n4383);
nand_5 g03998(new_n4383, new_n1080, new_n4384);
nand_5 g03999(new_n4384, new_n1075, new_n4385);
nand_5 g04000(new_n4385, new_n1070, new_n4386);
nand_5 g04001(new_n4386, new_n1143, new_n4387);
nand_5 g04002(new_n4387, new_n1148, new_n4388);
nand_5 g04003(new_n4388, new_n1065, new_n4389);
nand_5 g04004(new_n4389, new_n1062, new_n4390);
nand_5 g04005(new_n4390, new_n1156, new_n4391);
nand_5 g04006(new_n4391, new_n1057, new_n4392);
nand_5 g04007(new_n4392, new_n1053, new_n4393);
nand_5 g04008(new_n4393, new_n1050, new_n4394);
nand_5 g04009(new_n4394, new_n1045, new_n4395);
nand_5 g04010(new_n4395, new_n1040, new_n4396);
nand_5 g04011(new_n4396, new_n1036, new_n4397);
nand_5 g04012(new_n4397, new_n1033, new_n4398);
nand_5 g04013(new_n4398, new_n1028, new_n4399);
nand_5 g04014(new_n4399, new_n1026, new_n4400);
nand_5 g04015(new_n4400, new_n1021, new_n4401);
nand_5 g04016(new_n4401, new_n1017, new_n4402);
nand_5 g04017(new_n4402, new_n1012, new_n4403);
nand_5 g04018(new_n4403, n650, new_n4404);
nor_5  g04019(new_n4404, new_n1006, n3090);
not_4  g04020(new_n579, new_n4406);
not_4  g04021(new_n572, new_n4407);
nand_5 g04022(new_n1651, new_n4407, new_n4408);
nand_5 g04023(new_n4408, new_n1649, new_n4409);
nand_5 g04024(new_n4409, new_n1646, new_n4410);
nand_5 g04025(new_n4410, new_n1643, new_n4411);
nand_5 g04026(new_n4411, new_n1641, new_n4412);
nand_5 g04027(new_n4412, new_n1638, new_n4413);
nand_5 g04028(new_n4413, new_n1635, new_n4414);
nand_5 g04029(new_n4414, new_n1632, new_n4415);
nand_5 g04030(new_n4415, new_n1628, new_n4416);
nand_5 g04031(new_n4416, new_n1625, new_n4417);
nand_5 g04032(new_n4417, new_n1621, new_n4418);
nand_5 g04033(new_n4418, new_n1618, new_n4419);
nand_5 g04034(new_n4419, new_n1778, new_n4420);
nand_5 g04035(new_n4420, new_n1782, new_n4421);
nand_5 g04036(new_n4421, new_n1614, new_n4422);
nand_5 g04037(new_n4422, new_n1611, new_n4423);
nand_5 g04038(new_n4423, new_n1789, new_n4424);
nand_5 g04039(new_n4424, new_n1608, new_n4425);
nand_5 g04040(new_n4425, new_n1605, new_n4426);
nand_5 g04041(new_n4426, new_n1795, new_n4427);
nand_5 g04042(new_n4427, new_n1799, new_n4428);
nand_5 g04043(new_n4428, new_n1602, new_n4429);
nand_5 g04044(new_n4429, new_n1599, new_n4430);
nand_5 g04045(new_n4430, new_n1596, new_n4431);
nand_5 g04046(new_n4431, new_n1593, new_n4432);
nand_5 g04047(new_n4432, new_n1806, new_n4433);
nand_5 g04048(new_n4433, new_n1589, new_n4434);
nand_5 g04049(new_n4434, new_n1586, new_n4435);
nand_5 g04050(new_n4435, new_n1583, new_n4436);
nand_5 g04051(new_n4436, new_n1580, new_n4437_1);
nand_5 g04052(new_n4437_1, new_n1576, new_n4438);
nand_5 g04053(new_n4438, new_n1573, new_n4439);
nand_5 g04054(new_n4439, new_n1570, new_n4440);
nand_5 g04055(new_n4440, new_n1567, new_n4441);
nand_5 g04056(new_n4441, new_n1564, new_n4442);
nand_5 g04057(new_n4442, new_n1561, new_n4443);
nand_5 g04058(new_n4443, new_n1338, new_n4444);
nand_5 g04059(new_n4444, new_n1331, new_n4445);
nand_5 g04060(new_n4445, new_n1326, new_n4446);
nand_5 g04061(new_n4446, new_n1321, new_n4447);
nand_5 g04062(new_n4447, new_n1318, new_n4448);
nand_5 g04063(new_n4448, new_n1315, new_n4449);
nand_5 g04064(new_n4449, new_n1312, new_n4450);
nand_5 g04065(new_n4450, new_n1309, new_n4451);
nand_5 g04066(new_n4451, new_n1307, new_n4452);
nand_5 g04067(new_n4452, new_n1304, new_n4453);
nand_5 g04068(new_n4453, new_n1300, new_n4454);
nand_5 g04069(new_n4454, new_n1297, new_n4455);
nand_5 g04070(new_n4455, new_n1294, new_n4456);
nand_5 g04071(new_n4456, new_n1355, new_n4457);
nand_5 g04072(new_n4457, new_n1291, new_n4458);
nand_5 g04073(new_n4458, new_n1288, new_n4459);
nand_5 g04074(new_n4459, new_n1283, new_n4460);
nand_5 g04075(new_n4460, new_n1363, new_n4461);
nand_5 g04076(new_n4461, new_n1280, new_n4462);
nand_5 g04077(new_n4462, new_n1370, new_n4463);
nand_5 g04078(new_n4463, new_n1373, new_n4464);
nand_5 g04079(new_n4464, new_n1277, new_n4465);
nand_5 g04080(new_n4465, new_n1272, new_n4466);
nand_5 g04081(new_n4466, new_n1269, new_n4467);
nand_5 g04082(new_n4467, new_n1380, new_n4468);
nand_5 g04083(new_n4468, new_n1264, new_n4469);
nand_5 g04084(new_n4469, new_n1259, new_n4470);
nand_5 g04085(new_n4470, new_n1388, new_n4471);
nand_5 g04086(new_n4471, new_n1392, new_n4472);
nand_5 g04087(new_n4472, new_n1256, new_n4473);
nand_5 g04088(new_n4473, new_n1252, new_n4474);
nand_5 g04089(new_n4474, new_n1249, new_n4475);
nand_5 g04090(new_n4475, new_n1244, new_n4476);
nand_5 g04091(new_n4476, new_n1240, new_n4477);
nand_5 g04092(new_n4477, new_n1234, new_n4478);
nand_5 g04093(new_n4478, new_n1231, new_n4479);
nand_5 g04094(new_n4479, new_n1227, new_n4480);
nand_5 g04095(new_n4480, new_n1407, new_n4481);
nand_5 g04096(new_n4481, new_n1223, new_n4482);
nand_5 g04097(new_n4482, new_n1218, new_n4483);
nand_5 g04098(new_n4483, new_n1213, new_n4484);
nand_5 g04099(new_n4484, new_n1210, new_n4485);
nand_5 g04100(new_n4485, new_n1206, new_n4486);
nand_5 g04101(new_n4486, new_n1418, new_n4487);
nand_5 g04102(new_n4487, new_n1422, new_n4488);
nand_5 g04103(new_n4488, new_n1428, new_n4489);
nand_5 g04104(new_n4489, new_n1203, new_n4490);
nand_5 g04105(new_n4490, new_n1433, new_n4491);
nand_5 g04106(new_n4491, n6147, new_n4492);
nor_5  g04107(new_n4492, new_n4406, n3242);
nand_5 g04108(new_n496, new_n415, new_n4494);
nand_5 g04109(new_n445, new_n435, new_n4495);
nand_5 g04110(new_n516, new_n390, new_n4496);
nor_5  g04111(new_n4496, new_n4495, new_n4497);
nand_5 g04112(new_n2064, new_n1707, new_n4498);
nor_5  g04113(new_n4498, new_n1697, new_n4499);
nand_5 g04114(new_n4499, new_n4497, new_n4500);
nor_5  g04115(new_n4500, new_n4494, new_n4501);
nor_5  g04116(new_n1645, new_n1311, new_n4502);
nand_5 g04117(new_n476, new_n471, new_n4503);
nand_5 g04118(new_n1656, new_n1278, new_n4504);
nor_5  g04119(new_n4504, new_n4503, new_n4505);
nand_5 g04120(new_n4505, new_n4502, new_n4506);
nor_5  g04121(new_n4506, new_n999, new_n4507);
nand_5 g04122(new_n4507, new_n4501, new_n4508);
nor_5  g04123(new_n1258, new_n1251, new_n4509);
nand_5 g04124(new_n2053, new_n1720, new_n4510);
nor_5  g04125(new_n4510, new_n1687, new_n4511);
nand_5 g04126(new_n4511, new_n4509, new_n4512);
nor_5  g04127(new_n462_1, new_n421, new_n4513);
nand_5 g04128(new_n506, new_n410, new_n4514);
nand_5 g04129(new_n511, new_n405, new_n4515);
nor_5  g04130(new_n4515, new_n4514, new_n4516);
nand_5 g04131(new_n4516, new_n4513, new_n4517);
nor_5  g04132(new_n4517, new_n4512, new_n4518);
nor_5  g04133(new_n1325, new_n1222_1, new_n4519);
nand_5 g04134(new_n934, new_n915, new_n4520);
nand_5 g04135(new_n1587, new_n1082, new_n4521);
nor_5  g04136(new_n4521, new_n4520, new_n4522);
nand_5 g04137(new_n4522, new_n4519, new_n4523);
nand_5 g04138(new_n1048, new_n541, new_n4524);
nor_5  g04139(new_n4524, new_n552, new_n4525);
nand_5 g04140(new_n2024, new_n1619, new_n4526);
nor_5  g04141(new_n4526, new_n1598, new_n4527);
nand_5 g04142(new_n4527, new_n4525, new_n4528);
nor_5  g04143(new_n4528, new_n4523, new_n4529);
nand_5 g04144(new_n4529, new_n4518, new_n4530);
nor_5  g04145(new_n4530, new_n4508, new_n4531);
nor_5  g04146(new_n1061, new_n965, new_n4532);
nand_5 g04147(new_n4532, new_n1015, new_n4533);
nor_5  g04148(new_n1634, new_n1299, new_n4534);
nand_5 g04149(new_n486, new_n466, new_n4535);
nand_5 g04150(new_n1670, new_n1289, new_n4536);
nor_5  g04151(new_n4536, new_n4535, new_n4537);
nand_5 g04152(new_n4537, new_n4534, new_n4538);
nand_5 g04153(new_n946, new_n566, new_n4539);
nand_5 g04154(new_n1574, new_n1201, new_n4540);
nor_5  g04155(new_n4540, new_n4539, new_n4541_1);
nand_5 g04156(new_n1270, new_n1232, new_n4542);
nand_5 g04157(new_n1562, new_n1204, new_n4543);
nor_5  g04158(new_n4543, new_n4542, new_n4544);
nand_5 g04159(new_n4544, new_n4541_1, new_n4545);
nor_5  g04160(new_n4545, new_n4538, new_n4546);
nand_5 g04161(new_n1068, new_n979, new_n4547);
nand_5 g04162(new_n1031, new_n531, new_n4548);
nor_5  g04163(new_n4548, new_n562, new_n4549);
nand_5 g04164(new_n2037, new_n1612, new_n4550);
nor_5  g04165(new_n4550, new_n1604, new_n4551);
nand_5 g04166(new_n4551, new_n4549, new_n4552);
nor_5  g04167(new_n4552, new_n4547, new_n4553);
nand_5 g04168(new_n4553, new_n4546, new_n4554);
nor_5  g04169(new_n4554, new_n4533, new_n4555);
nand_5 g04170(new_n4555, new_n4531, n3340);
not_4  g04171(n6460, new_n4557);
nand_5 g04172(new_n2020, new_n4557, new_n4558);
nand_5 g04173(new_n4558, new_n435, new_n4559);
nand_5 g04174(new_n4559, new_n819, new_n4560);
nand_5 g04175(new_n4560, new_n432, new_n4561);
nand_5 g04176(new_n4561, new_n427_1, new_n4562);
nand_5 g04177(new_n4562, new_n422, new_n4563);
nand_5 g04178(new_n4563, new_n828, new_n4564);
nand_5 g04179(new_n4564, new_n834, new_n4565);
nand_5 g04180(new_n4565, new_n840, new_n4566);
nand_5 g04181(new_n4566, new_n417, new_n4567);
nand_5 g04182(new_n4567, new_n847, new_n4568);
nand_5 g04183(new_n4568, new_n853, new_n4569);
nand_5 g04184(new_n4569, new_n859, new_n4570);
nand_5 g04185(new_n4570, new_n412, new_n4571);
nand_5 g04186(new_n4571, new_n866, new_n4572);
nand_5 g04187(new_n4572, new_n872, new_n4573);
nand_5 g04188(new_n4573, new_n878, new_n4574);
nand_5 g04189(new_n4574, new_n407, new_n4575);
nand_5 g04190(new_n4575, new_n885, new_n4576);
nand_5 g04191(new_n4576, new_n402, new_n4577);
nand_5 g04192(new_n4577, new_n397, new_n4578);
nand_5 g04193(new_n4578, new_n392, new_n4579);
nand_5 g04194(new_n4579, new_n894, new_n4580);
nand_5 g04195(new_n4580, new_n1087, new_n4581);
nand_5 g04196(new_n4581, new_n1129, new_n4582);
nand_5 g04197(new_n4582, new_n1084, new_n4583);
nand_5 g04198(new_n4583, new_n1134, new_n4584);
nand_5 g04199(new_n4584, new_n1080, new_n4585);
nand_5 g04200(new_n4585, new_n1075, new_n4586);
nand_5 g04201(new_n4586, new_n1070, new_n4587);
nand_5 g04202(new_n4587, new_n1143, new_n4588);
nand_5 g04203(new_n4588, new_n1148, new_n4589);
nand_5 g04204(new_n4589, new_n1065, new_n4590);
nand_5 g04205(new_n4590, new_n1062, new_n4591);
nand_5 g04206(new_n4591, new_n1156, new_n4592);
nand_5 g04207(new_n4592, new_n1057, new_n4593);
nand_5 g04208(new_n4593, new_n1053, new_n4594);
nand_5 g04209(new_n4594, new_n1050, new_n4595);
nand_5 g04210(new_n4595, new_n1045, new_n4596);
nand_5 g04211(new_n4596, new_n1040, new_n4597);
nand_5 g04212(new_n4597, new_n1036, new_n4598);
nand_5 g04213(new_n4598, new_n1033, new_n4599);
nand_5 g04214(new_n4599, new_n1028, new_n4600);
nand_5 g04215(new_n4600, new_n1026, new_n4601);
nand_5 g04216(new_n4601, new_n1021, new_n4602);
nand_5 g04217(new_n4602, new_n1017, new_n4603);
nand_5 g04218(new_n4603, new_n1012, new_n4604_1);
nand_5 g04219(new_n4604_1, new_n1009, new_n4605);
nand_5 g04220(new_n4605, new_n1004, new_n4606);
nand_5 g04221(new_n4606, new_n1000, new_n4607);
nand_5 g04222(new_n4607, new_n995, new_n4608);
nand_5 g04223(new_n4608, new_n990, new_n4609);
nand_5 g04224(new_n4609, new_n985, new_n4610);
nand_5 g04225(new_n4610, new_n981, new_n4611);
nand_5 g04226(new_n4611, new_n1179, new_n4612);
nand_5 g04227(new_n4612, new_n976, new_n4613);
nand_5 g04228(new_n4613, new_n971, new_n4614);
nand_5 g04229(new_n4614, new_n966, new_n4615_1);
nand_5 g04230(new_n4615_1, new_n961, new_n4616);
nand_5 g04231(new_n4616, new_n957, new_n4617);
nand_5 g04232(new_n4617, new_n952, new_n4618);
nand_5 g04233(new_n4618, new_n948_1, new_n4619);
nand_5 g04234(new_n4619, new_n943, new_n4620);
nand_5 g04235(new_n4620, new_n941, new_n4621);
nand_5 g04236(new_n4621, new_n938, new_n4622);
nand_5 g04237(new_n4622, new_n936, new_n4623);
nand_5 g04238(new_n4623, new_n931, new_n4624);
nand_5 g04239(new_n4624, new_n927, new_n4625);
nand_5 g04240(new_n4625, new_n922, new_n4626);
nand_5 g04241(new_n4626, new_n917, new_n4627);
nand_5 g04242(new_n4627, new_n912, new_n4628);
nand_5 g04243(new_n4628, new_n907, new_n4629);
nand_5 g04244(new_n4629, new_n903, new_n4630);
nand_5 g04245(new_n4630, new_n2066, new_n4631);
nand_5 g04246(new_n4631, new_n2063, new_n4632);
nand_5 g04247(new_n4632, new_n2062, new_n4633);
nand_5 g04248(new_n4633, new_n2058, new_n4634);
nand_5 g04249(new_n4634, new_n2055, new_n4635);
nand_5 g04250(new_n4635, new_n2051, new_n4636);
nand_5 g04251(new_n4636, new_n2046, new_n4637);
nand_5 g04252(new_n4637, new_n2042, new_n4638);
nand_5 g04253(new_n4638, new_n2039, new_n4639);
nand_5 g04254(new_n4639, new_n2036, new_n4640);
nand_5 g04255(new_n4640, new_n2033, new_n4641);
nand_5 g04256(new_n4641, new_n2029, new_n4642);
nand_5 g04257(new_n4642, n3130, new_n4643);
nor_5  g04258(new_n4643, new_n2023, n3603);
nand_5 g04259(new_n1027_1, new_n531, new_n4645);
nand_5 g04260(new_n4645, new_n650_1, new_n4646);
nand_5 g04261(new_n4646, new_n528, new_n4647);
nand_5 g04262(new_n4647, new_n523, new_n4648);
nand_5 g04263(new_n4648, new_n518, new_n4649);
nand_5 g04264(new_n4649, new_n659, new_n4650);
nand_5 g04265(new_n4650, new_n665, new_n4651);
nand_5 g04266(new_n4651, new_n672, new_n4652);
nand_5 g04267(new_n4652, new_n513, new_n4653);
nand_5 g04268(new_n4653, new_n679, new_n4654);
nand_5 g04269(new_n4654, new_n685, new_n4655);
nand_5 g04270(new_n4655, new_n691, new_n4656);
nand_5 g04271(new_n4656, new_n508, new_n4657);
nand_5 g04272(new_n4657, new_n698, new_n4658);
nand_5 g04273(new_n4658, new_n503, new_n4659_1);
nand_5 g04274(new_n4659_1, new_n704, new_n4660);
nand_5 g04275(new_n4660, new_n498_1, new_n4661);
nand_5 g04276(new_n4661, new_n711, new_n4662);
nand_5 g04277(new_n4662, new_n493, new_n4663);
nand_5 g04278(new_n4663, new_n718, new_n4664);
nand_5 g04279(new_n4664, new_n488, new_n4665);
nand_5 g04280(new_n4665, new_n725, new_n4666);
nand_5 g04281(new_n4666, new_n483, new_n4667);
nand_5 g04282(new_n4667, new_n732, new_n4668);
nand_5 g04283(new_n4668, new_n478, new_n4669);
nand_5 g04284(new_n4669, new_n739, new_n4670);
nand_5 g04285(new_n4670, new_n745, new_n4671);
nand_5 g04286(new_n4671, new_n751, new_n4672_1);
nand_5 g04287(new_n4672_1, new_n473, new_n4673);
nand_5 g04288(new_n4673, new_n758, new_n4674);
nand_5 g04289(new_n4674, new_n764, new_n4675);
nand_5 g04290(new_n4675, new_n770, new_n4676);
nand_5 g04291(new_n4676, new_n468, new_n4677);
nand_5 g04292(new_n4677, new_n777, new_n4678);
nand_5 g04293(new_n4678, new_n783, new_n4679);
nand_5 g04294(new_n4679, new_n789, new_n4680);
nand_5 g04295(new_n4680, new_n463, new_n4681);
nand_5 g04296(new_n4681, new_n796, new_n4682);
nand_5 g04297(new_n4682, new_n458, new_n4683);
nand_5 g04298(new_n4683, new_n453, new_n4684);
nand_5 g04299(new_n4684, new_n447, new_n4685);
nand_5 g04300(new_n4685, new_n805, new_n4686);
nand_5 g04301(new_n4686, new_n811, new_n4687);
nand_5 g04302(new_n4687, new_n442, new_n4688);
nand_5 g04303(new_n4688, new_n437, new_n4689);
nand_5 g04304(new_n4689, new_n819, new_n4690);
nand_5 g04305(new_n4690, new_n432, new_n4691);
nand_5 g04306(new_n4691, new_n427_1, new_n4692);
nand_5 g04307(new_n4692, new_n422, new_n4693);
nand_5 g04308(new_n4693, new_n828, new_n4694);
nand_5 g04309(new_n4694, new_n834, new_n4695);
nand_5 g04310(new_n4695, new_n840, new_n4696);
nand_5 g04311(new_n4696, new_n417, new_n4697);
nand_5 g04312(new_n4697, new_n847, new_n4698);
nand_5 g04313(new_n4698, new_n853, new_n4699);
nand_5 g04314(new_n4699, new_n859, new_n4700);
nand_5 g04315(new_n4700, new_n412, new_n4701);
nand_5 g04316(new_n4701, new_n866, new_n4702);
nand_5 g04317(new_n4702, new_n872, new_n4703);
nand_5 g04318(new_n4703, new_n878, new_n4704);
nand_5 g04319(new_n4704, new_n407, new_n4705);
nand_5 g04320(new_n4705, new_n885, new_n4706);
nand_5 g04321(new_n4706, new_n402, new_n4707);
nand_5 g04322(new_n4707, new_n397, new_n4708);
nand_5 g04323(new_n4708, new_n392, new_n4709);
nand_5 g04324(new_n4709, new_n894, new_n4710);
nand_5 g04325(new_n4710, new_n1087, new_n4711);
nand_5 g04326(new_n4711, new_n1129, new_n4712);
nand_5 g04327(new_n4712, new_n1084, new_n4713);
nand_5 g04328(new_n4713, new_n1134, new_n4714);
nand_5 g04329(new_n4714, new_n1080, new_n4715);
nand_5 g04330(new_n4715, new_n1075, new_n4716);
nand_5 g04331(new_n4716, new_n1070, new_n4717);
nand_5 g04332(new_n4717, new_n1143, new_n4718);
nand_5 g04333(new_n4718, new_n1148, new_n4719);
nand_5 g04334(new_n4719, new_n1065, new_n4720);
nand_5 g04335(new_n4720, new_n1062, new_n4721);
nand_5 g04336(new_n4721, new_n1156, new_n4722);
nand_5 g04337(new_n4722, new_n1057, new_n4723);
nand_5 g04338(new_n4723, new_n1053, new_n4724);
nand_5 g04339(new_n4724, new_n1050, new_n4725);
nand_5 g04340(new_n4725, new_n1045, new_n4726);
nand_5 g04341(new_n4726, new_n1040, new_n4727);
nand_5 g04342(new_n4727, new_n1036, new_n4728);
nand_5 g04343(new_n4728, n3799, new_n4729);
nor_5  g04344(new_n4729, new_n1030, n3854);
nand_5 g04345(new_n1316, new_n731, new_n4731);
nand_5 g04346(new_n4731, new_n1315, new_n4732);
nand_5 g04347(new_n4732, new_n1312, new_n4733);
nand_5 g04348(new_n4733, new_n1309, new_n4734);
nand_5 g04349(new_n4734, new_n1307, new_n4735);
nand_5 g04350(new_n4735, new_n1304, new_n4736);
nand_5 g04351(new_n4736, new_n1300, new_n4737);
nand_5 g04352(new_n4737, new_n1297, new_n4738);
nand_5 g04353(new_n4738, new_n1294, new_n4739);
nand_5 g04354(new_n4739, new_n1355, new_n4740);
nand_5 g04355(new_n4740, new_n1291, new_n4741);
nand_5 g04356(new_n4741, new_n1288, new_n4742);
nand_5 g04357(new_n4742, new_n1283, new_n4743);
nand_5 g04358(new_n4743, new_n1363, new_n4744);
nand_5 g04359(new_n4744, new_n1280, new_n4745);
nand_5 g04360(new_n4745, new_n1370, new_n4746);
nand_5 g04361(new_n4746, new_n1373, new_n4747);
nand_5 g04362(new_n4747, new_n1277, new_n4748);
nand_5 g04363(new_n4748, new_n1272, new_n4749);
nand_5 g04364(new_n4749, new_n1269, new_n4750);
nand_5 g04365(new_n4750, new_n1380, new_n4751);
nand_5 g04366(new_n4751, new_n1264, new_n4752);
nand_5 g04367(new_n4752, new_n1259, new_n4753);
nand_5 g04368(new_n4753, new_n1388, new_n4754);
nand_5 g04369(new_n4754, new_n1392, new_n4755_1);
nand_5 g04370(new_n4755_1, new_n1256, new_n4756);
nand_5 g04371(new_n4756, new_n1252, new_n4757);
nand_5 g04372(new_n4757, new_n1249, new_n4758);
nand_5 g04373(new_n4758, new_n1244, new_n4759);
nand_5 g04374(new_n4759, new_n1240, new_n4760);
nand_5 g04375(new_n4760, new_n1234, new_n4761);
nand_5 g04376(new_n4761, new_n1231, new_n4762);
nand_5 g04377(new_n4762, new_n1227, new_n4763);
nand_5 g04378(new_n4763, new_n1407, new_n4764);
nand_5 g04379(new_n4764, new_n1223, new_n4765);
nand_5 g04380(new_n4765, new_n1218, new_n4766);
nand_5 g04381(new_n4766, new_n1213, new_n4767);
nand_5 g04382(new_n4767, new_n1210, new_n4768);
nand_5 g04383(new_n4768, new_n1206, new_n4769);
nand_5 g04384(new_n4769, new_n1418, new_n4770);
nand_5 g04385(new_n4770, new_n1422, new_n4771);
nand_5 g04386(new_n4771, new_n1428, new_n4772);
nand_5 g04387(new_n4772, new_n1203, new_n4773);
nand_5 g04388(new_n4773, new_n1433, new_n4774_1);
nand_5 g04389(new_n4774_1, new_n581, new_n4775);
nand_5 g04390(new_n4775, new_n574, new_n4776);
nand_5 g04391(new_n4776, new_n568, new_n4777);
nand_5 g04392(new_n4777, new_n589, new_n4778);
nand_5 g04393(new_n4778, new_n595, new_n4779);
nand_5 g04394(new_n4779, new_n601, new_n4780);
nand_5 g04395(new_n4780, new_n563, new_n4781);
nand_5 g04396(new_n4781, new_n608, new_n4782);
nand_5 g04397(new_n4782, new_n558, new_n4783);
nand_5 g04398(new_n4783, new_n615, new_n4784);
nand_5 g04399(new_n4784, new_n553, new_n4785_1);
nand_5 g04400(new_n4785_1, new_n622, new_n4786);
nand_5 g04401(new_n4786, new_n628, new_n4787);
nand_5 g04402(new_n4787, new_n548, new_n4788);
nand_5 g04403(new_n4788, new_n543_1, new_n4789);
nand_5 g04404(new_n4789, new_n636, new_n4790);
nand_5 g04405(new_n4790, new_n642, new_n4791);
nand_5 g04406(new_n4791, new_n538, new_n4792);
nand_5 g04407(new_n4792, new_n533, new_n4793);
nand_5 g04408(new_n4793, new_n650_1, new_n4794);
nand_5 g04409(new_n4794, new_n528, new_n4795);
nand_5 g04410(new_n4795, new_n523, new_n4796);
nand_5 g04411(new_n4796, new_n518, new_n4797);
nand_5 g04412(new_n4797, new_n659, new_n4798);
nand_5 g04413(new_n4798, new_n665, new_n4799);
nand_5 g04414(new_n4799, new_n672, new_n4800);
nand_5 g04415(new_n4800, new_n513, new_n4801);
nand_5 g04416(new_n4801, new_n679, new_n4802);
nand_5 g04417(new_n4802, new_n685, new_n4803);
nand_5 g04418(new_n4803, new_n691, new_n4804);
nand_5 g04419(new_n4804, new_n508, new_n4805);
nand_5 g04420(new_n4805, new_n698, new_n4806);
nand_5 g04421(new_n4806, new_n503, new_n4807);
nand_5 g04422(new_n4807, new_n704, new_n4808);
nand_5 g04423(new_n4808, new_n498_1, new_n4809);
nand_5 g04424(new_n4809, new_n711, new_n4810);
nand_5 g04425(new_n4810, new_n493, new_n4811);
nand_5 g04426(new_n4811, new_n718, new_n4812);
nand_5 g04427(new_n4812, new_n488, new_n4813);
nand_5 g04428(new_n4813, new_n725, new_n4814);
nand_5 g04429(new_n4814, n12573, new_n4815);
nor_5  g04430(new_n4815, new_n480, n3901);
nor_5  g04431(n12218, n9893, new_n4817);
not_4  g04432(new_n4817, new_n4818);
nand_5 g04433(new_n4818, new_n2062, new_n4819);
nand_5 g04434(new_n4819, new_n2058, new_n4820);
nand_5 g04435(new_n4820, new_n2055, new_n4821);
nand_5 g04436(new_n4821, new_n2051, new_n4822);
nand_5 g04437(new_n4822, new_n2046, new_n4823);
nand_5 g04438(new_n4823, new_n2042, new_n4824);
nand_5 g04439(new_n4824, new_n2039, new_n4825);
nand_5 g04440(new_n4825, new_n2036, new_n4826);
nand_5 g04441(new_n4826, new_n2033, new_n4827);
nand_5 g04442(new_n4827, new_n2029, new_n4828);
nand_5 g04443(new_n4828, new_n2026, new_n4829);
nand_5 g04444(new_n4829, new_n2022, new_n4830);
nand_5 g04445(new_n4830, new_n2018, new_n4831);
nand_5 g04446(new_n4831, new_n1726, new_n4832);
nand_5 g04447(new_n4832, new_n1722, new_n4833);
nand_5 g04448(new_n4833, new_n1718, new_n4834);
nand_5 g04449(new_n4834, new_n1713, new_n4835);
nand_5 g04450(new_n4835, new_n1737, new_n4836);
nand_5 g04451(new_n4836, new_n1709, new_n4837);
nand_5 g04452(new_n4837, new_n1742, new_n4838);
nand_5 g04453(new_n4838, new_n1704, new_n4839);
nand_5 g04454(new_n4839, new_n1702_1, new_n4840);
nand_5 g04455(new_n4840, new_n1698, new_n4841);
nand_5 g04456(new_n4841, new_n1695, new_n4842);
nand_5 g04457(new_n4842, new_n1692, new_n4843);
nand_5 g04458(new_n4843, new_n1752, new_n4844);
nand_5 g04459(new_n4844, new_n1688, new_n4845);
nand_5 g04460(new_n4845, new_n1685, new_n4846);
nand_5 g04461(new_n4846, new_n1680, new_n4847);
nand_5 g04462(new_n4847, new_n1676, new_n4848);
nand_5 g04463(new_n4848, new_n1672, new_n4849);
nand_5 g04464(new_n4849, new_n1669, new_n4850);
nand_5 g04465(new_n4850, new_n1666, new_n4851);
nand_5 g04466(new_n4851, new_n1663, new_n4852);
nand_5 g04467(new_n4852, new_n1658, new_n4853);
nand_5 g04468(new_n4853, new_n1653, new_n4854);
nand_5 g04469(new_n4854, new_n1651, new_n4855);
nand_5 g04470(new_n4855, new_n1649, new_n4856);
nand_5 g04471(new_n4856, new_n1646, new_n4857);
nand_5 g04472(new_n4857, new_n1643, new_n4858_1);
nand_5 g04473(new_n4858_1, new_n1641, new_n4859);
nand_5 g04474(new_n4859, new_n1638, new_n4860);
nand_5 g04475(new_n4860, new_n1635, new_n4861);
nand_5 g04476(new_n4861, new_n1632, new_n4862);
nand_5 g04477(new_n4862, new_n1628, new_n4863);
nand_5 g04478(new_n4863, new_n1625, new_n4864);
nand_5 g04479(new_n4864, new_n1621, new_n4865);
nand_5 g04480(new_n4865, new_n1618, new_n4866);
nand_5 g04481(new_n4866, new_n1778, new_n4867);
nand_5 g04482(new_n4867, new_n1782, new_n4868);
nand_5 g04483(new_n4868, new_n1614, new_n4869);
nand_5 g04484(new_n4869, new_n1611, new_n4870);
nand_5 g04485(new_n4870, new_n1789, new_n4871);
nand_5 g04486(new_n4871, new_n1608, new_n4872);
nand_5 g04487(new_n4872, new_n1605, new_n4873);
nand_5 g04488(new_n4873, new_n1795, new_n4874);
nand_5 g04489(new_n4874, new_n1799, new_n4875);
nand_5 g04490(new_n4875, new_n1602, new_n4876);
nand_5 g04491(new_n4876, new_n1599, new_n4877);
nand_5 g04492(new_n4877, new_n1596, new_n4878);
nand_5 g04493(new_n4878, new_n1593, new_n4879);
nand_5 g04494(new_n4879, new_n1806, new_n4880);
nand_5 g04495(new_n4880, new_n1589, new_n4881);
nand_5 g04496(new_n4881, new_n1586, new_n4882);
nand_5 g04497(new_n4882, new_n1583, new_n4883);
nand_5 g04498(new_n4883, new_n1580, new_n4884);
nand_5 g04499(new_n4884, new_n1576, new_n4885);
nand_5 g04500(new_n4885, new_n1573, new_n4886);
nand_5 g04501(new_n4886, new_n1570, new_n4887);
nand_5 g04502(new_n4887, new_n1567, new_n4888);
nand_5 g04503(new_n4888, new_n1564, new_n4889);
nand_5 g04504(new_n4889, new_n1561, new_n4890);
nand_5 g04505(new_n4890, new_n1338, new_n4891);
nand_5 g04506(new_n4891, new_n1331, new_n4892);
nand_5 g04507(new_n4892, new_n1326, new_n4893);
nand_5 g04508(new_n4893, new_n1321, new_n4894);
nand_5 g04509(new_n4894, new_n1318, new_n4895_1);
nand_5 g04510(new_n4895_1, new_n1315, new_n4896);
nand_5 g04511(new_n4896, new_n1312, new_n4897);
nand_5 g04512(new_n4897, new_n1309, new_n4898);
nand_5 g04513(new_n4898, new_n1307, new_n4899);
nand_5 g04514(new_n4899, new_n1304, new_n4900);
nand_5 g04515(new_n4900, new_n1300, new_n4901);
nand_5 g04516(new_n4901, new_n1297, new_n4902);
nand_5 g04517(new_n4902, n427, new_n4903);
nor_5  g04518(new_n4903, new_n767, n4125);
not_4  g04519(new_n737_1, new_n4905);
nand_5 g04520(new_n1312, new_n4905, new_n4906);
nand_5 g04521(new_n4906, new_n1309, new_n4907_1);
nand_5 g04522(new_n4907_1, new_n1307, new_n4908);
nand_5 g04523(new_n4908, new_n1304, new_n4909);
nand_5 g04524(new_n4909, new_n1300, new_n4910);
nand_5 g04525(new_n4910, new_n1297, new_n4911);
nand_5 g04526(new_n4911, new_n1294, new_n4912);
nand_5 g04527(new_n4912, new_n1355, new_n4913);
nand_5 g04528(new_n4913, new_n1291, new_n4914);
nand_5 g04529(new_n4914, new_n1288, new_n4915);
nand_5 g04530(new_n4915, new_n1283, new_n4916);
nand_5 g04531(new_n4916, new_n1363, new_n4917);
nand_5 g04532(new_n4917, new_n1280, new_n4918);
nand_5 g04533(new_n4918, new_n1370, new_n4919);
nand_5 g04534(new_n4919, new_n1373, new_n4920);
nand_5 g04535(new_n4920, new_n1277, new_n4921);
nand_5 g04536(new_n4921, new_n1272, new_n4922);
nand_5 g04537(new_n4922, new_n1269, new_n4923);
nand_5 g04538(new_n4923, new_n1380, new_n4924);
nand_5 g04539(new_n4924, new_n1264, new_n4925);
nand_5 g04540(new_n4925, new_n1259, new_n4926);
nand_5 g04541(new_n4926, new_n1388, new_n4927);
nand_5 g04542(new_n4927, new_n1392, new_n4928);
nand_5 g04543(new_n4928, new_n1256, new_n4929);
nand_5 g04544(new_n4929, new_n1252, new_n4930);
nand_5 g04545(new_n4930, new_n1249, new_n4931);
nand_5 g04546(new_n4931, new_n1244, new_n4932);
nand_5 g04547(new_n4932, new_n1240, new_n4933);
nand_5 g04548(new_n4933, new_n1234, new_n4934);
nand_5 g04549(new_n4934, new_n1231, new_n4935);
nand_5 g04550(new_n4935, new_n1227, new_n4936);
nand_5 g04551(new_n4936, new_n1407, new_n4937);
nand_5 g04552(new_n4937, new_n1223, new_n4938);
nand_5 g04553(new_n4938, new_n1218, new_n4939);
nand_5 g04554(new_n4939, new_n1213, new_n4940);
nand_5 g04555(new_n4940, new_n1210, new_n4941);
nand_5 g04556(new_n4941, new_n1206, new_n4942);
nand_5 g04557(new_n4942, new_n1418, new_n4943);
nand_5 g04558(new_n4943, new_n1422, new_n4944);
nand_5 g04559(new_n4944, new_n1428, new_n4945);
nand_5 g04560(new_n4945, new_n1203, new_n4946);
nand_5 g04561(new_n4946, new_n1433, new_n4947);
nand_5 g04562(new_n4947, new_n581, new_n4948);
nand_5 g04563(new_n4948, new_n574, new_n4949);
nand_5 g04564(new_n4949, new_n568, new_n4950);
nand_5 g04565(new_n4950, new_n589, new_n4951);
nand_5 g04566(new_n4951, new_n595, new_n4952);
nand_5 g04567(new_n4952, new_n601, new_n4953);
nand_5 g04568(new_n4953, new_n563, new_n4954);
nand_5 g04569(new_n4954, new_n608, new_n4955);
nand_5 g04570(new_n4955, new_n558, new_n4956);
nand_5 g04571(new_n4956, new_n615, new_n4957);
nand_5 g04572(new_n4957, new_n553, new_n4958);
nand_5 g04573(new_n4958, new_n622, new_n4959);
nand_5 g04574(new_n4959, new_n628, new_n4960);
nand_5 g04575(new_n4960, new_n548, new_n4961);
nand_5 g04576(new_n4961, new_n543_1, new_n4962);
nand_5 g04577(new_n4962, new_n636, new_n4963);
nand_5 g04578(new_n4963, new_n642, new_n4964);
nand_5 g04579(new_n4964, new_n538, new_n4965);
nand_5 g04580(new_n4965, new_n533, new_n4966);
nand_5 g04581(new_n4966, new_n650_1, new_n4967);
nand_5 g04582(new_n4967, new_n528, new_n4968);
nand_5 g04583(new_n4968, new_n523, new_n4969);
nand_5 g04584(new_n4969, new_n518, new_n4970);
nand_5 g04585(new_n4970, new_n659, new_n4971_1);
nand_5 g04586(new_n4971_1, new_n665, new_n4972);
nand_5 g04587(new_n4972, new_n672, new_n4973);
nand_5 g04588(new_n4973, new_n513, new_n4974);
nand_5 g04589(new_n4974, new_n679, new_n4975);
nand_5 g04590(new_n4975, new_n685, new_n4976);
nand_5 g04591(new_n4976, new_n691, new_n4977);
nand_5 g04592(new_n4977, new_n508, new_n4978);
nand_5 g04593(new_n4978, new_n698, new_n4979);
nand_5 g04594(new_n4979, new_n503, new_n4980);
nand_5 g04595(new_n4980, new_n704, new_n4981);
nand_5 g04596(new_n4981, new_n498_1, new_n4982);
nand_5 g04597(new_n4982, new_n711, new_n4983);
nand_5 g04598(new_n4983, new_n493, new_n4984);
nand_5 g04599(new_n4984, new_n718, new_n4985);
nand_5 g04600(new_n4985, new_n488, new_n4986);
nand_5 g04601(new_n4986, new_n725, new_n4987);
nand_5 g04602(new_n4987, new_n483, new_n4988);
nand_5 g04603(new_n4988, new_n732, new_n4989);
nand_5 g04604(new_n4989, n10736, new_n4990);
nor_5  g04605(new_n4990, new_n475, n4279);
nand_5 g04606(new_n1581, new_n690, new_n4992);
nand_5 g04607(new_n4992, new_n1580, new_n4993);
nand_5 g04608(new_n4993, new_n1576, new_n4994);
nand_5 g04609(new_n4994, new_n1573, new_n4995);
nand_5 g04610(new_n4995, new_n1570, new_n4996);
nand_5 g04611(new_n4996, new_n1567, new_n4997);
nand_5 g04612(new_n4997, new_n1564, new_n4998);
nand_5 g04613(new_n4998, new_n1561, new_n4999);
nand_5 g04614(new_n4999, new_n1338, new_n5000);
nand_5 g04615(new_n5000, new_n1331, new_n5001);
nand_5 g04616(new_n5001, new_n1326, new_n5002);
nand_5 g04617(new_n5002, new_n1321, new_n5003);
nand_5 g04618(new_n5003, new_n1318, new_n5004);
nand_5 g04619(new_n5004, new_n1315, new_n5005);
nand_5 g04620(new_n5005, new_n1312, new_n5006);
nand_5 g04621(new_n5006, new_n1309, new_n5007);
nand_5 g04622(new_n5007, new_n1307, new_n5008);
nand_5 g04623(new_n5008, new_n1304, new_n5009_1);
nand_5 g04624(new_n5009_1, new_n1300, new_n5010);
nand_5 g04625(new_n5010, new_n1297, new_n5011);
nand_5 g04626(new_n5011, new_n1294, new_n5012);
nand_5 g04627(new_n5012, new_n1355, new_n5013);
nand_5 g04628(new_n5013, new_n1291, new_n5014_1);
nand_5 g04629(new_n5014_1, new_n1288, new_n5015);
nand_5 g04630(new_n5015, new_n1283, new_n5016);
nand_5 g04631(new_n5016, new_n1363, new_n5017);
nand_5 g04632(new_n5017, new_n1280, new_n5018);
nand_5 g04633(new_n5018, new_n1370, new_n5019);
nand_5 g04634(new_n5019, new_n1373, new_n5020);
nand_5 g04635(new_n5020, new_n1277, new_n5021);
nand_5 g04636(new_n5021, new_n1272, new_n5022);
nand_5 g04637(new_n5022, new_n1269, new_n5023_1);
nand_5 g04638(new_n5023_1, new_n1380, new_n5024);
nand_5 g04639(new_n5024, new_n1264, new_n5025);
nand_5 g04640(new_n5025, new_n1259, new_n5026);
nand_5 g04641(new_n5026, new_n1388, new_n5027);
nand_5 g04642(new_n5027, new_n1392, new_n5028);
nand_5 g04643(new_n5028, new_n1256, new_n5029);
nand_5 g04644(new_n5029, new_n1252, new_n5030);
nand_5 g04645(new_n5030, new_n1249, new_n5031);
nand_5 g04646(new_n5031, new_n1244, new_n5032);
nand_5 g04647(new_n5032, new_n1240, new_n5033_1);
nand_5 g04648(new_n5033_1, new_n1234, new_n5034);
nand_5 g04649(new_n5034, new_n1231, new_n5035);
nand_5 g04650(new_n5035, new_n1227, new_n5036);
nand_5 g04651(new_n5036, new_n1407, new_n5037);
nand_5 g04652(new_n5037, new_n1223, new_n5038);
nand_5 g04653(new_n5038, new_n1218, new_n5039);
nand_5 g04654(new_n5039, new_n1213, new_n5040);
nand_5 g04655(new_n5040, new_n1210, new_n5041);
nand_5 g04656(new_n5041, new_n1206, new_n5042);
nand_5 g04657(new_n5042, new_n1418, new_n5043);
nand_5 g04658(new_n5043, new_n1422, new_n5044);
nand_5 g04659(new_n5044, new_n1428, new_n5045);
nand_5 g04660(new_n5045, new_n1203, new_n5046_1);
nand_5 g04661(new_n5046_1, new_n1433, new_n5047);
nand_5 g04662(new_n5047, new_n581, new_n5048);
nand_5 g04663(new_n5048, new_n574, new_n5049);
nand_5 g04664(new_n5049, new_n568, new_n5050);
nand_5 g04665(new_n5050, new_n589, new_n5051);
nand_5 g04666(new_n5051, new_n595, new_n5052);
nand_5 g04667(new_n5052, new_n601, new_n5053);
nand_5 g04668(new_n5053, new_n563, new_n5054);
nand_5 g04669(new_n5054, new_n608, new_n5055);
nand_5 g04670(new_n5055, new_n558, new_n5056);
nand_5 g04671(new_n5056, new_n615, new_n5057);
nand_5 g04672(new_n5057, new_n553, new_n5058);
nand_5 g04673(new_n5058, new_n622, new_n5059);
nand_5 g04674(new_n5059, new_n628, new_n5060);
nand_5 g04675(new_n5060, new_n548, new_n5061);
nand_5 g04676(new_n5061, new_n543_1, new_n5062);
nand_5 g04677(new_n5062, new_n636, new_n5063);
nand_5 g04678(new_n5063, new_n642, new_n5064);
nand_5 g04679(new_n5064, new_n538, new_n5065);
nand_5 g04680(new_n5065, new_n533, new_n5066);
nand_5 g04681(new_n5066, new_n650_1, new_n5067);
nand_5 g04682(new_n5067, new_n528, new_n5068);
nand_5 g04683(new_n5068, new_n523, new_n5069);
nand_5 g04684(new_n5069, new_n518, new_n5070);
nand_5 g04685(new_n5070, new_n659, new_n5071);
nand_5 g04686(new_n5071, new_n665, new_n5072);
nand_5 g04687(new_n5072, new_n672, new_n5073);
nand_5 g04688(new_n5073, new_n513, new_n5074);
nand_5 g04689(new_n5074, new_n679, new_n5075);
nand_5 g04690(new_n5075, n2454, new_n5076);
nor_5  g04691(new_n5076, new_n682_1, n4305);
nand_5 g04692(new_n1281, new_n788, new_n5078);
nand_5 g04693(new_n5078, new_n1363, new_n5079);
nand_5 g04694(new_n5079, new_n1280, new_n5080);
nand_5 g04695(new_n5080, new_n1370, new_n5081);
nand_5 g04696(new_n5081, new_n1373, new_n5082);
nand_5 g04697(new_n5082, new_n1277, new_n5083);
nand_5 g04698(new_n5083, new_n1272, new_n5084);
nand_5 g04699(new_n5084, new_n1269, new_n5085);
nand_5 g04700(new_n5085, new_n1380, new_n5086);
nand_5 g04701(new_n5086, new_n1264, new_n5087);
nand_5 g04702(new_n5087, new_n1259, new_n5088);
nand_5 g04703(new_n5088, new_n1388, new_n5089);
nand_5 g04704(new_n5089, new_n1392, new_n5090);
nand_5 g04705(new_n5090, new_n1256, new_n5091);
nand_5 g04706(new_n5091, new_n1252, new_n5092);
nand_5 g04707(new_n5092, new_n1249, new_n5093);
nand_5 g04708(new_n5093, new_n1244, new_n5094);
nand_5 g04709(new_n5094, new_n1240, new_n5095);
nand_5 g04710(new_n5095, new_n1234, new_n5096);
nand_5 g04711(new_n5096, new_n1231, new_n5097);
nand_5 g04712(new_n5097, new_n1227, new_n5098);
nand_5 g04713(new_n5098, new_n1407, new_n5099);
nand_5 g04714(new_n5099, new_n1223, new_n5100);
nand_5 g04715(new_n5100, new_n1218, new_n5101);
nand_5 g04716(new_n5101, new_n1213, new_n5102);
nand_5 g04717(new_n5102, new_n1210, new_n5103);
nand_5 g04718(new_n5103, new_n1206, new_n5104);
nand_5 g04719(new_n5104, new_n1418, new_n5105);
nand_5 g04720(new_n5105, new_n1422, new_n5106);
nand_5 g04721(new_n5106, new_n1428, new_n5107);
nand_5 g04722(new_n5107, new_n1203, new_n5108);
nand_5 g04723(new_n5108, new_n1433, new_n5109);
nand_5 g04724(new_n5109, new_n581, new_n5110);
nand_5 g04725(new_n5110, new_n574, new_n5111);
nand_5 g04726(new_n5111, new_n568, new_n5112);
nand_5 g04727(new_n5112, new_n589, new_n5113);
nand_5 g04728(new_n5113, new_n595, new_n5114);
nand_5 g04729(new_n5114, new_n601, new_n5115);
nand_5 g04730(new_n5115, new_n563, new_n5116);
nand_5 g04731(new_n5116, new_n608, new_n5117);
nand_5 g04732(new_n5117, new_n558, new_n5118);
nand_5 g04733(new_n5118, new_n615, new_n5119);
nand_5 g04734(new_n5119, new_n553, new_n5120);
nand_5 g04735(new_n5120, new_n622, new_n5121);
nand_5 g04736(new_n5121, new_n628, new_n5122);
nand_5 g04737(new_n5122, new_n548, new_n5123);
nand_5 g04738(new_n5123, new_n543_1, new_n5124);
nand_5 g04739(new_n5124, new_n636, new_n5125);
nand_5 g04740(new_n5125, new_n642, new_n5126);
nand_5 g04741(new_n5126, new_n538, new_n5127);
nand_5 g04742(new_n5127, new_n533, new_n5128);
nand_5 g04743(new_n5128, new_n650_1, new_n5129);
nand_5 g04744(new_n5129, new_n528, new_n5130);
nand_5 g04745(new_n5130, new_n523, new_n5131);
nand_5 g04746(new_n5131, new_n518, new_n5132);
nand_5 g04747(new_n5132, new_n659, new_n5133);
nand_5 g04748(new_n5133, new_n665, new_n5134);
nand_5 g04749(new_n5134, new_n672, new_n5135);
nand_5 g04750(new_n5135, new_n513, new_n5136);
nand_5 g04751(new_n5136, new_n679, new_n5137);
nand_5 g04752(new_n5137, new_n685, new_n5138);
nand_5 g04753(new_n5138, new_n691, new_n5139);
nand_5 g04754(new_n5139, new_n508, new_n5140);
nand_5 g04755(new_n5140, new_n698, new_n5141);
nand_5 g04756(new_n5141, new_n503, new_n5142);
nand_5 g04757(new_n5142, new_n704, new_n5143);
nand_5 g04758(new_n5143, new_n498_1, new_n5144);
nand_5 g04759(new_n5144, new_n711, new_n5145);
nand_5 g04760(new_n5145, new_n493, new_n5146);
nand_5 g04761(new_n5146, new_n718, new_n5147);
nand_5 g04762(new_n5147, new_n488, new_n5148);
nand_5 g04763(new_n5148, new_n725, new_n5149);
nand_5 g04764(new_n5149, new_n483, new_n5150);
nand_5 g04765(new_n5150, new_n732, new_n5151);
nand_5 g04766(new_n5151, new_n478, new_n5152);
nand_5 g04767(new_n5152, new_n739, new_n5153);
nand_5 g04768(new_n5153, new_n745, new_n5154);
nand_5 g04769(new_n5154, new_n751, new_n5155);
nand_5 g04770(new_n5155, new_n473, new_n5156);
nand_5 g04771(new_n5156, new_n758, new_n5157);
nand_5 g04772(new_n5157, new_n764, new_n5158);
nand_5 g04773(new_n5158, new_n770, new_n5159);
nand_5 g04774(new_n5159, new_n468, new_n5160);
nand_5 g04775(new_n5160, new_n777, new_n5161);
nand_5 g04776(new_n5161, n2615, new_n5162);
nor_5  g04777(new_n5162, new_n780, n4345);
not_4  g04778(new_n1177, new_n5164);
nand_5 g04779(new_n5164, new_n508, new_n5165);
nand_5 g04780(new_n5165, new_n698, new_n5166);
nand_5 g04781(new_n5166, new_n503, new_n5167);
nand_5 g04782(new_n5167, new_n704, new_n5168);
nand_5 g04783(new_n5168, new_n498_1, new_n5169);
nand_5 g04784(new_n5169, new_n711, new_n5170);
nand_5 g04785(new_n5170, new_n493, new_n5171);
nand_5 g04786(new_n5171, new_n718, new_n5172);
nand_5 g04787(new_n5172, new_n488, new_n5173);
nand_5 g04788(new_n5173, new_n725, new_n5174);
nand_5 g04789(new_n5174, new_n483, new_n5175);
nand_5 g04790(new_n5175, new_n732, new_n5176);
nand_5 g04791(new_n5176, new_n478, new_n5177);
nand_5 g04792(new_n5177, new_n739, new_n5178);
nand_5 g04793(new_n5178, new_n745, new_n5179);
nand_5 g04794(new_n5179, new_n751, new_n5180);
nand_5 g04795(new_n5180, new_n473, new_n5181);
nand_5 g04796(new_n5181, new_n758, new_n5182);
nand_5 g04797(new_n5182, new_n764, new_n5183);
nand_5 g04798(new_n5183, new_n770, new_n5184_1);
nand_5 g04799(new_n5184_1, new_n468, new_n5185_1);
nand_5 g04800(new_n5185_1, new_n777, new_n5186);
nand_5 g04801(new_n5186, new_n783, new_n5187);
nand_5 g04802(new_n5187, new_n789, new_n5188);
nand_5 g04803(new_n5188, new_n463, new_n5189);
nand_5 g04804(new_n5189, new_n796, new_n5190);
nand_5 g04805(new_n5190, new_n458, new_n5191);
nand_5 g04806(new_n5191, new_n453, new_n5192);
nand_5 g04807(new_n5192, new_n447, new_n5193);
nand_5 g04808(new_n5193, new_n805, new_n5194);
nand_5 g04809(new_n5194, new_n811, new_n5195);
nand_5 g04810(new_n5195, new_n442, new_n5196);
nand_5 g04811(new_n5196, new_n437, new_n5197);
nand_5 g04812(new_n5197, new_n819, new_n5198);
nand_5 g04813(new_n5198, new_n432, new_n5199);
nand_5 g04814(new_n5199, new_n427_1, new_n5200);
nand_5 g04815(new_n5200, new_n422, new_n5201);
nand_5 g04816(new_n5201, new_n828, new_n5202);
nand_5 g04817(new_n5202, new_n834, new_n5203);
nand_5 g04818(new_n5203, new_n840, new_n5204);
nand_5 g04819(new_n5204, new_n417, new_n5205);
nand_5 g04820(new_n5205, new_n847, new_n5206);
nand_5 g04821(new_n5206, new_n853, new_n5207);
nand_5 g04822(new_n5207, new_n859, new_n5208);
nand_5 g04823(new_n5208, new_n412, new_n5209);
nand_5 g04824(new_n5209, new_n866, new_n5210);
nand_5 g04825(new_n5210, new_n872, new_n5211);
nand_5 g04826(new_n5211, new_n878, new_n5212);
nand_5 g04827(new_n5212, new_n407, new_n5213);
nand_5 g04828(new_n5213, new_n885, new_n5214);
nand_5 g04829(new_n5214, new_n402, new_n5215);
nand_5 g04830(new_n5215, new_n397, new_n5216);
nand_5 g04831(new_n5216, new_n392, new_n5217);
nand_5 g04832(new_n5217, new_n894, new_n5218);
nand_5 g04833(new_n5218, new_n1087, new_n5219);
nand_5 g04834(new_n5219, new_n1129, new_n5220);
nand_5 g04835(new_n5220, new_n1084, new_n5221);
nand_5 g04836(new_n5221, new_n1134, new_n5222);
nand_5 g04837(new_n5222, new_n1080, new_n5223);
nand_5 g04838(new_n5223, new_n1075, new_n5224);
nand_5 g04839(new_n5224, new_n1070, new_n5225_1);
nand_5 g04840(new_n5225_1, new_n1143, new_n5226);
nand_5 g04841(new_n5226, new_n1148, new_n5227);
nand_5 g04842(new_n5227, new_n1065, new_n5228);
nand_5 g04843(new_n5228, new_n1062, new_n5229);
nand_5 g04844(new_n5229, new_n1156, new_n5230);
nand_5 g04845(new_n5230, new_n1057, new_n5231);
nand_5 g04846(new_n5231, new_n1053, new_n5232);
nand_5 g04847(new_n5232, new_n1050, new_n5233);
nand_5 g04848(new_n5233, new_n1045, new_n5234);
nand_5 g04849(new_n5234, new_n1040, new_n5235);
nand_5 g04850(new_n5235, new_n1036, new_n5236);
nand_5 g04851(new_n5236, new_n1033, new_n5237);
nand_5 g04852(new_n5237, new_n1028, new_n5238);
nand_5 g04853(new_n5238, new_n1026, new_n5239);
nand_5 g04854(new_n5239, new_n1021, new_n5240);
nand_5 g04855(new_n5240, new_n1017, new_n5241);
nand_5 g04856(new_n5241, new_n1012, new_n5242);
nand_5 g04857(new_n5242, new_n1009, new_n5243);
nand_5 g04858(new_n5243, new_n1004, new_n5244);
nand_5 g04859(new_n5244, new_n1000, new_n5245);
nand_5 g04860(new_n5245, new_n995, new_n5246);
nand_5 g04861(new_n5246, new_n990, new_n5247);
nand_5 g04862(new_n5247, new_n985, new_n5248);
nand_5 g04863(new_n5248, n8044, new_n5249);
nor_5  g04864(new_n5249, new_n978, n4437);
nor_5  g04865(n2895, n1568, new_n5251);
not_4  g04866(new_n5251, new_n5252);
nand_5 g04867(new_n5252, new_n503, new_n5253);
nand_5 g04868(new_n5253, new_n704, new_n5254);
nand_5 g04869(new_n5254, new_n498_1, new_n5255);
nand_5 g04870(new_n5255, new_n711, new_n5256);
nand_5 g04871(new_n5256, new_n493, new_n5257);
nand_5 g04872(new_n5257, new_n718, new_n5258);
nand_5 g04873(new_n5258, new_n488, new_n5259);
nand_5 g04874(new_n5259, new_n725, new_n5260);
nand_5 g04875(new_n5260, new_n483, new_n5261);
nand_5 g04876(new_n5261, new_n732, new_n5262);
nand_5 g04877(new_n5262, new_n478, new_n5263);
nand_5 g04878(new_n5263, new_n739, new_n5264);
nand_5 g04879(new_n5264, new_n745, new_n5265);
nand_5 g04880(new_n5265, new_n751, new_n5266);
nand_5 g04881(new_n5266, new_n473, new_n5267);
nand_5 g04882(new_n5267, new_n758, new_n5268);
nand_5 g04883(new_n5268, new_n764, new_n5269);
nand_5 g04884(new_n5269, new_n770, new_n5270);
nand_5 g04885(new_n5270, new_n468, new_n5271);
nand_5 g04886(new_n5271, new_n777, new_n5272);
nand_5 g04887(new_n5272, new_n783, new_n5273);
nand_5 g04888(new_n5273, new_n789, new_n5274);
nand_5 g04889(new_n5274, new_n463, new_n5275);
nand_5 g04890(new_n5275, new_n796, new_n5276);
nand_5 g04891(new_n5276, new_n458, new_n5277);
nand_5 g04892(new_n5277, new_n453, new_n5278);
nand_5 g04893(new_n5278, new_n447, new_n5279);
nand_5 g04894(new_n5279, new_n805, new_n5280);
nand_5 g04895(new_n5280, new_n811, new_n5281);
nand_5 g04896(new_n5281, new_n442, new_n5282);
nand_5 g04897(new_n5282, new_n437, new_n5283);
nand_5 g04898(new_n5283, new_n819, new_n5284);
nand_5 g04899(new_n5284, new_n432, new_n5285);
nand_5 g04900(new_n5285, new_n427_1, new_n5286);
nand_5 g04901(new_n5286, new_n422, new_n5287);
nand_5 g04902(new_n5287, new_n828, new_n5288);
nand_5 g04903(new_n5288, new_n834, new_n5289);
nand_5 g04904(new_n5289, new_n840, new_n5290);
nand_5 g04905(new_n5290, new_n417, new_n5291);
nand_5 g04906(new_n5291, new_n847, new_n5292);
nand_5 g04907(new_n5292, new_n853, new_n5293);
nand_5 g04908(new_n5293, new_n859, new_n5294);
nand_5 g04909(new_n5294, new_n412, new_n5295);
nand_5 g04910(new_n5295, new_n866, new_n5296);
nand_5 g04911(new_n5296, new_n872, new_n5297);
nand_5 g04912(new_n5297, new_n878, new_n5298);
nand_5 g04913(new_n5298, new_n407, new_n5299);
nand_5 g04914(new_n5299, new_n885, new_n5300);
nand_5 g04915(new_n5300, new_n402, new_n5301);
nand_5 g04916(new_n5301, new_n397, new_n5302);
nand_5 g04917(new_n5302, new_n392, new_n5303);
nand_5 g04918(new_n5303, new_n894, new_n5304);
nand_5 g04919(new_n5304, new_n1087, new_n5305);
nand_5 g04920(new_n5305, new_n1129, new_n5306);
nand_5 g04921(new_n5306, new_n1084, new_n5307);
nand_5 g04922(new_n5307, new_n1134, new_n5308);
nand_5 g04923(new_n5308, new_n1080, new_n5309);
nand_5 g04924(new_n5309, new_n1075, new_n5310);
nand_5 g04925(new_n5310, new_n1070, new_n5311);
nand_5 g04926(new_n5311, new_n1143, new_n5312);
nand_5 g04927(new_n5312, new_n1148, new_n5313);
nand_5 g04928(new_n5313, new_n1065, new_n5314);
nand_5 g04929(new_n5314, new_n1062, new_n5315);
nand_5 g04930(new_n5315, new_n1156, new_n5316);
nand_5 g04931(new_n5316, new_n1057, new_n5317);
nand_5 g04932(new_n5317, new_n1053, new_n5318);
nand_5 g04933(new_n5318, new_n1050, new_n5319);
nand_5 g04934(new_n5319, new_n1045, new_n5320);
nand_5 g04935(new_n5320, new_n1040, new_n5321);
nand_5 g04936(new_n5321, new_n1036, new_n5322);
nand_5 g04937(new_n5322, new_n1033, new_n5323);
nand_5 g04938(new_n5323, new_n1028, new_n5324);
nand_5 g04939(new_n5324, new_n1026, new_n5325);
nand_5 g04940(new_n5325, new_n1021, new_n5326);
nand_5 g04941(new_n5326, new_n1017, new_n5327);
nand_5 g04942(new_n5327, new_n1012, new_n5328);
nand_5 g04943(new_n5328, new_n1009, new_n5329);
nand_5 g04944(new_n5329, new_n1004, new_n5330);
nand_5 g04945(new_n5330, new_n1000, new_n5331);
nand_5 g04946(new_n5331, new_n995, new_n5332);
nand_5 g04947(new_n5332, new_n990, new_n5333);
nand_5 g04948(new_n5333, new_n985, new_n5334);
nand_5 g04949(new_n5334, new_n981, new_n5335);
nand_5 g04950(new_n5335, new_n1179, new_n5336);
nand_5 g04951(new_n5336, n5184, new_n5337);
nor_5  g04952(new_n5337, new_n973, n4541);
nand_5 g04953(new_n910, new_n1302, new_n5339);
nand_5 g04954(new_n5339, new_n471, new_n5340);
nand_5 g04955(new_n5340, new_n758, new_n5341);
nand_5 g04956(new_n5341, new_n764, new_n5342);
nand_5 g04957(new_n5342, new_n770, new_n5343);
nand_5 g04958(new_n5343, new_n468, new_n5344);
nand_5 g04959(new_n5344, new_n777, new_n5345);
nand_5 g04960(new_n5345, new_n783, new_n5346);
nand_5 g04961(new_n5346, new_n789, new_n5347);
nand_5 g04962(new_n5347, new_n463, new_n5348);
nand_5 g04963(new_n5348, new_n796, new_n5349);
nand_5 g04964(new_n5349, new_n458, new_n5350);
nand_5 g04965(new_n5350, new_n453, new_n5351);
nand_5 g04966(new_n5351, new_n447, new_n5352);
nand_5 g04967(new_n5352, new_n805, new_n5353);
nand_5 g04968(new_n5353, new_n811, new_n5354);
nand_5 g04969(new_n5354, new_n442, new_n5355);
nand_5 g04970(new_n5355, new_n437, new_n5356);
nand_5 g04971(new_n5356, new_n819, new_n5357);
nand_5 g04972(new_n5357, new_n432, new_n5358);
nand_5 g04973(new_n5358, new_n427_1, new_n5359);
nand_5 g04974(new_n5359, new_n422, new_n5360);
nand_5 g04975(new_n5360, new_n828, new_n5361);
nand_5 g04976(new_n5361, new_n834, new_n5362);
nand_5 g04977(new_n5362, new_n840, new_n5363);
nand_5 g04978(new_n5363, new_n417, new_n5364);
nand_5 g04979(new_n5364, new_n847, new_n5365);
nand_5 g04980(new_n5365, new_n853, new_n5366);
nand_5 g04981(new_n5366, new_n859, new_n5367);
nand_5 g04982(new_n5367, new_n412, new_n5368);
nand_5 g04983(new_n5368, new_n866, new_n5369);
nand_5 g04984(new_n5369, new_n872, new_n5370);
nand_5 g04985(new_n5370, new_n878, new_n5371);
nand_5 g04986(new_n5371, new_n407, new_n5372);
nand_5 g04987(new_n5372, new_n885, new_n5373);
nand_5 g04988(new_n5373, new_n402, new_n5374);
nand_5 g04989(new_n5374, new_n397, new_n5375);
nand_5 g04990(new_n5375, new_n392, new_n5376);
nand_5 g04991(new_n5376, new_n894, new_n5377);
nand_5 g04992(new_n5377, new_n1087, new_n5378);
nand_5 g04993(new_n5378, new_n1129, new_n5379);
nand_5 g04994(new_n5379, new_n1084, new_n5380);
nand_5 g04995(new_n5380, new_n1134, new_n5381);
nand_5 g04996(new_n5381, new_n1080, new_n5382);
nand_5 g04997(new_n5382, new_n1075, new_n5383);
nand_5 g04998(new_n5383, new_n1070, new_n5384);
nand_5 g04999(new_n5384, new_n1143, new_n5385);
nand_5 g05000(new_n5385, new_n1148, new_n5386);
nand_5 g05001(new_n5386, new_n1065, new_n5387);
nand_5 g05002(new_n5387, new_n1062, new_n5388);
nand_5 g05003(new_n5388, new_n1156, new_n5389);
nand_5 g05004(new_n5389, new_n1057, new_n5390);
nand_5 g05005(new_n5390, new_n1053, new_n5391);
nand_5 g05006(new_n5391, new_n1050, new_n5392);
nand_5 g05007(new_n5392, new_n1045, new_n5393);
nand_5 g05008(new_n5393, new_n1040, new_n5394);
nand_5 g05009(new_n5394, new_n1036, new_n5395);
nand_5 g05010(new_n5395, new_n1033, new_n5396);
nand_5 g05011(new_n5396, new_n1028, new_n5397);
nand_5 g05012(new_n5397, new_n1026, new_n5398);
nand_5 g05013(new_n5398, new_n1021, new_n5399);
nand_5 g05014(new_n5399, new_n1017, new_n5400);
nand_5 g05015(new_n5400, new_n1012, new_n5401);
nand_5 g05016(new_n5401, new_n1009, new_n5402);
nand_5 g05017(new_n5402, new_n1004, new_n5403);
nand_5 g05018(new_n5403, new_n1000, new_n5404);
nand_5 g05019(new_n5404, new_n995, new_n5405);
nand_5 g05020(new_n5405, new_n990, new_n5406);
nand_5 g05021(new_n5406, new_n985, new_n5407);
nand_5 g05022(new_n5407, new_n981, new_n5408);
nand_5 g05023(new_n5408, new_n1179, new_n5409);
nand_5 g05024(new_n5409, new_n976, new_n5410);
nand_5 g05025(new_n5410, new_n971, new_n5411);
nand_5 g05026(new_n5411, new_n966, new_n5412);
nand_5 g05027(new_n5412, new_n961, new_n5413);
nand_5 g05028(new_n5413, new_n957, new_n5414);
nand_5 g05029(new_n5414, new_n952, new_n5415);
nand_5 g05030(new_n5415, new_n948_1, new_n5416);
nand_5 g05031(new_n5416, new_n943, new_n5417);
nand_5 g05032(new_n5417, new_n941, new_n5418);
nand_5 g05033(new_n5418, new_n938, new_n5419);
nand_5 g05034(new_n5419, new_n936, new_n5420);
nand_5 g05035(new_n5420, new_n931, new_n5421);
nand_5 g05036(new_n5421, new_n927, new_n5422);
nand_5 g05037(new_n5422, new_n922, new_n5423);
nand_5 g05038(new_n5423, n8302, new_n5424);
nor_5  g05039(new_n5424, new_n914, n4604);
not_4  g05040(new_n1711, new_n5426);
nand_5 g05041(new_n1735, new_n1247, new_n5427);
nand_5 g05042(new_n5427, new_n832, new_n5428);
nand_5 g05043(new_n5428, new_n840, new_n5429);
nand_5 g05044(new_n5429, new_n417, new_n5430_1);
nand_5 g05045(new_n5430_1, new_n847, new_n5431);
nand_5 g05046(new_n5431, new_n853, new_n5432);
nand_5 g05047(new_n5432, new_n859, new_n5433);
nand_5 g05048(new_n5433, new_n412, new_n5434);
nand_5 g05049(new_n5434, new_n866, new_n5435);
nand_5 g05050(new_n5435, new_n872, new_n5436);
nand_5 g05051(new_n5436, new_n878, new_n5437);
nand_5 g05052(new_n5437, new_n407, new_n5438);
nand_5 g05053(new_n5438, new_n885, new_n5439);
nand_5 g05054(new_n5439, new_n402, new_n5440);
nand_5 g05055(new_n5440, new_n397, new_n5441);
nand_5 g05056(new_n5441, new_n392, new_n5442);
nand_5 g05057(new_n5442, new_n894, new_n5443);
nand_5 g05058(new_n5443, new_n1087, new_n5444);
nand_5 g05059(new_n5444, new_n1129, new_n5445);
nand_5 g05060(new_n5445, new_n1084, new_n5446);
nand_5 g05061(new_n5446, new_n1134, new_n5447);
nand_5 g05062(new_n5447, new_n1080, new_n5448);
nand_5 g05063(new_n5448, new_n1075, new_n5449_1);
nand_5 g05064(new_n5449_1, new_n1070, new_n5450);
nand_5 g05065(new_n5450, new_n1143, new_n5451);
nand_5 g05066(new_n5451, new_n1148, new_n5452);
nand_5 g05067(new_n5452, new_n1065, new_n5453);
nand_5 g05068(new_n5453, new_n1062, new_n5454);
nand_5 g05069(new_n5454, new_n1156, new_n5455);
nand_5 g05070(new_n5455, new_n1057, new_n5456);
nand_5 g05071(new_n5456, new_n1053, new_n5457);
nand_5 g05072(new_n5457, new_n1050, new_n5458);
nand_5 g05073(new_n5458, new_n1045, new_n5459);
nand_5 g05074(new_n5459, new_n1040, new_n5460);
nand_5 g05075(new_n5460, new_n1036, new_n5461);
nand_5 g05076(new_n5461, new_n1033, new_n5462);
nand_5 g05077(new_n5462, new_n1028, new_n5463);
nand_5 g05078(new_n5463, new_n1026, new_n5464);
nand_5 g05079(new_n5464, new_n1021, new_n5465);
nand_5 g05080(new_n5465, new_n1017, new_n5466);
nand_5 g05081(new_n5466, new_n1012, new_n5467_1);
nand_5 g05082(new_n5467_1, new_n1009, new_n5468);
nand_5 g05083(new_n5468, new_n1004, new_n5469);
nand_5 g05084(new_n5469, new_n1000, new_n5470);
nand_5 g05085(new_n5470, new_n995, new_n5471);
nand_5 g05086(new_n5471, new_n990, new_n5472);
nand_5 g05087(new_n5472, new_n985, new_n5473);
nand_5 g05088(new_n5473, new_n981, new_n5474);
nand_5 g05089(new_n5474, new_n1179, new_n5475);
nand_5 g05090(new_n5475, new_n976, new_n5476);
nand_5 g05091(new_n5476, new_n971, new_n5477);
nand_5 g05092(new_n5477, new_n966, new_n5478);
nand_5 g05093(new_n5478, new_n961, new_n5479_1);
nand_5 g05094(new_n5479_1, new_n957, new_n5480);
nand_5 g05095(new_n5480, new_n952, new_n5481);
nand_5 g05096(new_n5481, new_n948_1, new_n5482);
nand_5 g05097(new_n5482, new_n943, new_n5483);
nand_5 g05098(new_n5483, new_n941, new_n5484);
nand_5 g05099(new_n5484, new_n938, new_n5485);
nand_5 g05100(new_n5485, new_n936, new_n5486);
nand_5 g05101(new_n5486, new_n931, new_n5487);
nand_5 g05102(new_n5487, new_n927, new_n5488);
nand_5 g05103(new_n5488, new_n922, new_n5489);
nand_5 g05104(new_n5489, new_n917, new_n5490);
nand_5 g05105(new_n5490, new_n912, new_n5491);
nand_5 g05106(new_n5491, new_n907, new_n5492);
nand_5 g05107(new_n5492, new_n903, new_n5493);
nand_5 g05108(new_n5493, new_n2066, new_n5494);
nand_5 g05109(new_n5494, new_n2063, new_n5495);
nand_5 g05110(new_n5495, new_n2062, new_n5496);
nand_5 g05111(new_n5496, new_n2058, new_n5497);
nand_5 g05112(new_n5497, new_n2055, new_n5498);
nand_5 g05113(new_n5498, new_n2051, new_n5499);
nand_5 g05114(new_n5499, new_n2046, new_n5500);
nand_5 g05115(new_n5500, new_n2042, new_n5501);
nand_5 g05116(new_n5501, new_n2039, new_n5502_1);
nand_5 g05117(new_n5502_1, new_n2036, new_n5503);
nand_5 g05118(new_n5503, new_n2033, new_n5504);
nand_5 g05119(new_n5504, new_n2029, new_n5505);
nand_5 g05120(new_n5505, new_n2026, new_n5506);
nand_5 g05121(new_n5506, new_n2022, new_n5507);
nand_5 g05122(new_n5507, new_n2018, new_n5508);
nand_5 g05123(new_n5508, new_n1726, new_n5509);
nand_5 g05124(new_n5509, new_n1722, new_n5510);
nand_5 g05125(new_n5510, new_n1718, new_n5511);
nand_5 g05126(new_n5511, n12976, new_n5512);
nor_5  g05127(new_n5512, new_n5426, n4672);
nor_5  g05128(n13295, n760, new_n5514);
not_4  g05129(new_n5514, new_n5515);
nand_5 g05130(new_n5515, new_n1789, new_n5516);
nand_5 g05131(new_n5516, new_n1608, new_n5517);
nand_5 g05132(new_n5517, new_n1605, new_n5518);
nand_5 g05133(new_n5518, new_n1795, new_n5519);
nand_5 g05134(new_n5519, new_n1799, new_n5520);
nand_5 g05135(new_n5520, new_n1602, new_n5521);
nand_5 g05136(new_n5521, new_n1599, new_n5522);
nand_5 g05137(new_n5522, new_n1596, new_n5523);
nand_5 g05138(new_n5523, new_n1593, new_n5524);
nand_5 g05139(new_n5524, new_n1806, new_n5525);
nand_5 g05140(new_n5525, new_n1589, new_n5526);
nand_5 g05141(new_n5526, new_n1586, new_n5527);
nand_5 g05142(new_n5527, new_n1583, new_n5528);
nand_5 g05143(new_n5528, new_n1580, new_n5529);
nand_5 g05144(new_n5529, new_n1576, new_n5530);
nand_5 g05145(new_n5530, new_n1573, new_n5531);
nand_5 g05146(new_n5531, new_n1570, new_n5532);
nand_5 g05147(new_n5532, new_n1567, new_n5533);
nand_5 g05148(new_n5533, new_n1564, new_n5534);
nand_5 g05149(new_n5534, new_n1561, new_n5535);
nand_5 g05150(new_n5535, new_n1338, new_n5536);
nand_5 g05151(new_n5536, new_n1331, new_n5537);
nand_5 g05152(new_n5537, new_n1326, new_n5538);
nand_5 g05153(new_n5538, new_n1321, new_n5539);
nand_5 g05154(new_n5539, new_n1318, new_n5540);
nand_5 g05155(new_n5540, new_n1315, new_n5541);
nand_5 g05156(new_n5541, new_n1312, new_n5542);
nand_5 g05157(new_n5542, new_n1309, new_n5543);
nand_5 g05158(new_n5543, new_n1307, new_n5544);
nand_5 g05159(new_n5544, new_n1304, new_n5545);
nand_5 g05160(new_n5545, new_n1300, new_n5546);
nand_5 g05161(new_n5546, new_n1297, new_n5547);
nand_5 g05162(new_n5547, new_n1294, new_n5548);
nand_5 g05163(new_n5548, new_n1355, new_n5549);
nand_5 g05164(new_n5549, new_n1291, new_n5550_1);
nand_5 g05165(new_n5550_1, new_n1288, new_n5551);
nand_5 g05166(new_n5551, new_n1283, new_n5552);
nand_5 g05167(new_n5552, new_n1363, new_n5553);
nand_5 g05168(new_n5553, new_n1280, new_n5554);
nand_5 g05169(new_n5554, new_n1370, new_n5555);
nand_5 g05170(new_n5555, new_n1373, new_n5556);
nand_5 g05171(new_n5556, new_n1277, new_n5557);
nand_5 g05172(new_n5557, new_n1272, new_n5558);
nand_5 g05173(new_n5558, new_n1269, new_n5559);
nand_5 g05174(new_n5559, new_n1380, new_n5560);
nand_5 g05175(new_n5560, new_n1264, new_n5561);
nand_5 g05176(new_n5561, new_n1259, new_n5562);
nand_5 g05177(new_n5562, new_n1388, new_n5563);
nand_5 g05178(new_n5563, new_n1392, new_n5564);
nand_5 g05179(new_n5564, new_n1256, new_n5565);
nand_5 g05180(new_n5565, new_n1252, new_n5566);
nand_5 g05181(new_n5566, new_n1249, new_n5567);
nand_5 g05182(new_n5567, new_n1244, new_n5568);
nand_5 g05183(new_n5568, new_n1240, new_n5569);
nand_5 g05184(new_n5569, new_n1234, new_n5570);
nand_5 g05185(new_n5570, new_n1231, new_n5571);
nand_5 g05186(new_n5571, new_n1227, new_n5572);
nand_5 g05187(new_n5572, new_n1407, new_n5573);
nand_5 g05188(new_n5573, new_n1223, new_n5574);
nand_5 g05189(new_n5574, new_n1218, new_n5575);
nand_5 g05190(new_n5575, new_n1213, new_n5576);
nand_5 g05191(new_n5576, new_n1210, new_n5577);
nand_5 g05192(new_n5577, new_n1206, new_n5578);
nand_5 g05193(new_n5578, new_n1418, new_n5579);
nand_5 g05194(new_n5579, new_n1422, new_n5580);
nand_5 g05195(new_n5580, new_n1428, new_n5581);
nand_5 g05196(new_n5581, new_n1203, new_n5582);
nand_5 g05197(new_n5582, new_n1433, new_n5583);
nand_5 g05198(new_n5583, new_n581, new_n5584);
nand_5 g05199(new_n5584, new_n574, new_n5585);
nand_5 g05200(new_n5585, new_n568, new_n5586_1);
nand_5 g05201(new_n5586_1, new_n589, new_n5587);
nand_5 g05202(new_n5587, new_n595, new_n5588);
nand_5 g05203(new_n5588, new_n601, new_n5589);
nand_5 g05204(new_n5589, new_n563, new_n5590);
nand_5 g05205(new_n5590, new_n608, new_n5591);
nand_5 g05206(new_n5591, new_n558, new_n5592);
nand_5 g05207(new_n5592, new_n615, new_n5593);
nand_5 g05208(new_n5593, new_n553, new_n5594);
nand_5 g05209(new_n5594, new_n622, new_n5595);
nand_5 g05210(new_n5595, new_n628, new_n5596);
nand_5 g05211(new_n5596, new_n548, new_n5597);
nand_5 g05212(new_n5597, new_n543_1, new_n5598);
nand_5 g05213(new_n5598, new_n636, new_n5599);
nand_5 g05214(new_n5599, n3652, new_n5600);
nor_5  g05215(new_n5600, new_n639, n4858);
nand_5 g05216(new_n1648, new_n1078, new_n5602);
nand_5 g05217(new_n5602, new_n1075, new_n5603);
nand_5 g05218(new_n5603, new_n1070, new_n5604);
nand_5 g05219(new_n5604, new_n1143, new_n5605);
nand_5 g05220(new_n5605, new_n1148, new_n5606);
nand_5 g05221(new_n5606, new_n1065, new_n5607);
nand_5 g05222(new_n5607, new_n1062, new_n5608);
nand_5 g05223(new_n5608, new_n1156, new_n5609);
nand_5 g05224(new_n5609, new_n1057, new_n5610);
nand_5 g05225(new_n5610, new_n1053, new_n5611);
nand_5 g05226(new_n5611, new_n1050, new_n5612);
nand_5 g05227(new_n5612, new_n1045, new_n5613);
nand_5 g05228(new_n5613, new_n1040, new_n5614);
nand_5 g05229(new_n5614, new_n1036, new_n5615);
nand_5 g05230(new_n5615, new_n1033, new_n5616);
nand_5 g05231(new_n5616, new_n1028, new_n5617);
nand_5 g05232(new_n5617, new_n1026, new_n5618);
nand_5 g05233(new_n5618, new_n1021, new_n5619);
nand_5 g05234(new_n5619, new_n1017, new_n5620);
nand_5 g05235(new_n5620, new_n1012, new_n5621);
nand_5 g05236(new_n5621, new_n1009, new_n5622);
nand_5 g05237(new_n5622, new_n1004, new_n5623);
nand_5 g05238(new_n5623, new_n1000, new_n5624);
nand_5 g05239(new_n5624, new_n995, new_n5625);
nand_5 g05240(new_n5625, new_n990, new_n5626);
nand_5 g05241(new_n5626, new_n985, new_n5627);
nand_5 g05242(new_n5627, new_n981, new_n5628);
nand_5 g05243(new_n5628, new_n1179, new_n5629);
nand_5 g05244(new_n5629, new_n976, new_n5630);
nand_5 g05245(new_n5630, new_n971, new_n5631);
nand_5 g05246(new_n5631, new_n966, new_n5632);
nand_5 g05247(new_n5632, new_n961, new_n5633);
nand_5 g05248(new_n5633, new_n957, new_n5634);
nand_5 g05249(new_n5634, new_n952, new_n5635);
nand_5 g05250(new_n5635, new_n948_1, new_n5636);
nand_5 g05251(new_n5636, new_n943, new_n5637);
nand_5 g05252(new_n5637, new_n941, new_n5638);
nand_5 g05253(new_n5638, new_n938, new_n5639);
nand_5 g05254(new_n5639, new_n936, new_n5640);
nand_5 g05255(new_n5640, new_n931, new_n5641);
nand_5 g05256(new_n5641, new_n927, new_n5642);
nand_5 g05257(new_n5642, new_n922, new_n5643);
nand_5 g05258(new_n5643, new_n917, new_n5644);
nand_5 g05259(new_n5644, new_n912, new_n5645);
nand_5 g05260(new_n5645, new_n907, new_n5646);
nand_5 g05261(new_n5646, new_n903, new_n5647);
nand_5 g05262(new_n5647, new_n2066, new_n5648);
nand_5 g05263(new_n5648, new_n2063, new_n5649);
nand_5 g05264(new_n5649, new_n2062, new_n5650);
nand_5 g05265(new_n5650, new_n2058, new_n5651);
nand_5 g05266(new_n5651, new_n2055, new_n5652);
nand_5 g05267(new_n5652, new_n2051, new_n5653);
nand_5 g05268(new_n5653, new_n2046, new_n5654);
nand_5 g05269(new_n5654, new_n2042, new_n5655);
nand_5 g05270(new_n5655, new_n2039, new_n5656);
nand_5 g05271(new_n5656, new_n2036, new_n5657);
nand_5 g05272(new_n5657, new_n2033, new_n5658);
nand_5 g05273(new_n5658, new_n2029, new_n5659);
nand_5 g05274(new_n5659, new_n2026, new_n5660);
nand_5 g05275(new_n5660, new_n2022, new_n5661);
nand_5 g05276(new_n5661, new_n2018, new_n5662);
nand_5 g05277(new_n5662, new_n1726, new_n5663);
nand_5 g05278(new_n5663, new_n1722, new_n5664);
nand_5 g05279(new_n5664, new_n1718, new_n5665);
nand_5 g05280(new_n5665, new_n1713, new_n5666);
nand_5 g05281(new_n5666, new_n1737, new_n5667);
nand_5 g05282(new_n5667, new_n1709, new_n5668);
nand_5 g05283(new_n5668, new_n1742, new_n5669);
nand_5 g05284(new_n5669, new_n1704, new_n5670);
nand_5 g05285(new_n5670, new_n1702_1, new_n5671);
nand_5 g05286(new_n5671, new_n1698, new_n5672);
nand_5 g05287(new_n5672, new_n1695, new_n5673);
nand_5 g05288(new_n5673, new_n1692, new_n5674);
nand_5 g05289(new_n5674, new_n1752, new_n5675);
nand_5 g05290(new_n5675, new_n1688, new_n5676);
nand_5 g05291(new_n5676, new_n1685, new_n5677);
nand_5 g05292(new_n5677, new_n1680, new_n5678);
nand_5 g05293(new_n5678, new_n1676, new_n5679);
nand_5 g05294(new_n5679, new_n1672, new_n5680);
nand_5 g05295(new_n5680, new_n1669, new_n5681);
nand_5 g05296(new_n5681, new_n1666, new_n5682);
nand_5 g05297(new_n5682, new_n1663, new_n5683);
nand_5 g05298(new_n5683, new_n1658, new_n5684);
nand_5 g05299(new_n5684, new_n1653, new_n5685);
nand_5 g05300(new_n5685, n1222, new_n5686);
nor_5  g05301(new_n5686, new_n571, n4971);
not_4  g05302(new_n905, new_n5688);
nand_5 g05303(new_n902, new_n762, new_n5689);
nand_5 g05304(new_n5689, new_n770, new_n5690);
nand_5 g05305(new_n5690, new_n468, new_n5691);
nand_5 g05306(new_n5691, new_n777, new_n5692);
nand_5 g05307(new_n5692, new_n783, new_n5693);
nand_5 g05308(new_n5693, new_n789, new_n5694);
nand_5 g05309(new_n5694, new_n463, new_n5695);
nand_5 g05310(new_n5695, new_n796, new_n5696);
nand_5 g05311(new_n5696, new_n458, new_n5697);
nand_5 g05312(new_n5697, new_n453, new_n5698);
nand_5 g05313(new_n5698, new_n447, new_n5699);
nand_5 g05314(new_n5699, new_n805, new_n5700);
nand_5 g05315(new_n5700, new_n811, new_n5701);
nand_5 g05316(new_n5701, new_n442, new_n5702);
nand_5 g05317(new_n5702, new_n437, new_n5703);
nand_5 g05318(new_n5703, new_n819, new_n5704);
nand_5 g05319(new_n5704, new_n432, new_n5705);
nand_5 g05320(new_n5705, new_n427_1, new_n5706);
nand_5 g05321(new_n5706, new_n422, new_n5707);
nand_5 g05322(new_n5707, new_n828, new_n5708);
nand_5 g05323(new_n5708, new_n834, new_n5709);
nand_5 g05324(new_n5709, new_n840, new_n5710);
nand_5 g05325(new_n5710, new_n417, new_n5711);
nand_5 g05326(new_n5711, new_n847, new_n5712);
nand_5 g05327(new_n5712, new_n853, new_n5713);
nand_5 g05328(new_n5713, new_n859, new_n5714);
nand_5 g05329(new_n5714, new_n412, new_n5715);
nand_5 g05330(new_n5715, new_n866, new_n5716);
nand_5 g05331(new_n5716, new_n872, new_n5717);
nand_5 g05332(new_n5717, new_n878, new_n5718);
nand_5 g05333(new_n5718, new_n407, new_n5719);
nand_5 g05334(new_n5719, new_n885, new_n5720);
nand_5 g05335(new_n5720, new_n402, new_n5721);
nand_5 g05336(new_n5721, new_n397, new_n5722);
nand_5 g05337(new_n5722, new_n392, new_n5723);
nand_5 g05338(new_n5723, new_n894, new_n5724);
nand_5 g05339(new_n5724, new_n1087, new_n5725_1);
nand_5 g05340(new_n5725_1, new_n1129, new_n5726);
nand_5 g05341(new_n5726, new_n1084, new_n5727);
nand_5 g05342(new_n5727, new_n1134, new_n5728);
nand_5 g05343(new_n5728, new_n1080, new_n5729);
nand_5 g05344(new_n5729, new_n1075, new_n5730);
nand_5 g05345(new_n5730, new_n1070, new_n5731);
nand_5 g05346(new_n5731, new_n1143, new_n5732);
nand_5 g05347(new_n5732, new_n1148, new_n5733);
nand_5 g05348(new_n5733, new_n1065, new_n5734);
nand_5 g05349(new_n5734, new_n1062, new_n5735);
nand_5 g05350(new_n5735, new_n1156, new_n5736);
nand_5 g05351(new_n5736, new_n1057, new_n5737);
nand_5 g05352(new_n5737, new_n1053, new_n5738);
nand_5 g05353(new_n5738, new_n1050, new_n5739);
nand_5 g05354(new_n5739, new_n1045, new_n5740);
nand_5 g05355(new_n5740, new_n1040, new_n5741);
nand_5 g05356(new_n5741, new_n1036, new_n5742);
nand_5 g05357(new_n5742, new_n1033, new_n5743);
nand_5 g05358(new_n5743, new_n1028, new_n5744);
nand_5 g05359(new_n5744, new_n1026, new_n5745);
nand_5 g05360(new_n5745, new_n1021, new_n5746);
nand_5 g05361(new_n5746, new_n1017, new_n5747);
nand_5 g05362(new_n5747, new_n1012, new_n5748);
nand_5 g05363(new_n5748, new_n1009, new_n5749);
nand_5 g05364(new_n5749, new_n1004, new_n5750);
nand_5 g05365(new_n5750, new_n1000, new_n5751);
nand_5 g05366(new_n5751, new_n995, new_n5752);
nand_5 g05367(new_n5752, new_n990, new_n5753);
nand_5 g05368(new_n5753, new_n985, new_n5754);
nand_5 g05369(new_n5754, new_n981, new_n5755);
nand_5 g05370(new_n5755, new_n1179, new_n5756);
nand_5 g05371(new_n5756, new_n976, new_n5757);
nand_5 g05372(new_n5757, new_n971, new_n5758);
nand_5 g05373(new_n5758, new_n966, new_n5759);
nand_5 g05374(new_n5759, new_n961, new_n5760);
nand_5 g05375(new_n5760, new_n957, new_n5761);
nand_5 g05376(new_n5761, new_n952, new_n5762);
nand_5 g05377(new_n5762, new_n948_1, new_n5763);
nand_5 g05378(new_n5763, new_n943, new_n5764);
nand_5 g05379(new_n5764, new_n941, new_n5765);
nand_5 g05380(new_n5765, new_n938, new_n5766);
nand_5 g05381(new_n5766, new_n936, new_n5767);
nand_5 g05382(new_n5767, new_n931, new_n5768);
nand_5 g05383(new_n5768, new_n927, new_n5769);
nand_5 g05384(new_n5769, new_n922, new_n5770);
nand_5 g05385(new_n5770, new_n917, new_n5771);
nand_5 g05386(new_n5771, new_n912, new_n5772);
nand_5 g05387(new_n5772, n14072, new_n5773);
nor_5  g05388(new_n5773, new_n5688, n5479);
nand_5 g05389(new_n1670, new_n1417, new_n5775);
nand_5 g05390(new_n5775, new_n1669, new_n5776);
nand_5 g05391(new_n5776, new_n1666, new_n5777);
nand_5 g05392(new_n5777, new_n1663, new_n5778);
nand_5 g05393(new_n5778, new_n1658, new_n5779);
nand_5 g05394(new_n5779, new_n1653, new_n5780);
nand_5 g05395(new_n5780, new_n1651, new_n5781);
nand_5 g05396(new_n5781, new_n1649, new_n5782);
nand_5 g05397(new_n5782, new_n1646, new_n5783);
nand_5 g05398(new_n5783, new_n1643, new_n5784);
nand_5 g05399(new_n5784, new_n1641, new_n5785);
nand_5 g05400(new_n5785, new_n1638, new_n5786_1);
nand_5 g05401(new_n5786_1, new_n1635, new_n5787);
nand_5 g05402(new_n5787, new_n1632, new_n5788);
nand_5 g05403(new_n5788, new_n1628, new_n5789);
nand_5 g05404(new_n5789, new_n1625, new_n5790);
nand_5 g05405(new_n5790, new_n1621, new_n5791);
nand_5 g05406(new_n5791, new_n1618, new_n5792);
nand_5 g05407(new_n5792, new_n1778, new_n5793);
nand_5 g05408(new_n5793, new_n1782, new_n5794);
nand_5 g05409(new_n5794, new_n1614, new_n5795);
nand_5 g05410(new_n5795, new_n1611, new_n5796);
nand_5 g05411(new_n5796, new_n1789, new_n5797);
nand_5 g05412(new_n5797, new_n1608, new_n5798);
nand_5 g05413(new_n5798, new_n1605, new_n5799);
nand_5 g05414(new_n5799, new_n1795, new_n5800);
nand_5 g05415(new_n5800, new_n1799, new_n5801);
nand_5 g05416(new_n5801, new_n1602, new_n5802);
nand_5 g05417(new_n5802, new_n1599, new_n5803);
nand_5 g05418(new_n5803, new_n1596, new_n5804);
nand_5 g05419(new_n5804, new_n1593, new_n5805);
nand_5 g05420(new_n5805, new_n1806, new_n5806_1);
nand_5 g05421(new_n5806_1, new_n1589, new_n5807);
nand_5 g05422(new_n5807, new_n1586, new_n5808);
nand_5 g05423(new_n5808, new_n1583, new_n5809);
nand_5 g05424(new_n5809, new_n1580, new_n5810);
nand_5 g05425(new_n5810, new_n1576, new_n5811);
nand_5 g05426(new_n5811, new_n1573, new_n5812);
nand_5 g05427(new_n5812, new_n1570, new_n5813);
nand_5 g05428(new_n5813, new_n1567, new_n5814);
nand_5 g05429(new_n5814, new_n1564, new_n5815);
nand_5 g05430(new_n5815, new_n1561, new_n5816);
nand_5 g05431(new_n5816, new_n1338, new_n5817);
nand_5 g05432(new_n5817, new_n1331, new_n5818);
nand_5 g05433(new_n5818, new_n1326, new_n5819);
nand_5 g05434(new_n5819, new_n1321, new_n5820);
nand_5 g05435(new_n5820, new_n1318, new_n5821);
nand_5 g05436(new_n5821, new_n1315, new_n5822);
nand_5 g05437(new_n5822, new_n1312, new_n5823);
nand_5 g05438(new_n5823, new_n1309, new_n5824);
nand_5 g05439(new_n5824, new_n1307, new_n5825);
nand_5 g05440(new_n5825, new_n1304, new_n5826);
nand_5 g05441(new_n5826, new_n1300, new_n5827);
nand_5 g05442(new_n5827, new_n1297, new_n5828);
nand_5 g05443(new_n5828, new_n1294, new_n5829);
nand_5 g05444(new_n5829, new_n1355, new_n5830);
nand_5 g05445(new_n5830, new_n1291, new_n5831);
nand_5 g05446(new_n5831, new_n1288, new_n5832);
nand_5 g05447(new_n5832, new_n1283, new_n5833);
nand_5 g05448(new_n5833, new_n1363, new_n5834);
nand_5 g05449(new_n5834, new_n1280, new_n5835);
nand_5 g05450(new_n5835, new_n1370, new_n5836);
nand_5 g05451(new_n5836, new_n1373, new_n5837);
nand_5 g05452(new_n5837, new_n1277, new_n5838);
nand_5 g05453(new_n5838, new_n1272, new_n5839);
nand_5 g05454(new_n5839, new_n1269, new_n5840);
nand_5 g05455(new_n5840, new_n1380, new_n5841);
nand_5 g05456(new_n5841, new_n1264, new_n5842);
nand_5 g05457(new_n5842, new_n1259, new_n5843);
nand_5 g05458(new_n5843, new_n1388, new_n5844);
nand_5 g05459(new_n5844, new_n1392, new_n5845);
nand_5 g05460(new_n5845, new_n1256, new_n5846);
nand_5 g05461(new_n5846, new_n1252, new_n5847);
nand_5 g05462(new_n5847, new_n1249, new_n5848);
nand_5 g05463(new_n5848, new_n1244, new_n5849);
nand_5 g05464(new_n5849, new_n1240, new_n5850);
nand_5 g05465(new_n5850, new_n1234, new_n5851_1);
nand_5 g05466(new_n5851_1, new_n1231, new_n5852);
nand_5 g05467(new_n5852, new_n1227, new_n5853);
nand_5 g05468(new_n5853, new_n1407, new_n5854);
nand_5 g05469(new_n5854, new_n1223, new_n5855);
nand_5 g05470(new_n5855, new_n1218, new_n5856);
nand_5 g05471(new_n5856, new_n1213, new_n5857);
nand_5 g05472(new_n5857, new_n1210, new_n5858);
nand_5 g05473(new_n5858, n5046, new_n5859);
nor_5  g05474(new_n5859, new_n882, n5550);
not_4  g05475(new_n803, new_n5861);
nand_5 g05476(new_n1272, new_n5861, new_n5862);
nand_5 g05477(new_n5862, new_n1269, new_n5863);
nand_5 g05478(new_n5863, new_n1380, new_n5864);
nand_5 g05479(new_n5864, new_n1264, new_n5865);
nand_5 g05480(new_n5865, new_n1259, new_n5866);
nand_5 g05481(new_n5866, new_n1388, new_n5867);
nand_5 g05482(new_n5867, new_n1392, new_n5868);
nand_5 g05483(new_n5868, new_n1256, new_n5869);
nand_5 g05484(new_n5869, new_n1252, new_n5870);
nand_5 g05485(new_n5870, new_n1249, new_n5871);
nand_5 g05486(new_n5871, new_n1244, new_n5872);
nand_5 g05487(new_n5872, new_n1240, new_n5873);
nand_5 g05488(new_n5873, new_n1234, new_n5874);
nand_5 g05489(new_n5874, new_n1231, new_n5875);
nand_5 g05490(new_n5875, new_n1227, new_n5876);
nand_5 g05491(new_n5876, new_n1407, new_n5877);
nand_5 g05492(new_n5877, new_n1223, new_n5878);
nand_5 g05493(new_n5878, new_n1218, new_n5879);
nand_5 g05494(new_n5879, new_n1213, new_n5880);
nand_5 g05495(new_n5880, new_n1210, new_n5881);
nand_5 g05496(new_n5881, new_n1206, new_n5882);
nand_5 g05497(new_n5882, new_n1418, new_n5883);
nand_5 g05498(new_n5883, new_n1422, new_n5884);
nand_5 g05499(new_n5884, new_n1428, new_n5885);
nand_5 g05500(new_n5885, new_n1203, new_n5886);
nand_5 g05501(new_n5886, new_n1433, new_n5887);
nand_5 g05502(new_n5887, new_n581, new_n5888);
nand_5 g05503(new_n5888, new_n574, new_n5889);
nand_5 g05504(new_n5889, new_n568, new_n5890);
nand_5 g05505(new_n5890, new_n589, new_n5891);
nand_5 g05506(new_n5891, new_n595, new_n5892);
nand_5 g05507(new_n5892, new_n601, new_n5893);
nand_5 g05508(new_n5893, new_n563, new_n5894);
nand_5 g05509(new_n5894, new_n608, new_n5895);
nand_5 g05510(new_n5895, new_n558, new_n5896);
nand_5 g05511(new_n5896, new_n615, new_n5897);
nand_5 g05512(new_n5897, new_n553, new_n5898);
nand_5 g05513(new_n5898, new_n622, new_n5899);
nand_5 g05514(new_n5899, new_n628, new_n5900);
nand_5 g05515(new_n5900, new_n548, new_n5901);
nand_5 g05516(new_n5901, new_n543_1, new_n5902);
nand_5 g05517(new_n5902, new_n636, new_n5903);
nand_5 g05518(new_n5903, new_n642, new_n5904);
nand_5 g05519(new_n5904, new_n538, new_n5905);
nand_5 g05520(new_n5905, new_n533, new_n5906);
nand_5 g05521(new_n5906, new_n650_1, new_n5907);
nand_5 g05522(new_n5907, new_n528, new_n5908);
nand_5 g05523(new_n5908, new_n523, new_n5909);
nand_5 g05524(new_n5909, new_n518, new_n5910);
nand_5 g05525(new_n5910, new_n659, new_n5911);
nand_5 g05526(new_n5911, new_n665, new_n5912);
nand_5 g05527(new_n5912, new_n672, new_n5913);
nand_5 g05528(new_n5913, new_n513, new_n5914);
nand_5 g05529(new_n5914, new_n679, new_n5915);
nand_5 g05530(new_n5915, new_n685, new_n5916);
nand_5 g05531(new_n5916, new_n691, new_n5917);
nand_5 g05532(new_n5917, new_n508, new_n5918);
nand_5 g05533(new_n5918, new_n698, new_n5919);
nand_5 g05534(new_n5919, new_n503, new_n5920);
nand_5 g05535(new_n5920, new_n704, new_n5921);
nand_5 g05536(new_n5921, new_n498_1, new_n5922);
nand_5 g05537(new_n5922, new_n711, new_n5923);
nand_5 g05538(new_n5923, new_n493, new_n5924);
nand_5 g05539(new_n5924, new_n718, new_n5925);
nand_5 g05540(new_n5925, new_n488, new_n5926);
nand_5 g05541(new_n5926, new_n725, new_n5927);
nand_5 g05542(new_n5927, new_n483, new_n5928);
nand_5 g05543(new_n5928, new_n732, new_n5929);
nand_5 g05544(new_n5929, new_n478, new_n5930);
nand_5 g05545(new_n5930, new_n739, new_n5931);
nand_5 g05546(new_n5931, new_n745, new_n5932);
nand_5 g05547(new_n5932, new_n751, new_n5933);
nand_5 g05548(new_n5933, new_n473, new_n5934);
nand_5 g05549(new_n5934, new_n758, new_n5935);
nand_5 g05550(new_n5935, new_n764, new_n5936);
nand_5 g05551(new_n5936, new_n770, new_n5937);
nand_5 g05552(new_n5937, new_n468, new_n5938);
nand_5 g05553(new_n5938, new_n777, new_n5939);
nand_5 g05554(new_n5939, new_n783, new_n5940);
nand_5 g05555(new_n5940, new_n789, new_n5941);
nand_5 g05556(new_n5941, new_n463, new_n5942);
nand_5 g05557(new_n5942, new_n796, new_n5943_1);
nand_5 g05558(new_n5943_1, new_n458, new_n5944);
nand_5 g05559(new_n5944, new_n453, new_n5945);
nand_5 g05560(new_n5945, n8552, new_n5946);
nor_5  g05561(new_n5946, new_n444, n5586);
nand_5 g05562(new_n1601, new_n1007, new_n5948);
nand_5 g05563(new_n5948, new_n1004, new_n5949);
nand_5 g05564(new_n5949, new_n1000, new_n5950_1);
nand_5 g05565(new_n5950_1, new_n995, new_n5951);
nand_5 g05566(new_n5951, new_n990, new_n5952);
nand_5 g05567(new_n5952, new_n985, new_n5953);
nand_5 g05568(new_n5953, new_n981, new_n5954);
nand_5 g05569(new_n5954, new_n1179, new_n5955);
nand_5 g05570(new_n5955, new_n976, new_n5956);
nand_5 g05571(new_n5956, new_n971, new_n5957);
nand_5 g05572(new_n5957, new_n966, new_n5958);
nand_5 g05573(new_n5958, new_n961, new_n5959);
nand_5 g05574(new_n5959, new_n957, new_n5960_1);
nand_5 g05575(new_n5960_1, new_n952, new_n5961);
nand_5 g05576(new_n5961, new_n948_1, new_n5962);
nand_5 g05577(new_n5962, new_n943, new_n5963);
nand_5 g05578(new_n5963, new_n941, new_n5964);
nand_5 g05579(new_n5964, new_n938, new_n5965);
nand_5 g05580(new_n5965, new_n936, new_n5966);
nand_5 g05581(new_n5966, new_n931, new_n5967);
nand_5 g05582(new_n5967, new_n927, new_n5968);
nand_5 g05583(new_n5968, new_n922, new_n5969);
nand_5 g05584(new_n5969, new_n917, new_n5970);
nand_5 g05585(new_n5970, new_n912, new_n5971);
nand_5 g05586(new_n5971, new_n907, new_n5972);
nand_5 g05587(new_n5972, new_n903, new_n5973);
nand_5 g05588(new_n5973, new_n2066, new_n5974);
nand_5 g05589(new_n5974, new_n2063, new_n5975);
nand_5 g05590(new_n5975, new_n2062, new_n5976);
nand_5 g05591(new_n5976, new_n2058, new_n5977);
nand_5 g05592(new_n5977, new_n2055, new_n5978);
nand_5 g05593(new_n5978, new_n2051, new_n5979);
nand_5 g05594(new_n5979, new_n2046, new_n5980);
nand_5 g05595(new_n5980, new_n2042, new_n5981);
nand_5 g05596(new_n5981, new_n2039, new_n5982);
nand_5 g05597(new_n5982, new_n2036, new_n5983);
nand_5 g05598(new_n5983, new_n2033, new_n5984);
nand_5 g05599(new_n5984, new_n2029, new_n5985);
nand_5 g05600(new_n5985, new_n2026, new_n5986);
nand_5 g05601(new_n5986, new_n2022, new_n5987_1);
nand_5 g05602(new_n5987_1, new_n2018, new_n5988);
nand_5 g05603(new_n5988, new_n1726, new_n5989);
nand_5 g05604(new_n5989, new_n1722, new_n5990);
nand_5 g05605(new_n5990, new_n1718, new_n5991);
nand_5 g05606(new_n5991, new_n1713, new_n5992);
nand_5 g05607(new_n5992, new_n1737, new_n5993);
nand_5 g05608(new_n5993, new_n1709, new_n5994);
nand_5 g05609(new_n5994, new_n1742, new_n5995);
nand_5 g05610(new_n5995, new_n1704, new_n5996);
nand_5 g05611(new_n5996, new_n1702_1, new_n5997);
nand_5 g05612(new_n5997, new_n1698, new_n5998);
nand_5 g05613(new_n5998, new_n1695, new_n5999);
nand_5 g05614(new_n5999, new_n1692, new_n6000);
nand_5 g05615(new_n6000, new_n1752, new_n6001);
nand_5 g05616(new_n6001, new_n1688, new_n6002);
nand_5 g05617(new_n6002, new_n1685, new_n6003);
nand_5 g05618(new_n6003, new_n1680, new_n6004);
nand_5 g05619(new_n6004, new_n1676, new_n6005);
nand_5 g05620(new_n6005, new_n1672, new_n6006);
nand_5 g05621(new_n6006, new_n1669, new_n6007_1);
nand_5 g05622(new_n6007_1, new_n1666, new_n6008);
nand_5 g05623(new_n6008, new_n1663, new_n6009);
nand_5 g05624(new_n6009, new_n1658, new_n6010);
nand_5 g05625(new_n6010, new_n1653, new_n6011);
nand_5 g05626(new_n6011, new_n1651, new_n6012_1);
nand_5 g05627(new_n6012_1, new_n1649, new_n6013);
nand_5 g05628(new_n6013, new_n1646, new_n6014);
nand_5 g05629(new_n6014, new_n1643, new_n6015);
nand_5 g05630(new_n6015, new_n1641, new_n6016);
nand_5 g05631(new_n6016, new_n1638, new_n6017);
nand_5 g05632(new_n6017, new_n1635, new_n6018);
nand_5 g05633(new_n6018, new_n1632, new_n6019);
nand_5 g05634(new_n6019, new_n1628, new_n6020);
nand_5 g05635(new_n6020, new_n1625, new_n6021);
nand_5 g05636(new_n6021, new_n1621, new_n6022);
nand_5 g05637(new_n6022, new_n1618, new_n6023);
nand_5 g05638(new_n6023, new_n1778, new_n6024);
nand_5 g05639(new_n6024, new_n1782, new_n6025);
nand_5 g05640(new_n6025, new_n1614, new_n6026);
nand_5 g05641(new_n6026, new_n1611, new_n6027);
nand_5 g05642(new_n6027, new_n1789, new_n6028);
nand_5 g05643(new_n6028, new_n1608, new_n6029);
nand_5 g05644(new_n6029, new_n1605, new_n6030);
nand_5 g05645(new_n6030, new_n1795, new_n6031);
nand_5 g05646(new_n6031, n7652, new_n6032);
nor_5  g05647(new_n6032, new_n520, n5806);
nand_5 g05648(new_n1683, new_n1208, new_n6034);
nand_5 g05649(new_n6034, new_n405, new_n6035);
nand_5 g05650(new_n6035, new_n885, new_n6036);
nand_5 g05651(new_n6036, new_n402, new_n6037);
nand_5 g05652(new_n6037, new_n397, new_n6038);
nand_5 g05653(new_n6038, new_n392, new_n6039);
nand_5 g05654(new_n6039, new_n894, new_n6040);
nand_5 g05655(new_n6040, new_n1087, new_n6041);
nand_5 g05656(new_n6041, new_n1129, new_n6042);
nand_5 g05657(new_n6042, new_n1084, new_n6043);
nand_5 g05658(new_n6043, new_n1134, new_n6044);
nand_5 g05659(new_n6044, new_n1080, new_n6045);
nand_5 g05660(new_n6045, new_n1075, new_n6046);
nand_5 g05661(new_n6046, new_n1070, new_n6047);
nand_5 g05662(new_n6047, new_n1143, new_n6048);
nand_5 g05663(new_n6048, new_n1148, new_n6049);
nand_5 g05664(new_n6049, new_n1065, new_n6050);
nand_5 g05665(new_n6050, new_n1062, new_n6051);
nand_5 g05666(new_n6051, new_n1156, new_n6052);
nand_5 g05667(new_n6052, new_n1057, new_n6053);
nand_5 g05668(new_n6053, new_n1053, new_n6054_1);
nand_5 g05669(new_n6054_1, new_n1050, new_n6055);
nand_5 g05670(new_n6055, new_n1045, new_n6056);
nand_5 g05671(new_n6056, new_n1040, new_n6057);
nand_5 g05672(new_n6057, new_n1036, new_n6058);
nand_5 g05673(new_n6058, new_n1033, new_n6059);
nand_5 g05674(new_n6059, new_n1028, new_n6060);
nand_5 g05675(new_n6060, new_n1026, new_n6061);
nand_5 g05676(new_n6061, new_n1021, new_n6062);
nand_5 g05677(new_n6062, new_n1017, new_n6063);
nand_5 g05678(new_n6063, new_n1012, new_n6064);
nand_5 g05679(new_n6064, new_n1009, new_n6065);
nand_5 g05680(new_n6065, new_n1004, new_n6066);
nand_5 g05681(new_n6066, new_n1000, new_n6067);
nand_5 g05682(new_n6067, new_n995, new_n6068);
nand_5 g05683(new_n6068, new_n990, new_n6069);
nand_5 g05684(new_n6069, new_n985, new_n6070);
nand_5 g05685(new_n6070, new_n981, new_n6071);
nand_5 g05686(new_n6071, new_n1179, new_n6072);
nand_5 g05687(new_n6072, new_n976, new_n6073);
nand_5 g05688(new_n6073, new_n971, new_n6074);
nand_5 g05689(new_n6074, new_n966, new_n6075);
nand_5 g05690(new_n6075, new_n961, new_n6076);
nand_5 g05691(new_n6076, new_n957, new_n6077);
nand_5 g05692(new_n6077, new_n952, new_n6078);
nand_5 g05693(new_n6078, new_n948_1, new_n6079);
nand_5 g05694(new_n6079, new_n943, new_n6080);
nand_5 g05695(new_n6080, new_n941, new_n6081);
nand_5 g05696(new_n6081, new_n938, new_n6082);
nand_5 g05697(new_n6082, new_n936, new_n6083);
nand_5 g05698(new_n6083, new_n931, new_n6084);
nand_5 g05699(new_n6084, new_n927, new_n6085);
nand_5 g05700(new_n6085, new_n922, new_n6086);
nand_5 g05701(new_n6086, new_n917, new_n6087);
nand_5 g05702(new_n6087, new_n912, new_n6088);
nand_5 g05703(new_n6088, new_n907, new_n6089);
nand_5 g05704(new_n6089, new_n903, new_n6090);
nand_5 g05705(new_n6090, new_n2066, new_n6091);
nand_5 g05706(new_n6091, new_n2063, new_n6092);
nand_5 g05707(new_n6092, new_n2062, new_n6093);
nand_5 g05708(new_n6093, new_n2058, new_n6094);
nand_5 g05709(new_n6094, new_n2055, new_n6095);
nand_5 g05710(new_n6095, new_n2051, new_n6096);
nand_5 g05711(new_n6096, new_n2046, new_n6097);
nand_5 g05712(new_n6097, new_n2042, new_n6098);
nand_5 g05713(new_n6098, new_n2039, new_n6099);
nand_5 g05714(new_n6099, new_n2036, new_n6100);
nand_5 g05715(new_n6100, new_n2033, new_n6101);
nand_5 g05716(new_n6101, new_n2029, new_n6102);
nand_5 g05717(new_n6102, new_n2026, new_n6103);
nand_5 g05718(new_n6103, new_n2022, new_n6104);
nand_5 g05719(new_n6104, new_n2018, new_n6105);
nand_5 g05720(new_n6105, new_n1726, new_n6106);
nand_5 g05721(new_n6106, new_n1722, new_n6107);
nand_5 g05722(new_n6107, new_n1718, new_n6108);
nand_5 g05723(new_n6108, new_n1713, new_n6109);
nand_5 g05724(new_n6109, new_n1737, new_n6110);
nand_5 g05725(new_n6110, new_n1709, new_n6111);
nand_5 g05726(new_n6111, new_n1742, new_n6112);
nand_5 g05727(new_n6112, new_n1704, new_n6113);
nand_5 g05728(new_n6113, new_n1702_1, new_n6114_1);
nand_5 g05729(new_n6114_1, new_n1698, new_n6115);
nand_5 g05730(new_n6115, new_n1695, new_n6116);
nand_5 g05731(new_n6116, new_n1692, new_n6117);
nand_5 g05732(new_n6117, new_n1752, new_n6118);
nand_5 g05733(new_n6118, n13944, new_n6119);
nor_5  g05734(new_n6119, new_n1215, n5851);
not_4  g05735(new_n1319, new_n6121);
nand_5 g05736(new_n6121, new_n936, new_n6122);
nand_5 g05737(new_n6122, new_n931, new_n6123);
nand_5 g05738(new_n6123, new_n927, new_n6124);
nand_5 g05739(new_n6124, new_n922, new_n6125);
nand_5 g05740(new_n6125, new_n917, new_n6126);
nand_5 g05741(new_n6126, new_n912, new_n6127);
nand_5 g05742(new_n6127, new_n907, new_n6128);
nand_5 g05743(new_n6128, new_n903, new_n6129);
nand_5 g05744(new_n6129, new_n2066, new_n6130);
nand_5 g05745(new_n6130, new_n2063, new_n6131);
nand_5 g05746(new_n6131, new_n2062, new_n6132);
nand_5 g05747(new_n6132, new_n2058, new_n6133);
nand_5 g05748(new_n6133, new_n2055, new_n6134);
nand_5 g05749(new_n6134, new_n2051, new_n6135);
nand_5 g05750(new_n6135, new_n2046, new_n6136);
nand_5 g05751(new_n6136, new_n2042, new_n6137);
nand_5 g05752(new_n6137, new_n2039, new_n6138);
nand_5 g05753(new_n6138, new_n2036, new_n6139);
nand_5 g05754(new_n6139, new_n2033, new_n6140);
nand_5 g05755(new_n6140, new_n2029, new_n6141);
nand_5 g05756(new_n6141, new_n2026, new_n6142);
nand_5 g05757(new_n6142, new_n2022, new_n6143);
nand_5 g05758(new_n6143, new_n2018, new_n6144);
nand_5 g05759(new_n6144, new_n1726, new_n6145);
nand_5 g05760(new_n6145, new_n1722, new_n6146);
nand_5 g05761(new_n6146, new_n1718, new_n6147_1);
nand_5 g05762(new_n6147_1, new_n1713, new_n6148);
nand_5 g05763(new_n6148, new_n1737, new_n6149);
nand_5 g05764(new_n6149, new_n1709, new_n6150);
nand_5 g05765(new_n6150, new_n1742, new_n6151);
nand_5 g05766(new_n6151, new_n1704, new_n6152);
nand_5 g05767(new_n6152, new_n1702_1, new_n6153);
nand_5 g05768(new_n6153, new_n1698, new_n6154);
nand_5 g05769(new_n6154, new_n1695, new_n6155);
nand_5 g05770(new_n6155, new_n1692, new_n6156);
nand_5 g05771(new_n6156, new_n1752, new_n6157);
nand_5 g05772(new_n6157, new_n1688, new_n6158);
nand_5 g05773(new_n6158, new_n1685, new_n6159);
nand_5 g05774(new_n6159, new_n1680, new_n6160);
nand_5 g05775(new_n6160, new_n1676, new_n6161);
nand_5 g05776(new_n6161, new_n1672, new_n6162);
nand_5 g05777(new_n6162, new_n1669, new_n6163);
nand_5 g05778(new_n6163, new_n1666, new_n6164);
nand_5 g05779(new_n6164, new_n1663, new_n6165);
nand_5 g05780(new_n6165, new_n1658, new_n6166);
nand_5 g05781(new_n6166, new_n1653, new_n6167);
nand_5 g05782(new_n6167, new_n1651, new_n6168);
nand_5 g05783(new_n6168, new_n1649, new_n6169);
nand_5 g05784(new_n6169, new_n1646, new_n6170);
nand_5 g05785(new_n6170, new_n1643, new_n6171);
nand_5 g05786(new_n6171, new_n1641, new_n6172);
nand_5 g05787(new_n6172, new_n1638, new_n6173);
nand_5 g05788(new_n6173, new_n1635, new_n6174);
nand_5 g05789(new_n6174, new_n1632, new_n6175);
nand_5 g05790(new_n6175, new_n1628, new_n6176);
nand_5 g05791(new_n6176, new_n1625, new_n6177);
nand_5 g05792(new_n6177, new_n1621, new_n6178);
nand_5 g05793(new_n6178, new_n1618, new_n6179);
nand_5 g05794(new_n6179, new_n1778, new_n6180);
nand_5 g05795(new_n6180, new_n1782, new_n6181);
nand_5 g05796(new_n6181, new_n1614, new_n6182);
nand_5 g05797(new_n6182, new_n1611, new_n6183);
nand_5 g05798(new_n6183, new_n1789, new_n6184);
nand_5 g05799(new_n6184, new_n1608, new_n6185);
nand_5 g05800(new_n6185, new_n1605, new_n6186);
nand_5 g05801(new_n6186, new_n1795, new_n6187);
nand_5 g05802(new_n6187, new_n1799, new_n6188);
nand_5 g05803(new_n6188, new_n1602, new_n6189);
nand_5 g05804(new_n6189, new_n1599, new_n6190);
nand_5 g05805(new_n6190, new_n1596, new_n6191);
nand_5 g05806(new_n6191, new_n1593, new_n6192);
nand_5 g05807(new_n6192, new_n1806, new_n6193);
nand_5 g05808(new_n6193, new_n1589, new_n6194);
nand_5 g05809(new_n6194, new_n1586, new_n6195);
nand_5 g05810(new_n6195, new_n1583, new_n6196);
nand_5 g05811(new_n6196, new_n1580, new_n6197);
nand_5 g05812(new_n6197, new_n1576, new_n6198_1);
nand_5 g05813(new_n6198_1, new_n1573, new_n6199);
nand_5 g05814(new_n6199, new_n1570, new_n6200);
nand_5 g05815(new_n6200, new_n1567, new_n6201);
nand_5 g05816(new_n6201, new_n1564, new_n6202);
nand_5 g05817(new_n6202, new_n1561, new_n6203);
nand_5 g05818(new_n6203, new_n1338, new_n6204);
nand_5 g05819(new_n6204, new_n1331, new_n6205);
nand_5 g05820(new_n6205, n4659, new_n6206);
nor_5  g05821(new_n6206, new_n1323, n5987);
nand_5 g05822(new_n1621, new_n1622, new_n6208);
nand_5 g05823(new_n6208, new_n1618, new_n6209);
nand_5 g05824(new_n6209, new_n1778, new_n6210);
nand_5 g05825(new_n6210, new_n1782, new_n6211);
nand_5 g05826(new_n6211, new_n1614, new_n6212);
nand_5 g05827(new_n6212, new_n1611, new_n6213);
nand_5 g05828(new_n6213, new_n1789, new_n6214);
nand_5 g05829(new_n6214, new_n1608, new_n6215);
nand_5 g05830(new_n6215, new_n1605, new_n6216);
nand_5 g05831(new_n6216, new_n1795, new_n6217);
nand_5 g05832(new_n6217, new_n1799, new_n6218);
nand_5 g05833(new_n6218, new_n1602, new_n6219);
nand_5 g05834(new_n6219, new_n1599, new_n6220);
nand_5 g05835(new_n6220, new_n1596, new_n6221);
nand_5 g05836(new_n6221, new_n1593, new_n6222);
nand_5 g05837(new_n6222, new_n1806, new_n6223);
nand_5 g05838(new_n6223, new_n1589, new_n6224);
nand_5 g05839(new_n6224, new_n1586, new_n6225);
nand_5 g05840(new_n6225, new_n1583, new_n6226);
nand_5 g05841(new_n6226, new_n1580, new_n6227);
nand_5 g05842(new_n6227, new_n1576, new_n6228);
nand_5 g05843(new_n6228, new_n1573, new_n6229);
nand_5 g05844(new_n6229, new_n1570, new_n6230);
nand_5 g05845(new_n6230, new_n1567, new_n6231);
nand_5 g05846(new_n6231, new_n1564, new_n6232);
nand_5 g05847(new_n6232, new_n1561, new_n6233);
nand_5 g05848(new_n6233, new_n1338, new_n6234);
nand_5 g05849(new_n6234, new_n1331, new_n6235);
nand_5 g05850(new_n6235, new_n1326, new_n6236);
nand_5 g05851(new_n6236, new_n1321, new_n6237);
nand_5 g05852(new_n6237, new_n1318, new_n6238);
nand_5 g05853(new_n6238, new_n1315, new_n6239);
nand_5 g05854(new_n6239, new_n1312, new_n6240);
nand_5 g05855(new_n6240, new_n1309, new_n6241);
nand_5 g05856(new_n6241, new_n1307, new_n6242);
nand_5 g05857(new_n6242, new_n1304, new_n6243);
nand_5 g05858(new_n6243, new_n1300, new_n6244);
nand_5 g05859(new_n6244, new_n1297, new_n6245);
nand_5 g05860(new_n6245, new_n1294, new_n6246);
nand_5 g05861(new_n6246, new_n1355, new_n6247);
nand_5 g05862(new_n6247, new_n1291, new_n6248);
nand_5 g05863(new_n6248, new_n1288, new_n6249);
nand_5 g05864(new_n6249, new_n1283, new_n6250);
nand_5 g05865(new_n6250, new_n1363, new_n6251_1);
nand_5 g05866(new_n6251_1, new_n1280, new_n6252);
nand_5 g05867(new_n6252, new_n1370, new_n6253);
nand_5 g05868(new_n6253, new_n1373, new_n6254);
nand_5 g05869(new_n6254, new_n1277, new_n6255);
nand_5 g05870(new_n6255, new_n1272, new_n6256);
nand_5 g05871(new_n6256, new_n1269, new_n6257);
nand_5 g05872(new_n6257, new_n1380, new_n6258_1);
nand_5 g05873(new_n6258_1, new_n1264, new_n6259);
nand_5 g05874(new_n6259, new_n1259, new_n6260);
nand_5 g05875(new_n6260, new_n1388, new_n6261);
nand_5 g05876(new_n6261, new_n1392, new_n6262);
nand_5 g05877(new_n6262, new_n1256, new_n6263);
nand_5 g05878(new_n6263, new_n1252, new_n6264);
nand_5 g05879(new_n6264, new_n1249, new_n6265);
nand_5 g05880(new_n6265, new_n1244, new_n6266);
nand_5 g05881(new_n6266, new_n1240, new_n6267);
nand_5 g05882(new_n6267, new_n1234, new_n6268);
nand_5 g05883(new_n6268, new_n1231, new_n6269);
nand_5 g05884(new_n6269, new_n1227, new_n6270_1);
nand_5 g05885(new_n6270_1, new_n1407, new_n6271);
nand_5 g05886(new_n6271, new_n1223, new_n6272);
nand_5 g05887(new_n6272, new_n1218, new_n6273);
nand_5 g05888(new_n6273, new_n1213, new_n6274);
nand_5 g05889(new_n6274, new_n1210, new_n6275_1);
nand_5 g05890(new_n6275_1, new_n1206, new_n6276);
nand_5 g05891(new_n6276, new_n1418, new_n6277);
nand_5 g05892(new_n6277, new_n1422, new_n6278);
nand_5 g05893(new_n6278, new_n1428, new_n6279);
nand_5 g05894(new_n6279, new_n1203, new_n6280);
nand_5 g05895(new_n6280, new_n1433, new_n6281);
nand_5 g05896(new_n6281, new_n581, new_n6282);
nand_5 g05897(new_n6282, new_n574, new_n6283);
nand_5 g05898(new_n6283, new_n568, new_n6284);
nand_5 g05899(new_n6284, new_n589, new_n6285);
nand_5 g05900(new_n6285, new_n595, new_n6286);
nand_5 g05901(new_n6286, new_n601, new_n6287);
nand_5 g05902(new_n6287, new_n563, new_n6288);
nand_5 g05903(new_n6288, new_n608, new_n6289);
nand_5 g05904(new_n6289, new_n558, new_n6290);
nand_5 g05905(new_n6290, new_n615, new_n6291);
nand_5 g05906(new_n6291, n5225, new_n6292);
nor_5  g05907(new_n6292, new_n550, n6012);
nand_5 g05908(new_n1257, new_n818, new_n6294);
nand_5 g05909(new_n6294, new_n1388, new_n6295);
nand_5 g05910(new_n6295, new_n1392, new_n6296);
nand_5 g05911(new_n6296, new_n1256, new_n6297);
nand_5 g05912(new_n6297, new_n1252, new_n6298);
nand_5 g05913(new_n6298, new_n1249, new_n6299);
nand_5 g05914(new_n6299, new_n1244, new_n6300);
nand_5 g05915(new_n6300, new_n1240, new_n6301);
nand_5 g05916(new_n6301, new_n1234, new_n6302);
nand_5 g05917(new_n6302, new_n1231, new_n6303);
nand_5 g05918(new_n6303, new_n1227, new_n6304);
nand_5 g05919(new_n6304, new_n1407, new_n6305);
nand_5 g05920(new_n6305, new_n1223, new_n6306);
nand_5 g05921(new_n6306, new_n1218, new_n6307);
nand_5 g05922(new_n6307, new_n1213, new_n6308);
nand_5 g05923(new_n6308, new_n1210, new_n6309);
nand_5 g05924(new_n6309, new_n1206, new_n6310);
nand_5 g05925(new_n6310, new_n1418, new_n6311);
nand_5 g05926(new_n6311, new_n1422, new_n6312);
nand_5 g05927(new_n6312, new_n1428, new_n6313);
nand_5 g05928(new_n6313, new_n1203, new_n6314_1);
nand_5 g05929(new_n6314_1, new_n1433, new_n6315);
nand_5 g05930(new_n6315, new_n581, new_n6316);
nand_5 g05931(new_n6316, new_n574, new_n6317);
nand_5 g05932(new_n6317, new_n568, new_n6318);
nand_5 g05933(new_n6318, new_n589, new_n6319);
nand_5 g05934(new_n6319, new_n595, new_n6320);
nand_5 g05935(new_n6320, new_n601, new_n6321);
nand_5 g05936(new_n6321, new_n563, new_n6322);
nand_5 g05937(new_n6322, new_n608, new_n6323);
nand_5 g05938(new_n6323, new_n558, new_n6324);
nand_5 g05939(new_n6324, new_n615, new_n6325);
nand_5 g05940(new_n6325, new_n553, new_n6326);
nand_5 g05941(new_n6326, new_n622, new_n6327);
nand_5 g05942(new_n6327, new_n628, new_n6328);
nand_5 g05943(new_n6328, new_n548, new_n6329);
nand_5 g05944(new_n6329, new_n543_1, new_n6330);
nand_5 g05945(new_n6330, new_n636, new_n6331);
nand_5 g05946(new_n6331, new_n642, new_n6332);
nand_5 g05947(new_n6332, new_n538, new_n6333);
nand_5 g05948(new_n6333, new_n533, new_n6334);
nand_5 g05949(new_n6334, new_n650_1, new_n6335);
nand_5 g05950(new_n6335, new_n528, new_n6336);
nand_5 g05951(new_n6336, new_n523, new_n6337);
nand_5 g05952(new_n6337, new_n518, new_n6338);
nand_5 g05953(new_n6338, new_n659, new_n6339);
nand_5 g05954(new_n6339, new_n665, new_n6340);
nand_5 g05955(new_n6340, new_n672, new_n6341);
nand_5 g05956(new_n6341, new_n513, new_n6342);
nand_5 g05957(new_n6342, new_n679, new_n6343);
nand_5 g05958(new_n6343, new_n685, new_n6344);
nand_5 g05959(new_n6344, new_n691, new_n6345);
nand_5 g05960(new_n6345, new_n508, new_n6346);
nand_5 g05961(new_n6346, new_n698, new_n6347);
nand_5 g05962(new_n6347, new_n503, new_n6348);
nand_5 g05963(new_n6348, new_n704, new_n6349);
nand_5 g05964(new_n6349, new_n498_1, new_n6350);
nand_5 g05965(new_n6350, new_n711, new_n6351);
nand_5 g05966(new_n6351, new_n493, new_n6352);
nand_5 g05967(new_n6352, new_n718, new_n6353);
nand_5 g05968(new_n6353, new_n488, new_n6354);
nand_5 g05969(new_n6354, new_n725, new_n6355);
nand_5 g05970(new_n6355, new_n483, new_n6356);
nand_5 g05971(new_n6356, new_n732, new_n6357);
nand_5 g05972(new_n6357, new_n478, new_n6358);
nand_5 g05973(new_n6358, new_n739, new_n6359);
nand_5 g05974(new_n6359, new_n745, new_n6360);
nand_5 g05975(new_n6360, new_n751, new_n6361);
nand_5 g05976(new_n6361, new_n473, new_n6362_1);
nand_5 g05977(new_n6362_1, new_n758, new_n6363);
nand_5 g05978(new_n6363, new_n764, new_n6364);
nand_5 g05979(new_n6364, new_n770, new_n6365);
nand_5 g05980(new_n6365, new_n468, new_n6366);
nand_5 g05981(new_n6366, new_n777, new_n6367);
nand_5 g05982(new_n6367, new_n783, new_n6368);
nand_5 g05983(new_n6368, new_n789, new_n6369);
nand_5 g05984(new_n6369, new_n463, new_n6370);
nand_5 g05985(new_n6370, new_n796, new_n6371);
nand_5 g05986(new_n6371, new_n458, new_n6372);
nand_5 g05987(new_n6372, new_n453, new_n6373);
nand_5 g05988(new_n6373, new_n447, new_n6374);
nand_5 g05989(new_n6374, new_n805, new_n6375);
nand_5 g05990(new_n6375, new_n811, new_n6376);
nand_5 g05991(new_n6376, new_n442, new_n6377);
nand_5 g05992(new_n6377, n3673, new_n6378);
nor_5  g05993(new_n6378, new_n434, n6198);
nand_5 g05994(new_n1734, new_n1709, new_n6380);
nand_5 g05995(new_n6380, new_n1742, new_n6381);
nand_5 g05996(new_n6381, new_n1704, new_n6382);
nand_5 g05997(new_n6382, new_n1702_1, new_n6383);
nand_5 g05998(new_n6383, new_n1698, new_n6384);
nand_5 g05999(new_n6384, new_n1695, new_n6385);
nand_5 g06000(new_n6385, new_n1692, new_n6386);
nand_5 g06001(new_n6386, new_n1752, new_n6387);
nand_5 g06002(new_n6387, new_n1688, new_n6388);
nand_5 g06003(new_n6388, new_n1685, new_n6389);
nand_5 g06004(new_n6389, new_n1680, new_n6390);
nand_5 g06005(new_n6390, new_n1676, new_n6391);
nand_5 g06006(new_n6391, new_n1672, new_n6392);
nand_5 g06007(new_n6392, new_n1669, new_n6393);
nand_5 g06008(new_n6393, new_n1666, new_n6394);
nand_5 g06009(new_n6394, new_n1663, new_n6395);
nand_5 g06010(new_n6395, new_n1658, new_n6396);
nand_5 g06011(new_n6396, new_n1653, new_n6397);
nand_5 g06012(new_n6397, new_n1651, new_n6398);
nand_5 g06013(new_n6398, new_n1649, new_n6399);
nand_5 g06014(new_n6399, new_n1646, new_n6400);
nand_5 g06015(new_n6400, new_n1643, new_n6401);
nand_5 g06016(new_n6401, new_n1641, new_n6402);
nand_5 g06017(new_n6402, new_n1638, new_n6403);
nand_5 g06018(new_n6403, new_n1635, new_n6404);
nand_5 g06019(new_n6404, new_n1632, new_n6405);
nand_5 g06020(new_n6405, new_n1628, new_n6406);
nand_5 g06021(new_n6406, new_n1625, new_n6407);
nand_5 g06022(new_n6407, new_n1621, new_n6408);
nand_5 g06023(new_n6408, new_n1618, new_n6409);
nand_5 g06024(new_n6409, new_n1778, new_n6410);
nand_5 g06025(new_n6410, new_n1782, new_n6411);
nand_5 g06026(new_n6411, new_n1614, new_n6412);
nand_5 g06027(new_n6412, new_n1611, new_n6413);
nand_5 g06028(new_n6413, new_n1789, new_n6414);
nand_5 g06029(new_n6414, new_n1608, new_n6415);
nand_5 g06030(new_n6415, new_n1605, new_n6416);
nand_5 g06031(new_n6416, new_n1795, new_n6417);
nand_5 g06032(new_n6417, new_n1799, new_n6418);
nand_5 g06033(new_n6418, new_n1602, new_n6419);
nand_5 g06034(new_n6419, new_n1599, new_n6420);
nand_5 g06035(new_n6420, new_n1596, new_n6421);
nand_5 g06036(new_n6421, new_n1593, new_n6422);
nand_5 g06037(new_n6422, new_n1806, new_n6423);
nand_5 g06038(new_n6423, new_n1589, new_n6424);
nand_5 g06039(new_n6424, new_n1586, new_n6425);
nand_5 g06040(new_n6425, new_n1583, new_n6426);
nand_5 g06041(new_n6426, new_n1580, new_n6427);
nand_5 g06042(new_n6427, new_n1576, new_n6428);
nand_5 g06043(new_n6428, new_n1573, new_n6429);
nand_5 g06044(new_n6429, new_n1570, new_n6430);
nand_5 g06045(new_n6430, new_n1567, new_n6431);
nand_5 g06046(new_n6431, new_n1564, new_n6432);
nand_5 g06047(new_n6432, new_n1561, new_n6433);
nand_5 g06048(new_n6433, new_n1338, new_n6434);
nand_5 g06049(new_n6434, new_n1331, new_n6435);
nand_5 g06050(new_n6435, new_n1326, new_n6436_1);
nand_5 g06051(new_n6436_1, new_n1321, new_n6437);
nand_5 g06052(new_n6437, new_n1318, new_n6438);
nand_5 g06053(new_n6438, new_n1315, new_n6439);
nand_5 g06054(new_n6439, new_n1312, new_n6440);
nand_5 g06055(new_n6440, new_n1309, new_n6441);
nand_5 g06056(new_n6441, new_n1307, new_n6442);
nand_5 g06057(new_n6442, new_n1304, new_n6443);
nand_5 g06058(new_n6443, new_n1300, new_n6444);
nand_5 g06059(new_n6444, new_n1297, new_n6445);
nand_5 g06060(new_n6445, new_n1294, new_n6446);
nand_5 g06061(new_n6446, new_n1355, new_n6447);
nand_5 g06062(new_n6447, new_n1291, new_n6448);
nand_5 g06063(new_n6448, new_n1288, new_n6449);
nand_5 g06064(new_n6449, new_n1283, new_n6450);
nand_5 g06065(new_n6450, new_n1363, new_n6451);
nand_5 g06066(new_n6451, new_n1280, new_n6452);
nand_5 g06067(new_n6452, new_n1370, new_n6453);
nand_5 g06068(new_n6453, new_n1373, new_n6454);
nand_5 g06069(new_n6454, new_n1277, new_n6455);
nand_5 g06070(new_n6455, new_n1272, new_n6456);
nand_5 g06071(new_n6456, new_n1269, new_n6457);
nand_5 g06072(new_n6457, new_n1380, new_n6458);
nand_5 g06073(new_n6458, new_n1264, new_n6459);
nand_5 g06074(new_n6459, new_n1259, new_n6460_1);
nand_5 g06075(new_n6460_1, new_n1388, new_n6461);
nand_5 g06076(new_n6461, new_n1392, new_n6462);
nand_5 g06077(new_n6462, new_n1256, new_n6463);
nand_5 g06078(new_n6463, n666, new_n6464);
nor_5  g06079(new_n6464, new_n825, n6275);
not_4  g06080(new_n2060, new_n6466);
not_4  g06081(new_n2056, new_n6467);
nand_5 g06082(new_n6467, new_n783, new_n6468);
nand_5 g06083(new_n6468, new_n789, new_n6469);
nand_5 g06084(new_n6469, new_n463, new_n6470);
nand_5 g06085(new_n6470, new_n796, new_n6471);
nand_5 g06086(new_n6471, new_n458, new_n6472);
nand_5 g06087(new_n6472, new_n453, new_n6473);
nand_5 g06088(new_n6473, new_n447, new_n6474);
nand_5 g06089(new_n6474, new_n805, new_n6475);
nand_5 g06090(new_n6475, new_n811, new_n6476);
nand_5 g06091(new_n6476, new_n442, new_n6477);
nand_5 g06092(new_n6477, new_n437, new_n6478);
nand_5 g06093(new_n6478, new_n819, new_n6479);
nand_5 g06094(new_n6479, new_n432, new_n6480_1);
nand_5 g06095(new_n6480_1, new_n427_1, new_n6481);
nand_5 g06096(new_n6481, new_n422, new_n6482);
nand_5 g06097(new_n6482, new_n828, new_n6483);
nand_5 g06098(new_n6483, new_n834, new_n6484);
nand_5 g06099(new_n6484, new_n840, new_n6485);
nand_5 g06100(new_n6485, new_n417, new_n6486);
nand_5 g06101(new_n6486, new_n847, new_n6487);
nand_5 g06102(new_n6487, new_n853, new_n6488);
nand_5 g06103(new_n6488, new_n859, new_n6489);
nand_5 g06104(new_n6489, new_n412, new_n6490);
nand_5 g06105(new_n6490, new_n866, new_n6491);
nand_5 g06106(new_n6491, new_n872, new_n6492);
nand_5 g06107(new_n6492, new_n878, new_n6493);
nand_5 g06108(new_n6493, new_n407, new_n6494);
nand_5 g06109(new_n6494, new_n885, new_n6495);
nand_5 g06110(new_n6495, new_n402, new_n6496);
nand_5 g06111(new_n6496, new_n397, new_n6497);
nand_5 g06112(new_n6497, new_n392, new_n6498);
nand_5 g06113(new_n6498, new_n894, new_n6499);
nand_5 g06114(new_n6499, new_n1087, new_n6500);
nand_5 g06115(new_n6500, new_n1129, new_n6501);
nand_5 g06116(new_n6501, new_n1084, new_n6502);
nand_5 g06117(new_n6502, new_n1134, new_n6503);
nand_5 g06118(new_n6503, new_n1080, new_n6504);
nand_5 g06119(new_n6504, new_n1075, new_n6505);
nand_5 g06120(new_n6505, new_n1070, new_n6506);
nand_5 g06121(new_n6506, new_n1143, new_n6507);
nand_5 g06122(new_n6507, new_n1148, new_n6508);
nand_5 g06123(new_n6508, new_n1065, new_n6509);
nand_5 g06124(new_n6509, new_n1062, new_n6510);
nand_5 g06125(new_n6510, new_n1156, new_n6511);
nand_5 g06126(new_n6511, new_n1057, new_n6512);
nand_5 g06127(new_n6512, new_n1053, new_n6513);
nand_5 g06128(new_n6513, new_n1050, new_n6514);
nand_5 g06129(new_n6514, new_n1045, new_n6515);
nand_5 g06130(new_n6515, new_n1040, new_n6516);
nand_5 g06131(new_n6516, new_n1036, new_n6517_1);
nand_5 g06132(new_n6517_1, new_n1033, new_n6518);
nand_5 g06133(new_n6518, new_n1028, new_n6519);
nand_5 g06134(new_n6519, new_n1026, new_n6520);
nand_5 g06135(new_n6520, new_n1021, new_n6521);
nand_5 g06136(new_n6521, new_n1017, new_n6522);
nand_5 g06137(new_n6522, new_n1012, new_n6523);
nand_5 g06138(new_n6523, new_n1009, new_n6524);
nand_5 g06139(new_n6524, new_n1004, new_n6525);
nand_5 g06140(new_n6525, new_n1000, new_n6526);
nand_5 g06141(new_n6526, new_n995, new_n6527);
nand_5 g06142(new_n6527, new_n990, new_n6528);
nand_5 g06143(new_n6528, new_n985, new_n6529);
nand_5 g06144(new_n6529, new_n981, new_n6530);
nand_5 g06145(new_n6530, new_n1179, new_n6531);
nand_5 g06146(new_n6531, new_n976, new_n6532);
nand_5 g06147(new_n6532, new_n971, new_n6533);
nand_5 g06148(new_n6533, new_n966, new_n6534);
nand_5 g06149(new_n6534, new_n961, new_n6535);
nand_5 g06150(new_n6535, new_n957, new_n6536);
nand_5 g06151(new_n6536, new_n952, new_n6537);
nand_5 g06152(new_n6537, new_n948_1, new_n6538);
nand_5 g06153(new_n6538, new_n943, new_n6539);
nand_5 g06154(new_n6539, new_n941, new_n6540);
nand_5 g06155(new_n6540, new_n938, new_n6541);
nand_5 g06156(new_n6541, new_n936, new_n6542);
nand_5 g06157(new_n6542, new_n931, new_n6543);
nand_5 g06158(new_n6543, new_n927, new_n6544);
nand_5 g06159(new_n6544, new_n922, new_n6545);
nand_5 g06160(new_n6545, new_n917, new_n6546);
nand_5 g06161(new_n6546, new_n912, new_n6547);
nand_5 g06162(new_n6547, new_n907, new_n6548);
nand_5 g06163(new_n6548, new_n903, new_n6549);
nand_5 g06164(new_n6549, new_n2066, new_n6550);
nand_5 g06165(new_n6550, new_n2063, new_n6551);
nand_5 g06166(new_n6551, n6999, new_n6552);
nor_5  g06167(new_n6552, new_n6466, n6314);
nand_5 g06168(new_n1587, new_n678, new_n6554);
nand_5 g06169(new_n6554, new_n1586, new_n6555_1);
nand_5 g06170(new_n6555_1, new_n1583, new_n6556);
nand_5 g06171(new_n6556, new_n1580, new_n6557);
nand_5 g06172(new_n6557, new_n1576, new_n6558);
nand_5 g06173(new_n6558, new_n1573, new_n6559);
nand_5 g06174(new_n6559, new_n1570, new_n6560);
nand_5 g06175(new_n6560, new_n1567, new_n6561);
nand_5 g06176(new_n6561, new_n1564, new_n6562);
nand_5 g06177(new_n6562, new_n1561, new_n6563);
nand_5 g06178(new_n6563, new_n1338, new_n6564);
nand_5 g06179(new_n6564, new_n1331, new_n6565);
nand_5 g06180(new_n6565, new_n1326, new_n6566);
nand_5 g06181(new_n6566, new_n1321, new_n6567);
nand_5 g06182(new_n6567, new_n1318, new_n6568);
nand_5 g06183(new_n6568, new_n1315, new_n6569);
nand_5 g06184(new_n6569, new_n1312, new_n6570);
nand_5 g06185(new_n6570, new_n1309, new_n6571);
nand_5 g06186(new_n6571, new_n1307, new_n6572);
nand_5 g06187(new_n6572, new_n1304, new_n6573);
nand_5 g06188(new_n6573, new_n1300, new_n6574);
nand_5 g06189(new_n6574, new_n1297, new_n6575);
nand_5 g06190(new_n6575, new_n1294, new_n6576);
nand_5 g06191(new_n6576, new_n1355, new_n6577);
nand_5 g06192(new_n6577, new_n1291, new_n6578);
nand_5 g06193(new_n6578, new_n1288, new_n6579);
nand_5 g06194(new_n6579, new_n1283, new_n6580);
nand_5 g06195(new_n6580, new_n1363, new_n6581);
nand_5 g06196(new_n6581, new_n1280, new_n6582);
nand_5 g06197(new_n6582, new_n1370, new_n6583);
nand_5 g06198(new_n6583, new_n1373, new_n6584);
nand_5 g06199(new_n6584, new_n1277, new_n6585);
nand_5 g06200(new_n6585, new_n1272, new_n6586_1);
nand_5 g06201(new_n6586_1, new_n1269, new_n6587);
nand_5 g06202(new_n6587, new_n1380, new_n6588);
nand_5 g06203(new_n6588, new_n1264, new_n6589);
nand_5 g06204(new_n6589, new_n1259, new_n6590);
nand_5 g06205(new_n6590, new_n1388, new_n6591);
nand_5 g06206(new_n6591, new_n1392, new_n6592);
nand_5 g06207(new_n6592, new_n1256, new_n6593);
nand_5 g06208(new_n6593, new_n1252, new_n6594);
nand_5 g06209(new_n6594, new_n1249, new_n6595);
nand_5 g06210(new_n6595, new_n1244, new_n6596);
nand_5 g06211(new_n6596, new_n1240, new_n6597);
nand_5 g06212(new_n6597, new_n1234, new_n6598);
nand_5 g06213(new_n6598, new_n1231, new_n6599);
nand_5 g06214(new_n6599, new_n1227, new_n6600);
nand_5 g06215(new_n6600, new_n1407, new_n6601);
nand_5 g06216(new_n6601, new_n1223, new_n6602);
nand_5 g06217(new_n6602, new_n1218, new_n6603);
nand_5 g06218(new_n6603, new_n1213, new_n6604);
nand_5 g06219(new_n6604, new_n1210, new_n6605);
nand_5 g06220(new_n6605, new_n1206, new_n6606);
nand_5 g06221(new_n6606, new_n1418, new_n6607);
nand_5 g06222(new_n6607, new_n1422, new_n6608);
nand_5 g06223(new_n6608, new_n1428, new_n6609);
nand_5 g06224(new_n6609, new_n1203, new_n6610);
nand_5 g06225(new_n6610, new_n1433, new_n6611);
nand_5 g06226(new_n6611, new_n581, new_n6612);
nand_5 g06227(new_n6612, new_n574, new_n6613);
nand_5 g06228(new_n6613, new_n568, new_n6614);
nand_5 g06229(new_n6614, new_n589, new_n6615);
nand_5 g06230(new_n6615, new_n595, new_n6616);
nand_5 g06231(new_n6616, new_n601, new_n6617);
nand_5 g06232(new_n6617, new_n563, new_n6618);
nand_5 g06233(new_n6618, new_n608, new_n6619);
nand_5 g06234(new_n6619, new_n558, new_n6620);
nand_5 g06235(new_n6620, new_n615, new_n6621);
nand_5 g06236(new_n6621, new_n553, new_n6622);
nand_5 g06237(new_n6622, new_n622, new_n6623);
nand_5 g06238(new_n6623, new_n628, new_n6624);
nand_5 g06239(new_n6624, new_n548, new_n6625);
nand_5 g06240(new_n6625, new_n543_1, new_n6626);
nand_5 g06241(new_n6626, new_n636, new_n6627);
nand_5 g06242(new_n6627, new_n642, new_n6628);
nand_5 g06243(new_n6628, new_n538, new_n6629);
nand_5 g06244(new_n6629, new_n533, new_n6630);
nand_5 g06245(new_n6630, new_n650_1, new_n6631);
nand_5 g06246(new_n6631, new_n528, new_n6632);
nand_5 g06247(new_n6632, new_n523, new_n6633);
nand_5 g06248(new_n6633, new_n518, new_n6634);
nand_5 g06249(new_n6634, new_n659, new_n6635);
nand_5 g06250(new_n6635, new_n665, new_n6636);
nand_5 g06251(new_n6636, new_n672, new_n6637);
nand_5 g06252(new_n6637, n3506, new_n6638);
nor_5  g06253(new_n6638, new_n510, n6682);
nand_5 g06254(new_n1289, new_n776, new_n6640);
nand_5 g06255(new_n6640, new_n1288, new_n6641);
nand_5 g06256(new_n6641, new_n1283, new_n6642);
nand_5 g06257(new_n6642, new_n1363, new_n6643);
nand_5 g06258(new_n6643, new_n1280, new_n6644);
nand_5 g06259(new_n6644, new_n1370, new_n6645);
nand_5 g06260(new_n6645, new_n1373, new_n6646);
nand_5 g06261(new_n6646, new_n1277, new_n6647);
nand_5 g06262(new_n6647, new_n1272, new_n6648);
nand_5 g06263(new_n6648, new_n1269, new_n6649);
nand_5 g06264(new_n6649, new_n1380, new_n6650);
nand_5 g06265(new_n6650, new_n1264, new_n6651);
nand_5 g06266(new_n6651, new_n1259, new_n6652);
nand_5 g06267(new_n6652, new_n1388, new_n6653);
nand_5 g06268(new_n6653, new_n1392, new_n6654);
nand_5 g06269(new_n6654, new_n1256, new_n6655);
nand_5 g06270(new_n6655, new_n1252, new_n6656);
nand_5 g06271(new_n6656, new_n1249, new_n6657);
nand_5 g06272(new_n6657, new_n1244, new_n6658);
nand_5 g06273(new_n6658, new_n1240, new_n6659);
nand_5 g06274(new_n6659, new_n1234, new_n6660);
nand_5 g06275(new_n6660, new_n1231, new_n6661);
nand_5 g06276(new_n6661, new_n1227, new_n6662);
nand_5 g06277(new_n6662, new_n1407, new_n6663);
nand_5 g06278(new_n6663, new_n1223, new_n6664);
nand_5 g06279(new_n6664, new_n1218, new_n6665);
nand_5 g06280(new_n6665, new_n1213, new_n6666);
nand_5 g06281(new_n6666, new_n1210, new_n6667);
nand_5 g06282(new_n6667, new_n1206, new_n6668);
nand_5 g06283(new_n6668, new_n1418, new_n6669);
nand_5 g06284(new_n6669, new_n1422, new_n6670);
nand_5 g06285(new_n6670, new_n1428, new_n6671);
nand_5 g06286(new_n6671, new_n1203, new_n6672);
nand_5 g06287(new_n6672, new_n1433, new_n6673);
nand_5 g06288(new_n6673, new_n581, new_n6674);
nand_5 g06289(new_n6674, new_n574, new_n6675);
nand_5 g06290(new_n6675, new_n568, new_n6676);
nand_5 g06291(new_n6676, new_n589, new_n6677);
nand_5 g06292(new_n6677, new_n595, new_n6678);
nand_5 g06293(new_n6678, new_n601, new_n6679);
nand_5 g06294(new_n6679, new_n563, new_n6680_1);
nand_5 g06295(new_n6680_1, new_n608, new_n6681);
nand_5 g06296(new_n6681, new_n558, new_n6682_1);
nand_5 g06297(new_n6682_1, new_n615, new_n6683);
nand_5 g06298(new_n6683, new_n553, new_n6684);
nand_5 g06299(new_n6684, new_n622, new_n6685);
nand_5 g06300(new_n6685, new_n628, new_n6686);
nand_5 g06301(new_n6686, new_n548, new_n6687);
nand_5 g06302(new_n6687, new_n543_1, new_n6688);
nand_5 g06303(new_n6688, new_n636, new_n6689);
nand_5 g06304(new_n6689, new_n642, new_n6690);
nand_5 g06305(new_n6690, new_n538, new_n6691);
nand_5 g06306(new_n6691, new_n533, new_n6692);
nand_5 g06307(new_n6692, new_n650_1, new_n6693_1);
nand_5 g06308(new_n6693_1, new_n528, new_n6694);
nand_5 g06309(new_n6694, new_n523, new_n6695);
nand_5 g06310(new_n6695, new_n518, new_n6696_1);
nand_5 g06311(new_n6696_1, new_n659, new_n6697);
nand_5 g06312(new_n6697, new_n665, new_n6698);
nand_5 g06313(new_n6698, new_n672, new_n6699);
nand_5 g06314(new_n6699, new_n513, new_n6700);
nand_5 g06315(new_n6700, new_n679, new_n6701);
nand_5 g06316(new_n6701, new_n685, new_n6702);
nand_5 g06317(new_n6702, new_n691, new_n6703_1);
nand_5 g06318(new_n6703_1, new_n508, new_n6704);
nand_5 g06319(new_n6704, new_n698, new_n6705);
nand_5 g06320(new_n6705, new_n503, new_n6706);
nand_5 g06321(new_n6706, new_n704, new_n6707);
nand_5 g06322(new_n6707, new_n498_1, new_n6708);
nand_5 g06323(new_n6708, new_n711, new_n6709);
nand_5 g06324(new_n6709, new_n493, new_n6710);
nand_5 g06325(new_n6710, new_n718, new_n6711);
nand_5 g06326(new_n6711, new_n488, new_n6712);
nand_5 g06327(new_n6712, new_n725, new_n6713);
nand_5 g06328(new_n6713, new_n483, new_n6714);
nand_5 g06329(new_n6714, new_n732, new_n6715);
nand_5 g06330(new_n6715, new_n478, new_n6716);
nand_5 g06331(new_n6716, new_n739, new_n6717);
nand_5 g06332(new_n6717, new_n745, new_n6718);
nand_5 g06333(new_n6718, new_n751, new_n6719);
nand_5 g06334(new_n6719, new_n473, new_n6720);
nand_5 g06335(new_n6720, new_n758, new_n6721);
nand_5 g06336(new_n6721, new_n764, new_n6722);
nand_5 g06337(new_n6722, new_n770, new_n6723);
nand_5 g06338(new_n6723, n6517, new_n6724);
nor_5  g06339(new_n6724, new_n465, n6696);
nand_5 g06340(new_n1566, new_n955, new_n6726);
nand_5 g06341(new_n6726, new_n952, new_n6727);
nand_5 g06342(new_n6727, new_n948_1, new_n6728);
nand_5 g06343(new_n6728, new_n943, new_n6729);
nand_5 g06344(new_n6729, new_n941, new_n6730);
nand_5 g06345(new_n6730, new_n938, new_n6731);
nand_5 g06346(new_n6731, new_n936, new_n6732);
nand_5 g06347(new_n6732, new_n931, new_n6733);
nand_5 g06348(new_n6733, new_n927, new_n6734);
nand_5 g06349(new_n6734, new_n922, new_n6735);
nand_5 g06350(new_n6735, new_n917, new_n6736);
nand_5 g06351(new_n6736, new_n912, new_n6737);
nand_5 g06352(new_n6737, new_n907, new_n6738);
nand_5 g06353(new_n6738, new_n903, new_n6739);
nand_5 g06354(new_n6739, new_n2066, new_n6740);
nand_5 g06355(new_n6740, new_n2063, new_n6741);
nand_5 g06356(new_n6741, new_n2062, new_n6742);
nand_5 g06357(new_n6742, new_n2058, new_n6743);
nand_5 g06358(new_n6743, new_n2055, new_n6744);
nand_5 g06359(new_n6744, new_n2051, new_n6745);
nand_5 g06360(new_n6745, new_n2046, new_n6746);
nand_5 g06361(new_n6746, new_n2042, new_n6747);
nand_5 g06362(new_n6747, new_n2039, new_n6748);
nand_5 g06363(new_n6748, new_n2036, new_n6749);
nand_5 g06364(new_n6749, new_n2033, new_n6750);
nand_5 g06365(new_n6750, new_n2029, new_n6751);
nand_5 g06366(new_n6751, new_n2026, new_n6752);
nand_5 g06367(new_n6752, new_n2022, new_n6753);
nand_5 g06368(new_n6753, new_n2018, new_n6754);
nand_5 g06369(new_n6754, new_n1726, new_n6755);
nand_5 g06370(new_n6755, new_n1722, new_n6756);
nand_5 g06371(new_n6756, new_n1718, new_n6757);
nand_5 g06372(new_n6757, new_n1713, new_n6758_1);
nand_5 g06373(new_n6758_1, new_n1737, new_n6759);
nand_5 g06374(new_n6759, new_n1709, new_n6760);
nand_5 g06375(new_n6760, new_n1742, new_n6761);
nand_5 g06376(new_n6761, new_n1704, new_n6762);
nand_5 g06377(new_n6762, new_n1702_1, new_n6763);
nand_5 g06378(new_n6763, new_n1698, new_n6764);
nand_5 g06379(new_n6764, new_n1695, new_n6765);
nand_5 g06380(new_n6765, new_n1692, new_n6766);
nand_5 g06381(new_n6766, new_n1752, new_n6767);
nand_5 g06382(new_n6767, new_n1688, new_n6768);
nand_5 g06383(new_n6768, new_n1685, new_n6769);
nand_5 g06384(new_n6769, new_n1680, new_n6770);
nand_5 g06385(new_n6770, new_n1676, new_n6771);
nand_5 g06386(new_n6771, new_n1672, new_n6772);
nand_5 g06387(new_n6772, new_n1669, new_n6773);
nand_5 g06388(new_n6773, new_n1666, new_n6774);
nand_5 g06389(new_n6774, new_n1663, new_n6775);
nand_5 g06390(new_n6775, new_n1658, new_n6776);
nand_5 g06391(new_n6776, new_n1653, new_n6777);
nand_5 g06392(new_n6777, new_n1651, new_n6778);
nand_5 g06393(new_n6778, new_n1649, new_n6779);
nand_5 g06394(new_n6779, new_n1646, new_n6780);
nand_5 g06395(new_n6780, new_n1643, new_n6781);
nand_5 g06396(new_n6781, new_n1641, new_n6782);
nand_5 g06397(new_n6782, new_n1638, new_n6783);
nand_5 g06398(new_n6783, new_n1635, new_n6784);
nand_5 g06399(new_n6784, new_n1632, new_n6785);
nand_5 g06400(new_n6785, new_n1628, new_n6786_1);
nand_5 g06401(new_n6786_1, new_n1625, new_n6787);
nand_5 g06402(new_n6787, new_n1621, new_n6788);
nand_5 g06403(new_n6788, new_n1618, new_n6789);
nand_5 g06404(new_n6789, new_n1778, new_n6790);
nand_5 g06405(new_n6790, new_n1782, new_n6791_1);
nand_5 g06406(new_n6791_1, new_n1614, new_n6792);
nand_5 g06407(new_n6792, new_n1611, new_n6793);
nand_5 g06408(new_n6793, new_n1789, new_n6794);
nand_5 g06409(new_n6794, new_n1608, new_n6795);
nand_5 g06410(new_n6795, new_n1605, new_n6796);
nand_5 g06411(new_n6796, new_n1795, new_n6797);
nand_5 g06412(new_n6797, new_n1799, new_n6798);
nand_5 g06413(new_n6798, new_n1602, new_n6799);
nand_5 g06414(new_n6799, new_n1599, new_n6800);
nand_5 g06415(new_n6800, new_n1596, new_n6801);
nand_5 g06416(new_n6801, new_n1593, new_n6802);
nand_5 g06417(new_n6802, new_n1806, new_n6803);
nand_5 g06418(new_n6803, new_n1589, new_n6804);
nand_5 g06419(new_n6804, new_n1586, new_n6805);
nand_5 g06420(new_n6805, new_n1583, new_n6806);
nand_5 g06421(new_n6806, new_n1580, new_n6807);
nand_5 g06422(new_n6807, new_n1576, new_n6808);
nand_5 g06423(new_n6808, new_n1573, new_n6809);
nand_5 g06424(new_n6809, n11875, new_n6810_1);
nor_5  g06425(new_n6810_1, new_n701, n6786);
nand_5 g06426(new_n2035, new_n445, new_n6812);
nand_5 g06427(new_n6812, new_n805, new_n6813);
nand_5 g06428(new_n6813, new_n811, new_n6814);
nand_5 g06429(new_n6814, new_n442, new_n6815);
nand_5 g06430(new_n6815, new_n437, new_n6816);
nand_5 g06431(new_n6816, new_n819, new_n6817);
nand_5 g06432(new_n6817, new_n432, new_n6818);
nand_5 g06433(new_n6818, new_n427_1, new_n6819);
nand_5 g06434(new_n6819, new_n422, new_n6820);
nand_5 g06435(new_n6820, new_n828, new_n6821);
nand_5 g06436(new_n6821, new_n834, new_n6822);
nand_5 g06437(new_n6822, new_n840, new_n6823);
nand_5 g06438(new_n6823, new_n417, new_n6824);
nand_5 g06439(new_n6824, new_n847, new_n6825);
nand_5 g06440(new_n6825, new_n853, new_n6826);
nand_5 g06441(new_n6826, new_n859, new_n6827);
nand_5 g06442(new_n6827, new_n412, new_n6828);
nand_5 g06443(new_n6828, new_n866, new_n6829);
nand_5 g06444(new_n6829, new_n872, new_n6830);
nand_5 g06445(new_n6830, new_n878, new_n6831);
nand_5 g06446(new_n6831, new_n407, new_n6832);
nand_5 g06447(new_n6832, new_n885, new_n6833);
nand_5 g06448(new_n6833, new_n402, new_n6834);
nand_5 g06449(new_n6834, new_n397, new_n6835);
nand_5 g06450(new_n6835, new_n392, new_n6836);
nand_5 g06451(new_n6836, new_n894, new_n6837);
nand_5 g06452(new_n6837, new_n1087, new_n6838);
nand_5 g06453(new_n6838, new_n1129, new_n6839);
nand_5 g06454(new_n6839, new_n1084, new_n6840);
nand_5 g06455(new_n6840, new_n1134, new_n6841);
nand_5 g06456(new_n6841, new_n1080, new_n6842);
nand_5 g06457(new_n6842, new_n1075, new_n6843);
nand_5 g06458(new_n6843, new_n1070, new_n6844);
nand_5 g06459(new_n6844, new_n1143, new_n6845);
nand_5 g06460(new_n6845, new_n1148, new_n6846);
nand_5 g06461(new_n6846, new_n1065, new_n6847);
nand_5 g06462(new_n6847, new_n1062, new_n6848);
nand_5 g06463(new_n6848, new_n1156, new_n6849);
nand_5 g06464(new_n6849, new_n1057, new_n6850);
nand_5 g06465(new_n6850, new_n1053, new_n6851);
nand_5 g06466(new_n6851, new_n1050, new_n6852);
nand_5 g06467(new_n6852, new_n1045, new_n6853_1);
nand_5 g06468(new_n6853_1, new_n1040, new_n6854);
nand_5 g06469(new_n6854, new_n1036, new_n6855);
nand_5 g06470(new_n6855, new_n1033, new_n6856);
nand_5 g06471(new_n6856, new_n1028, new_n6857);
nand_5 g06472(new_n6857, new_n1026, new_n6858);
nand_5 g06473(new_n6858, new_n1021, new_n6859);
nand_5 g06474(new_n6859, new_n1017, new_n6860);
nand_5 g06475(new_n6860, new_n1012, new_n6861);
nand_5 g06476(new_n6861, new_n1009, new_n6862);
nand_5 g06477(new_n6862, new_n1004, new_n6863);
nand_5 g06478(new_n6863, new_n1000, new_n6864);
nand_5 g06479(new_n6864, new_n995, new_n6865);
nand_5 g06480(new_n6865, new_n990, new_n6866);
nand_5 g06481(new_n6866, new_n985, new_n6867);
nand_5 g06482(new_n6867, new_n981, new_n6868);
nand_5 g06483(new_n6868, new_n1179, new_n6869);
nand_5 g06484(new_n6869, new_n976, new_n6870);
nand_5 g06485(new_n6870, new_n971, new_n6871);
nand_5 g06486(new_n6871, new_n966, new_n6872);
nand_5 g06487(new_n6872, new_n961, new_n6873_1);
nand_5 g06488(new_n6873_1, new_n957, new_n6874);
nand_5 g06489(new_n6874, new_n952, new_n6875);
nand_5 g06490(new_n6875, new_n948_1, new_n6876);
nand_5 g06491(new_n6876, new_n943, new_n6877);
nand_5 g06492(new_n6877, new_n941, new_n6878);
nand_5 g06493(new_n6878, new_n938, new_n6879);
nand_5 g06494(new_n6879, new_n936, new_n6880);
nand_5 g06495(new_n6880, new_n931, new_n6881);
nand_5 g06496(new_n6881, new_n927, new_n6882);
nand_5 g06497(new_n6882, new_n922, new_n6883);
nand_5 g06498(new_n6883, new_n917, new_n6884);
nand_5 g06499(new_n6884, new_n912, new_n6885);
nand_5 g06500(new_n6885, new_n907, new_n6886);
nand_5 g06501(new_n6886, new_n903, new_n6887);
nand_5 g06502(new_n6887, new_n2066, new_n6888);
nand_5 g06503(new_n6888, new_n2063, new_n6889);
nand_5 g06504(new_n6889, new_n2062, new_n6890);
nand_5 g06505(new_n6890, new_n2058, new_n6891);
nand_5 g06506(new_n6891, new_n2055, new_n6892);
nand_5 g06507(new_n6892, new_n2051, new_n6893);
nand_5 g06508(new_n6893, new_n2046, new_n6894);
nand_5 g06509(new_n6894, new_n2042, new_n6895);
nand_5 g06510(new_n6895, n11345, new_n6896);
nor_5  g06511(new_n6896, new_n1367, n6853);
nand_5 g06512(new_n1628, new_n1629, new_n6898);
nand_5 g06513(new_n6898, new_n1625, new_n6899);
nand_5 g06514(new_n6899, new_n1621, new_n6900);
nand_5 g06515(new_n6900, new_n1618, new_n6901);
nand_5 g06516(new_n6901, new_n1778, new_n6902);
nand_5 g06517(new_n6902, new_n1782, new_n6903);
nand_5 g06518(new_n6903, new_n1614, new_n6904);
nand_5 g06519(new_n6904, new_n1611, new_n6905);
nand_5 g06520(new_n6905, new_n1789, new_n6906);
nand_5 g06521(new_n6906, new_n1608, new_n6907);
nand_5 g06522(new_n6907, new_n1605, new_n6908);
nand_5 g06523(new_n6908, new_n1795, new_n6909);
nand_5 g06524(new_n6909, new_n1799, new_n6910);
nand_5 g06525(new_n6910, new_n1602, new_n6911);
nand_5 g06526(new_n6911, new_n1599, new_n6912);
nand_5 g06527(new_n6912, new_n1596, new_n6913);
nand_5 g06528(new_n6913, new_n1593, new_n6914);
nand_5 g06529(new_n6914, new_n1806, new_n6915);
nand_5 g06530(new_n6915, new_n1589, new_n6916);
nand_5 g06531(new_n6916, new_n1586, new_n6917);
nand_5 g06532(new_n6917, new_n1583, new_n6918);
nand_5 g06533(new_n6918, new_n1580, new_n6919);
nand_5 g06534(new_n6919, new_n1576, new_n6920);
nand_5 g06535(new_n6920, new_n1573, new_n6921);
nand_5 g06536(new_n6921, new_n1570, new_n6922);
nand_5 g06537(new_n6922, new_n1567, new_n6923);
nand_5 g06538(new_n6923, new_n1564, new_n6924);
nand_5 g06539(new_n6924, new_n1561, new_n6925);
nand_5 g06540(new_n6925, new_n1338, new_n6926);
nand_5 g06541(new_n6926, new_n1331, new_n6927);
nand_5 g06542(new_n6927, new_n1326, new_n6928);
nand_5 g06543(new_n6928, new_n1321, new_n6929);
nand_5 g06544(new_n6929, new_n1318, new_n6930);
nand_5 g06545(new_n6930, new_n1315, new_n6931);
nand_5 g06546(new_n6931, new_n1312, new_n6932);
nand_5 g06547(new_n6932, new_n1309, new_n6933);
nand_5 g06548(new_n6933, new_n1307, new_n6934);
nand_5 g06549(new_n6934, new_n1304, new_n6935);
nand_5 g06550(new_n6935, new_n1300, new_n6936);
nand_5 g06551(new_n6936, new_n1297, new_n6937);
nand_5 g06552(new_n6937, new_n1294, new_n6938);
nand_5 g06553(new_n6938, new_n1355, new_n6939);
nand_5 g06554(new_n6939, new_n1291, new_n6940);
nand_5 g06555(new_n6940, new_n1288, new_n6941);
nand_5 g06556(new_n6941, new_n1283, new_n6942);
nand_5 g06557(new_n6942, new_n1363, new_n6943);
nand_5 g06558(new_n6943, new_n1280, new_n6944);
nand_5 g06559(new_n6944, new_n1370, new_n6945);
nand_5 g06560(new_n6945, new_n1373, new_n6946_1);
nand_5 g06561(new_n6946_1, new_n1277, new_n6947);
nand_5 g06562(new_n6947, new_n1272, new_n6948);
nand_5 g06563(new_n6948, new_n1269, new_n6949);
nand_5 g06564(new_n6949, new_n1380, new_n6950);
nand_5 g06565(new_n6950, new_n1264, new_n6951);
nand_5 g06566(new_n6951, new_n1259, new_n6952_1);
nand_5 g06567(new_n6952_1, new_n1388, new_n6953);
nand_5 g06568(new_n6953, new_n1392, new_n6954);
nand_5 g06569(new_n6954, new_n1256, new_n6955);
nand_5 g06570(new_n6955, new_n1252, new_n6956);
nand_5 g06571(new_n6956, new_n1249, new_n6957);
nand_5 g06572(new_n6957, new_n1244, new_n6958);
nand_5 g06573(new_n6958, new_n1240, new_n6959);
nand_5 g06574(new_n6959, new_n1234, new_n6960);
nand_5 g06575(new_n6960, new_n1231, new_n6961);
nand_5 g06576(new_n6961, new_n1227, new_n6962);
nand_5 g06577(new_n6962, new_n1407, new_n6963);
nand_5 g06578(new_n6963, new_n1223, new_n6964);
nand_5 g06579(new_n6964, new_n1218, new_n6965);
nand_5 g06580(new_n6965, new_n1213, new_n6966);
nand_5 g06581(new_n6966, new_n1210, new_n6967);
nand_5 g06582(new_n6967, new_n1206, new_n6968);
nand_5 g06583(new_n6968, new_n1418, new_n6969);
nand_5 g06584(new_n6969, new_n1422, new_n6970);
nand_5 g06585(new_n6970, new_n1428, new_n6971);
nand_5 g06586(new_n6971, new_n1203, new_n6972);
nand_5 g06587(new_n6972, new_n1433, new_n6973);
nand_5 g06588(new_n6973, new_n581, new_n6974);
nand_5 g06589(new_n6974, new_n574, new_n6975);
nand_5 g06590(new_n6975, new_n568, new_n6976);
nand_5 g06591(new_n6976, new_n589, new_n6977);
nand_5 g06592(new_n6977, new_n595, new_n6978);
nand_5 g06593(new_n6978, new_n601, new_n6979_1);
nand_5 g06594(new_n6979_1, new_n563, new_n6980);
nand_5 g06595(new_n6980, new_n608, new_n6981);
nand_5 g06596(new_n6981, n13109, new_n6982);
nor_5  g06597(new_n6982, new_n555, n6952);
nand_5 g06598(new_n968, new_n966, new_n6984);
nand_5 g06599(new_n6984, new_n961, new_n6985);
nand_5 g06600(new_n6985, new_n957, new_n6986);
nand_5 g06601(new_n6986, new_n952, new_n6987);
nand_5 g06602(new_n6987, new_n948_1, new_n6988);
nand_5 g06603(new_n6988, new_n943, new_n6989);
nand_5 g06604(new_n6989, new_n941, new_n6990);
nand_5 g06605(new_n6990, new_n938, new_n6991);
nand_5 g06606(new_n6991, new_n936, new_n6992);
nand_5 g06607(new_n6992, new_n931, new_n6993);
nand_5 g06608(new_n6993, new_n927, new_n6994);
nand_5 g06609(new_n6994, new_n922, new_n6995);
nand_5 g06610(new_n6995, new_n917, new_n6996);
nand_5 g06611(new_n6996, new_n912, new_n6997);
nand_5 g06612(new_n6997, new_n907, new_n6998);
nand_5 g06613(new_n6998, new_n903, new_n6999_1);
nand_5 g06614(new_n6999_1, new_n2066, new_n7000);
nand_5 g06615(new_n7000, new_n2063, new_n7001);
nand_5 g06616(new_n7001, new_n2062, new_n7002);
nand_5 g06617(new_n7002, new_n2058, new_n7003);
nand_5 g06618(new_n7003, new_n2055, new_n7004);
nand_5 g06619(new_n7004, new_n2051, new_n7005);
nand_5 g06620(new_n7005, new_n2046, new_n7006);
nand_5 g06621(new_n7006, new_n2042, new_n7007);
nand_5 g06622(new_n7007, new_n2039, new_n7008);
nand_5 g06623(new_n7008, new_n2036, new_n7009);
nand_5 g06624(new_n7009, new_n2033, new_n7010);
nand_5 g06625(new_n7010, new_n2029, new_n7011);
nand_5 g06626(new_n7011, new_n2026, new_n7012);
nand_5 g06627(new_n7012, new_n2022, new_n7013);
nand_5 g06628(new_n7013, new_n2018, new_n7014);
nand_5 g06629(new_n7014, new_n1726, new_n7015);
nand_5 g06630(new_n7015, new_n1722, new_n7016);
nand_5 g06631(new_n7016, new_n1718, new_n7017);
nand_5 g06632(new_n7017, new_n1713, new_n7018);
nand_5 g06633(new_n7018, new_n1737, new_n7019);
nand_5 g06634(new_n7019, new_n1709, new_n7020);
nand_5 g06635(new_n7020, new_n1742, new_n7021);
nand_5 g06636(new_n7021, new_n1704, new_n7022);
nand_5 g06637(new_n7022, new_n1702_1, new_n7023);
nand_5 g06638(new_n7023, new_n1698, new_n7024);
nand_5 g06639(new_n7024, new_n1695, new_n7025);
nand_5 g06640(new_n7025, new_n1692, new_n7026);
nand_5 g06641(new_n7026, new_n1752, new_n7027);
nand_5 g06642(new_n7027, new_n1688, new_n7028);
nand_5 g06643(new_n7028, new_n1685, new_n7029);
nand_5 g06644(new_n7029, new_n1680, new_n7030);
nand_5 g06645(new_n7030, new_n1676, new_n7031);
nand_5 g06646(new_n7031, new_n1672, new_n7032);
nand_5 g06647(new_n7032, new_n1669, new_n7033);
nand_5 g06648(new_n7033, new_n1666, new_n7034);
nand_5 g06649(new_n7034, new_n1663, new_n7035);
nand_5 g06650(new_n7035, new_n1658, new_n7036);
nand_5 g06651(new_n7036, new_n1653, new_n7037);
nand_5 g06652(new_n7037, new_n1651, new_n7038);
nand_5 g06653(new_n7038, new_n1649, new_n7039);
nand_5 g06654(new_n7039, new_n1646, new_n7040);
nand_5 g06655(new_n7040, new_n1643, new_n7041);
nand_5 g06656(new_n7041, new_n1641, new_n7042);
nand_5 g06657(new_n7042, new_n1638, new_n7043);
nand_5 g06658(new_n7043, new_n1635, new_n7044);
nand_5 g06659(new_n7044, new_n1632, new_n7045);
nand_5 g06660(new_n7045, new_n1628, new_n7046);
nand_5 g06661(new_n7046, new_n1625, new_n7047);
nand_5 g06662(new_n7047, new_n1621, new_n7048);
nand_5 g06663(new_n7048, new_n1618, new_n7049);
nand_5 g06664(new_n7049, new_n1778, new_n7050);
nand_5 g06665(new_n7050, new_n1782, new_n7051);
nand_5 g06666(new_n7051, new_n1614, new_n7052);
nand_5 g06667(new_n7052, new_n1611, new_n7053);
nand_5 g06668(new_n7053, new_n1789, new_n7054);
nand_5 g06669(new_n7054, new_n1608, new_n7055);
nand_5 g06670(new_n7055, new_n1605, new_n7056);
nand_5 g06671(new_n7056, new_n1795, new_n7057);
nand_5 g06672(new_n7057, new_n1799, new_n7058);
nand_5 g06673(new_n7058, new_n1602, new_n7059);
nand_5 g06674(new_n7059, new_n1599, new_n7060);
nand_5 g06675(new_n7060, new_n1596, new_n7061);
nand_5 g06676(new_n7061, new_n1593, new_n7062);
nand_5 g06677(new_n7062, new_n1806, new_n7063);
nand_5 g06678(new_n7063, new_n1589, new_n7064);
nand_5 g06679(new_n7064, new_n1586, new_n7065);
nand_5 g06680(new_n7065, new_n1583, new_n7066);
nand_5 g06681(new_n7066, new_n1580, new_n7067);
nand_5 g06682(new_n7067, n8635, new_n7068);
nor_5  g06683(new_n7068, new_n695, n6979);
nand_5 g06684(new_n1720, new_n1387, new_n7070);
nand_5 g06685(new_n7070, new_n1718, new_n7071_1);
nand_5 g06686(new_n7071_1, new_n1713, new_n7072);
nand_5 g06687(new_n7072, new_n1737, new_n7073_1);
nand_5 g06688(new_n7073_1, new_n1709, new_n7074);
nand_5 g06689(new_n7074, new_n1742, new_n7075);
nand_5 g06690(new_n7075, new_n1704, new_n7076);
nand_5 g06691(new_n7076, new_n1702_1, new_n7077);
nand_5 g06692(new_n7077, new_n1698, new_n7078);
nand_5 g06693(new_n7078, new_n1695, new_n7079);
nand_5 g06694(new_n7079, new_n1692, new_n7080);
nand_5 g06695(new_n7080, new_n1752, new_n7081);
nand_5 g06696(new_n7081, new_n1688, new_n7082);
nand_5 g06697(new_n7082, new_n1685, new_n7083);
nand_5 g06698(new_n7083, new_n1680, new_n7084);
nand_5 g06699(new_n7084, new_n1676, new_n7085);
nand_5 g06700(new_n7085, new_n1672, new_n7086);
nand_5 g06701(new_n7086, new_n1669, new_n7087);
nand_5 g06702(new_n7087, new_n1666, new_n7088);
nand_5 g06703(new_n7088, new_n1663, new_n7089);
nand_5 g06704(new_n7089, new_n1658, new_n7090);
nand_5 g06705(new_n7090, new_n1653, new_n7091);
nand_5 g06706(new_n7091, new_n1651, new_n7092);
nand_5 g06707(new_n7092, new_n1649, new_n7093);
nand_5 g06708(new_n7093, new_n1646, new_n7094);
nand_5 g06709(new_n7094, new_n1643, new_n7095);
nand_5 g06710(new_n7095, new_n1641, new_n7096);
nand_5 g06711(new_n7096, new_n1638, new_n7097);
nand_5 g06712(new_n7097, new_n1635, new_n7098);
nand_5 g06713(new_n7098, new_n1632, new_n7099);
nand_5 g06714(new_n7099, new_n1628, new_n7100);
nand_5 g06715(new_n7100, new_n1625, new_n7101);
nand_5 g06716(new_n7101, new_n1621, new_n7102);
nand_5 g06717(new_n7102, new_n1618, new_n7103);
nand_5 g06718(new_n7103, new_n1778, new_n7104_1);
nand_5 g06719(new_n7104_1, new_n1782, new_n7105);
nand_5 g06720(new_n7105, new_n1614, new_n7106);
nand_5 g06721(new_n7106, new_n1611, new_n7107);
nand_5 g06722(new_n7107, new_n1789, new_n7108);
nand_5 g06723(new_n7108, new_n1608, new_n7109);
nand_5 g06724(new_n7109, new_n1605, new_n7110);
nand_5 g06725(new_n7110, new_n1795, new_n7111);
nand_5 g06726(new_n7111, new_n1799, new_n7112);
nand_5 g06727(new_n7112, new_n1602, new_n7113);
nand_5 g06728(new_n7113, new_n1599, new_n7114);
nand_5 g06729(new_n7114, new_n1596, new_n7115);
nand_5 g06730(new_n7115, new_n1593, new_n7116);
nand_5 g06731(new_n7116, new_n1806, new_n7117);
nand_5 g06732(new_n7117, new_n1589, new_n7118);
nand_5 g06733(new_n7118, new_n1586, new_n7119);
nand_5 g06734(new_n7119, new_n1583, new_n7120);
nand_5 g06735(new_n7120, new_n1580, new_n7121);
nand_5 g06736(new_n7121, new_n1576, new_n7122);
nand_5 g06737(new_n7122, new_n1573, new_n7123);
nand_5 g06738(new_n7123, new_n1570, new_n7124);
nand_5 g06739(new_n7124, new_n1567, new_n7125);
nand_5 g06740(new_n7125, new_n1564, new_n7126);
nand_5 g06741(new_n7126, new_n1561, new_n7127);
nand_5 g06742(new_n7127, new_n1338, new_n7128);
nand_5 g06743(new_n7128, new_n1331, new_n7129);
nand_5 g06744(new_n7129, new_n1326, new_n7130);
nand_5 g06745(new_n7130, new_n1321, new_n7131);
nand_5 g06746(new_n7131, new_n1318, new_n7132_1);
nand_5 g06747(new_n7132_1, new_n1315, new_n7133);
nand_5 g06748(new_n7133, new_n1312, new_n7134);
nand_5 g06749(new_n7134, new_n1309, new_n7135);
nand_5 g06750(new_n7135, new_n1307, new_n7136);
nand_5 g06751(new_n7136, new_n1304, new_n7137);
nand_5 g06752(new_n7137, new_n1300, new_n7138);
nand_5 g06753(new_n7138, new_n1297, new_n7139);
nand_5 g06754(new_n7139, new_n1294, new_n7140);
nand_5 g06755(new_n7140, new_n1355, new_n7141);
nand_5 g06756(new_n7141, new_n1291, new_n7142);
nand_5 g06757(new_n7142, new_n1288, new_n7143);
nand_5 g06758(new_n7143, new_n1283, new_n7144);
nand_5 g06759(new_n7144, new_n1363, new_n7145);
nand_5 g06760(new_n7145, new_n1280, new_n7146);
nand_5 g06761(new_n7146, new_n1370, new_n7147);
nand_5 g06762(new_n7147, new_n1373, new_n7148);
nand_5 g06763(new_n7148, new_n1277, new_n7149);
nand_5 g06764(new_n7149, new_n1272, new_n7150);
nand_5 g06765(new_n7150, new_n1269, new_n7151);
nand_5 g06766(new_n7151, new_n1380, new_n7152_1);
nand_5 g06767(new_n7152_1, new_n1264, new_n7153);
nand_5 g06768(new_n7153, n14408, new_n7154);
nor_5  g06769(new_n7154, new_n816, n7071);
nand_5 g06770(new_n1725, new_n430, new_n7156);
nand_5 g06771(new_n7156, new_n427_1, new_n7157);
nand_5 g06772(new_n7157, new_n422, new_n7158);
nand_5 g06773(new_n7158, new_n828, new_n7159);
nand_5 g06774(new_n7159, new_n834, new_n7160);
nand_5 g06775(new_n7160, new_n840, new_n7161);
nand_5 g06776(new_n7161, new_n417, new_n7162);
nand_5 g06777(new_n7162, new_n847, new_n7163);
nand_5 g06778(new_n7163, new_n853, new_n7164);
nand_5 g06779(new_n7164, new_n859, new_n7165);
nand_5 g06780(new_n7165, new_n412, new_n7166);
nand_5 g06781(new_n7166, new_n866, new_n7167);
nand_5 g06782(new_n7167, new_n872, new_n7168);
nand_5 g06783(new_n7168, new_n878, new_n7169);
nand_5 g06784(new_n7169, new_n407, new_n7170);
nand_5 g06785(new_n7170, new_n885, new_n7171);
nand_5 g06786(new_n7171, new_n402, new_n7172);
nand_5 g06787(new_n7172, new_n397, new_n7173);
nand_5 g06788(new_n7173, new_n392, new_n7174);
nand_5 g06789(new_n7174, new_n894, new_n7175);
nand_5 g06790(new_n7175, new_n1087, new_n7176);
nand_5 g06791(new_n7176, new_n1129, new_n7177);
nand_5 g06792(new_n7177, new_n1084, new_n7178);
nand_5 g06793(new_n7178, new_n1134, new_n7179);
nand_5 g06794(new_n7179, new_n1080, new_n7180);
nand_5 g06795(new_n7180, new_n1075, new_n7181);
nand_5 g06796(new_n7181, new_n1070, new_n7182);
nand_5 g06797(new_n7182, new_n1143, new_n7183);
nand_5 g06798(new_n7183, new_n1148, new_n7184);
nand_5 g06799(new_n7184, new_n1065, new_n7185);
nand_5 g06800(new_n7185, new_n1062, new_n7186);
nand_5 g06801(new_n7186, new_n1156, new_n7187);
nand_5 g06802(new_n7187, new_n1057, new_n7188);
nand_5 g06803(new_n7188, new_n1053, new_n7189);
nand_5 g06804(new_n7189, new_n1050, new_n7190);
nand_5 g06805(new_n7190, new_n1045, new_n7191);
nand_5 g06806(new_n7191, new_n1040, new_n7192);
nand_5 g06807(new_n7192, new_n1036, new_n7193);
nand_5 g06808(new_n7193, new_n1033, new_n7194);
nand_5 g06809(new_n7194, new_n1028, new_n7195);
nand_5 g06810(new_n7195, new_n1026, new_n7196);
nand_5 g06811(new_n7196, new_n1021, new_n7197);
nand_5 g06812(new_n7197, new_n1017, new_n7198);
nand_5 g06813(new_n7198, new_n1012, new_n7199);
nand_5 g06814(new_n7199, new_n1009, new_n7200);
nand_5 g06815(new_n7200, new_n1004, new_n7201);
nand_5 g06816(new_n7201, new_n1000, new_n7202);
nand_5 g06817(new_n7202, new_n995, new_n7203);
nand_5 g06818(new_n7203, new_n990, new_n7204);
nand_5 g06819(new_n7204, new_n985, new_n7205);
nand_5 g06820(new_n7205, new_n981, new_n7206);
nand_5 g06821(new_n7206, new_n1179, new_n7207);
nand_5 g06822(new_n7207, new_n976, new_n7208);
nand_5 g06823(new_n7208, new_n971, new_n7209);
nand_5 g06824(new_n7209, new_n966, new_n7210);
nand_5 g06825(new_n7210, new_n961, new_n7211);
nand_5 g06826(new_n7211, new_n957, new_n7212);
nand_5 g06827(new_n7212, new_n952, new_n7213);
nand_5 g06828(new_n7213, new_n948_1, new_n7214);
nand_5 g06829(new_n7214, new_n943, new_n7215);
nand_5 g06830(new_n7215, new_n941, new_n7216);
nand_5 g06831(new_n7216, new_n938, new_n7217);
nand_5 g06832(new_n7217, new_n936, new_n7218);
nand_5 g06833(new_n7218, new_n931, new_n7219);
nand_5 g06834(new_n7219, new_n927, new_n7220);
nand_5 g06835(new_n7220, new_n922, new_n7221);
nand_5 g06836(new_n7221, new_n917, new_n7222);
nand_5 g06837(new_n7222, new_n912, new_n7223);
nand_5 g06838(new_n7223, new_n907, new_n7224);
nand_5 g06839(new_n7224, new_n903, new_n7225);
nand_5 g06840(new_n7225, new_n2066, new_n7226);
nand_5 g06841(new_n7226, new_n2063, new_n7227);
nand_5 g06842(new_n7227, new_n2062, new_n7228);
nand_5 g06843(new_n7228, new_n2058, new_n7229);
nand_5 g06844(new_n7229, new_n2055, new_n7230);
nand_5 g06845(new_n7230, new_n2051, new_n7231);
nand_5 g06846(new_n7231, new_n2046, new_n7232);
nand_5 g06847(new_n7232, new_n2042, new_n7233);
nand_5 g06848(new_n7233, new_n2039, new_n7234);
nand_5 g06849(new_n7234, new_n2036, new_n7235);
nand_5 g06850(new_n7235, new_n2033, new_n7236);
nand_5 g06851(new_n7236, new_n2029, new_n7237);
nand_5 g06852(new_n7237, new_n2026, new_n7238);
nand_5 g06853(new_n7238, new_n2022, new_n7239);
nand_5 g06854(new_n7239, n5023, new_n7240);
nor_5  g06855(new_n7240, new_n1261, n7073);
not_4  g06856(new_n1336, new_n7242);
nor_5  g06857(n13992, n5014, new_n7243);
not_4  g06858(new_n7243, new_n7244);
nand_5 g06859(new_n7244, new_n941, new_n7245);
nand_5 g06860(new_n7245, new_n938, new_n7246_1);
nand_5 g06861(new_n7246_1, new_n936, new_n7247);
nand_5 g06862(new_n7247, new_n931, new_n7248);
nand_5 g06863(new_n7248, new_n927, new_n7249);
nand_5 g06864(new_n7249, new_n922, new_n7250);
nand_5 g06865(new_n7250, new_n917, new_n7251);
nand_5 g06866(new_n7251, new_n912, new_n7252);
nand_5 g06867(new_n7252, new_n907, new_n7253);
nand_5 g06868(new_n7253, new_n903, new_n7254);
nand_5 g06869(new_n7254, new_n2066, new_n7255);
nand_5 g06870(new_n7255, new_n2063, new_n7256);
nand_5 g06871(new_n7256, new_n2062, new_n7257);
nand_5 g06872(new_n7257, new_n2058, new_n7258);
nand_5 g06873(new_n7258, new_n2055, new_n7259);
nand_5 g06874(new_n7259, new_n2051, new_n7260);
nand_5 g06875(new_n7260, new_n2046, new_n7261);
nand_5 g06876(new_n7261, new_n2042, new_n7262);
nand_5 g06877(new_n7262, new_n2039, new_n7263);
nand_5 g06878(new_n7263, new_n2036, new_n7264);
nand_5 g06879(new_n7264, new_n2033, new_n7265_1);
nand_5 g06880(new_n7265_1, new_n2029, new_n7266);
nand_5 g06881(new_n7266, new_n2026, new_n7267);
nand_5 g06882(new_n7267, new_n2022, new_n7268);
nand_5 g06883(new_n7268, new_n2018, new_n7269);
nand_5 g06884(new_n7269, new_n1726, new_n7270);
nand_5 g06885(new_n7270, new_n1722, new_n7271);
nand_5 g06886(new_n7271, new_n1718, new_n7272_1);
nand_5 g06887(new_n7272_1, new_n1713, new_n7273);
nand_5 g06888(new_n7273, new_n1737, new_n7274);
nand_5 g06889(new_n7274, new_n1709, new_n7275);
nand_5 g06890(new_n7275, new_n1742, new_n7276);
nand_5 g06891(new_n7276, new_n1704, new_n7277);
nand_5 g06892(new_n7277, new_n1702_1, new_n7278);
nand_5 g06893(new_n7278, new_n1698, new_n7279);
nand_5 g06894(new_n7279, new_n1695, new_n7280);
nand_5 g06895(new_n7280, new_n1692, new_n7281);
nand_5 g06896(new_n7281, new_n1752, new_n7282_1);
nand_5 g06897(new_n7282_1, new_n1688, new_n7283);
nand_5 g06898(new_n7283, new_n1685, new_n7284);
nand_5 g06899(new_n7284, new_n1680, new_n7285);
nand_5 g06900(new_n7285, new_n1676, new_n7286);
nand_5 g06901(new_n7286, new_n1672, new_n7287);
nand_5 g06902(new_n7287, new_n1669, new_n7288);
nand_5 g06903(new_n7288, new_n1666, new_n7289);
nand_5 g06904(new_n7289, new_n1663, new_n7290);
nand_5 g06905(new_n7290, new_n1658, new_n7291);
nand_5 g06906(new_n7291, new_n1653, new_n7292);
nand_5 g06907(new_n7292, new_n1651, new_n7293);
nand_5 g06908(new_n7293, new_n1649, new_n7294);
nand_5 g06909(new_n7294, new_n1646, new_n7295);
nand_5 g06910(new_n7295, new_n1643, new_n7296);
nand_5 g06911(new_n7296, new_n1641, new_n7297);
nand_5 g06912(new_n7297, new_n1638, new_n7298);
nand_5 g06913(new_n7298, new_n1635, new_n7299);
nand_5 g06914(new_n7299, new_n1632, new_n7300);
nand_5 g06915(new_n7300, new_n1628, new_n7301);
nand_5 g06916(new_n7301, new_n1625, new_n7302);
nand_5 g06917(new_n7302, new_n1621, new_n7303);
nand_5 g06918(new_n7303, new_n1618, new_n7304);
nand_5 g06919(new_n7304, new_n1778, new_n7305);
nand_5 g06920(new_n7305, new_n1782, new_n7306);
nand_5 g06921(new_n7306, new_n1614, new_n7307);
nand_5 g06922(new_n7307, new_n1611, new_n7308);
nand_5 g06923(new_n7308, new_n1789, new_n7309);
nand_5 g06924(new_n7309, new_n1608, new_n7310);
nand_5 g06925(new_n7310, new_n1605, new_n7311);
nand_5 g06926(new_n7311, new_n1795, new_n7312);
nand_5 g06927(new_n7312, new_n1799, new_n7313);
nand_5 g06928(new_n7313, new_n1602, new_n7314);
nand_5 g06929(new_n7314, new_n1599, new_n7315);
nand_5 g06930(new_n7315, new_n1596, new_n7316);
nand_5 g06931(new_n7316, new_n1593, new_n7317);
nand_5 g06932(new_n7317, new_n1806, new_n7318);
nand_5 g06933(new_n7318, new_n1589, new_n7319);
nand_5 g06934(new_n7319, new_n1586, new_n7320);
nand_5 g06935(new_n7320, new_n1583, new_n7321);
nand_5 g06936(new_n7321, new_n1580, new_n7322);
nand_5 g06937(new_n7322, new_n1576, new_n7323);
nand_5 g06938(new_n7323, new_n1573, new_n7324);
nand_5 g06939(new_n7324, new_n1570, new_n7325);
nand_5 g06940(new_n7325, new_n1567, new_n7326);
nand_5 g06941(new_n7326, new_n1564, new_n7327);
nand_5 g06942(new_n7327, new_n1561, new_n7328);
nand_5 g06943(new_n7328, n11590, new_n7329);
nor_5  g06944(new_n7329, new_n7242, n7132);
nand_5 g06945(new_n1305, new_n750, new_n7331);
nand_5 g06946(new_n7331, new_n1304, new_n7332);
nand_5 g06947(new_n7332, new_n1300, new_n7333);
nand_5 g06948(new_n7333, new_n1297, new_n7334);
nand_5 g06949(new_n7334, new_n1294, new_n7335);
nand_5 g06950(new_n7335, new_n1355, new_n7336);
nand_5 g06951(new_n7336, new_n1291, new_n7337);
nand_5 g06952(new_n7337, new_n1288, new_n7338);
nand_5 g06953(new_n7338, new_n1283, new_n7339);
nand_5 g06954(new_n7339, new_n1363, new_n7340);
nand_5 g06955(new_n7340, new_n1280, new_n7341);
nand_5 g06956(new_n7341, new_n1370, new_n7342);
nand_5 g06957(new_n7342, new_n1373, new_n7343);
nand_5 g06958(new_n7343, new_n1277, new_n7344);
nand_5 g06959(new_n7344, new_n1272, new_n7345);
nand_5 g06960(new_n7345, new_n1269, new_n7346);
nand_5 g06961(new_n7346, new_n1380, new_n7347);
nand_5 g06962(new_n7347, new_n1264, new_n7348);
nand_5 g06963(new_n7348, new_n1259, new_n7349);
nand_5 g06964(new_n7349, new_n1388, new_n7350);
nand_5 g06965(new_n7350, new_n1392, new_n7351);
nand_5 g06966(new_n7351, new_n1256, new_n7352);
nand_5 g06967(new_n7352, new_n1252, new_n7353);
nand_5 g06968(new_n7353, new_n1249, new_n7354_1);
nand_5 g06969(new_n7354_1, new_n1244, new_n7355);
nand_5 g06970(new_n7355, new_n1240, new_n7356);
nand_5 g06971(new_n7356, new_n1234, new_n7357);
nand_5 g06972(new_n7357, new_n1231, new_n7358);
nand_5 g06973(new_n7358, new_n1227, new_n7359);
nand_5 g06974(new_n7359, new_n1407, new_n7360);
nand_5 g06975(new_n7360, new_n1223, new_n7361);
nand_5 g06976(new_n7361, new_n1218, new_n7362);
nand_5 g06977(new_n7362, new_n1213, new_n7363);
nand_5 g06978(new_n7363, new_n1210, new_n7364);
nand_5 g06979(new_n7364, new_n1206, new_n7365);
nand_5 g06980(new_n7365, new_n1418, new_n7366);
nand_5 g06981(new_n7366, new_n1422, new_n7367);
nand_5 g06982(new_n7367, new_n1428, new_n7368);
nand_5 g06983(new_n7368, new_n1203, new_n7369);
nand_5 g06984(new_n7369, new_n1433, new_n7370);
nand_5 g06985(new_n7370, new_n581, new_n7371);
nand_5 g06986(new_n7371, new_n574, new_n7372);
nand_5 g06987(new_n7372, new_n568, new_n7373);
nand_5 g06988(new_n7373, new_n589, new_n7374);
nand_5 g06989(new_n7374, new_n595, new_n7375);
nand_5 g06990(new_n7375, new_n601, new_n7376);
nand_5 g06991(new_n7376, new_n563, new_n7377);
nand_5 g06992(new_n7377, new_n608, new_n7378);
nand_5 g06993(new_n7378, new_n558, new_n7379);
nand_5 g06994(new_n7379, new_n615, new_n7380);
nand_5 g06995(new_n7380, new_n553, new_n7381);
nand_5 g06996(new_n7381, new_n622, new_n7382_1);
nand_5 g06997(new_n7382_1, new_n628, new_n7383);
nand_5 g06998(new_n7383, new_n548, new_n7384);
nand_5 g06999(new_n7384, new_n543_1, new_n7385);
nand_5 g07000(new_n7385, new_n636, new_n7386);
nand_5 g07001(new_n7386, new_n642, new_n7387);
nand_5 g07002(new_n7387, new_n538, new_n7388);
nand_5 g07003(new_n7388, new_n533, new_n7389);
nand_5 g07004(new_n7389, new_n650_1, new_n7390);
nand_5 g07005(new_n7390, new_n528, new_n7391);
nand_5 g07006(new_n7391, new_n523, new_n7392);
nand_5 g07007(new_n7392, new_n518, new_n7393);
nand_5 g07008(new_n7393, new_n659, new_n7394);
nand_5 g07009(new_n7394, new_n665, new_n7395);
nand_5 g07010(new_n7395, new_n672, new_n7396);
nand_5 g07011(new_n7396, new_n513, new_n7397);
nand_5 g07012(new_n7397, new_n679, new_n7398);
nand_5 g07013(new_n7398, new_n685, new_n7399);
nand_5 g07014(new_n7399, new_n691, new_n7400);
nand_5 g07015(new_n7400, new_n508, new_n7401);
nand_5 g07016(new_n7401, new_n698, new_n7402);
nand_5 g07017(new_n7402, new_n503, new_n7403);
nand_5 g07018(new_n7403, new_n704, new_n7404);
nand_5 g07019(new_n7404, new_n498_1, new_n7405);
nand_5 g07020(new_n7405, new_n711, new_n7406);
nand_5 g07021(new_n7406, new_n493, new_n7407);
nand_5 g07022(new_n7407, new_n718, new_n7408);
nand_5 g07023(new_n7408, new_n488, new_n7409);
nand_5 g07024(new_n7409, new_n725, new_n7410);
nand_5 g07025(new_n7410, new_n483, new_n7411);
nand_5 g07026(new_n7411, new_n732, new_n7412);
nand_5 g07027(new_n7412, new_n478, new_n7413);
nand_5 g07028(new_n7413, new_n739, new_n7414);
nand_5 g07029(new_n7414, n9830, new_n7415);
nor_5  g07030(new_n7415, new_n742, n7152);
nand_5 g07031(new_n1597, new_n658, new_n7417);
nand_5 g07032(new_n7417, new_n1596, new_n7418);
nand_5 g07033(new_n7418, new_n1593, new_n7419);
nand_5 g07034(new_n7419, new_n1806, new_n7420);
nand_5 g07035(new_n7420, new_n1589, new_n7421);
nand_5 g07036(new_n7421, new_n1586, new_n7422);
nand_5 g07037(new_n7422, new_n1583, new_n7423);
nand_5 g07038(new_n7423, new_n1580, new_n7424);
nand_5 g07039(new_n7424, new_n1576, new_n7425);
nand_5 g07040(new_n7425, new_n1573, new_n7426);
nand_5 g07041(new_n7426, new_n1570, new_n7427);
nand_5 g07042(new_n7427, new_n1567, new_n7428);
nand_5 g07043(new_n7428, new_n1564, new_n7429);
nand_5 g07044(new_n7429, new_n1561, new_n7430);
nand_5 g07045(new_n7430, new_n1338, new_n7431);
nand_5 g07046(new_n7431, new_n1331, new_n7432);
nand_5 g07047(new_n7432, new_n1326, new_n7433);
nand_5 g07048(new_n7433, new_n1321, new_n7434);
nand_5 g07049(new_n7434, new_n1318, new_n7435);
nand_5 g07050(new_n7435, new_n1315, new_n7436);
nand_5 g07051(new_n7436, new_n1312, new_n7437);
nand_5 g07052(new_n7437, new_n1309, new_n7438);
nand_5 g07053(new_n7438, new_n1307, new_n7439);
nand_5 g07054(new_n7439, new_n1304, new_n7440);
nand_5 g07055(new_n7440, new_n1300, new_n7441);
nand_5 g07056(new_n7441, new_n1297, new_n7442);
nand_5 g07057(new_n7442, new_n1294, new_n7443);
nand_5 g07058(new_n7443, new_n1355, new_n7444);
nand_5 g07059(new_n7444, new_n1291, new_n7445);
nand_5 g07060(new_n7445, new_n1288, new_n7446);
nand_5 g07061(new_n7446, new_n1283, new_n7447);
nand_5 g07062(new_n7447, new_n1363, new_n7448);
nand_5 g07063(new_n7448, new_n1280, new_n7449);
nand_5 g07064(new_n7449, new_n1370, new_n7450_1);
nand_5 g07065(new_n7450_1, new_n1373, new_n7451);
nand_5 g07066(new_n7451, new_n1277, new_n7452);
nand_5 g07067(new_n7452, new_n1272, new_n7453);
nand_5 g07068(new_n7453, new_n1269, new_n7454);
nand_5 g07069(new_n7454, new_n1380, new_n7455);
nand_5 g07070(new_n7455, new_n1264, new_n7456);
nand_5 g07071(new_n7456, new_n1259, new_n7457);
nand_5 g07072(new_n7457, new_n1388, new_n7458);
nand_5 g07073(new_n7458, new_n1392, new_n7459);
nand_5 g07074(new_n7459, new_n1256, new_n7460);
nand_5 g07075(new_n7460, new_n1252, new_n7461);
nand_5 g07076(new_n7461, new_n1249, new_n7462);
nand_5 g07077(new_n7462, new_n1244, new_n7463);
nand_5 g07078(new_n7463, new_n1240, new_n7464);
nand_5 g07079(new_n7464, new_n1234, new_n7465);
nand_5 g07080(new_n7465, new_n1231, new_n7466);
nand_5 g07081(new_n7466, new_n1227, new_n7467);
nand_5 g07082(new_n7467, new_n1407, new_n7468);
nand_5 g07083(new_n7468, new_n1223, new_n7469);
nand_5 g07084(new_n7469, new_n1218, new_n7470);
nand_5 g07085(new_n7470, new_n1213, new_n7471);
nand_5 g07086(new_n7471, new_n1210, new_n7472);
nand_5 g07087(new_n7472, new_n1206, new_n7473);
nand_5 g07088(new_n7473, new_n1418, new_n7474);
nand_5 g07089(new_n7474, new_n1422, new_n7475);
nand_5 g07090(new_n7475, new_n1428, new_n7476);
nand_5 g07091(new_n7476, new_n1203, new_n7477);
nand_5 g07092(new_n7477, new_n1433, new_n7478);
nand_5 g07093(new_n7478, new_n581, new_n7479);
nand_5 g07094(new_n7479, new_n574, new_n7480);
nand_5 g07095(new_n7480, new_n568, new_n7481);
nand_5 g07096(new_n7481, new_n589, new_n7482);
nand_5 g07097(new_n7482, new_n595, new_n7483);
nand_5 g07098(new_n7483, new_n601, new_n7484);
nand_5 g07099(new_n7484, new_n563, new_n7485);
nand_5 g07100(new_n7485, new_n608, new_n7486);
nand_5 g07101(new_n7486, new_n558, new_n7487);
nand_5 g07102(new_n7487, new_n615, new_n7488);
nand_5 g07103(new_n7488, new_n553, new_n7489);
nand_5 g07104(new_n7489, new_n622, new_n7490);
nand_5 g07105(new_n7490, new_n628, new_n7491);
nand_5 g07106(new_n7491, new_n548, new_n7492);
nand_5 g07107(new_n7492, new_n543_1, new_n7493);
nand_5 g07108(new_n7493, new_n636, new_n7494);
nand_5 g07109(new_n7494, new_n642, new_n7495);
nand_5 g07110(new_n7495, new_n538, new_n7496);
nand_5 g07111(new_n7496, new_n533, new_n7497);
nand_5 g07112(new_n7497, new_n650_1, new_n7498);
nand_5 g07113(new_n7498, new_n528, new_n7499);
nand_5 g07114(new_n7499, new_n523, new_n7500);
nand_5 g07115(new_n7500, n13093, new_n7501);
nor_5  g07116(new_n7501, new_n515, n7246);
not_4  g07117(n10573, new_n7503);
nand_5 g07118(new_n1073, new_n7503, new_n7504);
nand_5 g07119(new_n7504, new_n593, new_n7505);
nand_5 g07120(new_n7505, new_n601, new_n7506);
nand_5 g07121(new_n7506, new_n563, new_n7507);
nand_5 g07122(new_n7507, new_n608, new_n7508);
nand_5 g07123(new_n7508, new_n558, new_n7509);
nand_5 g07124(new_n7509, new_n615, new_n7510);
nand_5 g07125(new_n7510, new_n553, new_n7511);
nand_5 g07126(new_n7511, new_n622, new_n7512);
nand_5 g07127(new_n7512, new_n628, new_n7513);
nand_5 g07128(new_n7513, new_n548, new_n7514);
nand_5 g07129(new_n7514, new_n543_1, new_n7515);
nand_5 g07130(new_n7515, new_n636, new_n7516);
nand_5 g07131(new_n7516, new_n642, new_n7517);
nand_5 g07132(new_n7517, new_n538, new_n7518);
nand_5 g07133(new_n7518, new_n533, new_n7519);
nand_5 g07134(new_n7519, new_n650_1, new_n7520);
nand_5 g07135(new_n7520, new_n528, new_n7521);
nand_5 g07136(new_n7521, new_n523, new_n7522);
nand_5 g07137(new_n7522, new_n518, new_n7523);
nand_5 g07138(new_n7523, new_n659, new_n7524);
nand_5 g07139(new_n7524, new_n665, new_n7525);
nand_5 g07140(new_n7525, new_n672, new_n7526);
nand_5 g07141(new_n7526, new_n513, new_n7527);
nand_5 g07142(new_n7527, new_n679, new_n7528);
nand_5 g07143(new_n7528, new_n685, new_n7529);
nand_5 g07144(new_n7529, new_n691, new_n7530);
nand_5 g07145(new_n7530, new_n508, new_n7531);
nand_5 g07146(new_n7531, new_n698, new_n7532);
nand_5 g07147(new_n7532, new_n503, new_n7533);
nand_5 g07148(new_n7533, new_n704, new_n7534);
nand_5 g07149(new_n7534, new_n498_1, new_n7535);
nand_5 g07150(new_n7535, new_n711, new_n7536);
nand_5 g07151(new_n7536, new_n493, new_n7537);
nand_5 g07152(new_n7537, new_n718, new_n7538);
nand_5 g07153(new_n7538, new_n488, new_n7539);
nand_5 g07154(new_n7539, new_n725, new_n7540);
nand_5 g07155(new_n7540, new_n483, new_n7541);
nand_5 g07156(new_n7541, new_n732, new_n7542);
nand_5 g07157(new_n7542, new_n478, new_n7543);
nand_5 g07158(new_n7543, new_n739, new_n7544);
nand_5 g07159(new_n7544, new_n745, new_n7545);
nand_5 g07160(new_n7545, new_n751, new_n7546);
nand_5 g07161(new_n7546, new_n473, new_n7547);
nand_5 g07162(new_n7547, new_n758, new_n7548);
nand_5 g07163(new_n7548, new_n764, new_n7549);
nand_5 g07164(new_n7549, new_n770, new_n7550);
nand_5 g07165(new_n7550, new_n468, new_n7551);
nand_5 g07166(new_n7551, new_n777, new_n7552);
nand_5 g07167(new_n7552, new_n783, new_n7553);
nand_5 g07168(new_n7553, new_n789, new_n7554);
nand_5 g07169(new_n7554, new_n463, new_n7555);
nand_5 g07170(new_n7555, new_n796, new_n7556);
nand_5 g07171(new_n7556, new_n458, new_n7557);
nand_5 g07172(new_n7557, new_n453, new_n7558);
nand_5 g07173(new_n7558, new_n447, new_n7559);
nand_5 g07174(new_n7559, new_n805, new_n7560);
nand_5 g07175(new_n7560, new_n811, new_n7561);
nand_5 g07176(new_n7561, new_n442, new_n7562);
nand_5 g07177(new_n7562, new_n437, new_n7563);
nand_5 g07178(new_n7563, new_n819, new_n7564);
nand_5 g07179(new_n7564, new_n432, new_n7565);
nand_5 g07180(new_n7565, new_n427_1, new_n7566);
nand_5 g07181(new_n7566, new_n422, new_n7567);
nand_5 g07182(new_n7567, new_n828, new_n7568);
nand_5 g07183(new_n7568, new_n834, new_n7569);
nand_5 g07184(new_n7569, new_n840, new_n7570);
nand_5 g07185(new_n7570, new_n417, new_n7571);
nand_5 g07186(new_n7571, new_n847, new_n7572);
nand_5 g07187(new_n7572, new_n853, new_n7573);
nand_5 g07188(new_n7573, new_n859, new_n7574);
nand_5 g07189(new_n7574, new_n412, new_n7575);
nand_5 g07190(new_n7575, new_n866, new_n7576);
nand_5 g07191(new_n7576, new_n872, new_n7577);
nand_5 g07192(new_n7577, new_n878, new_n7578);
nand_5 g07193(new_n7578, new_n407, new_n7579);
nand_5 g07194(new_n7579, new_n885, new_n7580);
nand_5 g07195(new_n7580, new_n402, new_n7581);
nand_5 g07196(new_n7581, new_n397, new_n7582);
nand_5 g07197(new_n7582, new_n392, new_n7583);
nand_5 g07198(new_n7583, new_n894, new_n7584);
nand_5 g07199(new_n7584, new_n1087, new_n7585);
nand_5 g07200(new_n7585, new_n1129, new_n7586);
nand_5 g07201(new_n7586, new_n1084, new_n7587);
nand_5 g07202(new_n7587, new_n1134, new_n7588);
nand_5 g07203(new_n7588, n1776, new_n7589);
nor_5  g07204(new_n7589, new_n1077, n7265);
nand_5 g07205(new_n1403, new_n1223, new_n7591);
nand_5 g07206(new_n7591, new_n1218, new_n7592);
nand_5 g07207(new_n7592, new_n1213, new_n7593);
nand_5 g07208(new_n7593, new_n1210, new_n7594);
nand_5 g07209(new_n7594, new_n1206, new_n7595);
nand_5 g07210(new_n7595, new_n1418, new_n7596);
nand_5 g07211(new_n7596, new_n1422, new_n7597);
nand_5 g07212(new_n7597, new_n1428, new_n7598);
nand_5 g07213(new_n7598, new_n1203, new_n7599);
nand_5 g07214(new_n7599, new_n1433, new_n7600);
nand_5 g07215(new_n7600, new_n581, new_n7601);
nand_5 g07216(new_n7601, new_n574, new_n7602);
nand_5 g07217(new_n7602, new_n568, new_n7603);
nand_5 g07218(new_n7603, new_n589, new_n7604);
nand_5 g07219(new_n7604, new_n595, new_n7605);
nand_5 g07220(new_n7605, new_n601, new_n7606);
nand_5 g07221(new_n7606, new_n563, new_n7607);
nand_5 g07222(new_n7607, new_n608, new_n7608);
nand_5 g07223(new_n7608, new_n558, new_n7609);
nand_5 g07224(new_n7609, new_n615, new_n7610);
nand_5 g07225(new_n7610, new_n553, new_n7611);
nand_5 g07226(new_n7611, new_n622, new_n7612);
nand_5 g07227(new_n7612, new_n628, new_n7613);
nand_5 g07228(new_n7613, new_n548, new_n7614);
nand_5 g07229(new_n7614, new_n543_1, new_n7615);
nand_5 g07230(new_n7615, new_n636, new_n7616);
nand_5 g07231(new_n7616, new_n642, new_n7617);
nand_5 g07232(new_n7617, new_n538, new_n7618);
nand_5 g07233(new_n7618, new_n533, new_n7619);
nand_5 g07234(new_n7619, new_n650_1, new_n7620);
nand_5 g07235(new_n7620, new_n528, new_n7621);
nand_5 g07236(new_n7621, new_n523, new_n7622);
nand_5 g07237(new_n7622, new_n518, new_n7623);
nand_5 g07238(new_n7623, new_n659, new_n7624);
nand_5 g07239(new_n7624, new_n665, new_n7625);
nand_5 g07240(new_n7625, new_n672, new_n7626);
nand_5 g07241(new_n7626, new_n513, new_n7627);
nand_5 g07242(new_n7627, new_n679, new_n7628);
nand_5 g07243(new_n7628, new_n685, new_n7629);
nand_5 g07244(new_n7629, new_n691, new_n7630);
nand_5 g07245(new_n7630, new_n508, new_n7631);
nand_5 g07246(new_n7631, new_n698, new_n7632);
nand_5 g07247(new_n7632, new_n503, new_n7633);
nand_5 g07248(new_n7633, new_n704, new_n7634);
nand_5 g07249(new_n7634, new_n498_1, new_n7635);
nand_5 g07250(new_n7635, new_n711, new_n7636);
nand_5 g07251(new_n7636, new_n493, new_n7637);
nand_5 g07252(new_n7637, new_n718, new_n7638);
nand_5 g07253(new_n7638, new_n488, new_n7639);
nand_5 g07254(new_n7639, new_n725, new_n7640);
nand_5 g07255(new_n7640, new_n483, new_n7641);
nand_5 g07256(new_n7641, new_n732, new_n7642);
nand_5 g07257(new_n7642, new_n478, new_n7643);
nand_5 g07258(new_n7643, new_n739, new_n7644);
nand_5 g07259(new_n7644, new_n745, new_n7645);
nand_5 g07260(new_n7645, new_n751, new_n7646);
nand_5 g07261(new_n7646, new_n473, new_n7647);
nand_5 g07262(new_n7647, new_n758, new_n7648);
nand_5 g07263(new_n7648, new_n764, new_n7649);
nand_5 g07264(new_n7649, new_n770, new_n7650);
nand_5 g07265(new_n7650, new_n468, new_n7651);
nand_5 g07266(new_n7651, new_n777, new_n7652_1);
nand_5 g07267(new_n7652_1, new_n783, new_n7653);
nand_5 g07268(new_n7653, new_n789, new_n7654);
nand_5 g07269(new_n7654, new_n463, new_n7655_1);
nand_5 g07270(new_n7655_1, new_n796, new_n7656);
nand_5 g07271(new_n7656, new_n458, new_n7657);
nand_5 g07272(new_n7657, new_n453, new_n7658);
nand_5 g07273(new_n7658, new_n447, new_n7659);
nand_5 g07274(new_n7659, new_n805, new_n7660);
nand_5 g07275(new_n7660, new_n811, new_n7661);
nand_5 g07276(new_n7661, new_n442, new_n7662);
nand_5 g07277(new_n7662, new_n437, new_n7663);
nand_5 g07278(new_n7663, new_n819, new_n7664);
nand_5 g07279(new_n7664, new_n432, new_n7665);
nand_5 g07280(new_n7665, new_n427_1, new_n7666);
nand_5 g07281(new_n7666, new_n422, new_n7667_1);
nand_5 g07282(new_n7667_1, new_n828, new_n7668);
nand_5 g07283(new_n7668, new_n834, new_n7669);
nand_5 g07284(new_n7669, new_n840, new_n7670);
nand_5 g07285(new_n7670, new_n417, new_n7671);
nand_5 g07286(new_n7671, new_n847, new_n7672);
nand_5 g07287(new_n7672, new_n853, new_n7673);
nand_5 g07288(new_n7673, new_n859, new_n7674);
nand_5 g07289(new_n7674, n844, new_n7675);
nor_5  g07290(new_n7675, new_n409, n7382);
not_4  g07291(new_n1793, new_n7677);
nand_5 g07292(new_n7677, new_n1017, new_n7678);
nand_5 g07293(new_n7678, new_n1012, new_n7679);
nand_5 g07294(new_n7679, new_n1009, new_n7680);
nand_5 g07295(new_n7680, new_n1004, new_n7681);
nand_5 g07296(new_n7681, new_n1000, new_n7682);
nand_5 g07297(new_n7682, new_n995, new_n7683);
nand_5 g07298(new_n7683, new_n990, new_n7684);
nand_5 g07299(new_n7684, new_n985, new_n7685);
nand_5 g07300(new_n7685, new_n981, new_n7686);
nand_5 g07301(new_n7686, new_n1179, new_n7687);
nand_5 g07302(new_n7687, new_n976, new_n7688);
nand_5 g07303(new_n7688, new_n971, new_n7689);
nand_5 g07304(new_n7689, new_n966, new_n7690);
nand_5 g07305(new_n7690, new_n961, new_n7691);
nand_5 g07306(new_n7691, new_n957, new_n7692);
nand_5 g07307(new_n7692, new_n952, new_n7693);
nand_5 g07308(new_n7693, new_n948_1, new_n7694);
nand_5 g07309(new_n7694, new_n943, new_n7695);
nand_5 g07310(new_n7695, new_n941, new_n7696);
nand_5 g07311(new_n7696, new_n938, new_n7697);
nand_5 g07312(new_n7697, new_n936, new_n7698);
nand_5 g07313(new_n7698, new_n931, new_n7699);
nand_5 g07314(new_n7699, new_n927, new_n7700);
nand_5 g07315(new_n7700, new_n922, new_n7701);
nand_5 g07316(new_n7701, new_n917, new_n7702);
nand_5 g07317(new_n7702, new_n912, new_n7703);
nand_5 g07318(new_n7703, new_n907, new_n7704);
nand_5 g07319(new_n7704, new_n903, new_n7705);
nand_5 g07320(new_n7705, new_n2066, new_n7706);
nand_5 g07321(new_n7706, new_n2063, new_n7707);
nand_5 g07322(new_n7707, new_n2062, new_n7708);
nand_5 g07323(new_n7708, new_n2058, new_n7709);
nand_5 g07324(new_n7709, new_n2055, new_n7710);
nand_5 g07325(new_n7710, new_n2051, new_n7711);
nand_5 g07326(new_n7711, new_n2046, new_n7712);
nand_5 g07327(new_n7712, new_n2042, new_n7713);
nand_5 g07328(new_n7713, new_n2039, new_n7714);
nand_5 g07329(new_n7714, new_n2036, new_n7715);
nand_5 g07330(new_n7715, new_n2033, new_n7716);
nand_5 g07331(new_n7716, new_n2029, new_n7717);
nand_5 g07332(new_n7717, new_n2026, new_n7718);
nand_5 g07333(new_n7718, new_n2022, new_n7719);
nand_5 g07334(new_n7719, new_n2018, new_n7720);
nand_5 g07335(new_n7720, new_n1726, new_n7721);
nand_5 g07336(new_n7721, new_n1722, new_n7722);
nand_5 g07337(new_n7722, new_n1718, new_n7723);
nand_5 g07338(new_n7723, new_n1713, new_n7724);
nand_5 g07339(new_n7724, new_n1737, new_n7725);
nand_5 g07340(new_n7725, new_n1709, new_n7726);
nand_5 g07341(new_n7726, new_n1742, new_n7727);
nand_5 g07342(new_n7727, new_n1704, new_n7728);
nand_5 g07343(new_n7728, new_n1702_1, new_n7729);
nand_5 g07344(new_n7729, new_n1698, new_n7730);
nand_5 g07345(new_n7730, new_n1695, new_n7731);
nand_5 g07346(new_n7731, new_n1692, new_n7732);
nand_5 g07347(new_n7732, new_n1752, new_n7733);
nand_5 g07348(new_n7733, new_n1688, new_n7734);
nand_5 g07349(new_n7734, new_n1685, new_n7735);
nand_5 g07350(new_n7735, new_n1680, new_n7736);
nand_5 g07351(new_n7736, new_n1676, new_n7737);
nand_5 g07352(new_n7737, new_n1672, new_n7738);
nand_5 g07353(new_n7738, new_n1669, new_n7739);
nand_5 g07354(new_n7739, new_n1666, new_n7740);
nand_5 g07355(new_n7740, new_n1663, new_n7741);
nand_5 g07356(new_n7741, new_n1658, new_n7742);
nand_5 g07357(new_n7742, new_n1653, new_n7743);
nand_5 g07358(new_n7743, new_n1651, new_n7744);
nand_5 g07359(new_n7744, new_n1649, new_n7745);
nand_5 g07360(new_n7745, new_n1646, new_n7746);
nand_5 g07361(new_n7746, new_n1643, new_n7747);
nand_5 g07362(new_n7747, new_n1641, new_n7748_1);
nand_5 g07363(new_n7748_1, new_n1638, new_n7749);
nand_5 g07364(new_n7749, new_n1635, new_n7750);
nand_5 g07365(new_n7750, new_n1632, new_n7751);
nand_5 g07366(new_n7751, new_n1628, new_n7752);
nand_5 g07367(new_n7752, new_n1625, new_n7753);
nand_5 g07368(new_n7753, new_n1621, new_n7754);
nand_5 g07369(new_n7754, new_n1618, new_n7755);
nand_5 g07370(new_n7755, new_n1778, new_n7756);
nand_5 g07371(new_n7756, new_n1782, new_n7757);
nand_5 g07372(new_n7757, new_n1614, new_n7758);
nand_5 g07373(new_n7758, new_n1611, new_n7759);
nand_5 g07374(new_n7759, new_n1789, new_n7760);
nand_5 g07375(new_n7760, new_n1608, new_n7761);
nand_5 g07376(new_n7761, n13882, new_n7762);
nor_5  g07377(new_n7762, new_n647, n7655);
nand_5 g07378(new_n1148, new_n1140, new_n7764);
nand_5 g07379(new_n7764, new_n1065, new_n7765);
nand_5 g07380(new_n7765, new_n1062, new_n7766);
nand_5 g07381(new_n7766, new_n1156, new_n7767);
nand_5 g07382(new_n7767, new_n1057, new_n7768);
nand_5 g07383(new_n7768, new_n1053, new_n7769);
nand_5 g07384(new_n7769, new_n1050, new_n7770);
nand_5 g07385(new_n7770, new_n1045, new_n7771_1);
nand_5 g07386(new_n7771_1, new_n1040, new_n7772);
nand_5 g07387(new_n7772, new_n1036, new_n7773);
nand_5 g07388(new_n7773, new_n1033, new_n7774);
nand_5 g07389(new_n7774, new_n1028, new_n7775);
nand_5 g07390(new_n7775, new_n1026, new_n7776);
nand_5 g07391(new_n7776, new_n1021, new_n7777);
nand_5 g07392(new_n7777, new_n1017, new_n7778);
nand_5 g07393(new_n7778, new_n1012, new_n7779);
nand_5 g07394(new_n7779, new_n1009, new_n7780);
nand_5 g07395(new_n7780, new_n1004, new_n7781);
nand_5 g07396(new_n7781, new_n1000, new_n7782);
nand_5 g07397(new_n7782, new_n995, new_n7783);
nand_5 g07398(new_n7783, new_n990, new_n7784);
nand_5 g07399(new_n7784, new_n985, new_n7785);
nand_5 g07400(new_n7785, new_n981, new_n7786);
nand_5 g07401(new_n7786, new_n1179, new_n7787);
nand_5 g07402(new_n7787, new_n976, new_n7788);
nand_5 g07403(new_n7788, new_n971, new_n7789);
nand_5 g07404(new_n7789, new_n966, new_n7790);
nand_5 g07405(new_n7790, new_n961, new_n7791);
nand_5 g07406(new_n7791, new_n957, new_n7792);
nand_5 g07407(new_n7792, new_n952, new_n7793);
nand_5 g07408(new_n7793, new_n948_1, new_n7794);
nand_5 g07409(new_n7794, new_n943, new_n7795);
nand_5 g07410(new_n7795, new_n941, new_n7796);
nand_5 g07411(new_n7796, new_n938, new_n7797);
nand_5 g07412(new_n7797, new_n936, new_n7798);
nand_5 g07413(new_n7798, new_n931, new_n7799);
nand_5 g07414(new_n7799, new_n927, new_n7800);
nand_5 g07415(new_n7800, new_n922, new_n7801);
nand_5 g07416(new_n7801, new_n917, new_n7802);
nand_5 g07417(new_n7802, new_n912, new_n7803);
nand_5 g07418(new_n7803, new_n907, new_n7804);
nand_5 g07419(new_n7804, new_n903, new_n7805);
nand_5 g07420(new_n7805, new_n2066, new_n7806);
nand_5 g07421(new_n7806, new_n2063, new_n7807);
nand_5 g07422(new_n7807, new_n2062, new_n7808);
nand_5 g07423(new_n7808, new_n2058, new_n7809);
nand_5 g07424(new_n7809, new_n2055, new_n7810);
nand_5 g07425(new_n7810, new_n2051, new_n7811);
nand_5 g07426(new_n7811, new_n2046, new_n7812);
nand_5 g07427(new_n7812, new_n2042, new_n7813);
nand_5 g07428(new_n7813, new_n2039, new_n7814);
nand_5 g07429(new_n7814, new_n2036, new_n7815);
nand_5 g07430(new_n7815, new_n2033, new_n7816);
nand_5 g07431(new_n7816, new_n2029, new_n7817);
nand_5 g07432(new_n7817, new_n2026, new_n7818);
nand_5 g07433(new_n7818, new_n2022, new_n7819);
nand_5 g07434(new_n7819, new_n2018, new_n7820);
nand_5 g07435(new_n7820, new_n1726, new_n7821);
nand_5 g07436(new_n7821, new_n1722, new_n7822);
nand_5 g07437(new_n7822, new_n1718, new_n7823);
nand_5 g07438(new_n7823, new_n1713, new_n7824);
nand_5 g07439(new_n7824, new_n1737, new_n7825_1);
nand_5 g07440(new_n7825_1, new_n1709, new_n7826);
nand_5 g07441(new_n7826, new_n1742, new_n7827);
nand_5 g07442(new_n7827, new_n1704, new_n7828);
nand_5 g07443(new_n7828, new_n1702_1, new_n7829);
nand_5 g07444(new_n7829, new_n1698, new_n7830);
nand_5 g07445(new_n7830, new_n1695, new_n7831);
nand_5 g07446(new_n7831, new_n1692, new_n7832_1);
nand_5 g07447(new_n7832_1, new_n1752, new_n7833);
nand_5 g07448(new_n7833, new_n1688, new_n7834);
nand_5 g07449(new_n7834, new_n1685, new_n7835);
nand_5 g07450(new_n7835, new_n1680, new_n7836);
nand_5 g07451(new_n7836, new_n1676, new_n7837);
nand_5 g07452(new_n7837, new_n1672, new_n7838);
nand_5 g07453(new_n7838, new_n1669, new_n7839);
nand_5 g07454(new_n7839, new_n1666, new_n7840);
nand_5 g07455(new_n7840, new_n1663, new_n7841);
nand_5 g07456(new_n7841, new_n1658, new_n7842);
nand_5 g07457(new_n7842, new_n1653, new_n7843);
nand_5 g07458(new_n7843, new_n1651, new_n7844);
nand_5 g07459(new_n7844, new_n1649, new_n7845);
nand_5 g07460(new_n7845, new_n1646, new_n7846);
nand_5 g07461(new_n7846, new_n1643, new_n7847);
nand_5 g07462(new_n7847, n1763, new_n7848);
nor_5  g07463(new_n7848, new_n598, n7771);
nand_5 g07464(new_n2024, new_n1268_1, new_n7850);
nand_5 g07465(new_n7850, new_n2022, new_n7851);
nand_5 g07466(new_n7851, new_n2018, new_n7852);
nand_5 g07467(new_n7852, new_n1726, new_n7853);
nand_5 g07468(new_n7853, new_n1722, new_n7854);
nand_5 g07469(new_n7854, new_n1718, new_n7855);
nand_5 g07470(new_n7855, new_n1713, new_n7856);
nand_5 g07471(new_n7856, new_n1737, new_n7857);
nand_5 g07472(new_n7857, new_n1709, new_n7858);
nand_5 g07473(new_n7858, new_n1742, new_n7859);
nand_5 g07474(new_n7859, new_n1704, new_n7860);
nand_5 g07475(new_n7860, new_n1702_1, new_n7861);
nand_5 g07476(new_n7861, new_n1698, new_n7862);
nand_5 g07477(new_n7862, new_n1695, new_n7863);
nand_5 g07478(new_n7863, new_n1692, new_n7864);
nand_5 g07479(new_n7864, new_n1752, new_n7865);
nand_5 g07480(new_n7865, new_n1688, new_n7866);
nand_5 g07481(new_n7866, new_n1685, new_n7867);
nand_5 g07482(new_n7867, new_n1680, new_n7868);
nand_5 g07483(new_n7868, new_n1676, new_n7869);
nand_5 g07484(new_n7869, new_n1672, new_n7870);
nand_5 g07485(new_n7870, new_n1669, new_n7871);
nand_5 g07486(new_n7871, new_n1666, new_n7872);
nand_5 g07487(new_n7872, new_n1663, new_n7873);
nand_5 g07488(new_n7873, new_n1658, new_n7874);
nand_5 g07489(new_n7874, new_n1653, new_n7875);
nand_5 g07490(new_n7875, new_n1651, new_n7876);
nand_5 g07491(new_n7876, new_n1649, new_n7877);
nand_5 g07492(new_n7877, new_n1646, new_n7878);
nand_5 g07493(new_n7878, new_n1643, new_n7879);
nand_5 g07494(new_n7879, new_n1641, new_n7880);
nand_5 g07495(new_n7880, new_n1638, new_n7881);
nand_5 g07496(new_n7881, new_n1635, new_n7882);
nand_5 g07497(new_n7882, new_n1632, new_n7883);
nand_5 g07498(new_n7883, new_n1628, new_n7884);
nand_5 g07499(new_n7884, new_n1625, new_n7885);
nand_5 g07500(new_n7885, new_n1621, new_n7886);
nand_5 g07501(new_n7886, new_n1618, new_n7887);
nand_5 g07502(new_n7887, new_n1778, new_n7888);
nand_5 g07503(new_n7888, new_n1782, new_n7889);
nand_5 g07504(new_n7889, new_n1614, new_n7890);
nand_5 g07505(new_n7890, new_n1611, new_n7891);
nand_5 g07506(new_n7891, new_n1789, new_n7892);
nand_5 g07507(new_n7892, new_n1608, new_n7893);
nand_5 g07508(new_n7893, new_n1605, new_n7894);
nand_5 g07509(new_n7894, new_n1795, new_n7895);
nand_5 g07510(new_n7895, new_n1799, new_n7896);
nand_5 g07511(new_n7896, new_n1602, new_n7897);
nand_5 g07512(new_n7897, new_n1599, new_n7898);
nand_5 g07513(new_n7898, new_n1596, new_n7899);
nand_5 g07514(new_n7899, new_n1593, new_n7900);
nand_5 g07515(new_n7900, new_n1806, new_n7901);
nand_5 g07516(new_n7901, new_n1589, new_n7902);
nand_5 g07517(new_n7902, new_n1586, new_n7903);
nand_5 g07518(new_n7903, new_n1583, new_n7904);
nand_5 g07519(new_n7904, new_n1580, new_n7905);
nand_5 g07520(new_n7905, new_n1576, new_n7906);
nand_5 g07521(new_n7906, new_n1573, new_n7907);
nand_5 g07522(new_n7907, new_n1570, new_n7908);
nand_5 g07523(new_n7908, new_n1567, new_n7909);
nand_5 g07524(new_n7909, new_n1564, new_n7910);
nand_5 g07525(new_n7910, new_n1561, new_n7911);
nand_5 g07526(new_n7911, new_n1338, new_n7912);
nand_5 g07527(new_n7912, new_n1331, new_n7913);
nand_5 g07528(new_n7913, new_n1326, new_n7914);
nand_5 g07529(new_n7914, new_n1321, new_n7915);
nand_5 g07530(new_n7915, new_n1318, new_n7916);
nand_5 g07531(new_n7916, new_n1315, new_n7917);
nand_5 g07532(new_n7917, new_n1312, new_n7918);
nand_5 g07533(new_n7918, new_n1309, new_n7919);
nand_5 g07534(new_n7919, new_n1307, new_n7920);
nand_5 g07535(new_n7920, new_n1304, new_n7921);
nand_5 g07536(new_n7921, new_n1300, new_n7922);
nand_5 g07537(new_n7922, new_n1297, new_n7923);
nand_5 g07538(new_n7923, new_n1294, new_n7924);
nand_5 g07539(new_n7924, new_n1355, new_n7925);
nand_5 g07540(new_n7925, new_n1291, new_n7926);
nand_5 g07541(new_n7926, new_n1288, new_n7927);
nand_5 g07542(new_n7927, new_n1283, new_n7928);
nand_5 g07543(new_n7928, new_n1363, new_n7929);
nand_5 g07544(new_n7929, new_n1280, new_n7930);
nand_5 g07545(new_n7930, new_n1370, new_n7931);
nand_5 g07546(new_n7931, new_n1373, new_n7932);
nand_5 g07547(new_n7932, new_n1277, new_n7933);
nand_5 g07548(new_n7933, n11404, new_n7934);
nor_5  g07549(new_n7934, new_n802, n7825);
not_4  g07550(n12009, new_n7936);
nand_5 g07551(new_n1141, new_n7936, new_n7937);
nand_5 g07552(new_n7937, new_n561, new_n7938);
nand_5 g07553(new_n7938, new_n608, new_n7939);
nand_5 g07554(new_n7939, new_n558, new_n7940);
nand_5 g07555(new_n7940, new_n615, new_n7941_1);
nand_5 g07556(new_n7941_1, new_n553, new_n7942);
nand_5 g07557(new_n7942, new_n622, new_n7943);
nand_5 g07558(new_n7943, new_n628, new_n7944);
nand_5 g07559(new_n7944, new_n548, new_n7945);
nand_5 g07560(new_n7945, new_n543_1, new_n7946);
nand_5 g07561(new_n7946, new_n636, new_n7947);
nand_5 g07562(new_n7947, new_n642, new_n7948);
nand_5 g07563(new_n7948, new_n538, new_n7949);
nand_5 g07564(new_n7949, new_n533, new_n7950);
nand_5 g07565(new_n7950, new_n650_1, new_n7951);
nand_5 g07566(new_n7951, new_n528, new_n7952);
nand_5 g07567(new_n7952, new_n523, new_n7953);
nand_5 g07568(new_n7953, new_n518, new_n7954);
nand_5 g07569(new_n7954, new_n659, new_n7955);
nand_5 g07570(new_n7955, new_n665, new_n7956);
nand_5 g07571(new_n7956, new_n672, new_n7957);
nand_5 g07572(new_n7957, new_n513, new_n7958);
nand_5 g07573(new_n7958, new_n679, new_n7959);
nand_5 g07574(new_n7959, new_n685, new_n7960);
nand_5 g07575(new_n7960, new_n691, new_n7961);
nand_5 g07576(new_n7961, new_n508, new_n7962);
nand_5 g07577(new_n7962, new_n698, new_n7963);
nand_5 g07578(new_n7963, new_n503, new_n7964);
nand_5 g07579(new_n7964, new_n704, new_n7965);
nand_5 g07580(new_n7965, new_n498_1, new_n7966);
nand_5 g07581(new_n7966, new_n711, new_n7967);
nand_5 g07582(new_n7967, new_n493, new_n7968);
nand_5 g07583(new_n7968, new_n718, new_n7969);
nand_5 g07584(new_n7969, new_n488, new_n7970);
nand_5 g07585(new_n7970, new_n725, new_n7971);
nand_5 g07586(new_n7971, new_n483, new_n7972_1);
nand_5 g07587(new_n7972_1, new_n732, new_n7973);
nand_5 g07588(new_n7973, new_n478, new_n7974);
nand_5 g07589(new_n7974, new_n739, new_n7975);
nand_5 g07590(new_n7975, new_n745, new_n7976);
nand_5 g07591(new_n7976, new_n751, new_n7977);
nand_5 g07592(new_n7977, new_n473, new_n7978);
nand_5 g07593(new_n7978, new_n758, new_n7979);
nand_5 g07594(new_n7979, new_n764, new_n7980);
nand_5 g07595(new_n7980, new_n770, new_n7981);
nand_5 g07596(new_n7981, new_n468, new_n7982);
nand_5 g07597(new_n7982, new_n777, new_n7983);
nand_5 g07598(new_n7983, new_n783, new_n7984);
nand_5 g07599(new_n7984, new_n789, new_n7985);
nand_5 g07600(new_n7985, new_n463, new_n7986);
nand_5 g07601(new_n7986, new_n796, new_n7987);
nand_5 g07602(new_n7987, new_n458, new_n7988_1);
nand_5 g07603(new_n7988_1, new_n453, new_n7989);
nand_5 g07604(new_n7989, new_n447, new_n7990);
nand_5 g07605(new_n7990, new_n805, new_n7991);
nand_5 g07606(new_n7991, new_n811, new_n7992);
nand_5 g07607(new_n7992, new_n442, new_n7993);
nand_5 g07608(new_n7993, new_n437, new_n7994);
nand_5 g07609(new_n7994, new_n819, new_n7995);
nand_5 g07610(new_n7995, new_n432, new_n7996);
nand_5 g07611(new_n7996, new_n427_1, new_n7997);
nand_5 g07612(new_n7997, new_n422, new_n7998);
nand_5 g07613(new_n7998, new_n828, new_n7999);
nand_5 g07614(new_n7999, new_n834, new_n8000);
nand_5 g07615(new_n8000, new_n840, new_n8001);
nand_5 g07616(new_n8001, new_n417, new_n8002_1);
nand_5 g07617(new_n8002_1, new_n847, new_n8003);
nand_5 g07618(new_n8003, new_n853, new_n8004);
nand_5 g07619(new_n8004, new_n859, new_n8005);
nand_5 g07620(new_n8005, new_n412, new_n8006);
nand_5 g07621(new_n8006, new_n866, new_n8007);
nand_5 g07622(new_n8007, new_n872, new_n8008);
nand_5 g07623(new_n8008, new_n878, new_n8009);
nand_5 g07624(new_n8009, new_n407, new_n8010);
nand_5 g07625(new_n8010, new_n885, new_n8011);
nand_5 g07626(new_n8011, new_n402, new_n8012);
nand_5 g07627(new_n8012, new_n397, new_n8013);
nand_5 g07628(new_n8013, new_n392, new_n8014);
nand_5 g07629(new_n8014, new_n894, new_n8015);
nand_5 g07630(new_n8015, new_n1087, new_n8016);
nand_5 g07631(new_n8016, new_n1129, new_n8017);
nand_5 g07632(new_n8017, new_n1084, new_n8018);
nand_5 g07633(new_n8018, new_n1134, new_n8019);
nand_5 g07634(new_n8019, new_n1080, new_n8020);
nand_5 g07635(new_n8020, new_n1075, new_n8021);
nand_5 g07636(new_n8021, n13363, new_n8022);
nor_5  g07637(new_n8022, new_n1067, n8068);
nand_5 g07638(new_n1579, new_n974, new_n8024);
nand_5 g07639(new_n8024, new_n971, new_n8025);
nand_5 g07640(new_n8025, new_n966, new_n8026);
nand_5 g07641(new_n8026, new_n961, new_n8027);
nand_5 g07642(new_n8027, new_n957, new_n8028);
nand_5 g07643(new_n8028, new_n952, new_n8029);
nand_5 g07644(new_n8029, new_n948_1, new_n8030);
nand_5 g07645(new_n8030, new_n943, new_n8031);
nand_5 g07646(new_n8031, new_n941, new_n8032);
nand_5 g07647(new_n8032, new_n938, new_n8033);
nand_5 g07648(new_n8033, new_n936, new_n8034);
nand_5 g07649(new_n8034, new_n931, new_n8035);
nand_5 g07650(new_n8035, new_n927, new_n8036);
nand_5 g07651(new_n8036, new_n922, new_n8037);
nand_5 g07652(new_n8037, new_n917, new_n8038);
nand_5 g07653(new_n8038, new_n912, new_n8039);
nand_5 g07654(new_n8039, new_n907, new_n8040);
nand_5 g07655(new_n8040, new_n903, new_n8041);
nand_5 g07656(new_n8041, new_n2066, new_n8042);
nand_5 g07657(new_n8042, new_n2063, new_n8043);
nand_5 g07658(new_n8043, new_n2062, new_n8044_1);
nand_5 g07659(new_n8044_1, new_n2058, new_n8045);
nand_5 g07660(new_n8045, new_n2055, new_n8046);
nand_5 g07661(new_n8046, new_n2051, new_n8047);
nand_5 g07662(new_n8047, new_n2046, new_n8048);
nand_5 g07663(new_n8048, new_n2042, new_n8049);
nand_5 g07664(new_n8049, new_n2039, new_n8050);
nand_5 g07665(new_n8050, new_n2036, new_n8051);
nand_5 g07666(new_n8051, new_n2033, new_n8052);
nand_5 g07667(new_n8052, new_n2029, new_n8053);
nand_5 g07668(new_n8053, new_n2026, new_n8054);
nand_5 g07669(new_n8054, new_n2022, new_n8055);
nand_5 g07670(new_n8055, new_n2018, new_n8056);
nand_5 g07671(new_n8056, new_n1726, new_n8057);
nand_5 g07672(new_n8057, new_n1722, new_n8058);
nand_5 g07673(new_n8058, new_n1718, new_n8059);
nand_5 g07674(new_n8059, new_n1713, new_n8060);
nand_5 g07675(new_n8060, new_n1737, new_n8061);
nand_5 g07676(new_n8061, new_n1709, new_n8062);
nand_5 g07677(new_n8062, new_n1742, new_n8063);
nand_5 g07678(new_n8063, new_n1704, new_n8064);
nand_5 g07679(new_n8064, new_n1702_1, new_n8065);
nand_5 g07680(new_n8065, new_n1698, new_n8066);
nand_5 g07681(new_n8066, new_n1695, new_n8067);
nand_5 g07682(new_n8067, new_n1692, new_n8068_1);
nand_5 g07683(new_n8068_1, new_n1752, new_n8069);
nand_5 g07684(new_n8069, new_n1688, new_n8070);
nand_5 g07685(new_n8070, new_n1685, new_n8071);
nand_5 g07686(new_n8071, new_n1680, new_n8072);
nand_5 g07687(new_n8072, new_n1676, new_n8073_1);
nand_5 g07688(new_n8073_1, new_n1672, new_n8074);
nand_5 g07689(new_n8074, new_n1669, new_n8075);
nand_5 g07690(new_n8075, new_n1666, new_n8076);
nand_5 g07691(new_n8076, new_n1663, new_n8077);
nand_5 g07692(new_n8077, new_n1658, new_n8078);
nand_5 g07693(new_n8078, new_n1653, new_n8079);
nand_5 g07694(new_n8079, new_n1651, new_n8080);
nand_5 g07695(new_n8080, new_n1649, new_n8081);
nand_5 g07696(new_n8081, new_n1646, new_n8082);
nand_5 g07697(new_n8082, new_n1643, new_n8083);
nand_5 g07698(new_n8083, new_n1641, new_n8084);
nand_5 g07699(new_n8084, new_n1638, new_n8085_1);
nand_5 g07700(new_n8085_1, new_n1635, new_n8086);
nand_5 g07701(new_n8086, new_n1632, new_n8087);
nand_5 g07702(new_n8087, new_n1628, new_n8088);
nand_5 g07703(new_n8088, new_n1625, new_n8089);
nand_5 g07704(new_n8089, new_n1621, new_n8090);
nand_5 g07705(new_n8090, new_n1618, new_n8091);
nand_5 g07706(new_n8091, new_n1778, new_n8092);
nand_5 g07707(new_n8092, new_n1782, new_n8093);
nand_5 g07708(new_n8093, new_n1614, new_n8094);
nand_5 g07709(new_n8094, new_n1611, new_n8095);
nand_5 g07710(new_n8095, new_n1789, new_n8096);
nand_5 g07711(new_n8096, new_n1608, new_n8097);
nand_5 g07712(new_n8097, new_n1605, new_n8098);
nand_5 g07713(new_n8098, new_n1795, new_n8099);
nand_5 g07714(new_n8099, new_n1799, new_n8100);
nand_5 g07715(new_n8100, new_n1602, new_n8101);
nand_5 g07716(new_n8101, new_n1599, new_n8102);
nand_5 g07717(new_n8102, new_n1596, new_n8103);
nand_5 g07718(new_n8103, new_n1593, new_n8104);
nand_5 g07719(new_n8104, new_n1806, new_n8105);
nand_5 g07720(new_n8105, new_n1589, new_n8106);
nand_5 g07721(new_n8106, new_n1586, new_n8107);
nand_5 g07722(new_n8107, n8800, new_n8108);
nor_5  g07723(new_n8108, new_n688, n8085);
nand_5 g07724(new_n1560, new_n946, new_n8110);
nand_5 g07725(new_n8110, new_n943, new_n8111);
nand_5 g07726(new_n8111, new_n941, new_n8112);
nand_5 g07727(new_n8112, new_n938, new_n8113);
nand_5 g07728(new_n8113, new_n936, new_n8114);
nand_5 g07729(new_n8114, new_n931, new_n8115);
nand_5 g07730(new_n8115, new_n927, new_n8116);
nand_5 g07731(new_n8116, new_n922, new_n8117);
nand_5 g07732(new_n8117, new_n917, new_n8118);
nand_5 g07733(new_n8118, new_n912, new_n8119);
nand_5 g07734(new_n8119, new_n907, new_n8120);
nand_5 g07735(new_n8120, new_n903, new_n8121);
nand_5 g07736(new_n8121, new_n2066, new_n8122);
nand_5 g07737(new_n8122, new_n2063, new_n8123);
nand_5 g07738(new_n8123, new_n2062, new_n8124_1);
nand_5 g07739(new_n8124_1, new_n2058, new_n8125);
nand_5 g07740(new_n8125, new_n2055, new_n8126);
nand_5 g07741(new_n8126, new_n2051, new_n8127);
nand_5 g07742(new_n8127, new_n2046, new_n8128);
nand_5 g07743(new_n8128, new_n2042, new_n8129);
nand_5 g07744(new_n8129, new_n2039, new_n8130);
nand_5 g07745(new_n8130, new_n2036, new_n8131);
nand_5 g07746(new_n8131, new_n2033, new_n8132);
nand_5 g07747(new_n8132, new_n2029, new_n8133);
nand_5 g07748(new_n8133, new_n2026, new_n8134);
nand_5 g07749(new_n8134, new_n2022, new_n8135);
nand_5 g07750(new_n8135, new_n2018, new_n8136);
nand_5 g07751(new_n8136, new_n1726, new_n8137);
nand_5 g07752(new_n8137, new_n1722, new_n8138);
nand_5 g07753(new_n8138, new_n1718, new_n8139);
nand_5 g07754(new_n8139, new_n1713, new_n8140);
nand_5 g07755(new_n8140, new_n1737, new_n8141);
nand_5 g07756(new_n8141, new_n1709, new_n8142);
nand_5 g07757(new_n8142, new_n1742, new_n8143);
nand_5 g07758(new_n8143, new_n1704, new_n8144_1);
nand_5 g07759(new_n8144_1, new_n1702_1, new_n8145);
nand_5 g07760(new_n8145, new_n1698, new_n8146);
nand_5 g07761(new_n8146, new_n1695, new_n8147);
nand_5 g07762(new_n8147, new_n1692, new_n8148);
nand_5 g07763(new_n8148, new_n1752, new_n8149);
nand_5 g07764(new_n8149, new_n1688, new_n8150);
nand_5 g07765(new_n8150, new_n1685, new_n8151);
nand_5 g07766(new_n8151, new_n1680, new_n8152);
nand_5 g07767(new_n8152, new_n1676, new_n8153);
nand_5 g07768(new_n8153, new_n1672, new_n8154);
nand_5 g07769(new_n8154, new_n1669, new_n8155);
nand_5 g07770(new_n8155, new_n1666, new_n8156);
nand_5 g07771(new_n8156, new_n1663, new_n8157);
nand_5 g07772(new_n8157, new_n1658, new_n8158);
nand_5 g07773(new_n8158, new_n1653, new_n8159);
nand_5 g07774(new_n8159, new_n1651, new_n8160);
nand_5 g07775(new_n8160, new_n1649, new_n8161);
nand_5 g07776(new_n8161, new_n1646, new_n8162);
nand_5 g07777(new_n8162, new_n1643, new_n8163);
nand_5 g07778(new_n8163, new_n1641, new_n8164);
nand_5 g07779(new_n8164, new_n1638, new_n8165);
nand_5 g07780(new_n8165, new_n1635, new_n8166);
nand_5 g07781(new_n8166, new_n1632, new_n8167);
nand_5 g07782(new_n8167, new_n1628, new_n8168);
nand_5 g07783(new_n8168, new_n1625, new_n8169);
nand_5 g07784(new_n8169, new_n1621, new_n8170);
nand_5 g07785(new_n8170, new_n1618, new_n8171);
nand_5 g07786(new_n8171, new_n1778, new_n8172);
nand_5 g07787(new_n8172, new_n1782, new_n8173);
nand_5 g07788(new_n8173, new_n1614, new_n8174);
nand_5 g07789(new_n8174, new_n1611, new_n8175);
nand_5 g07790(new_n8175, new_n1789, new_n8176);
nand_5 g07791(new_n8176, new_n1608, new_n8177);
nand_5 g07792(new_n8177, new_n1605, new_n8178);
nand_5 g07793(new_n8178, new_n1795, new_n8179);
nand_5 g07794(new_n8179, new_n1799, new_n8180);
nand_5 g07795(new_n8180, new_n1602, new_n8181);
nand_5 g07796(new_n8181, new_n1599, new_n8182);
nand_5 g07797(new_n8182, new_n1596, new_n8183);
nand_5 g07798(new_n8183, new_n1593, new_n8184);
nand_5 g07799(new_n8184, new_n1806, new_n8185);
nand_5 g07800(new_n8185, new_n1589, new_n8186);
nand_5 g07801(new_n8186, new_n1586, new_n8187);
nand_5 g07802(new_n8187, new_n1583, new_n8188);
nand_5 g07803(new_n8188, new_n1580, new_n8189);
nand_5 g07804(new_n8189, new_n1576, new_n8190);
nand_5 g07805(new_n8190, new_n1573, new_n8191);
nand_5 g07806(new_n8191, new_n1570, new_n8192);
nand_5 g07807(new_n8192, new_n1567, new_n8193);
nand_5 g07808(new_n8193, n9154, new_n8194);
nor_5  g07809(new_n8194, new_n708, n8124);
not_4  g07810(new_n892, new_n8196);
nand_5 g07811(new_n1203, new_n8196, new_n8197);
nand_5 g07812(new_n8197, new_n1433, new_n8198);
nand_5 g07813(new_n8198, new_n581, new_n8199);
nand_5 g07814(new_n8199, new_n574, new_n8200);
nand_5 g07815(new_n8200, new_n568, new_n8201);
nand_5 g07816(new_n8201, new_n589, new_n8202);
nand_5 g07817(new_n8202, new_n595, new_n8203);
nand_5 g07818(new_n8203, new_n601, new_n8204_1);
nand_5 g07819(new_n8204_1, new_n563, new_n8205);
nand_5 g07820(new_n8205, new_n608, new_n8206);
nand_5 g07821(new_n8206, new_n558, new_n8207);
nand_5 g07822(new_n8207, new_n615, new_n8208);
nand_5 g07823(new_n8208, new_n553, new_n8209);
nand_5 g07824(new_n8209, new_n622, new_n8210);
nand_5 g07825(new_n8210, new_n628, new_n8211);
nand_5 g07826(new_n8211, new_n548, new_n8212);
nand_5 g07827(new_n8212, new_n543_1, new_n8213);
nand_5 g07828(new_n8213, new_n636, new_n8214);
nand_5 g07829(new_n8214, new_n642, new_n8215_1);
nand_5 g07830(new_n8215_1, new_n538, new_n8216);
nand_5 g07831(new_n8216, new_n533, new_n8217);
nand_5 g07832(new_n8217, new_n650_1, new_n8218);
nand_5 g07833(new_n8218, new_n528, new_n8219);
nand_5 g07834(new_n8219, new_n523, new_n8220);
nand_5 g07835(new_n8220, new_n518, new_n8221);
nand_5 g07836(new_n8221, new_n659, new_n8222);
nand_5 g07837(new_n8222, new_n665, new_n8223);
nand_5 g07838(new_n8223, new_n672, new_n8224);
nand_5 g07839(new_n8224, new_n513, new_n8225);
nand_5 g07840(new_n8225, new_n679, new_n8226);
nand_5 g07841(new_n8226, new_n685, new_n8227);
nand_5 g07842(new_n8227, new_n691, new_n8228);
nand_5 g07843(new_n8228, new_n508, new_n8229);
nand_5 g07844(new_n8229, new_n698, new_n8230);
nand_5 g07845(new_n8230, new_n503, new_n8231);
nand_5 g07846(new_n8231, new_n704, new_n8232);
nand_5 g07847(new_n8232, new_n498_1, new_n8233);
nand_5 g07848(new_n8233, new_n711, new_n8234);
nand_5 g07849(new_n8234, new_n493, new_n8235);
nand_5 g07850(new_n8235, new_n718, new_n8236);
nand_5 g07851(new_n8236, new_n488, new_n8237);
nand_5 g07852(new_n8237, new_n725, new_n8238);
nand_5 g07853(new_n8238, new_n483, new_n8239);
nand_5 g07854(new_n8239, new_n732, new_n8240);
nand_5 g07855(new_n8240, new_n478, new_n8241);
nand_5 g07856(new_n8241, new_n739, new_n8242);
nand_5 g07857(new_n8242, new_n745, new_n8243);
nand_5 g07858(new_n8243, new_n751, new_n8244);
nand_5 g07859(new_n8244, new_n473, new_n8245);
nand_5 g07860(new_n8245, new_n758, new_n8246);
nand_5 g07861(new_n8246, new_n764, new_n8247);
nand_5 g07862(new_n8247, new_n770, new_n8248);
nand_5 g07863(new_n8248, new_n468, new_n8249);
nand_5 g07864(new_n8249, new_n777, new_n8250);
nand_5 g07865(new_n8250, new_n783, new_n8251);
nand_5 g07866(new_n8251, new_n789, new_n8252);
nand_5 g07867(new_n8252, new_n463, new_n8253);
nand_5 g07868(new_n8253, new_n796, new_n8254);
nand_5 g07869(new_n8254, new_n458, new_n8255);
nand_5 g07870(new_n8255, new_n453, new_n8256);
nand_5 g07871(new_n8256, new_n447, new_n8257);
nand_5 g07872(new_n8257, new_n805, new_n8258);
nand_5 g07873(new_n8258, new_n811, new_n8259);
nand_5 g07874(new_n8259, new_n442, new_n8260);
nand_5 g07875(new_n8260, new_n437, new_n8261);
nand_5 g07876(new_n8261, new_n819, new_n8262_1);
nand_5 g07877(new_n8262_1, new_n432, new_n8263);
nand_5 g07878(new_n8263, new_n427_1, new_n8264);
nand_5 g07879(new_n8264, new_n422, new_n8265);
nand_5 g07880(new_n8265, new_n828, new_n8266);
nand_5 g07881(new_n8266, new_n834, new_n8267);
nand_5 g07882(new_n8267, new_n840, new_n8268);
nand_5 g07883(new_n8268, new_n417, new_n8269);
nand_5 g07884(new_n8269, new_n847, new_n8270);
nand_5 g07885(new_n8270, new_n853, new_n8271);
nand_5 g07886(new_n8271, new_n859, new_n8272);
nand_5 g07887(new_n8272, new_n412, new_n8273);
nand_5 g07888(new_n8273, new_n866, new_n8274);
nand_5 g07889(new_n8274, new_n872, new_n8275);
nand_5 g07890(new_n8275, new_n878, new_n8276);
nand_5 g07891(new_n8276, new_n407, new_n8277);
nand_5 g07892(new_n8277, new_n885, new_n8278);
nand_5 g07893(new_n8278, new_n402, new_n8279);
nand_5 g07894(new_n8279, new_n397, new_n8280);
nand_5 g07895(new_n8280, n8780, new_n8281);
nor_5  g07896(new_n8281, new_n389_1, n8144);
not_4  g07897(new_n939, new_n8283);
nand_5 g07898(new_n937, new_n481, new_n8284);
nand_5 g07899(new_n8284, new_n732, new_n8285);
nand_5 g07900(new_n8285, new_n478, new_n8286);
nand_5 g07901(new_n8286, new_n739, new_n8287);
nand_5 g07902(new_n8287, new_n745, new_n8288);
nand_5 g07903(new_n8288, new_n751, new_n8289);
nand_5 g07904(new_n8289, new_n473, new_n8290);
nand_5 g07905(new_n8290, new_n758, new_n8291);
nand_5 g07906(new_n8291, new_n764, new_n8292);
nand_5 g07907(new_n8292, new_n770, new_n8293);
nand_5 g07908(new_n8293, new_n468, new_n8294);
nand_5 g07909(new_n8294, new_n777, new_n8295);
nand_5 g07910(new_n8295, new_n783, new_n8296);
nand_5 g07911(new_n8296, new_n789, new_n8297);
nand_5 g07912(new_n8297, new_n463, new_n8298);
nand_5 g07913(new_n8298, new_n796, new_n8299);
nand_5 g07914(new_n8299, new_n458, new_n8300);
nand_5 g07915(new_n8300, new_n453, new_n8301);
nand_5 g07916(new_n8301, new_n447, new_n8302_1);
nand_5 g07917(new_n8302_1, new_n805, new_n8303);
nand_5 g07918(new_n8303, new_n811, new_n8304);
nand_5 g07919(new_n8304, new_n442, new_n8305);
nand_5 g07920(new_n8305, new_n437, new_n8306_1);
nand_5 g07921(new_n8306_1, new_n819, new_n8307);
nand_5 g07922(new_n8307, new_n432, new_n8308);
nand_5 g07923(new_n8308, new_n427_1, new_n8309);
nand_5 g07924(new_n8309, new_n422, new_n8310);
nand_5 g07925(new_n8310, new_n828, new_n8311);
nand_5 g07926(new_n8311, new_n834, new_n8312);
nand_5 g07927(new_n8312, new_n840, new_n8313);
nand_5 g07928(new_n8313, new_n417, new_n8314);
nand_5 g07929(new_n8314, new_n847, new_n8315_1);
nand_5 g07930(new_n8315_1, new_n853, new_n8316);
nand_5 g07931(new_n8316, new_n859, new_n8317);
nand_5 g07932(new_n8317, new_n412, new_n8318);
nand_5 g07933(new_n8318, new_n866, new_n8319);
nand_5 g07934(new_n8319, new_n872, new_n8320);
nand_5 g07935(new_n8320, new_n878, new_n8321);
nand_5 g07936(new_n8321, new_n407, new_n8322);
nand_5 g07937(new_n8322, new_n885, new_n8323);
nand_5 g07938(new_n8323, new_n402, new_n8324);
nand_5 g07939(new_n8324, new_n397, new_n8325);
nand_5 g07940(new_n8325, new_n392, new_n8326);
nand_5 g07941(new_n8326, new_n894, new_n8327);
nand_5 g07942(new_n8327, new_n1087, new_n8328);
nand_5 g07943(new_n8328, new_n1129, new_n8329);
nand_5 g07944(new_n8329, new_n1084, new_n8330);
nand_5 g07945(new_n8330, new_n1134, new_n8331);
nand_5 g07946(new_n8331, new_n1080, new_n8332);
nand_5 g07947(new_n8332, new_n1075, new_n8333);
nand_5 g07948(new_n8333, new_n1070, new_n8334);
nand_5 g07949(new_n8334, new_n1143, new_n8335);
nand_5 g07950(new_n8335, new_n1148, new_n8336);
nand_5 g07951(new_n8336, new_n1065, new_n8337);
nand_5 g07952(new_n8337, new_n1062, new_n8338);
nand_5 g07953(new_n8338, new_n1156, new_n8339);
nand_5 g07954(new_n8339, new_n1057, new_n8340);
nand_5 g07955(new_n8340, new_n1053, new_n8341);
nand_5 g07956(new_n8341, new_n1050, new_n8342);
nand_5 g07957(new_n8342, new_n1045, new_n8343);
nand_5 g07958(new_n8343, new_n1040, new_n8344);
nand_5 g07959(new_n8344, new_n1036, new_n8345);
nand_5 g07960(new_n8345, new_n1033, new_n8346);
nand_5 g07961(new_n8346, new_n1028, new_n8347);
nand_5 g07962(new_n8347, new_n1026, new_n8348);
nand_5 g07963(new_n8348, new_n1021, new_n8349);
nand_5 g07964(new_n8349, new_n1017, new_n8350);
nand_5 g07965(new_n8350, new_n1012, new_n8351);
nand_5 g07966(new_n8351, new_n1009, new_n8352);
nand_5 g07967(new_n8352, new_n1004, new_n8353);
nand_5 g07968(new_n8353, new_n1000, new_n8354);
nand_5 g07969(new_n8354, new_n995, new_n8355);
nand_5 g07970(new_n8355, new_n990, new_n8356);
nand_5 g07971(new_n8356, new_n985, new_n8357);
nand_5 g07972(new_n8357, new_n981, new_n8358);
nand_5 g07973(new_n8358, new_n1179, new_n8359);
nand_5 g07974(new_n8359, new_n976, new_n8360);
nand_5 g07975(new_n8360, new_n971, new_n8361);
nand_5 g07976(new_n8361, new_n966, new_n8362);
nand_5 g07977(new_n8362, new_n961, new_n8363);
nand_5 g07978(new_n8363, new_n957, new_n8364);
nand_5 g07979(new_n8364, new_n952, new_n8365);
nand_5 g07980(new_n8365, new_n948_1, new_n8366);
nand_5 g07981(new_n8366, new_n943, new_n8367);
nand_5 g07982(new_n8367, n10407, new_n8368);
nor_5  g07983(new_n8368, new_n8283, n8215);
not_4  g07984(n656, new_n8370);
nand_5 g07985(new_n1286, new_n8370, new_n8371);
nand_5 g07986(new_n8371, new_n2053, new_n8372);
nand_5 g07987(new_n8372, new_n2051, new_n8373);
nand_5 g07988(new_n8373, new_n2046, new_n8374);
nand_5 g07989(new_n8374, new_n2042, new_n8375);
nand_5 g07990(new_n8375, new_n2039, new_n8376);
nand_5 g07991(new_n8376, new_n2036, new_n8377);
nand_5 g07992(new_n8377, new_n2033, new_n8378);
nand_5 g07993(new_n8378, new_n2029, new_n8379);
nand_5 g07994(new_n8379, new_n2026, new_n8380);
nand_5 g07995(new_n8380, new_n2022, new_n8381);
nand_5 g07996(new_n8381, new_n2018, new_n8382);
nand_5 g07997(new_n8382, new_n1726, new_n8383);
nand_5 g07998(new_n8383, new_n1722, new_n8384);
nand_5 g07999(new_n8384, new_n1718, new_n8385);
nand_5 g08000(new_n8385, new_n1713, new_n8386);
nand_5 g08001(new_n8386, new_n1737, new_n8387);
nand_5 g08002(new_n8387, new_n1709, new_n8388);
nand_5 g08003(new_n8388, new_n1742, new_n8389);
nand_5 g08004(new_n8389, new_n1704, new_n8390);
nand_5 g08005(new_n8390, new_n1702_1, new_n8391);
nand_5 g08006(new_n8391, new_n1698, new_n8392);
nand_5 g08007(new_n8392, new_n1695, new_n8393);
nand_5 g08008(new_n8393, new_n1692, new_n8394);
nand_5 g08009(new_n8394, new_n1752, new_n8395);
nand_5 g08010(new_n8395, new_n1688, new_n8396);
nand_5 g08011(new_n8396, new_n1685, new_n8397_1);
nand_5 g08012(new_n8397_1, new_n1680, new_n8398);
nand_5 g08013(new_n8398, new_n1676, new_n8399);
nand_5 g08014(new_n8399, new_n1672, new_n8400);
nand_5 g08015(new_n8400, new_n1669, new_n8401);
nand_5 g08016(new_n8401, new_n1666, new_n8402);
nand_5 g08017(new_n8402, new_n1663, new_n8403);
nand_5 g08018(new_n8403, new_n1658, new_n8404);
nand_5 g08019(new_n8404, new_n1653, new_n8405);
nand_5 g08020(new_n8405, new_n1651, new_n8406);
nand_5 g08021(new_n8406, new_n1649, new_n8407);
nand_5 g08022(new_n8407, new_n1646, new_n8408);
nand_5 g08023(new_n8408, new_n1643, new_n8409);
nand_5 g08024(new_n8409, new_n1641, new_n8410);
nand_5 g08025(new_n8410, new_n1638, new_n8411);
nand_5 g08026(new_n8411, new_n1635, new_n8412);
nand_5 g08027(new_n8412, new_n1632, new_n8413);
nand_5 g08028(new_n8413, new_n1628, new_n8414);
nand_5 g08029(new_n8414, new_n1625, new_n8415);
nand_5 g08030(new_n8415, new_n1621, new_n8416);
nand_5 g08031(new_n8416, new_n1618, new_n8417);
nand_5 g08032(new_n8417, new_n1778, new_n8418);
nand_5 g08033(new_n8418, new_n1782, new_n8419);
nand_5 g08034(new_n8419, new_n1614, new_n8420);
nand_5 g08035(new_n8420, new_n1611, new_n8421);
nand_5 g08036(new_n8421, new_n1789, new_n8422);
nand_5 g08037(new_n8422, new_n1608, new_n8423);
nand_5 g08038(new_n8423, new_n1605, new_n8424);
nand_5 g08039(new_n8424, new_n1795, new_n8425);
nand_5 g08040(new_n8425, new_n1799, new_n8426);
nand_5 g08041(new_n8426, new_n1602, new_n8427);
nand_5 g08042(new_n8427, new_n1599, new_n8428);
nand_5 g08043(new_n8428, new_n1596, new_n8429);
nand_5 g08044(new_n8429, new_n1593, new_n8430);
nand_5 g08045(new_n8430, new_n1806, new_n8431);
nand_5 g08046(new_n8431, new_n1589, new_n8432);
nand_5 g08047(new_n8432, new_n1586, new_n8433);
nand_5 g08048(new_n8433, new_n1583, new_n8434);
nand_5 g08049(new_n8434, new_n1580, new_n8435);
nand_5 g08050(new_n8435, new_n1576, new_n8436);
nand_5 g08051(new_n8436, new_n1573, new_n8437);
nand_5 g08052(new_n8437, new_n1570, new_n8438);
nand_5 g08053(new_n8438, new_n1567, new_n8439_1);
nand_5 g08054(new_n8439_1, new_n1564, new_n8440);
nand_5 g08055(new_n8440, new_n1561, new_n8441);
nand_5 g08056(new_n8441, new_n1338, new_n8442);
nand_5 g08057(new_n8442, new_n1331, new_n8443);
nand_5 g08058(new_n8443, new_n1326, new_n8444);
nand_5 g08059(new_n8444, new_n1321, new_n8445);
nand_5 g08060(new_n8445, new_n1318, new_n8446);
nand_5 g08061(new_n8446, new_n1315, new_n8447);
nand_5 g08062(new_n8447, new_n1312, new_n8448);
nand_5 g08063(new_n8448, new_n1309, new_n8449);
nand_5 g08064(new_n8449, new_n1307, new_n8450);
nand_5 g08065(new_n8450, new_n1304, new_n8451);
nand_5 g08066(new_n8451, new_n1300, new_n8452);
nand_5 g08067(new_n8452, new_n1297, new_n8453);
nand_5 g08068(new_n8453, new_n1294, new_n8454);
nand_5 g08069(new_n8454, new_n1355, new_n8455);
nand_5 g08070(new_n8455, n1093, new_n8456);
nor_5  g08071(new_n8456, new_n774, n8306);
nand_5 g08072(new_n1298, new_n757, new_n8458);
nand_5 g08073(new_n8458, new_n1297, new_n8459);
nand_5 g08074(new_n8459, new_n1294, new_n8460);
nand_5 g08075(new_n8460, new_n1355, new_n8461);
nand_5 g08076(new_n8461, new_n1291, new_n8462);
nand_5 g08077(new_n8462, new_n1288, new_n8463_1);
nand_5 g08078(new_n8463_1, new_n1283, new_n8464);
nand_5 g08079(new_n8464, new_n1363, new_n8465);
nand_5 g08080(new_n8465, new_n1280, new_n8466);
nand_5 g08081(new_n8466, new_n1370, new_n8467);
nand_5 g08082(new_n8467, new_n1373, new_n8468);
nand_5 g08083(new_n8468, new_n1277, new_n8469);
nand_5 g08084(new_n8469, new_n1272, new_n8470);
nand_5 g08085(new_n8470, new_n1269, new_n8471_1);
nand_5 g08086(new_n8471_1, new_n1380, new_n8472);
nand_5 g08087(new_n8472, new_n1264, new_n8473);
nand_5 g08088(new_n8473, new_n1259, new_n8474);
nand_5 g08089(new_n8474, new_n1388, new_n8475);
nand_5 g08090(new_n8475, new_n1392, new_n8476);
nand_5 g08091(new_n8476, new_n1256, new_n8477);
nand_5 g08092(new_n8477, new_n1252, new_n8478);
nand_5 g08093(new_n8478, new_n1249, new_n8479);
nand_5 g08094(new_n8479, new_n1244, new_n8480);
nand_5 g08095(new_n8480, new_n1240, new_n8481);
nand_5 g08096(new_n8481, new_n1234, new_n8482);
nand_5 g08097(new_n8482, new_n1231, new_n8483);
nand_5 g08098(new_n8483, new_n1227, new_n8484);
nand_5 g08099(new_n8484, new_n1407, new_n8485);
nand_5 g08100(new_n8485, new_n1223, new_n8486_1);
nand_5 g08101(new_n8486_1, new_n1218, new_n8487);
nand_5 g08102(new_n8487, new_n1213, new_n8488);
nand_5 g08103(new_n8488, new_n1210, new_n8489);
nand_5 g08104(new_n8489, new_n1206, new_n8490);
nand_5 g08105(new_n8490, new_n1418, new_n8491);
nand_5 g08106(new_n8491, new_n1422, new_n8492);
nand_5 g08107(new_n8492, new_n1428, new_n8493);
nand_5 g08108(new_n8493, new_n1203, new_n8494);
nand_5 g08109(new_n8494, new_n1433, new_n8495);
nand_5 g08110(new_n8495, new_n581, new_n8496);
nand_5 g08111(new_n8496, new_n574, new_n8497);
nand_5 g08112(new_n8497, new_n568, new_n8498);
nand_5 g08113(new_n8498, new_n589, new_n8499);
nand_5 g08114(new_n8499, new_n595, new_n8500);
nand_5 g08115(new_n8500, new_n601, new_n8501);
nand_5 g08116(new_n8501, new_n563, new_n8502);
nand_5 g08117(new_n8502, new_n608, new_n8503);
nand_5 g08118(new_n8503, new_n558, new_n8504);
nand_5 g08119(new_n8504, new_n615, new_n8505);
nand_5 g08120(new_n8505, new_n553, new_n8506);
nand_5 g08121(new_n8506, new_n622, new_n8507);
nand_5 g08122(new_n8507, new_n628, new_n8508);
nand_5 g08123(new_n8508, new_n548, new_n8509);
nand_5 g08124(new_n8509, new_n543_1, new_n8510);
nand_5 g08125(new_n8510, new_n636, new_n8511);
nand_5 g08126(new_n8511, new_n642, new_n8512);
nand_5 g08127(new_n8512, new_n538, new_n8513);
nand_5 g08128(new_n8513, new_n533, new_n8514);
nand_5 g08129(new_n8514, new_n650_1, new_n8515);
nand_5 g08130(new_n8515, new_n528, new_n8516);
nand_5 g08131(new_n8516, new_n523, new_n8517);
nand_5 g08132(new_n8517, new_n518, new_n8518);
nand_5 g08133(new_n8518, new_n659, new_n8519);
nand_5 g08134(new_n8519, new_n665, new_n8520);
nand_5 g08135(new_n8520, new_n672, new_n8521);
nand_5 g08136(new_n8521, new_n513, new_n8522);
nand_5 g08137(new_n8522, new_n679, new_n8523);
nand_5 g08138(new_n8523, new_n685, new_n8524);
nand_5 g08139(new_n8524, new_n691, new_n8525);
nand_5 g08140(new_n8525, new_n508, new_n8526);
nand_5 g08141(new_n8526, new_n698, new_n8527);
nand_5 g08142(new_n8527, new_n503, new_n8528);
nand_5 g08143(new_n8528, new_n704, new_n8529);
nand_5 g08144(new_n8529, new_n498_1, new_n8530);
nand_5 g08145(new_n8530, new_n711, new_n8531);
nand_5 g08146(new_n8531, new_n493, new_n8532);
nand_5 g08147(new_n8532, new_n718, new_n8533);
nand_5 g08148(new_n8533, new_n488, new_n8534);
nand_5 g08149(new_n8534, new_n725, new_n8535);
nand_5 g08150(new_n8535, new_n483, new_n8536);
nand_5 g08151(new_n8536, new_n732, new_n8537);
nand_5 g08152(new_n8537, new_n478, new_n8538);
nand_5 g08153(new_n8538, new_n739, new_n8539);
nand_5 g08154(new_n8539, new_n745, new_n8540);
nand_5 g08155(new_n8540, new_n751, new_n8541);
nand_5 g08156(new_n8541, n9544, new_n8542);
nor_5  g08157(new_n8542, new_n470, n8471);
nand_5 g08158(new_n2031, new_n1276, new_n8544);
nand_5 g08159(new_n8544, new_n2029, new_n8545);
nand_5 g08160(new_n8545, new_n2026, new_n8546);
nand_5 g08161(new_n8546, new_n2022, new_n8547);
nand_5 g08162(new_n8547, new_n2018, new_n8548);
nand_5 g08163(new_n8548, new_n1726, new_n8549);
nand_5 g08164(new_n8549, new_n1722, new_n8550_1);
nand_5 g08165(new_n8550_1, new_n1718, new_n8551);
nand_5 g08166(new_n8551, new_n1713, new_n8552_1);
nand_5 g08167(new_n8552_1, new_n1737, new_n8553);
nand_5 g08168(new_n8553, new_n1709, new_n8554);
nand_5 g08169(new_n8554, new_n1742, new_n8555);
nand_5 g08170(new_n8555, new_n1704, new_n8556);
nand_5 g08171(new_n8556, new_n1702_1, new_n8557);
nand_5 g08172(new_n8557, new_n1698, new_n8558);
nand_5 g08173(new_n8558, new_n1695, new_n8559);
nand_5 g08174(new_n8559, new_n1692, new_n8560);
nand_5 g08175(new_n8560, new_n1752, new_n8561);
nand_5 g08176(new_n8561, new_n1688, new_n8562);
nand_5 g08177(new_n8562, new_n1685, new_n8563);
nand_5 g08178(new_n8563, new_n1680, new_n8564);
nand_5 g08179(new_n8564, new_n1676, new_n8565);
nand_5 g08180(new_n8565, new_n1672, new_n8566);
nand_5 g08181(new_n8566, new_n1669, new_n8567);
nand_5 g08182(new_n8567, new_n1666, new_n8568);
nand_5 g08183(new_n8568, new_n1663, new_n8569);
nand_5 g08184(new_n8569, new_n1658, new_n8570);
nand_5 g08185(new_n8570, new_n1653, new_n8571);
nand_5 g08186(new_n8571, new_n1651, new_n8572);
nand_5 g08187(new_n8572, new_n1649, new_n8573);
nand_5 g08188(new_n8573, new_n1646, new_n8574);
nand_5 g08189(new_n8574, new_n1643, new_n8575);
nand_5 g08190(new_n8575, new_n1641, new_n8576);
nand_5 g08191(new_n8576, new_n1638, new_n8577);
nand_5 g08192(new_n8577, new_n1635, new_n8578);
nand_5 g08193(new_n8578, new_n1632, new_n8579);
nand_5 g08194(new_n8579, new_n1628, new_n8580);
nand_5 g08195(new_n8580, new_n1625, new_n8581);
nand_5 g08196(new_n8581, new_n1621, new_n8582);
nand_5 g08197(new_n8582, new_n1618, new_n8583);
nand_5 g08198(new_n8583, new_n1778, new_n8584);
nand_5 g08199(new_n8584, new_n1782, new_n8585);
nand_5 g08200(new_n8585, new_n1614, new_n8586);
nand_5 g08201(new_n8586, new_n1611, new_n8587);
nand_5 g08202(new_n8587, new_n1789, new_n8588);
nand_5 g08203(new_n8588, new_n1608, new_n8589);
nand_5 g08204(new_n8589, new_n1605, new_n8590);
nand_5 g08205(new_n8590, new_n1795, new_n8591);
nand_5 g08206(new_n8591, new_n1799, new_n8592);
nand_5 g08207(new_n8592, new_n1602, new_n8593);
nand_5 g08208(new_n8593, new_n1599, new_n8594);
nand_5 g08209(new_n8594, new_n1596, new_n8595);
nand_5 g08210(new_n8595, new_n1593, new_n8596);
nand_5 g08211(new_n8596, new_n1806, new_n8597);
nand_5 g08212(new_n8597, new_n1589, new_n8598_1);
nand_5 g08213(new_n8598_1, new_n1586, new_n8599);
nand_5 g08214(new_n8599, new_n1583, new_n8600);
nand_5 g08215(new_n8600, new_n1580, new_n8601);
nand_5 g08216(new_n8601, new_n1576, new_n8602);
nand_5 g08217(new_n8602, new_n1573, new_n8603);
nand_5 g08218(new_n8603, new_n1570, new_n8604_1);
nand_5 g08219(new_n8604_1, new_n1567, new_n8605);
nand_5 g08220(new_n8605, new_n1564, new_n8606);
nand_5 g08221(new_n8606, new_n1561, new_n8607);
nand_5 g08222(new_n8607, new_n1338, new_n8608);
nand_5 g08223(new_n8608, new_n1331, new_n8609);
nand_5 g08224(new_n8609, new_n1326, new_n8610);
nand_5 g08225(new_n8610, new_n1321, new_n8611);
nand_5 g08226(new_n8611, new_n1318, new_n8612);
nand_5 g08227(new_n8612, new_n1315, new_n8613);
nand_5 g08228(new_n8613, new_n1312, new_n8614);
nand_5 g08229(new_n8614, new_n1309, new_n8615);
nand_5 g08230(new_n8615, new_n1307, new_n8616);
nand_5 g08231(new_n8616, new_n1304, new_n8617);
nand_5 g08232(new_n8617, new_n1300, new_n8618);
nand_5 g08233(new_n8618, new_n1297, new_n8619);
nand_5 g08234(new_n8619, new_n1294, new_n8620);
nand_5 g08235(new_n8620, new_n1355, new_n8621);
nand_5 g08236(new_n8621, new_n1291, new_n8622);
nand_5 g08237(new_n8622, new_n1288, new_n8623);
nand_5 g08238(new_n8623, new_n1283, new_n8624);
nand_5 g08239(new_n8624, new_n1363, new_n8625);
nand_5 g08240(new_n8625, new_n1280, new_n8626);
nand_5 g08241(new_n8626, new_n1370, new_n8627);
nand_5 g08242(new_n8627, n5786, new_n8628);
nor_5  g08243(new_n8628, new_n451_1, n8604);
nand_5 g08244(new_n2028, new_n809, new_n8630);
nand_5 g08245(new_n8630, new_n442, new_n8631);
nand_5 g08246(new_n8631, new_n437, new_n8632);
nand_5 g08247(new_n8632, new_n819, new_n8633);
nand_5 g08248(new_n8633, new_n432, new_n8634);
nand_5 g08249(new_n8634, new_n427_1, new_n8635_1);
nand_5 g08250(new_n8635_1, new_n422, new_n8636);
nand_5 g08251(new_n8636, new_n828, new_n8637);
nand_5 g08252(new_n8637, new_n834, new_n8638);
nand_5 g08253(new_n8638, new_n840, new_n8639);
nand_5 g08254(new_n8639, new_n417, new_n8640);
nand_5 g08255(new_n8640, new_n847, new_n8641);
nand_5 g08256(new_n8641, new_n853, new_n8642);
nand_5 g08257(new_n8642, new_n859, new_n8643);
nand_5 g08258(new_n8643, new_n412, new_n8644);
nand_5 g08259(new_n8644, new_n866, new_n8645);
nand_5 g08260(new_n8645, new_n872, new_n8646);
nand_5 g08261(new_n8646, new_n878, new_n8647);
nand_5 g08262(new_n8647, new_n407, new_n8648);
nand_5 g08263(new_n8648, new_n885, new_n8649_1);
nand_5 g08264(new_n8649_1, new_n402, new_n8650);
nand_5 g08265(new_n8650, new_n397, new_n8651);
nand_5 g08266(new_n8651, new_n392, new_n8652);
nand_5 g08267(new_n8652, new_n894, new_n8653);
nand_5 g08268(new_n8653, new_n1087, new_n8654);
nand_5 g08269(new_n8654, new_n1129, new_n8655);
nand_5 g08270(new_n8655, new_n1084, new_n8656);
nand_5 g08271(new_n8656, new_n1134, new_n8657);
nand_5 g08272(new_n8657, new_n1080, new_n8658);
nand_5 g08273(new_n8658, new_n1075, new_n8659);
nand_5 g08274(new_n8659, new_n1070, new_n8660);
nand_5 g08275(new_n8660, new_n1143, new_n8661);
nand_5 g08276(new_n8661, new_n1148, new_n8662);
nand_5 g08277(new_n8662, new_n1065, new_n8663);
nand_5 g08278(new_n8663, new_n1062, new_n8664);
nand_5 g08279(new_n8664, new_n1156, new_n8665);
nand_5 g08280(new_n8665, new_n1057, new_n8666);
nand_5 g08281(new_n8666, new_n1053, new_n8667);
nand_5 g08282(new_n8667, new_n1050, new_n8668);
nand_5 g08283(new_n8668, new_n1045, new_n8669);
nand_5 g08284(new_n8669, new_n1040, new_n8670);
nand_5 g08285(new_n8670, new_n1036, new_n8671);
nand_5 g08286(new_n8671, new_n1033, new_n8672);
nand_5 g08287(new_n8672, new_n1028, new_n8673);
nand_5 g08288(new_n8673, new_n1026, new_n8674);
nand_5 g08289(new_n8674, new_n1021, new_n8675);
nand_5 g08290(new_n8675, new_n1017, new_n8676);
nand_5 g08291(new_n8676, new_n1012, new_n8677);
nand_5 g08292(new_n8677, new_n1009, new_n8678);
nand_5 g08293(new_n8678, new_n1004, new_n8679);
nand_5 g08294(new_n8679, new_n1000, new_n8680);
nand_5 g08295(new_n8680, new_n995, new_n8681);
nand_5 g08296(new_n8681, new_n990, new_n8682);
nand_5 g08297(new_n8682, new_n985, new_n8683);
nand_5 g08298(new_n8683, new_n981, new_n8684);
nand_5 g08299(new_n8684, new_n1179, new_n8685);
nand_5 g08300(new_n8685, new_n976, new_n8686);
nand_5 g08301(new_n8686, new_n971, new_n8687);
nand_5 g08302(new_n8687, new_n966, new_n8688);
nand_5 g08303(new_n8688, new_n961, new_n8689);
nand_5 g08304(new_n8689, new_n957, new_n8690);
nand_5 g08305(new_n8690, new_n952, new_n8691);
nand_5 g08306(new_n8691, new_n948_1, new_n8692);
nand_5 g08307(new_n8692, new_n943, new_n8693);
nand_5 g08308(new_n8693, new_n941, new_n8694);
nand_5 g08309(new_n8694, new_n938, new_n8695);
nand_5 g08310(new_n8695, new_n936, new_n8696);
nand_5 g08311(new_n8696, new_n931, new_n8697);
nand_5 g08312(new_n8697, new_n927, new_n8698);
nand_5 g08313(new_n8698, new_n922, new_n8699);
nand_5 g08314(new_n8699, new_n917, new_n8700);
nand_5 g08315(new_n8700, new_n912, new_n8701);
nand_5 g08316(new_n8701, new_n907, new_n8702);
nand_5 g08317(new_n8702, new_n903, new_n8703);
nand_5 g08318(new_n8703, new_n2066, new_n8704);
nand_5 g08319(new_n8704, new_n2063, new_n8705);
nand_5 g08320(new_n8705, new_n2062, new_n8706);
nand_5 g08321(new_n8706, new_n2058, new_n8707);
nand_5 g08322(new_n8707, new_n2055, new_n8708);
nand_5 g08323(new_n8708, new_n2051, new_n8709);
nand_5 g08324(new_n8709, new_n2046, new_n8710);
nand_5 g08325(new_n8710, new_n2042, new_n8711);
nand_5 g08326(new_n8711, new_n2039, new_n8712);
nand_5 g08327(new_n8712, new_n2036, new_n8713);
nand_5 g08328(new_n8713, n9589, new_n8714);
nor_5  g08329(new_n8714, new_n2030, n8909);
not_4  g08330(new_n521, new_n8716);
nand_5 g08331(new_n1799, new_n8716, new_n8717);
nand_5 g08332(new_n8717, new_n1602, new_n8718);
nand_5 g08333(new_n8718, new_n1599, new_n8719);
nand_5 g08334(new_n8719, new_n1596, new_n8720);
nand_5 g08335(new_n8720, new_n1593, new_n8721);
nand_5 g08336(new_n8721, new_n1806, new_n8722);
nand_5 g08337(new_n8722, new_n1589, new_n8723);
nand_5 g08338(new_n8723, new_n1586, new_n8724);
nand_5 g08339(new_n8724, new_n1583, new_n8725);
nand_5 g08340(new_n8725, new_n1580, new_n8726);
nand_5 g08341(new_n8726, new_n1576, new_n8727);
nand_5 g08342(new_n8727, new_n1573, new_n8728);
nand_5 g08343(new_n8728, new_n1570, new_n8729);
nand_5 g08344(new_n8729, new_n1567, new_n8730);
nand_5 g08345(new_n8730, new_n1564, new_n8731);
nand_5 g08346(new_n8731, new_n1561, new_n8732);
nand_5 g08347(new_n8732, new_n1338, new_n8733);
nand_5 g08348(new_n8733, new_n1331, new_n8734);
nand_5 g08349(new_n8734, new_n1326, new_n8735);
nand_5 g08350(new_n8735, new_n1321, new_n8736);
nand_5 g08351(new_n8736, new_n1318, new_n8737_1);
nand_5 g08352(new_n8737_1, new_n1315, new_n8738);
nand_5 g08353(new_n8738, new_n1312, new_n8739);
nand_5 g08354(new_n8739, new_n1309, new_n8740);
nand_5 g08355(new_n8740, new_n1307, new_n8741);
nand_5 g08356(new_n8741, new_n1304, new_n8742);
nand_5 g08357(new_n8742, new_n1300, new_n8743);
nand_5 g08358(new_n8743, new_n1297, new_n8744);
nand_5 g08359(new_n8744, new_n1294, new_n8745);
nand_5 g08360(new_n8745, new_n1355, new_n8746_1);
nand_5 g08361(new_n8746_1, new_n1291, new_n8747);
nand_5 g08362(new_n8747, new_n1288, new_n8748);
nand_5 g08363(new_n8748, new_n1283, new_n8749);
nand_5 g08364(new_n8749, new_n1363, new_n8750);
nand_5 g08365(new_n8750, new_n1280, new_n8751);
nand_5 g08366(new_n8751, new_n1370, new_n8752);
nand_5 g08367(new_n8752, new_n1373, new_n8753);
nand_5 g08368(new_n8753, new_n1277, new_n8754);
nand_5 g08369(new_n8754, new_n1272, new_n8755);
nand_5 g08370(new_n8755, new_n1269, new_n8756);
nand_5 g08371(new_n8756, new_n1380, new_n8757);
nand_5 g08372(new_n8757, new_n1264, new_n8758);
nand_5 g08373(new_n8758, new_n1259, new_n8759);
nand_5 g08374(new_n8759, new_n1388, new_n8760);
nand_5 g08375(new_n8760, new_n1392, new_n8761);
nand_5 g08376(new_n8761, new_n1256, new_n8762);
nand_5 g08377(new_n8762, new_n1252, new_n8763);
nand_5 g08378(new_n8763, new_n1249, new_n8764);
nand_5 g08379(new_n8764, new_n1244, new_n8765);
nand_5 g08380(new_n8765, new_n1240, new_n8766);
nand_5 g08381(new_n8766, new_n1234, new_n8767);
nand_5 g08382(new_n8767, new_n1231, new_n8768);
nand_5 g08383(new_n8768, new_n1227, new_n8769);
nand_5 g08384(new_n8769, new_n1407, new_n8770);
nand_5 g08385(new_n8770, new_n1223, new_n8771);
nand_5 g08386(new_n8771, new_n1218, new_n8772);
nand_5 g08387(new_n8772, new_n1213, new_n8773);
nand_5 g08388(new_n8773, new_n1210, new_n8774);
nand_5 g08389(new_n8774, new_n1206, new_n8775);
nand_5 g08390(new_n8775, new_n1418, new_n8776);
nand_5 g08391(new_n8776, new_n1422, new_n8777);
nand_5 g08392(new_n8777, new_n1428, new_n8778);
nand_5 g08393(new_n8778, new_n1203, new_n8779);
nand_5 g08394(new_n8779, new_n1433, new_n8780_1);
nand_5 g08395(new_n8780_1, new_n581, new_n8781);
nand_5 g08396(new_n8781, new_n574, new_n8782);
nand_5 g08397(new_n8782, new_n568, new_n8783);
nand_5 g08398(new_n8783, new_n589, new_n8784);
nand_5 g08399(new_n8784, new_n595, new_n8785);
nand_5 g08400(new_n8785, new_n601, new_n8786);
nand_5 g08401(new_n8786, new_n563, new_n8787);
nand_5 g08402(new_n8787, new_n608, new_n8788);
nand_5 g08403(new_n8788, new_n558, new_n8789);
nand_5 g08404(new_n8789, new_n615, new_n8790);
nand_5 g08405(new_n8790, new_n553, new_n8791);
nand_5 g08406(new_n8791, new_n622, new_n8792);
nand_5 g08407(new_n8792, new_n628, new_n8793);
nand_5 g08408(new_n8793, new_n548, new_n8794);
nand_5 g08409(new_n8794, new_n543_1, new_n8795);
nand_5 g08410(new_n8795, new_n636, new_n8796);
nand_5 g08411(new_n8796, new_n642, new_n8797);
nand_5 g08412(new_n8797, new_n538, new_n8798);
nand_5 g08413(new_n8798, new_n533, new_n8799_1);
nand_5 g08414(new_n8799_1, new_n650_1, new_n8800_1);
nand_5 g08415(new_n8800_1, n6680, new_n8801);
nor_5  g08416(new_n8801, new_n525, n9096);
nand_5 g08417(new_n1405, new_n864, new_n8803);
nand_5 g08418(new_n8803, new_n1690, new_n8804);
nand_5 g08419(new_n8804, new_n1752, new_n8805);
nand_5 g08420(new_n8805, new_n1688, new_n8806);
nand_5 g08421(new_n8806, new_n1685, new_n8807);
nand_5 g08422(new_n8807, new_n1680, new_n8808);
nand_5 g08423(new_n8808, new_n1676, new_n8809);
nand_5 g08424(new_n8809, new_n1672, new_n8810);
nand_5 g08425(new_n8810, new_n1669, new_n8811);
nand_5 g08426(new_n8811, new_n1666, new_n8812);
nand_5 g08427(new_n8812, new_n1663, new_n8813);
nand_5 g08428(new_n8813, new_n1658, new_n8814);
nand_5 g08429(new_n8814, new_n1653, new_n8815);
nand_5 g08430(new_n8815, new_n1651, new_n8816);
nand_5 g08431(new_n8816, new_n1649, new_n8817);
nand_5 g08432(new_n8817, new_n1646, new_n8818);
nand_5 g08433(new_n8818, new_n1643, new_n8819);
nand_5 g08434(new_n8819, new_n1641, new_n8820);
nand_5 g08435(new_n8820, new_n1638, new_n8821);
nand_5 g08436(new_n8821, new_n1635, new_n8822);
nand_5 g08437(new_n8822, new_n1632, new_n8823);
nand_5 g08438(new_n8823, new_n1628, new_n8824);
nand_5 g08439(new_n8824, new_n1625, new_n8825);
nand_5 g08440(new_n8825, new_n1621, new_n8826);
nand_5 g08441(new_n8826, new_n1618, new_n8827);
nand_5 g08442(new_n8827, new_n1778, new_n8828);
nand_5 g08443(new_n8828, new_n1782, new_n8829);
nand_5 g08444(new_n8829, new_n1614, new_n8830);
nand_5 g08445(new_n8830, new_n1611, new_n8831);
nand_5 g08446(new_n8831, new_n1789, new_n8832);
nand_5 g08447(new_n8832, new_n1608, new_n8833);
nand_5 g08448(new_n8833, new_n1605, new_n8834);
nand_5 g08449(new_n8834, new_n1795, new_n8835);
nand_5 g08450(new_n8835, new_n1799, new_n8836);
nand_5 g08451(new_n8836, new_n1602, new_n8837);
nand_5 g08452(new_n8837, new_n1599, new_n8838);
nand_5 g08453(new_n8838, new_n1596, new_n8839);
nand_5 g08454(new_n8839, new_n1593, new_n8840);
nand_5 g08455(new_n8840, new_n1806, new_n8841);
nand_5 g08456(new_n8841, new_n1589, new_n8842);
nand_5 g08457(new_n8842, new_n1586, new_n8843);
nand_5 g08458(new_n8843, new_n1583, new_n8844);
nand_5 g08459(new_n8844, new_n1580, new_n8845);
nand_5 g08460(new_n8845, new_n1576, new_n8846);
nand_5 g08461(new_n8846, new_n1573, new_n8847);
nand_5 g08462(new_n8847, new_n1570, new_n8848);
nand_5 g08463(new_n8848, new_n1567, new_n8849);
nand_5 g08464(new_n8849, new_n1564, new_n8850);
nand_5 g08465(new_n8850, new_n1561, new_n8851);
nand_5 g08466(new_n8851, new_n1338, new_n8852);
nand_5 g08467(new_n8852, new_n1331, new_n8853);
nand_5 g08468(new_n8853, new_n1326, new_n8854);
nand_5 g08469(new_n8854, new_n1321, new_n8855);
nand_5 g08470(new_n8855, new_n1318, new_n8856);
nand_5 g08471(new_n8856, new_n1315, new_n8857);
nand_5 g08472(new_n8857, new_n1312, new_n8858);
nand_5 g08473(new_n8858, new_n1309, new_n8859);
nand_5 g08474(new_n8859, new_n1307, new_n8860);
nand_5 g08475(new_n8860, new_n1304, new_n8861);
nand_5 g08476(new_n8861, new_n1300, new_n8862);
nand_5 g08477(new_n8862, new_n1297, new_n8863);
nand_5 g08478(new_n8863, new_n1294, new_n8864);
nand_5 g08479(new_n8864, new_n1355, new_n8865);
nand_5 g08480(new_n8865, new_n1291, new_n8866);
nand_5 g08481(new_n8866, new_n1288, new_n8867);
nand_5 g08482(new_n8867, new_n1283, new_n8868);
nand_5 g08483(new_n8868, new_n1363, new_n8869);
nand_5 g08484(new_n8869, new_n1280, new_n8870);
nand_5 g08485(new_n8870, new_n1370, new_n8871);
nand_5 g08486(new_n8871, new_n1373, new_n8872);
nand_5 g08487(new_n8872, new_n1277, new_n8873_1);
nand_5 g08488(new_n8873_1, new_n1272, new_n8874);
nand_5 g08489(new_n8874, new_n1269, new_n8875);
nand_5 g08490(new_n8875, new_n1380, new_n8876);
nand_5 g08491(new_n8876, new_n1264, new_n8877);
nand_5 g08492(new_n8877, new_n1259, new_n8878);
nand_5 g08493(new_n8878, new_n1388, new_n8879);
nand_5 g08494(new_n8879, new_n1392, new_n8880);
nand_5 g08495(new_n8880, new_n1256, new_n8881);
nand_5 g08496(new_n8881, new_n1252, new_n8882);
nand_5 g08497(new_n8882, new_n1249, new_n8883);
nand_5 g08498(new_n8883, new_n1244, new_n8884);
nand_5 g08499(new_n8884, new_n1240, new_n8885);
nand_5 g08500(new_n8885, new_n1234, new_n8886);
nand_5 g08501(new_n8886, new_n1231, new_n8887);
nand_5 g08502(new_n8887, n8439, new_n8888);
nor_5  g08503(new_n8888, new_n1224, n9342);
nand_5 g08504(new_n670, new_n993, new_n8890);
nand_5 g08505(new_n8890, new_n1591, new_n8891);
nand_5 g08506(new_n8891, new_n1806, new_n8892_1);
nand_5 g08507(new_n8892_1, new_n1589, new_n8893);
nand_5 g08508(new_n8893, new_n1586, new_n8894);
nand_5 g08509(new_n8894, new_n1583, new_n8895);
nand_5 g08510(new_n8895, new_n1580, new_n8896);
nand_5 g08511(new_n8896, new_n1576, new_n8897);
nand_5 g08512(new_n8897, new_n1573, new_n8898);
nand_5 g08513(new_n8898, new_n1570, new_n8899);
nand_5 g08514(new_n8899, new_n1567, new_n8900);
nand_5 g08515(new_n8900, new_n1564, new_n8901);
nand_5 g08516(new_n8901, new_n1561, new_n8902);
nand_5 g08517(new_n8902, new_n1338, new_n8903);
nand_5 g08518(new_n8903, new_n1331, new_n8904);
nand_5 g08519(new_n8904, new_n1326, new_n8905);
nand_5 g08520(new_n8905, new_n1321, new_n8906);
nand_5 g08521(new_n8906, new_n1318, new_n8907);
nand_5 g08522(new_n8907, new_n1315, new_n8908);
nand_5 g08523(new_n8908, new_n1312, new_n8909_1);
nand_5 g08524(new_n8909_1, new_n1309, new_n8910);
nand_5 g08525(new_n8910, new_n1307, new_n8911);
nand_5 g08526(new_n8911, new_n1304, new_n8912);
nand_5 g08527(new_n8912, new_n1300, new_n8913);
nand_5 g08528(new_n8913, new_n1297, new_n8914);
nand_5 g08529(new_n8914, new_n1294, new_n8915);
nand_5 g08530(new_n8915, new_n1355, new_n8916);
nand_5 g08531(new_n8916, new_n1291, new_n8917);
nand_5 g08532(new_n8917, new_n1288, new_n8918);
nand_5 g08533(new_n8918, new_n1283, new_n8919);
nand_5 g08534(new_n8919, new_n1363, new_n8920);
nand_5 g08535(new_n8920, new_n1280, new_n8921);
nand_5 g08536(new_n8921, new_n1370, new_n8922);
nand_5 g08537(new_n8922, new_n1373, new_n8923);
nand_5 g08538(new_n8923, new_n1277, new_n8924);
nand_5 g08539(new_n8924, new_n1272, new_n8925);
nand_5 g08540(new_n8925, new_n1269, new_n8926_1);
nand_5 g08541(new_n8926_1, new_n1380, new_n8927);
nand_5 g08542(new_n8927, new_n1264, new_n8928);
nand_5 g08543(new_n8928, new_n1259, new_n8929);
nand_5 g08544(new_n8929, new_n1388, new_n8930);
nand_5 g08545(new_n8930, new_n1392, new_n8931);
nand_5 g08546(new_n8931, new_n1256, new_n8932);
nand_5 g08547(new_n8932, new_n1252, new_n8933);
nand_5 g08548(new_n8933, new_n1249, new_n8934);
nand_5 g08549(new_n8934, new_n1244, new_n8935);
nand_5 g08550(new_n8935, new_n1240, new_n8936);
nand_5 g08551(new_n8936, new_n1234, new_n8937);
nand_5 g08552(new_n8937, new_n1231, new_n8938);
nand_5 g08553(new_n8938, new_n1227, new_n8939);
nand_5 g08554(new_n8939, new_n1407, new_n8940);
nand_5 g08555(new_n8940, new_n1223, new_n8941);
nand_5 g08556(new_n8941, new_n1218, new_n8942);
nand_5 g08557(new_n8942, new_n1213, new_n8943);
nand_5 g08558(new_n8943, new_n1210, new_n8944);
nand_5 g08559(new_n8944, new_n1206, new_n8945);
nand_5 g08560(new_n8945, new_n1418, new_n8946);
nand_5 g08561(new_n8946, new_n1422, new_n8947);
nand_5 g08562(new_n8947, new_n1428, new_n8948);
nand_5 g08563(new_n8948, new_n1203, new_n8949);
nand_5 g08564(new_n8949, new_n1433, new_n8950);
nand_5 g08565(new_n8950, new_n581, new_n8951);
nand_5 g08566(new_n8951, new_n574, new_n8952);
nand_5 g08567(new_n8952, new_n568, new_n8953);
nand_5 g08568(new_n8953, new_n589, new_n8954);
nand_5 g08569(new_n8954, new_n595, new_n8955);
nand_5 g08570(new_n8955, new_n601, new_n8956);
nand_5 g08571(new_n8956, new_n563, new_n8957);
nand_5 g08572(new_n8957, new_n608, new_n8958);
nand_5 g08573(new_n8958, new_n558, new_n8959);
nand_5 g08574(new_n8959, new_n615, new_n8960);
nand_5 g08575(new_n8960, new_n553, new_n8961);
nand_5 g08576(new_n8961, new_n622, new_n8962);
nand_5 g08577(new_n8962, new_n628, new_n8963);
nand_5 g08578(new_n8963, new_n548, new_n8964);
nand_5 g08579(new_n8964, new_n543_1, new_n8965);
nand_5 g08580(new_n8965, new_n636, new_n8966);
nand_5 g08581(new_n8966, new_n642, new_n8967);
nand_5 g08582(new_n8967, new_n538, new_n8968);
nand_5 g08583(new_n8968, new_n533, new_n8969);
nand_5 g08584(new_n8969, new_n650_1, new_n8970);
nand_5 g08585(new_n8970, new_n528, new_n8971);
nand_5 g08586(new_n8971, new_n523, new_n8972);
nand_5 g08587(new_n8972, new_n518, new_n8973);
nand_5 g08588(new_n8973, new_n659, new_n8974);
nand_5 g08589(new_n8974, n12614, new_n8975);
nor_5  g08590(new_n8975, new_n662, n9437);
nand_5 g08591(new_n1696, new_n1230, new_n8977);
nand_5 g08592(new_n8977, new_n1695, new_n8978);
nand_5 g08593(new_n8978, new_n1692, new_n8979);
nand_5 g08594(new_n8979, new_n1752, new_n8980);
nand_5 g08595(new_n8980, new_n1688, new_n8981);
nand_5 g08596(new_n8981, new_n1685, new_n8982);
nand_5 g08597(new_n8982, new_n1680, new_n8983);
nand_5 g08598(new_n8983, new_n1676, new_n8984);
nand_5 g08599(new_n8984, new_n1672, new_n8985);
nand_5 g08600(new_n8985, new_n1669, new_n8986);
nand_5 g08601(new_n8986, new_n1666, new_n8987);
nand_5 g08602(new_n8987, new_n1663, new_n8988);
nand_5 g08603(new_n8988, new_n1658, new_n8989);
nand_5 g08604(new_n8989, new_n1653, new_n8990);
nand_5 g08605(new_n8990, new_n1651, new_n8991);
nand_5 g08606(new_n8991, new_n1649, new_n8992);
nand_5 g08607(new_n8992, new_n1646, new_n8993);
nand_5 g08608(new_n8993, new_n1643, new_n8994);
nand_5 g08609(new_n8994, new_n1641, new_n8995);
nand_5 g08610(new_n8995, new_n1638, new_n8996);
nand_5 g08611(new_n8996, new_n1635, new_n8997_1);
nand_5 g08612(new_n8997_1, new_n1632, new_n8998);
nand_5 g08613(new_n8998, new_n1628, new_n8999);
nand_5 g08614(new_n8999, new_n1625, new_n9000);
nand_5 g08615(new_n9000, new_n1621, new_n9001);
nand_5 g08616(new_n9001, new_n1618, new_n9002);
nand_5 g08617(new_n9002, new_n1778, new_n9003);
nand_5 g08618(new_n9003, new_n1782, new_n9004);
nand_5 g08619(new_n9004, new_n1614, new_n9005);
nand_5 g08620(new_n9005, new_n1611, new_n9006);
nand_5 g08621(new_n9006, new_n1789, new_n9007);
nand_5 g08622(new_n9007, new_n1608, new_n9008);
nand_5 g08623(new_n9008, new_n1605, new_n9009);
nand_5 g08624(new_n9009, new_n1795, new_n9010);
nand_5 g08625(new_n9010, new_n1799, new_n9011);
nand_5 g08626(new_n9011, new_n1602, new_n9012);
nand_5 g08627(new_n9012, new_n1599, new_n9013);
nand_5 g08628(new_n9013, new_n1596, new_n9014);
nand_5 g08629(new_n9014, new_n1593, new_n9015);
nand_5 g08630(new_n9015, new_n1806, new_n9016);
nand_5 g08631(new_n9016, new_n1589, new_n9017);
nand_5 g08632(new_n9017, new_n1586, new_n9018);
nand_5 g08633(new_n9018, new_n1583, new_n9019);
nand_5 g08634(new_n9019, new_n1580, new_n9020);
nand_5 g08635(new_n9020, new_n1576, new_n9021);
nand_5 g08636(new_n9021, new_n1573, new_n9022);
nand_5 g08637(new_n9022, new_n1570, new_n9023);
nand_5 g08638(new_n9023, new_n1567, new_n9024);
nand_5 g08639(new_n9024, new_n1564, new_n9025);
nand_5 g08640(new_n9025, new_n1561, new_n9026_1);
nand_5 g08641(new_n9026_1, new_n1338, new_n9027);
nand_5 g08642(new_n9027, new_n1331, new_n9028);
nand_5 g08643(new_n9028, new_n1326, new_n9029);
nand_5 g08644(new_n9029, new_n1321, new_n9030);
nand_5 g08645(new_n9030, new_n1318, new_n9031);
nand_5 g08646(new_n9031, new_n1315, new_n9032);
nand_5 g08647(new_n9032, new_n1312, new_n9033);
nand_5 g08648(new_n9033, new_n1309, new_n9034);
nand_5 g08649(new_n9034, new_n1307, new_n9035);
nand_5 g08650(new_n9035, new_n1304, new_n9036);
nand_5 g08651(new_n9036, new_n1300, new_n9037);
nand_5 g08652(new_n9037, new_n1297, new_n9038);
nand_5 g08653(new_n9038, new_n1294, new_n9039);
nand_5 g08654(new_n9039, new_n1355, new_n9040);
nand_5 g08655(new_n9040, new_n1291, new_n9041);
nand_5 g08656(new_n9041, new_n1288, new_n9042);
nand_5 g08657(new_n9042, new_n1283, new_n9043);
nand_5 g08658(new_n9043, new_n1363, new_n9044);
nand_5 g08659(new_n9044, new_n1280, new_n9045);
nand_5 g08660(new_n9045, new_n1370, new_n9046);
nand_5 g08661(new_n9046, new_n1373, new_n9047);
nand_5 g08662(new_n9047, new_n1277, new_n9048);
nand_5 g08663(new_n9048, new_n1272, new_n9049);
nand_5 g08664(new_n9049, new_n1269, new_n9050);
nand_5 g08665(new_n9050, new_n1380, new_n9051);
nand_5 g08666(new_n9051, new_n1264, new_n9052);
nand_5 g08667(new_n9052, new_n1259, new_n9053);
nand_5 g08668(new_n9053, new_n1388, new_n9054);
nand_5 g08669(new_n9054, new_n1392, new_n9055);
nand_5 g08670(new_n9055, new_n1256, new_n9056);
nand_5 g08671(new_n9056, new_n1252, new_n9057);
nand_5 g08672(new_n9057, new_n1249, new_n9058);
nand_5 g08673(new_n9058, new_n1244, new_n9059);
nand_5 g08674(new_n9059, new_n1240, new_n9060);
nand_5 g08675(new_n9060, n12782, new_n9061);
nor_5  g08676(new_n9061, new_n844_1, n9447);
not_4  g08677(new_n1063, new_n9063);
nand_5 g08678(new_n9063, new_n558, new_n9064);
nand_5 g08679(new_n9064, new_n615, new_n9065);
nand_5 g08680(new_n9065, new_n553, new_n9066);
nand_5 g08681(new_n9066, new_n622, new_n9067);
nand_5 g08682(new_n9067, new_n628, new_n9068);
nand_5 g08683(new_n9068, new_n548, new_n9069);
nand_5 g08684(new_n9069, new_n543_1, new_n9070);
nand_5 g08685(new_n9070, new_n636, new_n9071);
nand_5 g08686(new_n9071, new_n642, new_n9072);
nand_5 g08687(new_n9072, new_n538, new_n9073);
nand_5 g08688(new_n9073, new_n533, new_n9074);
nand_5 g08689(new_n9074, new_n650_1, new_n9075);
nand_5 g08690(new_n9075, new_n528, new_n9076);
nand_5 g08691(new_n9076, new_n523, new_n9077);
nand_5 g08692(new_n9077, new_n518, new_n9078);
nand_5 g08693(new_n9078, new_n659, new_n9079);
nand_5 g08694(new_n9079, new_n665, new_n9080);
nand_5 g08695(new_n9080, new_n672, new_n9081);
nand_5 g08696(new_n9081, new_n513, new_n9082);
nand_5 g08697(new_n9082, new_n679, new_n9083);
nand_5 g08698(new_n9083, new_n685, new_n9084);
nand_5 g08699(new_n9084, new_n691, new_n9085);
nand_5 g08700(new_n9085, new_n508, new_n9086);
nand_5 g08701(new_n9086, new_n698, new_n9087);
nand_5 g08702(new_n9087, new_n503, new_n9088);
nand_5 g08703(new_n9088, new_n704, new_n9089);
nand_5 g08704(new_n9089, new_n498_1, new_n9090);
nand_5 g08705(new_n9090, new_n711, new_n9091);
nand_5 g08706(new_n9091, new_n493, new_n9092);
nand_5 g08707(new_n9092, new_n718, new_n9093);
nand_5 g08708(new_n9093, new_n488, new_n9094);
nand_5 g08709(new_n9094, new_n725, new_n9095);
nand_5 g08710(new_n9095, new_n483, new_n9096_1);
nand_5 g08711(new_n9096_1, new_n732, new_n9097);
nand_5 g08712(new_n9097, new_n478, new_n9098);
nand_5 g08713(new_n9098, new_n739, new_n9099);
nand_5 g08714(new_n9099, new_n745, new_n9100);
nand_5 g08715(new_n9100, new_n751, new_n9101);
nand_5 g08716(new_n9101, new_n473, new_n9102);
nand_5 g08717(new_n9102, new_n758, new_n9103);
nand_5 g08718(new_n9103, new_n764, new_n9104);
nand_5 g08719(new_n9104, new_n770, new_n9105);
nand_5 g08720(new_n9105, new_n468, new_n9106);
nand_5 g08721(new_n9106, new_n777, new_n9107);
nand_5 g08722(new_n9107, new_n783, new_n9108);
nand_5 g08723(new_n9108, new_n789, new_n9109);
nand_5 g08724(new_n9109, new_n463, new_n9110_1);
nand_5 g08725(new_n9110_1, new_n796, new_n9111);
nand_5 g08726(new_n9111, new_n458, new_n9112);
nand_5 g08727(new_n9112, new_n453, new_n9113);
nand_5 g08728(new_n9113, new_n447, new_n9114);
nand_5 g08729(new_n9114, new_n805, new_n9115);
nand_5 g08730(new_n9115, new_n811, new_n9116);
nand_5 g08731(new_n9116, new_n442, new_n9117);
nand_5 g08732(new_n9117, new_n437, new_n9118);
nand_5 g08733(new_n9118, new_n819, new_n9119);
nand_5 g08734(new_n9119, new_n432, new_n9120);
nand_5 g08735(new_n9120, new_n427_1, new_n9121);
nand_5 g08736(new_n9121, new_n422, new_n9122);
nand_5 g08737(new_n9122, new_n828, new_n9123);
nand_5 g08738(new_n9123, new_n834, new_n9124);
nand_5 g08739(new_n9124, new_n840, new_n9125);
nand_5 g08740(new_n9125, new_n417, new_n9126);
nand_5 g08741(new_n9126, new_n847, new_n9127);
nand_5 g08742(new_n9127, new_n853, new_n9128);
nand_5 g08743(new_n9128, new_n859, new_n9129);
nand_5 g08744(new_n9129, new_n412, new_n9130);
nand_5 g08745(new_n9130, new_n866, new_n9131);
nand_5 g08746(new_n9131, new_n872, new_n9132);
nand_5 g08747(new_n9132, new_n878, new_n9133);
nand_5 g08748(new_n9133, new_n407, new_n9134);
nand_5 g08749(new_n9134, new_n885, new_n9135);
nand_5 g08750(new_n9135, new_n402, new_n9136);
nand_5 g08751(new_n9136, new_n397, new_n9137);
nand_5 g08752(new_n9137, new_n392, new_n9138);
nand_5 g08753(new_n9138, new_n894, new_n9139);
nand_5 g08754(new_n9139, new_n1087, new_n9140);
nand_5 g08755(new_n9140, new_n1129, new_n9141);
nand_5 g08756(new_n9141, new_n1084, new_n9142);
nand_5 g08757(new_n9142, new_n1134, new_n9143);
nand_5 g08758(new_n9143, new_n1080, new_n9144);
nand_5 g08759(new_n9144, new_n1075, new_n9145);
nand_5 g08760(new_n9145, new_n1070, new_n9146);
nand_5 g08761(new_n9146, new_n1143, new_n9147);
nand_5 g08762(new_n9147, n4172, new_n9148);
nor_5  g08763(new_n9148, new_n1636, n9570);
nand_5 g08764(new_n1246, new_n1244, new_n9150);
nand_5 g08765(new_n9150, new_n1240, new_n9151);
nand_5 g08766(new_n9151, new_n1234, new_n9152);
nand_5 g08767(new_n9152, new_n1231, new_n9153);
nand_5 g08768(new_n9153, new_n1227, new_n9154_1);
nand_5 g08769(new_n9154_1, new_n1407, new_n9155);
nand_5 g08770(new_n9155, new_n1223, new_n9156);
nand_5 g08771(new_n9156, new_n1218, new_n9157);
nand_5 g08772(new_n9157, new_n1213, new_n9158);
nand_5 g08773(new_n9158, new_n1210, new_n9159);
nand_5 g08774(new_n9159, new_n1206, new_n9160);
nand_5 g08775(new_n9160, new_n1418, new_n9161);
nand_5 g08776(new_n9161, new_n1422, new_n9162);
nand_5 g08777(new_n9162, new_n1428, new_n9163);
nand_5 g08778(new_n9163, new_n1203, new_n9164);
nand_5 g08779(new_n9164, new_n1433, new_n9165);
nand_5 g08780(new_n9165, new_n581, new_n9166);
nand_5 g08781(new_n9166, new_n574, new_n9167);
nand_5 g08782(new_n9167, new_n568, new_n9168);
nand_5 g08783(new_n9168, new_n589, new_n9169);
nand_5 g08784(new_n9169, new_n595, new_n9170);
nand_5 g08785(new_n9170, new_n601, new_n9171);
nand_5 g08786(new_n9171, new_n563, new_n9172);
nand_5 g08787(new_n9172, new_n608, new_n9173);
nand_5 g08788(new_n9173, new_n558, new_n9174);
nand_5 g08789(new_n9174, new_n615, new_n9175);
nand_5 g08790(new_n9175, new_n553, new_n9176);
nand_5 g08791(new_n9176, new_n622, new_n9177);
nand_5 g08792(new_n9177, new_n628, new_n9178);
nand_5 g08793(new_n9178, new_n548, new_n9179);
nand_5 g08794(new_n9179, new_n543_1, new_n9180);
nand_5 g08795(new_n9180, new_n636, new_n9181);
nand_5 g08796(new_n9181, new_n642, new_n9182);
nand_5 g08797(new_n9182, new_n538, new_n9183);
nand_5 g08798(new_n9183, new_n533, new_n9184);
nand_5 g08799(new_n9184, new_n650_1, new_n9185);
nand_5 g08800(new_n9185, new_n528, new_n9186_1);
nand_5 g08801(new_n9186_1, new_n523, new_n9187);
nand_5 g08802(new_n9187, new_n518, new_n9188);
nand_5 g08803(new_n9188, new_n659, new_n9189);
nand_5 g08804(new_n9189, new_n665, new_n9190);
nand_5 g08805(new_n9190, new_n672, new_n9191);
nand_5 g08806(new_n9191, new_n513, new_n9192);
nand_5 g08807(new_n9192, new_n679, new_n9193);
nand_5 g08808(new_n9193, new_n685, new_n9194);
nand_5 g08809(new_n9194, new_n691, new_n9195);
nand_5 g08810(new_n9195, new_n508, new_n9196);
nand_5 g08811(new_n9196, new_n698, new_n9197);
nand_5 g08812(new_n9197, new_n503, new_n9198);
nand_5 g08813(new_n9198, new_n704, new_n9199);
nand_5 g08814(new_n9199, new_n498_1, new_n9200);
nand_5 g08815(new_n9200, new_n711, new_n9201);
nand_5 g08816(new_n9201, new_n493, new_n9202);
nand_5 g08817(new_n9202, new_n718, new_n9203);
nand_5 g08818(new_n9203, new_n488, new_n9204);
nand_5 g08819(new_n9204, new_n725, new_n9205);
nand_5 g08820(new_n9205, new_n483, new_n9206);
nand_5 g08821(new_n9206, new_n732, new_n9207);
nand_5 g08822(new_n9207, new_n478, new_n9208);
nand_5 g08823(new_n9208, new_n739, new_n9209);
nand_5 g08824(new_n9209, new_n745, new_n9210);
nand_5 g08825(new_n9210, new_n751, new_n9211);
nand_5 g08826(new_n9211, new_n473, new_n9212);
nand_5 g08827(new_n9212, new_n758, new_n9213);
nand_5 g08828(new_n9213, new_n764, new_n9214);
nand_5 g08829(new_n9214, new_n770, new_n9215);
nand_5 g08830(new_n9215, new_n468, new_n9216);
nand_5 g08831(new_n9216, new_n777, new_n9217);
nand_5 g08832(new_n9217, new_n783, new_n9218);
nand_5 g08833(new_n9218, new_n789, new_n9219);
nand_5 g08834(new_n9219, new_n463, new_n9220);
nand_5 g08835(new_n9220, new_n796, new_n9221);
nand_5 g08836(new_n9221, new_n458, new_n9222);
nand_5 g08837(new_n9222, new_n453, new_n9223);
nand_5 g08838(new_n9223, new_n447, new_n9224);
nand_5 g08839(new_n9224, new_n805, new_n9225);
nand_5 g08840(new_n9225, new_n811, new_n9226);
nand_5 g08841(new_n9226, new_n442, new_n9227);
nand_5 g08842(new_n9227, new_n437, new_n9228);
nand_5 g08843(new_n9228, new_n819, new_n9229);
nand_5 g08844(new_n9229, new_n432, new_n9230);
nand_5 g08845(new_n9230, new_n427_1, new_n9231);
nand_5 g08846(new_n9231, new_n422, new_n9232);
nand_5 g08847(new_n9232, new_n828, new_n9233);
nand_5 g08848(new_n9233, n13511, new_n9234);
nor_5  g08849(new_n9234, new_n831, n9665);
nand_5 g08850(new_n1035, new_n640, new_n9236);
nand_5 g08851(new_n9236, new_n538, new_n9237);
nand_5 g08852(new_n9237, new_n533, new_n9238);
nand_5 g08853(new_n9238, new_n650_1, new_n9239);
nand_5 g08854(new_n9239, new_n528, new_n9240);
nand_5 g08855(new_n9240, new_n523, new_n9241);
nand_5 g08856(new_n9241, new_n518, new_n9242);
nand_5 g08857(new_n9242, new_n659, new_n9243);
nand_5 g08858(new_n9243, new_n665, new_n9244);
nand_5 g08859(new_n9244, new_n672, new_n9245);
nand_5 g08860(new_n9245, new_n513, new_n9246);
nand_5 g08861(new_n9246, new_n679, new_n9247);
nand_5 g08862(new_n9247, new_n685, new_n9248);
nand_5 g08863(new_n9248, new_n691, new_n9249);
nand_5 g08864(new_n9249, new_n508, new_n9250);
nand_5 g08865(new_n9250, new_n698, new_n9251);
nand_5 g08866(new_n9251, new_n503, new_n9252_1);
nand_5 g08867(new_n9252_1, new_n704, new_n9253);
nand_5 g08868(new_n9253, new_n498_1, new_n9254);
nand_5 g08869(new_n9254, new_n711, new_n9255);
nand_5 g08870(new_n9255, new_n493, new_n9256);
nand_5 g08871(new_n9256, new_n718, new_n9257);
nand_5 g08872(new_n9257, new_n488, new_n9258);
nand_5 g08873(new_n9258, new_n725, new_n9259);
nand_5 g08874(new_n9259, new_n483, new_n9260);
nand_5 g08875(new_n9260, new_n732, new_n9261);
nand_5 g08876(new_n9261, new_n478, new_n9262);
nand_5 g08877(new_n9262, new_n739, new_n9263);
nand_5 g08878(new_n9263, new_n745, new_n9264);
nand_5 g08879(new_n9264, new_n751, new_n9265);
nand_5 g08880(new_n9265, new_n473, new_n9266);
nand_5 g08881(new_n9266, new_n758, new_n9267);
nand_5 g08882(new_n9267, new_n764, new_n9268);
nand_5 g08883(new_n9268, new_n770, new_n9269);
nand_5 g08884(new_n9269, new_n468, new_n9270);
nand_5 g08885(new_n9270, new_n777, new_n9271);
nand_5 g08886(new_n9271, new_n783, new_n9272);
nand_5 g08887(new_n9272, new_n789, new_n9273);
nand_5 g08888(new_n9273, new_n463, new_n9274);
nand_5 g08889(new_n9274, new_n796, new_n9275);
nand_5 g08890(new_n9275, new_n458, new_n9276);
nand_5 g08891(new_n9276, new_n453, new_n9277);
nand_5 g08892(new_n9277, new_n447, new_n9278);
nand_5 g08893(new_n9278, new_n805, new_n9279);
nand_5 g08894(new_n9279, new_n811, new_n9280);
nand_5 g08895(new_n9280, new_n442, new_n9281);
nand_5 g08896(new_n9281, new_n437, new_n9282);
nand_5 g08897(new_n9282, new_n819, new_n9283);
nand_5 g08898(new_n9283, new_n432, new_n9284);
nand_5 g08899(new_n9284, new_n427_1, new_n9285);
nand_5 g08900(new_n9285, new_n422, new_n9286);
nand_5 g08901(new_n9286, new_n828, new_n9287);
nand_5 g08902(new_n9287, new_n834, new_n9288);
nand_5 g08903(new_n9288, new_n840, new_n9289);
nand_5 g08904(new_n9289, new_n417, new_n9290);
nand_5 g08905(new_n9290, new_n847, new_n9291);
nand_5 g08906(new_n9291, new_n853, new_n9292);
nand_5 g08907(new_n9292, new_n859, new_n9293);
nand_5 g08908(new_n9293, new_n412, new_n9294);
nand_5 g08909(new_n9294, new_n866, new_n9295);
nand_5 g08910(new_n9295, new_n872, new_n9296);
nand_5 g08911(new_n9296, new_n878, new_n9297);
nand_5 g08912(new_n9297, new_n407, new_n9298);
nand_5 g08913(new_n9298, new_n885, new_n9299);
nand_5 g08914(new_n9299, new_n402, new_n9300);
nand_5 g08915(new_n9300, new_n397, new_n9301);
nand_5 g08916(new_n9301, new_n392, new_n9302);
nand_5 g08917(new_n9302, new_n894, new_n9303);
nand_5 g08918(new_n9303, new_n1087, new_n9304);
nand_5 g08919(new_n9304, new_n1129, new_n9305);
nand_5 g08920(new_n9305, new_n1084, new_n9306);
nand_5 g08921(new_n9306, new_n1134, new_n9307);
nand_5 g08922(new_n9307, new_n1080, new_n9308);
nand_5 g08923(new_n9308, new_n1075, new_n9309);
nand_5 g08924(new_n9309, new_n1070, new_n9310);
nand_5 g08925(new_n9310, new_n1143, new_n9311);
nand_5 g08926(new_n9311, new_n1148, new_n9312);
nand_5 g08927(new_n9312, new_n1065, new_n9313);
nand_5 g08928(new_n9313, new_n1062, new_n9314_1);
nand_5 g08929(new_n9314_1, new_n1156, new_n9315);
nand_5 g08930(new_n9315, new_n1057, new_n9316);
nand_5 g08931(new_n9316, new_n1053, new_n9317);
nand_5 g08932(new_n9317, new_n1050, new_n9318);
nand_5 g08933(new_n9318, new_n1045, new_n9319);
nand_5 g08934(new_n9319, n6873, new_n9320);
nor_5  g08935(new_n9320, new_n1780, n9717);
nand_5 g08936(new_n1805, new_n988, new_n9322);
nand_5 g08937(new_n9322, new_n985, new_n9323);
nand_5 g08938(new_n9323, new_n981, new_n9324);
nand_5 g08939(new_n9324, new_n1179, new_n9325);
nand_5 g08940(new_n9325, new_n976, new_n9326);
nand_5 g08941(new_n9326, new_n971, new_n9327);
nand_5 g08942(new_n9327, new_n966, new_n9328);
nand_5 g08943(new_n9328, new_n961, new_n9329);
nand_5 g08944(new_n9329, new_n957, new_n9330);
nand_5 g08945(new_n9330, new_n952, new_n9331);
nand_5 g08946(new_n9331, new_n948_1, new_n9332);
nand_5 g08947(new_n9332, new_n943, new_n9333);
nand_5 g08948(new_n9333, new_n941, new_n9334);
nand_5 g08949(new_n9334, new_n938, new_n9335);
nand_5 g08950(new_n9335, new_n936, new_n9336);
nand_5 g08951(new_n9336, new_n931, new_n9337);
nand_5 g08952(new_n9337, new_n927, new_n9338);
nand_5 g08953(new_n9338, new_n922, new_n9339);
nand_5 g08954(new_n9339, new_n917, new_n9340);
nand_5 g08955(new_n9340, new_n912, new_n9341);
nand_5 g08956(new_n9341, new_n907, new_n9342_1);
nand_5 g08957(new_n9342_1, new_n903, new_n9343);
nand_5 g08958(new_n9343, new_n2066, new_n9344);
nand_5 g08959(new_n9344, new_n2063, new_n9345);
nand_5 g08960(new_n9345, new_n2062, new_n9346);
nand_5 g08961(new_n9346, new_n2058, new_n9347);
nand_5 g08962(new_n9347, new_n2055, new_n9348);
nand_5 g08963(new_n9348, new_n2051, new_n9349);
nand_5 g08964(new_n9349, new_n2046, new_n9350);
nand_5 g08965(new_n9350, new_n2042, new_n9351);
nand_5 g08966(new_n9351, new_n2039, new_n9352);
nand_5 g08967(new_n9352, new_n2036, new_n9353);
nand_5 g08968(new_n9353, new_n2033, new_n9354);
nand_5 g08969(new_n9354, new_n2029, new_n9355);
nand_5 g08970(new_n9355, new_n2026, new_n9356);
nand_5 g08971(new_n9356, new_n2022, new_n9357);
nand_5 g08972(new_n9357, new_n2018, new_n9358);
nand_5 g08973(new_n9358, new_n1726, new_n9359);
nand_5 g08974(new_n9359, new_n1722, new_n9360);
nand_5 g08975(new_n9360, new_n1718, new_n9361);
nand_5 g08976(new_n9361, new_n1713, new_n9362);
nand_5 g08977(new_n9362, new_n1737, new_n9363);
nand_5 g08978(new_n9363, new_n1709, new_n9364);
nand_5 g08979(new_n9364, new_n1742, new_n9365);
nand_5 g08980(new_n9365, new_n1704, new_n9366);
nand_5 g08981(new_n9366, new_n1702_1, new_n9367);
nand_5 g08982(new_n9367, new_n1698, new_n9368);
nand_5 g08983(new_n9368, new_n1695, new_n9369);
nand_5 g08984(new_n9369, new_n1692, new_n9370);
nand_5 g08985(new_n9370, new_n1752, new_n9371);
nand_5 g08986(new_n9371, new_n1688, new_n9372);
nand_5 g08987(new_n9372, new_n1685, new_n9373);
nand_5 g08988(new_n9373, new_n1680, new_n9374);
nand_5 g08989(new_n9374, new_n1676, new_n9375);
nand_5 g08990(new_n9375, new_n1672, new_n9376);
nand_5 g08991(new_n9376, new_n1669, new_n9377);
nand_5 g08992(new_n9377, new_n1666, new_n9378);
nand_5 g08993(new_n9378, new_n1663, new_n9379);
nand_5 g08994(new_n9379, new_n1658, new_n9380);
nand_5 g08995(new_n9380, new_n1653, new_n9381);
nand_5 g08996(new_n9381, new_n1651, new_n9382);
nand_5 g08997(new_n9382, new_n1649, new_n9383);
nand_5 g08998(new_n9383, new_n1646, new_n9384);
nand_5 g08999(new_n9384, new_n1643, new_n9385);
nand_5 g09000(new_n9385, new_n1641, new_n9386);
nand_5 g09001(new_n9386, new_n1638, new_n9387);
nand_5 g09002(new_n9387, new_n1635, new_n9388);
nand_5 g09003(new_n9388, new_n1632, new_n9389);
nand_5 g09004(new_n9389, new_n1628, new_n9390);
nand_5 g09005(new_n9390, new_n1625, new_n9391);
nand_5 g09006(new_n9391, new_n1621, new_n9392);
nand_5 g09007(new_n9392, new_n1618, new_n9393);
nand_5 g09008(new_n9393, new_n1778, new_n9394);
nand_5 g09009(new_n9394, new_n1782, new_n9395);
nand_5 g09010(new_n9395, new_n1614, new_n9396);
nand_5 g09011(new_n9396, new_n1611, new_n9397);
nand_5 g09012(new_n9397, new_n1789, new_n9398);
nand_5 g09013(new_n9398, new_n1608, new_n9399);
nand_5 g09014(new_n9399, new_n1605, new_n9400);
nand_5 g09015(new_n9400, new_n1795, new_n9401);
nand_5 g09016(new_n9401, new_n1799, new_n9402);
nand_5 g09017(new_n9402, new_n1602, new_n9403);
nand_5 g09018(new_n9403, new_n1599, new_n9404);
nand_5 g09019(new_n9404, new_n1596, new_n9405);
nand_5 g09020(new_n9405, n4154, new_n9406);
nor_5  g09021(new_n9406, new_n1590, n10515);
nand_5 g09022(new_n872, new_n863, new_n9408);
nand_5 g09023(new_n9408, new_n878, new_n9409);
nand_5 g09024(new_n9409, new_n407, new_n9410);
nand_5 g09025(new_n9410, new_n885, new_n9411);
nand_5 g09026(new_n9411, new_n402, new_n9412);
nand_5 g09027(new_n9412, new_n397, new_n9413);
nand_5 g09028(new_n9413, new_n392, new_n9414);
nand_5 g09029(new_n9414, new_n894, new_n9415);
nand_5 g09030(new_n9415, new_n1087, new_n9416);
nand_5 g09031(new_n9416, new_n1129, new_n9417);
nand_5 g09032(new_n9417, new_n1084, new_n9418);
nand_5 g09033(new_n9418, new_n1134, new_n9419);
nand_5 g09034(new_n9419, new_n1080, new_n9420);
nand_5 g09035(new_n9420, new_n1075, new_n9421);
nand_5 g09036(new_n9421, new_n1070, new_n9422);
nand_5 g09037(new_n9422, new_n1143, new_n9423);
nand_5 g09038(new_n9423, new_n1148, new_n9424);
nand_5 g09039(new_n9424, new_n1065, new_n9425);
nand_5 g09040(new_n9425, new_n1062, new_n9426);
nand_5 g09041(new_n9426, new_n1156, new_n9427);
nand_5 g09042(new_n9427, new_n1057, new_n9428);
nand_5 g09043(new_n9428, new_n1053, new_n9429);
nand_5 g09044(new_n9429, new_n1050, new_n9430);
nand_5 g09045(new_n9430, new_n1045, new_n9431);
nand_5 g09046(new_n9431, new_n1040, new_n9432);
nand_5 g09047(new_n9432, new_n1036, new_n9433);
nand_5 g09048(new_n9433, new_n1033, new_n9434);
nand_5 g09049(new_n9434, new_n1028, new_n9435);
nand_5 g09050(new_n9435, new_n1026, new_n9436);
nand_5 g09051(new_n9436, new_n1021, new_n9437_1);
nand_5 g09052(new_n9437_1, new_n1017, new_n9438);
nand_5 g09053(new_n9438, new_n1012, new_n9439);
nand_5 g09054(new_n9439, new_n1009, new_n9440);
nand_5 g09055(new_n9440, new_n1004, new_n9441);
nand_5 g09056(new_n9441, new_n1000, new_n9442);
nand_5 g09057(new_n9442, new_n995, new_n9443);
nand_5 g09058(new_n9443, new_n990, new_n9444);
nand_5 g09059(new_n9444, new_n985, new_n9445);
nand_5 g09060(new_n9445, new_n981, new_n9446);
nand_5 g09061(new_n9446, new_n1179, new_n9447_1);
nand_5 g09062(new_n9447_1, new_n976, new_n9448);
nand_5 g09063(new_n9448, new_n971, new_n9449);
nand_5 g09064(new_n9449, new_n966, new_n9450);
nand_5 g09065(new_n9450, new_n961, new_n9451);
nand_5 g09066(new_n9451, new_n957, new_n9452);
nand_5 g09067(new_n9452, new_n952, new_n9453);
nand_5 g09068(new_n9453, new_n948_1, new_n9454);
nand_5 g09069(new_n9454, new_n943, new_n9455);
nand_5 g09070(new_n9455, new_n941, new_n9456);
nand_5 g09071(new_n9456, new_n938, new_n9457);
nand_5 g09072(new_n9457, new_n936, new_n9458);
nand_5 g09073(new_n9458, new_n931, new_n9459);
nand_5 g09074(new_n9459, new_n927, new_n9460);
nand_5 g09075(new_n9460, new_n922, new_n9461);
nand_5 g09076(new_n9461, new_n917, new_n9462);
nand_5 g09077(new_n9462, new_n912, new_n9463);
nand_5 g09078(new_n9463, new_n907, new_n9464);
nand_5 g09079(new_n9464, new_n903, new_n9465);
nand_5 g09080(new_n9465, new_n2066, new_n9466);
nand_5 g09081(new_n9466, new_n2063, new_n9467);
nand_5 g09082(new_n9467, new_n2062, new_n9468);
nand_5 g09083(new_n9468, new_n2058, new_n9469);
nand_5 g09084(new_n9469, new_n2055, new_n9470);
nand_5 g09085(new_n9470, new_n2051, new_n9471);
nand_5 g09086(new_n9471, new_n2046, new_n9472);
nand_5 g09087(new_n9472, new_n2042, new_n9473);
nand_5 g09088(new_n9473, new_n2039, new_n9474);
nand_5 g09089(new_n9474, new_n2036, new_n9475);
nand_5 g09090(new_n9475, new_n2033, new_n9476);
nand_5 g09091(new_n9476, new_n2029, new_n9477);
nand_5 g09092(new_n9477, new_n2026, new_n9478);
nand_5 g09093(new_n9478, new_n2022, new_n9479);
nand_5 g09094(new_n9479, new_n2018, new_n9480);
nand_5 g09095(new_n9480, new_n1726, new_n9481);
nand_5 g09096(new_n9481, new_n1722, new_n9482);
nand_5 g09097(new_n9482, new_n1718, new_n9483);
nand_5 g09098(new_n9483, new_n1713, new_n9484);
nand_5 g09099(new_n9484, new_n1737, new_n9485);
nand_5 g09100(new_n9485, new_n1709, new_n9486);
nand_5 g09101(new_n9486, new_n1742, new_n9487);
nand_5 g09102(new_n9487, new_n1704, new_n9488);
nand_5 g09103(new_n9488, new_n1702_1, new_n9489);
nand_5 g09104(new_n9489, new_n1698, new_n9490);
nand_5 g09105(new_n9490, new_n1695, new_n9491);
nand_5 g09106(new_n9491, n3910, new_n9492);
nor_5  g09107(new_n9492, new_n1689, n10591);
nand_5 g09108(new_n1292, new_n769, new_n9494);
nand_5 g09109(new_n9494, new_n1355, new_n9495);
nand_5 g09110(new_n9495, new_n1291, new_n9496);
nand_5 g09111(new_n9496, new_n1288, new_n9497);
nand_5 g09112(new_n9497, new_n1283, new_n9498);
nand_5 g09113(new_n9498, new_n1363, new_n9499);
nand_5 g09114(new_n9499, new_n1280, new_n9500);
nand_5 g09115(new_n9500, new_n1370, new_n9501);
nand_5 g09116(new_n9501, new_n1373, new_n9502);
nand_5 g09117(new_n9502, new_n1277, new_n9503);
nand_5 g09118(new_n9503, new_n1272, new_n9504);
nand_5 g09119(new_n9504, new_n1269, new_n9505);
nand_5 g09120(new_n9505, new_n1380, new_n9506);
nand_5 g09121(new_n9506, new_n1264, new_n9507);
nand_5 g09122(new_n9507, new_n1259, new_n9508);
nand_5 g09123(new_n9508, new_n1388, new_n9509);
nand_5 g09124(new_n9509, new_n1392, new_n9510);
nand_5 g09125(new_n9510, new_n1256, new_n9511);
nand_5 g09126(new_n9511, new_n1252, new_n9512);
nand_5 g09127(new_n9512, new_n1249, new_n9513);
nand_5 g09128(new_n9513, new_n1244, new_n9514);
nand_5 g09129(new_n9514, new_n1240, new_n9515);
nand_5 g09130(new_n9515, new_n1234, new_n9516);
nand_5 g09131(new_n9516, new_n1231, new_n9517);
nand_5 g09132(new_n9517, new_n1227, new_n9518);
nand_5 g09133(new_n9518, new_n1407, new_n9519);
nand_5 g09134(new_n9519, new_n1223, new_n9520);
nand_5 g09135(new_n9520, new_n1218, new_n9521);
nand_5 g09136(new_n9521, new_n1213, new_n9522);
nand_5 g09137(new_n9522, new_n1210, new_n9523);
nand_5 g09138(new_n9523, new_n1206, new_n9524);
nand_5 g09139(new_n9524, new_n1418, new_n9525);
nand_5 g09140(new_n9525, new_n1422, new_n9526);
nand_5 g09141(new_n9526, new_n1428, new_n9527);
nand_5 g09142(new_n9527, new_n1203, new_n9528);
nand_5 g09143(new_n9528, new_n1433, new_n9529);
nand_5 g09144(new_n9529, new_n581, new_n9530);
nand_5 g09145(new_n9530, new_n574, new_n9531);
nand_5 g09146(new_n9531, new_n568, new_n9532);
nand_5 g09147(new_n9532, new_n589, new_n9533);
nand_5 g09148(new_n9533, new_n595, new_n9534);
nand_5 g09149(new_n9534, new_n601, new_n9535);
nand_5 g09150(new_n9535, new_n563, new_n9536);
nand_5 g09151(new_n9536, new_n608, new_n9537);
nand_5 g09152(new_n9537, new_n558, new_n9538);
nand_5 g09153(new_n9538, new_n615, new_n9539);
nand_5 g09154(new_n9539, new_n553, new_n9540);
nand_5 g09155(new_n9540, new_n622, new_n9541);
nand_5 g09156(new_n9541, new_n628, new_n9542);
nand_5 g09157(new_n9542, new_n548, new_n9543_1);
nand_5 g09158(new_n9543_1, new_n543_1, new_n9544_1);
nand_5 g09159(new_n9544_1, new_n636, new_n9545);
nand_5 g09160(new_n9545, new_n642, new_n9546);
nand_5 g09161(new_n9546, new_n538, new_n9547);
nand_5 g09162(new_n9547, new_n533, new_n9548);
nand_5 g09163(new_n9548, new_n650_1, new_n9549);
nand_5 g09164(new_n9549, new_n528, new_n9550);
nand_5 g09165(new_n9550, new_n523, new_n9551);
nand_5 g09166(new_n9551, new_n518, new_n9552);
nand_5 g09167(new_n9552, new_n659, new_n9553);
nand_5 g09168(new_n9553, new_n665, new_n9554);
nand_5 g09169(new_n9554, new_n672, new_n9555_1);
nand_5 g09170(new_n9555_1, new_n513, new_n9556);
nand_5 g09171(new_n9556, new_n679, new_n9557);
nand_5 g09172(new_n9557, new_n685, new_n9558);
nand_5 g09173(new_n9558, new_n691, new_n9559);
nand_5 g09174(new_n9559, new_n508, new_n9560);
nand_5 g09175(new_n9560, new_n698, new_n9561);
nand_5 g09176(new_n9561, new_n503, new_n9562);
nand_5 g09177(new_n9562, new_n704, new_n9563);
nand_5 g09178(new_n9563, new_n498_1, new_n9564);
nand_5 g09179(new_n9564, new_n711, new_n9565);
nand_5 g09180(new_n9565, new_n493, new_n9566);
nand_5 g09181(new_n9566, new_n718, new_n9567);
nand_5 g09182(new_n9567, new_n488, new_n9568);
nand_5 g09183(new_n9568, new_n725, new_n9569);
nand_5 g09184(new_n9569, new_n483, new_n9570_1);
nand_5 g09185(new_n9570_1, new_n732, new_n9571);
nand_5 g09186(new_n9571, new_n478, new_n9572);
nand_5 g09187(new_n9572, new_n739, new_n9573);
nand_5 g09188(new_n9573, new_n745, new_n9574);
nand_5 g09189(new_n9574, new_n751, new_n9575);
nand_5 g09190(new_n9575, new_n473, new_n9576);
nand_5 g09191(new_n9576, new_n758, new_n9577);
nand_5 g09192(new_n9577, n10378, new_n9578);
nor_5  g09193(new_n9578, new_n761, n10791);
nand_5 g09194(new_n1694, new_n410, new_n9580);
nand_5 g09195(new_n9580, new_n866, new_n9581);
nand_5 g09196(new_n9581, new_n872, new_n9582);
nand_5 g09197(new_n9582, new_n878, new_n9583);
nand_5 g09198(new_n9583, new_n407, new_n9584);
nand_5 g09199(new_n9584, new_n885, new_n9585);
nand_5 g09200(new_n9585, new_n402, new_n9586);
nand_5 g09201(new_n9586, new_n397, new_n9587);
nand_5 g09202(new_n9587, new_n392, new_n9588);
nand_5 g09203(new_n9588, new_n894, new_n9589_1);
nand_5 g09204(new_n9589_1, new_n1087, new_n9590);
nand_5 g09205(new_n9590, new_n1129, new_n9591);
nand_5 g09206(new_n9591, new_n1084, new_n9592);
nand_5 g09207(new_n9592, new_n1134, new_n9593);
nand_5 g09208(new_n9593, new_n1080, new_n9594);
nand_5 g09209(new_n9594, new_n1075, new_n9595);
nand_5 g09210(new_n9595, new_n1070, new_n9596);
nand_5 g09211(new_n9596, new_n1143, new_n9597);
nand_5 g09212(new_n9597, new_n1148, new_n9598);
nand_5 g09213(new_n9598, new_n1065, new_n9599);
nand_5 g09214(new_n9599, new_n1062, new_n9600);
nand_5 g09215(new_n9600, new_n1156, new_n9601);
nand_5 g09216(new_n9601, new_n1057, new_n9602);
nand_5 g09217(new_n9602, new_n1053, new_n9603);
nand_5 g09218(new_n9603, new_n1050, new_n9604);
nand_5 g09219(new_n9604, new_n1045, new_n9605);
nand_5 g09220(new_n9605, new_n1040, new_n9606);
nand_5 g09221(new_n9606, new_n1036, new_n9607);
nand_5 g09222(new_n9607, new_n1033, new_n9608);
nand_5 g09223(new_n9608, new_n1028, new_n9609);
nand_5 g09224(new_n9609, new_n1026, new_n9610);
nand_5 g09225(new_n9610, new_n1021, new_n9611);
nand_5 g09226(new_n9611, new_n1017, new_n9612);
nand_5 g09227(new_n9612, new_n1012, new_n9613);
nand_5 g09228(new_n9613, new_n1009, new_n9614);
nand_5 g09229(new_n9614, new_n1004, new_n9615);
nand_5 g09230(new_n9615, new_n1000, new_n9616);
nand_5 g09231(new_n9616, new_n995, new_n9617);
nand_5 g09232(new_n9617, new_n990, new_n9618);
nand_5 g09233(new_n9618, new_n985, new_n9619);
nand_5 g09234(new_n9619, new_n981, new_n9620);
nand_5 g09235(new_n9620, new_n1179, new_n9621);
nand_5 g09236(new_n9621, new_n976, new_n9622);
nand_5 g09237(new_n9622, new_n971, new_n9623);
nand_5 g09238(new_n9623, new_n966, new_n9624);
nand_5 g09239(new_n9624, new_n961, new_n9625);
nand_5 g09240(new_n9625, new_n957, new_n9626);
nand_5 g09241(new_n9626, new_n952, new_n9627);
nand_5 g09242(new_n9627, new_n948_1, new_n9628);
nand_5 g09243(new_n9628, new_n943, new_n9629);
nand_5 g09244(new_n9629, new_n941, new_n9630);
nand_5 g09245(new_n9630, new_n938, new_n9631);
nand_5 g09246(new_n9631, new_n936, new_n9632);
nand_5 g09247(new_n9632, new_n931, new_n9633);
nand_5 g09248(new_n9633, new_n927, new_n9634);
nand_5 g09249(new_n9634, new_n922, new_n9635);
nand_5 g09250(new_n9635, new_n917, new_n9636);
nand_5 g09251(new_n9636, new_n912, new_n9637);
nand_5 g09252(new_n9637, new_n907, new_n9638);
nand_5 g09253(new_n9638, new_n903, new_n9639);
nand_5 g09254(new_n9639, new_n2066, new_n9640);
nand_5 g09255(new_n9640, new_n2063, new_n9641);
nand_5 g09256(new_n9641, new_n2062, new_n9642);
nand_5 g09257(new_n9642, new_n2058, new_n9643);
nand_5 g09258(new_n9643, new_n2055, new_n9644);
nand_5 g09259(new_n9644, new_n2051, new_n9645);
nand_5 g09260(new_n9645, new_n2046, new_n9646);
nand_5 g09261(new_n9646, new_n2042, new_n9647);
nand_5 g09262(new_n9647, new_n2039, new_n9648);
nand_5 g09263(new_n9648, new_n2036, new_n9649);
nand_5 g09264(new_n9649, new_n2033, new_n9650);
nand_5 g09265(new_n9650, new_n2029, new_n9651);
nand_5 g09266(new_n9651, new_n2026, new_n9652);
nand_5 g09267(new_n9652, new_n2022, new_n9653);
nand_5 g09268(new_n9653, new_n2018, new_n9654);
nand_5 g09269(new_n9654, new_n1726, new_n9655);
nand_5 g09270(new_n9655, new_n1722, new_n9656);
nand_5 g09271(new_n9656, new_n1718, new_n9657);
nand_5 g09272(new_n9657, new_n1713, new_n9658);
nand_5 g09273(new_n9658, new_n1737, new_n9659);
nand_5 g09274(new_n9659, new_n1709, new_n9660);
nand_5 g09275(new_n9660, new_n1742, new_n9661);
nand_5 g09276(new_n9661, new_n1704, new_n9662);
nand_5 g09277(new_n9662, new_n1702_1, new_n9663);
nand_5 g09278(new_n9663, n13186, new_n9664);
nor_5  g09279(new_n9664, new_n1228, n10802);
nand_5 g09280(new_n1716, new_n1254, new_n9666);
nand_5 g09281(new_n9666, new_n420, new_n9667);
nand_5 g09282(new_n9667, new_n828, new_n9668);
nand_5 g09283(new_n9668, new_n834, new_n9669);
nand_5 g09284(new_n9669, new_n840, new_n9670);
nand_5 g09285(new_n9670, new_n417, new_n9671);
nand_5 g09286(new_n9671, new_n847, new_n9672);
nand_5 g09287(new_n9672, new_n853, new_n9673);
nand_5 g09288(new_n9673, new_n859, new_n9674);
nand_5 g09289(new_n9674, new_n412, new_n9675);
nand_5 g09290(new_n9675, new_n866, new_n9676);
nand_5 g09291(new_n9676, new_n872, new_n9677);
nand_5 g09292(new_n9677, new_n878, new_n9678);
nand_5 g09293(new_n9678, new_n407, new_n9679);
nand_5 g09294(new_n9679, new_n885, new_n9680);
nand_5 g09295(new_n9680, new_n402, new_n9681);
nand_5 g09296(new_n9681, new_n397, new_n9682);
nand_5 g09297(new_n9682, new_n392, new_n9683);
nand_5 g09298(new_n9683, new_n894, new_n9684);
nand_5 g09299(new_n9684, new_n1087, new_n9685);
nand_5 g09300(new_n9685, new_n1129, new_n9686);
nand_5 g09301(new_n9686, new_n1084, new_n9687);
nand_5 g09302(new_n9687, new_n1134, new_n9688);
nand_5 g09303(new_n9688, new_n1080, new_n9689);
nand_5 g09304(new_n9689, new_n1075, new_n9690);
nand_5 g09305(new_n9690, new_n1070, new_n9691);
nand_5 g09306(new_n9691, new_n1143, new_n9692);
nand_5 g09307(new_n9692, new_n1148, new_n9693);
nand_5 g09308(new_n9693, new_n1065, new_n9694);
nand_5 g09309(new_n9694, new_n1062, new_n9695);
nand_5 g09310(new_n9695, new_n1156, new_n9696);
nand_5 g09311(new_n9696, new_n1057, new_n9697);
nand_5 g09312(new_n9697, new_n1053, new_n9698);
nand_5 g09313(new_n9698, new_n1050, new_n9699);
nand_5 g09314(new_n9699, new_n1045, new_n9700);
nand_5 g09315(new_n9700, new_n1040, new_n9701);
nand_5 g09316(new_n9701, new_n1036, new_n9702);
nand_5 g09317(new_n9702, new_n1033, new_n9703);
nand_5 g09318(new_n9703, new_n1028, new_n9704);
nand_5 g09319(new_n9704, new_n1026, new_n9705);
nand_5 g09320(new_n9705, new_n1021, new_n9706);
nand_5 g09321(new_n9706, new_n1017, new_n9707);
nand_5 g09322(new_n9707, new_n1012, new_n9708);
nand_5 g09323(new_n9708, new_n1009, new_n9709);
nand_5 g09324(new_n9709, new_n1004, new_n9710);
nand_5 g09325(new_n9710, new_n1000, new_n9711);
nand_5 g09326(new_n9711, new_n995, new_n9712);
nand_5 g09327(new_n9712, new_n990, new_n9713);
nand_5 g09328(new_n9713, new_n985, new_n9714);
nand_5 g09329(new_n9714, new_n981, new_n9715);
nand_5 g09330(new_n9715, new_n1179, new_n9716);
nand_5 g09331(new_n9716, new_n976, new_n9717_1);
nand_5 g09332(new_n9717_1, new_n971, new_n9718);
nand_5 g09333(new_n9718, new_n966, new_n9719);
nand_5 g09334(new_n9719, new_n961, new_n9720);
nand_5 g09335(new_n9720, new_n957, new_n9721);
nand_5 g09336(new_n9721, new_n952, new_n9722);
nand_5 g09337(new_n9722, new_n948_1, new_n9723);
nand_5 g09338(new_n9723, new_n943, new_n9724);
nand_5 g09339(new_n9724, new_n941, new_n9725);
nand_5 g09340(new_n9725, new_n938, new_n9726);
nand_5 g09341(new_n9726, new_n936, new_n9727);
nand_5 g09342(new_n9727, new_n931, new_n9728);
nand_5 g09343(new_n9728, new_n927, new_n9729);
nand_5 g09344(new_n9729, new_n922, new_n9730);
nand_5 g09345(new_n9730, new_n917, new_n9731);
nand_5 g09346(new_n9731, new_n912, new_n9732);
nand_5 g09347(new_n9732, new_n907, new_n9733);
nand_5 g09348(new_n9733, new_n903, new_n9734);
nand_5 g09349(new_n9734, new_n2066, new_n9735);
nand_5 g09350(new_n9735, new_n2063, new_n9736);
nand_5 g09351(new_n9736, new_n2062, new_n9737);
nand_5 g09352(new_n9737, new_n2058, new_n9738);
nand_5 g09353(new_n9738, new_n2055, new_n9739);
nand_5 g09354(new_n9739, new_n2051, new_n9740);
nand_5 g09355(new_n9740, new_n2046, new_n9741);
nand_5 g09356(new_n9741, new_n2042, new_n9742);
nand_5 g09357(new_n9742, new_n2039, new_n9743);
nand_5 g09358(new_n9743, new_n2036, new_n9744);
nand_5 g09359(new_n9744, new_n2033, new_n9745);
nand_5 g09360(new_n9745, new_n2029, new_n9746);
nand_5 g09361(new_n9746, new_n2026, new_n9747);
nand_5 g09362(new_n9747, new_n2022, new_n9748);
nand_5 g09363(new_n9748, new_n2018, new_n9749);
nand_5 g09364(new_n9749, new_n1726, new_n9750);
nand_5 g09365(new_n9750, n7667, new_n9751);
nor_5  g09366(new_n9751, new_n1719, n10915);
nand_5 g09367(new_n1682, new_n1680, new_n9753);
nand_5 g09368(new_n9753, new_n1676, new_n9754);
nand_5 g09369(new_n9754, new_n1672, new_n9755);
nand_5 g09370(new_n9755, new_n1669, new_n9756);
nand_5 g09371(new_n9756, new_n1666, new_n9757);
nand_5 g09372(new_n9757, new_n1663, new_n9758);
nand_5 g09373(new_n9758, new_n1658, new_n9759);
nand_5 g09374(new_n9759, new_n1653, new_n9760);
nand_5 g09375(new_n9760, new_n1651, new_n9761);
nand_5 g09376(new_n9761, new_n1649, new_n9762);
nand_5 g09377(new_n9762, new_n1646, new_n9763);
nand_5 g09378(new_n9763, new_n1643, new_n9764);
nand_5 g09379(new_n9764, new_n1641, new_n9765);
nand_5 g09380(new_n9765, new_n1638, new_n9766);
nand_5 g09381(new_n9766, new_n1635, new_n9767);
nand_5 g09382(new_n9767, new_n1632, new_n9768);
nand_5 g09383(new_n9768, new_n1628, new_n9769);
nand_5 g09384(new_n9769, new_n1625, new_n9770);
nand_5 g09385(new_n9770, new_n1621, new_n9771);
nand_5 g09386(new_n9771, new_n1618, new_n9772);
nand_5 g09387(new_n9772, new_n1778, new_n9773);
nand_5 g09388(new_n9773, new_n1782, new_n9774);
nand_5 g09389(new_n9774, new_n1614, new_n9775);
nand_5 g09390(new_n9775, new_n1611, new_n9776);
nand_5 g09391(new_n9776, new_n1789, new_n9777);
nand_5 g09392(new_n9777, new_n1608, new_n9778);
nand_5 g09393(new_n9778, new_n1605, new_n9779);
nand_5 g09394(new_n9779, new_n1795, new_n9780);
nand_5 g09395(new_n9780, new_n1799, new_n9781);
nand_5 g09396(new_n9781, new_n1602, new_n9782);
nand_5 g09397(new_n9782, new_n1599, new_n9783);
nand_5 g09398(new_n9783, new_n1596, new_n9784);
nand_5 g09399(new_n9784, new_n1593, new_n9785);
nand_5 g09400(new_n9785, new_n1806, new_n9786);
nand_5 g09401(new_n9786, new_n1589, new_n9787);
nand_5 g09402(new_n9787, new_n1586, new_n9788);
nand_5 g09403(new_n9788, new_n1583, new_n9789);
nand_5 g09404(new_n9789, new_n1580, new_n9790);
nand_5 g09405(new_n9790, new_n1576, new_n9791);
nand_5 g09406(new_n9791, new_n1573, new_n9792);
nand_5 g09407(new_n9792, new_n1570, new_n9793);
nand_5 g09408(new_n9793, new_n1567, new_n9794);
nand_5 g09409(new_n9794, new_n1564, new_n9795);
nand_5 g09410(new_n9795, new_n1561, new_n9796);
nand_5 g09411(new_n9796, new_n1338, new_n9797);
nand_5 g09412(new_n9797, new_n1331, new_n9798);
nand_5 g09413(new_n9798, new_n1326, new_n9799);
nand_5 g09414(new_n9799, new_n1321, new_n9800);
nand_5 g09415(new_n9800, new_n1318, new_n9801);
nand_5 g09416(new_n9801, new_n1315, new_n9802);
nand_5 g09417(new_n9802, new_n1312, new_n9803);
nand_5 g09418(new_n9803, new_n1309, new_n9804);
nand_5 g09419(new_n9804, new_n1307, new_n9805);
nand_5 g09420(new_n9805, new_n1304, new_n9806);
nand_5 g09421(new_n9806, new_n1300, new_n9807);
nand_5 g09422(new_n9807, new_n1297, new_n9808);
nand_5 g09423(new_n9808, new_n1294, new_n9809);
nand_5 g09424(new_n9809, new_n1355, new_n9810);
nand_5 g09425(new_n9810, new_n1291, new_n9811);
nand_5 g09426(new_n9811, new_n1288, new_n9812);
nand_5 g09427(new_n9812, new_n1283, new_n9813);
nand_5 g09428(new_n9813, new_n1363, new_n9814);
nand_5 g09429(new_n9814, new_n1280, new_n9815);
nand_5 g09430(new_n9815, new_n1370, new_n9816);
nand_5 g09431(new_n9816, new_n1373, new_n9817);
nand_5 g09432(new_n9817, new_n1277, new_n9818);
nand_5 g09433(new_n9818, new_n1272, new_n9819);
nand_5 g09434(new_n9819, new_n1269, new_n9820);
nand_5 g09435(new_n9820, new_n1380, new_n9821);
nand_5 g09436(new_n9821, new_n1264, new_n9822);
nand_5 g09437(new_n9822, new_n1259, new_n9823);
nand_5 g09438(new_n9823, new_n1388, new_n9824);
nand_5 g09439(new_n9824, new_n1392, new_n9825);
nand_5 g09440(new_n9825, new_n1256, new_n9826);
nand_5 g09441(new_n9826, new_n1252, new_n9827);
nand_5 g09442(new_n9827, new_n1249, new_n9828);
nand_5 g09443(new_n9828, new_n1244, new_n9829);
nand_5 g09444(new_n9829, new_n1240, new_n9830_1);
nand_5 g09445(new_n9830_1, new_n1234, new_n9831);
nand_5 g09446(new_n9831, new_n1231, new_n9832);
nand_5 g09447(new_n9832, new_n1227, new_n9833);
nand_5 g09448(new_n9833, new_n1407, new_n9834);
nand_5 g09449(new_n9834, new_n1223, new_n9835);
nand_5 g09450(new_n9835, new_n1218, new_n9836);
nand_5 g09451(new_n9836, n8649, new_n9837);
nor_5  g09452(new_n9837, new_n875, n11122);
nand_5 g09453(new_n1225, new_n858, new_n9839);
nand_5 g09454(new_n9839, new_n1407, new_n9840);
nand_5 g09455(new_n9840, new_n1223, new_n9841);
nand_5 g09456(new_n9841, new_n1218, new_n9842);
nand_5 g09457(new_n9842, new_n1213, new_n9843);
nand_5 g09458(new_n9843, new_n1210, new_n9844);
nand_5 g09459(new_n9844, new_n1206, new_n9845);
nand_5 g09460(new_n9845, new_n1418, new_n9846);
nand_5 g09461(new_n9846, new_n1422, new_n9847);
nand_5 g09462(new_n9847, new_n1428, new_n9848);
nand_5 g09463(new_n9848, new_n1203, new_n9849);
nand_5 g09464(new_n9849, new_n1433, new_n9850);
nand_5 g09465(new_n9850, new_n581, new_n9851);
nand_5 g09466(new_n9851, new_n574, new_n9852);
nand_5 g09467(new_n9852, new_n568, new_n9853);
nand_5 g09468(new_n9853, new_n589, new_n9854);
nand_5 g09469(new_n9854, new_n595, new_n9855);
nand_5 g09470(new_n9855, new_n601, new_n9856);
nand_5 g09471(new_n9856, new_n563, new_n9857);
nand_5 g09472(new_n9857, new_n608, new_n9858);
nand_5 g09473(new_n9858, new_n558, new_n9859);
nand_5 g09474(new_n9859, new_n615, new_n9860);
nand_5 g09475(new_n9860, new_n553, new_n9861);
nand_5 g09476(new_n9861, new_n622, new_n9862);
nand_5 g09477(new_n9862, new_n628, new_n9863);
nand_5 g09478(new_n9863, new_n548, new_n9864);
nand_5 g09479(new_n9864, new_n543_1, new_n9865);
nand_5 g09480(new_n9865, new_n636, new_n9866);
nand_5 g09481(new_n9866, new_n642, new_n9867);
nand_5 g09482(new_n9867, new_n538, new_n9868);
nand_5 g09483(new_n9868, new_n533, new_n9869);
nand_5 g09484(new_n9869, new_n650_1, new_n9870);
nand_5 g09485(new_n9870, new_n528, new_n9871);
nand_5 g09486(new_n9871, new_n523, new_n9872);
nand_5 g09487(new_n9872, new_n518, new_n9873);
nand_5 g09488(new_n9873, new_n659, new_n9874);
nand_5 g09489(new_n9874, new_n665, new_n9875);
nand_5 g09490(new_n9875, new_n672, new_n9876);
nand_5 g09491(new_n9876, new_n513, new_n9877);
nand_5 g09492(new_n9877, new_n679, new_n9878);
nand_5 g09493(new_n9878, new_n685, new_n9879);
nand_5 g09494(new_n9879, new_n691, new_n9880);
nand_5 g09495(new_n9880, new_n508, new_n9881);
nand_5 g09496(new_n9881, new_n698, new_n9882);
nand_5 g09497(new_n9882, new_n503, new_n9883);
nand_5 g09498(new_n9883, new_n704, new_n9884);
nand_5 g09499(new_n9884, new_n498_1, new_n9885);
nand_5 g09500(new_n9885, new_n711, new_n9886);
nand_5 g09501(new_n9886, new_n493, new_n9887);
nand_5 g09502(new_n9887, new_n718, new_n9888);
nand_5 g09503(new_n9888, new_n488, new_n9889);
nand_5 g09504(new_n9889, new_n725, new_n9890);
nand_5 g09505(new_n9890, new_n483, new_n9891);
nand_5 g09506(new_n9891, new_n732, new_n9892);
nand_5 g09507(new_n9892, new_n478, new_n9893_1);
nand_5 g09508(new_n9893_1, new_n739, new_n9894);
nand_5 g09509(new_n9894, new_n745, new_n9895);
nand_5 g09510(new_n9895, new_n751, new_n9896);
nand_5 g09511(new_n9896, new_n473, new_n9897);
nand_5 g09512(new_n9897, new_n758, new_n9898);
nand_5 g09513(new_n9898, new_n764, new_n9899);
nand_5 g09514(new_n9899, new_n770, new_n9900);
nand_5 g09515(new_n9900, new_n468, new_n9901);
nand_5 g09516(new_n9901, new_n777, new_n9902);
nand_5 g09517(new_n9902, new_n783, new_n9903);
nand_5 g09518(new_n9903, new_n789, new_n9904);
nand_5 g09519(new_n9904, new_n463, new_n9905);
nand_5 g09520(new_n9905, new_n796, new_n9906);
nand_5 g09521(new_n9906, new_n458, new_n9907);
nand_5 g09522(new_n9907, new_n453, new_n9908);
nand_5 g09523(new_n9908, new_n447, new_n9909);
nand_5 g09524(new_n9909, new_n805, new_n9910);
nand_5 g09525(new_n9910, new_n811, new_n9911);
nand_5 g09526(new_n9911, new_n442, new_n9912);
nand_5 g09527(new_n9912, new_n437, new_n9913);
nand_5 g09528(new_n9913, new_n819, new_n9914);
nand_5 g09529(new_n9914, new_n432, new_n9915);
nand_5 g09530(new_n9915, new_n427_1, new_n9916);
nand_5 g09531(new_n9916, new_n422, new_n9917);
nand_5 g09532(new_n9917, new_n828, new_n9918);
nand_5 g09533(new_n9918, new_n834, new_n9919);
nand_5 g09534(new_n9919, new_n840, new_n9920);
nand_5 g09535(new_n9920, new_n417, new_n9921_1);
nand_5 g09536(new_n9921_1, new_n847, new_n9922);
nand_5 g09537(new_n9922, n7748, new_n9923);
nor_5  g09538(new_n9923, new_n1699, n11393);
nand_5 g09539(new_n837, new_n417, new_n9925);
nand_5 g09540(new_n9925, new_n847, new_n9926);
nand_5 g09541(new_n9926, new_n853, new_n9927);
nand_5 g09542(new_n9927, new_n859, new_n9928);
nand_5 g09543(new_n9928, new_n412, new_n9929);
nand_5 g09544(new_n9929, new_n866, new_n9930);
nand_5 g09545(new_n9930, new_n872, new_n9931);
nand_5 g09546(new_n9931, new_n878, new_n9932);
nand_5 g09547(new_n9932, new_n407, new_n9933);
nand_5 g09548(new_n9933, new_n885, new_n9934);
nand_5 g09549(new_n9934, new_n402, new_n9935);
nand_5 g09550(new_n9935, new_n397, new_n9936_1);
nand_5 g09551(new_n9936_1, new_n392, new_n9937);
nand_5 g09552(new_n9937, new_n894, new_n9938);
nand_5 g09553(new_n9938, new_n1087, new_n9939);
nand_5 g09554(new_n9939, new_n1129, new_n9940);
nand_5 g09555(new_n9940, new_n1084, new_n9941);
nand_5 g09556(new_n9941, new_n1134, new_n9942);
nand_5 g09557(new_n9942, new_n1080, new_n9943);
nand_5 g09558(new_n9943, new_n1075, new_n9944);
nand_5 g09559(new_n9944, new_n1070, new_n9945);
nand_5 g09560(new_n9945, new_n1143, new_n9946);
nand_5 g09561(new_n9946, new_n1148, new_n9947);
nand_5 g09562(new_n9947, new_n1065, new_n9948);
nand_5 g09563(new_n9948, new_n1062, new_n9949);
nand_5 g09564(new_n9949, new_n1156, new_n9950);
nand_5 g09565(new_n9950, new_n1057, new_n9951);
nand_5 g09566(new_n9951, new_n1053, new_n9952);
nand_5 g09567(new_n9952, new_n1050, new_n9953);
nand_5 g09568(new_n9953, new_n1045, new_n9954);
nand_5 g09569(new_n9954, new_n1040, new_n9955);
nand_5 g09570(new_n9955, new_n1036, new_n9956);
nand_5 g09571(new_n9956, new_n1033, new_n9957);
nand_5 g09572(new_n9957, new_n1028, new_n9958);
nand_5 g09573(new_n9958, new_n1026, new_n9959);
nand_5 g09574(new_n9959, new_n1021, new_n9960);
nand_5 g09575(new_n9960, new_n1017, new_n9961);
nand_5 g09576(new_n9961, new_n1012, new_n9962);
nand_5 g09577(new_n9962, new_n1009, new_n9963);
nand_5 g09578(new_n9963, new_n1004, new_n9964);
nand_5 g09579(new_n9964, new_n1000, new_n9965);
nand_5 g09580(new_n9965, new_n995, new_n9966);
nand_5 g09581(new_n9966, new_n990, new_n9967);
nand_5 g09582(new_n9967, new_n985, new_n9968);
nand_5 g09583(new_n9968, new_n981, new_n9969);
nand_5 g09584(new_n9969, new_n1179, new_n9970);
nand_5 g09585(new_n9970, new_n976, new_n9971);
nand_5 g09586(new_n9971, new_n971, new_n9972);
nand_5 g09587(new_n9972, new_n966, new_n9973);
nand_5 g09588(new_n9973, new_n961, new_n9974);
nand_5 g09589(new_n9974, new_n957, new_n9975);
nand_5 g09590(new_n9975, new_n952, new_n9976);
nand_5 g09591(new_n9976, new_n948_1, new_n9977_1);
nand_5 g09592(new_n9977_1, new_n943, new_n9978);
nand_5 g09593(new_n9978, new_n941, new_n9979);
nand_5 g09594(new_n9979, new_n938, new_n9980);
nand_5 g09595(new_n9980, new_n936, new_n9981);
nand_5 g09596(new_n9981, new_n931, new_n9982);
nand_5 g09597(new_n9982, new_n927, new_n9983);
nand_5 g09598(new_n9983, new_n922, new_n9984);
nand_5 g09599(new_n9984, new_n917, new_n9985);
nand_5 g09600(new_n9985, new_n912, new_n9986);
nand_5 g09601(new_n9986, new_n907, new_n9987);
nand_5 g09602(new_n9987, new_n903, new_n9988);
nand_5 g09603(new_n9988, new_n2066, new_n9989);
nand_5 g09604(new_n9989, new_n2063, new_n9990);
nand_5 g09605(new_n9990, new_n2062, new_n9991);
nand_5 g09606(new_n9991, new_n2058, new_n9992);
nand_5 g09607(new_n9992, new_n2055, new_n9993);
nand_5 g09608(new_n9993, new_n2051, new_n9994);
nand_5 g09609(new_n9994, new_n2046, new_n9995);
nand_5 g09610(new_n9995, new_n2042, new_n9996);
nand_5 g09611(new_n9996, new_n2039, new_n9997);
nand_5 g09612(new_n9997, new_n2036, new_n9998);
nand_5 g09613(new_n9998, new_n2033, new_n9999);
nand_5 g09614(new_n9999, new_n2029, new_n10000);
nand_5 g09615(new_n10000, new_n2026, new_n10001);
nand_5 g09616(new_n10001, new_n2022, new_n10002);
nand_5 g09617(new_n10002, new_n2018, new_n10003);
nand_5 g09618(new_n10003, new_n1726, new_n10004);
nand_5 g09619(new_n10004, new_n1722, new_n10005);
nand_5 g09620(new_n10005, new_n1718, new_n10006);
nand_5 g09621(new_n10006, new_n1713, new_n10007);
nand_5 g09622(new_n10007, new_n1737, new_n10008);
nand_5 g09623(new_n10008, n13364, new_n10009);
nor_5  g09624(new_n10009, new_n1706, n11463);
nand_5 g09625(new_n942, new_n486, new_n10011);
nand_5 g09626(new_n10011, new_n725, new_n10012);
nand_5 g09627(new_n10012, new_n483, new_n10013);
nand_5 g09628(new_n10013, new_n732, new_n10014);
nand_5 g09629(new_n10014, new_n478, new_n10015);
nand_5 g09630(new_n10015, new_n739, new_n10016);
nand_5 g09631(new_n10016, new_n745, new_n10017);
nand_5 g09632(new_n10017, new_n751, new_n10018);
nand_5 g09633(new_n10018, new_n473, new_n10019);
nand_5 g09634(new_n10019, new_n758, new_n10020);
nand_5 g09635(new_n10020, new_n764, new_n10021);
nand_5 g09636(new_n10021, new_n770, new_n10022);
nand_5 g09637(new_n10022, new_n468, new_n10023);
nand_5 g09638(new_n10023, new_n777, new_n10024);
nand_5 g09639(new_n10024, new_n783, new_n10025);
nand_5 g09640(new_n10025, new_n789, new_n10026);
nand_5 g09641(new_n10026, new_n463, new_n10027);
nand_5 g09642(new_n10027, new_n796, new_n10028);
nand_5 g09643(new_n10028, new_n458, new_n10029);
nand_5 g09644(new_n10029, new_n453, new_n10030);
nand_5 g09645(new_n10030, new_n447, new_n10031);
nand_5 g09646(new_n10031, new_n805, new_n10032);
nand_5 g09647(new_n10032, new_n811, new_n10033);
nand_5 g09648(new_n10033, new_n442, new_n10034);
nand_5 g09649(new_n10034, new_n437, new_n10035);
nand_5 g09650(new_n10035, new_n819, new_n10036);
nand_5 g09651(new_n10036, new_n432, new_n10037);
nand_5 g09652(new_n10037, new_n427_1, new_n10038);
nand_5 g09653(new_n10038, new_n422, new_n10039);
nand_5 g09654(new_n10039, new_n828, new_n10040);
nand_5 g09655(new_n10040, new_n834, new_n10041);
nand_5 g09656(new_n10041, new_n840, new_n10042);
nand_5 g09657(new_n10042, new_n417, new_n10043);
nand_5 g09658(new_n10043, new_n847, new_n10044);
nand_5 g09659(new_n10044, new_n853, new_n10045);
nand_5 g09660(new_n10045, new_n859, new_n10046);
nand_5 g09661(new_n10046, new_n412, new_n10047);
nand_5 g09662(new_n10047, new_n866, new_n10048);
nand_5 g09663(new_n10048, new_n872, new_n10049);
nand_5 g09664(new_n10049, new_n878, new_n10050_1);
nand_5 g09665(new_n10050_1, new_n407, new_n10051_1);
nand_5 g09666(new_n10051_1, new_n885, new_n10052);
nand_5 g09667(new_n10052, new_n402, new_n10053);
nand_5 g09668(new_n10053, new_n397, new_n10054);
nand_5 g09669(new_n10054, new_n392, new_n10055);
nand_5 g09670(new_n10055, new_n894, new_n10056);
nand_5 g09671(new_n10056, new_n1087, new_n10057);
nand_5 g09672(new_n10057, new_n1129, new_n10058);
nand_5 g09673(new_n10058, new_n1084, new_n10059);
nand_5 g09674(new_n10059, new_n1134, new_n10060);
nand_5 g09675(new_n10060, new_n1080, new_n10061_1);
nand_5 g09676(new_n10061_1, new_n1075, new_n10062);
nand_5 g09677(new_n10062, new_n1070, new_n10063);
nand_5 g09678(new_n10063, new_n1143, new_n10064);
nand_5 g09679(new_n10064, new_n1148, new_n10065);
nand_5 g09680(new_n10065, new_n1065, new_n10066);
nand_5 g09681(new_n10066, new_n1062, new_n10067);
nand_5 g09682(new_n10067, new_n1156, new_n10068);
nand_5 g09683(new_n10068, new_n1057, new_n10069);
nand_5 g09684(new_n10069, new_n1053, new_n10070);
nand_5 g09685(new_n10070, new_n1050, new_n10071);
nand_5 g09686(new_n10071, new_n1045, new_n10072);
nand_5 g09687(new_n10072, new_n1040, new_n10073);
nand_5 g09688(new_n10073, new_n1036, new_n10074);
nand_5 g09689(new_n10074, new_n1033, new_n10075);
nand_5 g09690(new_n10075, new_n1028, new_n10076);
nand_5 g09691(new_n10076, new_n1026, new_n10077);
nand_5 g09692(new_n10077, new_n1021, new_n10078);
nand_5 g09693(new_n10078, new_n1017, new_n10079);
nand_5 g09694(new_n10079, new_n1012, new_n10080_1);
nand_5 g09695(new_n10080_1, new_n1009, new_n10081);
nand_5 g09696(new_n10081, new_n1004, new_n10082);
nand_5 g09697(new_n10082, new_n1000, new_n10083);
nand_5 g09698(new_n10083, new_n995, new_n10084);
nand_5 g09699(new_n10084, new_n990, new_n10085);
nand_5 g09700(new_n10085, new_n985, new_n10086);
nand_5 g09701(new_n10086, new_n981, new_n10087);
nand_5 g09702(new_n10087, new_n1179, new_n10088);
nand_5 g09703(new_n10088, new_n976, new_n10089);
nand_5 g09704(new_n10089, new_n971, new_n10090);
nand_5 g09705(new_n10090, new_n966, new_n10091);
nand_5 g09706(new_n10091, new_n961, new_n10092);
nand_5 g09707(new_n10092, new_n957, new_n10093);
nand_5 g09708(new_n10093, new_n952, new_n10094);
nand_5 g09709(new_n10094, n6436, new_n10095);
nor_5  g09710(new_n10095, new_n945, n11534);
nand_5 g09711(new_n1232, new_n846, new_n10097);
nand_5 g09712(new_n10097, new_n1231, new_n10098);
nand_5 g09713(new_n10098, new_n1227, new_n10099);
nand_5 g09714(new_n10099, new_n1407, new_n10100);
nand_5 g09715(new_n10100, new_n1223, new_n10101);
nand_5 g09716(new_n10101, new_n1218, new_n10102);
nand_5 g09717(new_n10102, new_n1213, new_n10103);
nand_5 g09718(new_n10103, new_n1210, new_n10104);
nand_5 g09719(new_n10104, new_n1206, new_n10105);
nand_5 g09720(new_n10105, new_n1418, new_n10106);
nand_5 g09721(new_n10106, new_n1422, new_n10107);
nand_5 g09722(new_n10107, new_n1428, new_n10108);
nand_5 g09723(new_n10108, new_n1203, new_n10109);
nand_5 g09724(new_n10109, new_n1433, new_n10110);
nand_5 g09725(new_n10110, new_n581, new_n10111);
nand_5 g09726(new_n10111, new_n574, new_n10112_1);
nand_5 g09727(new_n10112_1, new_n568, new_n10113);
nand_5 g09728(new_n10113, new_n589, new_n10114);
nand_5 g09729(new_n10114, new_n595, new_n10115);
nand_5 g09730(new_n10115, new_n601, new_n10116);
nand_5 g09731(new_n10116, new_n563, new_n10117);
nand_5 g09732(new_n10117, new_n608, new_n10118);
nand_5 g09733(new_n10118, new_n558, new_n10119);
nand_5 g09734(new_n10119, new_n615, new_n10120);
nand_5 g09735(new_n10120, new_n553, new_n10121);
nand_5 g09736(new_n10121, new_n622, new_n10122);
nand_5 g09737(new_n10122, new_n628, new_n10123);
nand_5 g09738(new_n10123, new_n548, new_n10124);
nand_5 g09739(new_n10124, new_n543_1, new_n10125);
nand_5 g09740(new_n10125, new_n636, new_n10126);
nand_5 g09741(new_n10126, new_n642, new_n10127);
nand_5 g09742(new_n10127, new_n538, new_n10128);
nand_5 g09743(new_n10128, new_n533, new_n10129);
nand_5 g09744(new_n10129, new_n650_1, new_n10130);
nand_5 g09745(new_n10130, new_n528, new_n10131);
nand_5 g09746(new_n10131, new_n523, new_n10132);
nand_5 g09747(new_n10132, new_n518, new_n10133);
nand_5 g09748(new_n10133, new_n659, new_n10134);
nand_5 g09749(new_n10134, new_n665, new_n10135);
nand_5 g09750(new_n10135, new_n672, new_n10136);
nand_5 g09751(new_n10136, new_n513, new_n10137);
nand_5 g09752(new_n10137, new_n679, new_n10138);
nand_5 g09753(new_n10138, new_n685, new_n10139);
nand_5 g09754(new_n10139, new_n691, new_n10140);
nand_5 g09755(new_n10140, new_n508, new_n10141);
nand_5 g09756(new_n10141, new_n698, new_n10142);
nand_5 g09757(new_n10142, new_n503, new_n10143);
nand_5 g09758(new_n10143, new_n704, new_n10144);
nand_5 g09759(new_n10144, new_n498_1, new_n10145);
nand_5 g09760(new_n10145, new_n711, new_n10146);
nand_5 g09761(new_n10146, new_n493, new_n10147_1);
nand_5 g09762(new_n10147_1, new_n718, new_n10148);
nand_5 g09763(new_n10148, new_n488, new_n10149);
nand_5 g09764(new_n10149, new_n725, new_n10150);
nand_5 g09765(new_n10150, new_n483, new_n10151);
nand_5 g09766(new_n10151, new_n732, new_n10152);
nand_5 g09767(new_n10152, new_n478, new_n10153);
nand_5 g09768(new_n10153, new_n739, new_n10154);
nand_5 g09769(new_n10154, new_n745, new_n10155);
nand_5 g09770(new_n10155, new_n751, new_n10156);
nand_5 g09771(new_n10156, new_n473, new_n10157);
nand_5 g09772(new_n10157, new_n758, new_n10158);
nand_5 g09773(new_n10158, new_n764, new_n10159);
nand_5 g09774(new_n10159, new_n770, new_n10160);
nand_5 g09775(new_n10160, new_n468, new_n10161);
nand_5 g09776(new_n10161, new_n777, new_n10162);
nand_5 g09777(new_n10162, new_n783, new_n10163);
nand_5 g09778(new_n10163, new_n789, new_n10164);
nand_5 g09779(new_n10164, new_n463, new_n10165);
nand_5 g09780(new_n10165, new_n796, new_n10166);
nand_5 g09781(new_n10166, new_n458, new_n10167);
nand_5 g09782(new_n10167, new_n453, new_n10168);
nand_5 g09783(new_n10168, new_n447, new_n10169);
nand_5 g09784(new_n10169, new_n805, new_n10170);
nand_5 g09785(new_n10170, new_n811, new_n10171);
nand_5 g09786(new_n10171, new_n442, new_n10172);
nand_5 g09787(new_n10172, new_n437, new_n10173);
nand_5 g09788(new_n10173, new_n819, new_n10174);
nand_5 g09789(new_n10174, new_n432, new_n10175);
nand_5 g09790(new_n10175, new_n427_1, new_n10176);
nand_5 g09791(new_n10176, new_n422, new_n10177);
nand_5 g09792(new_n10177, new_n828, new_n10178);
nand_5 g09793(new_n10178, new_n834, new_n10179);
nand_5 g09794(new_n10179, new_n840, new_n10180);
nand_5 g09795(new_n10180, n9186, new_n10181);
nor_5  g09796(new_n10181, new_n414, n11627);
not_4  g09797(new_n501, new_n10183);
nand_5 g09798(new_n1568_1, new_n703, new_n10184);
nand_5 g09799(new_n10184, new_n1567, new_n10185);
nand_5 g09800(new_n10185, new_n1564, new_n10186);
nand_5 g09801(new_n10186, new_n1561, new_n10187);
nand_5 g09802(new_n10187, new_n1338, new_n10188);
nand_5 g09803(new_n10188, new_n1331, new_n10189);
nand_5 g09804(new_n10189, new_n1326, new_n10190);
nand_5 g09805(new_n10190, new_n1321, new_n10191);
nand_5 g09806(new_n10191, new_n1318, new_n10192);
nand_5 g09807(new_n10192, new_n1315, new_n10193);
nand_5 g09808(new_n10193, new_n1312, new_n10194);
nand_5 g09809(new_n10194, new_n1309, new_n10195);
nand_5 g09810(new_n10195, new_n1307, new_n10196);
nand_5 g09811(new_n10196, new_n1304, new_n10197);
nand_5 g09812(new_n10197, new_n1300, new_n10198);
nand_5 g09813(new_n10198, new_n1297, new_n10199);
nand_5 g09814(new_n10199, new_n1294, new_n10200);
nand_5 g09815(new_n10200, new_n1355, new_n10201);
nand_5 g09816(new_n10201, new_n1291, new_n10202);
nand_5 g09817(new_n10202, new_n1288, new_n10203);
nand_5 g09818(new_n10203, new_n1283, new_n10204);
nand_5 g09819(new_n10204, new_n1363, new_n10205);
nand_5 g09820(new_n10205, new_n1280, new_n10206);
nand_5 g09821(new_n10206, new_n1370, new_n10207);
nand_5 g09822(new_n10207, new_n1373, new_n10208);
nand_5 g09823(new_n10208, new_n1277, new_n10209);
nand_5 g09824(new_n10209, new_n1272, new_n10210);
nand_5 g09825(new_n10210, new_n1269, new_n10211);
nand_5 g09826(new_n10211, new_n1380, new_n10212);
nand_5 g09827(new_n10212, new_n1264, new_n10213);
nand_5 g09828(new_n10213, new_n1259, new_n10214);
nand_5 g09829(new_n10214, new_n1388, new_n10215);
nand_5 g09830(new_n10215, new_n1392, new_n10216);
nand_5 g09831(new_n10216, new_n1256, new_n10217);
nand_5 g09832(new_n10217, new_n1252, new_n10218);
nand_5 g09833(new_n10218, new_n1249, new_n10219);
nand_5 g09834(new_n10219, new_n1244, new_n10220);
nand_5 g09835(new_n10220, new_n1240, new_n10221);
nand_5 g09836(new_n10221, new_n1234, new_n10222);
nand_5 g09837(new_n10222, new_n1231, new_n10223);
nand_5 g09838(new_n10223, new_n1227, new_n10224);
nand_5 g09839(new_n10224, new_n1407, new_n10225);
nand_5 g09840(new_n10225, new_n1223, new_n10226);
nand_5 g09841(new_n10226, new_n1218, new_n10227);
nand_5 g09842(new_n10227, new_n1213, new_n10228);
nand_5 g09843(new_n10228, new_n1210, new_n10229);
nand_5 g09844(new_n10229, new_n1206, new_n10230);
nand_5 g09845(new_n10230, new_n1418, new_n10231);
nand_5 g09846(new_n10231, new_n1422, new_n10232);
nand_5 g09847(new_n10232, new_n1428, new_n10233);
nand_5 g09848(new_n10233, new_n1203, new_n10234);
nand_5 g09849(new_n10234, new_n1433, new_n10235);
nand_5 g09850(new_n10235, new_n581, new_n10236);
nand_5 g09851(new_n10236, new_n574, new_n10237);
nand_5 g09852(new_n10237, new_n568, new_n10238);
nand_5 g09853(new_n10238, new_n589, new_n10239);
nand_5 g09854(new_n10239, new_n595, new_n10240);
nand_5 g09855(new_n10240, new_n601, new_n10241);
nand_5 g09856(new_n10241, new_n563, new_n10242);
nand_5 g09857(new_n10242, new_n608, new_n10243);
nand_5 g09858(new_n10243, new_n558, new_n10244);
nand_5 g09859(new_n10244, new_n615, new_n10245);
nand_5 g09860(new_n10245, new_n553, new_n10246);
nand_5 g09861(new_n10246, new_n622, new_n10247);
nand_5 g09862(new_n10247, new_n628, new_n10248);
nand_5 g09863(new_n10248, new_n548, new_n10249);
nand_5 g09864(new_n10249, new_n543_1, new_n10250);
nand_5 g09865(new_n10250, new_n636, new_n10251);
nand_5 g09866(new_n10251, new_n642, new_n10252);
nand_5 g09867(new_n10252, new_n538, new_n10253);
nand_5 g09868(new_n10253, new_n533, new_n10254);
nand_5 g09869(new_n10254, new_n650_1, new_n10255_1);
nand_5 g09870(new_n10255_1, new_n528, new_n10256);
nand_5 g09871(new_n10256, new_n523, new_n10257);
nand_5 g09872(new_n10257, new_n518, new_n10258);
nand_5 g09873(new_n10258, new_n659, new_n10259);
nand_5 g09874(new_n10259, new_n665, new_n10260);
nand_5 g09875(new_n10260, new_n672, new_n10261);
nand_5 g09876(new_n10261, new_n513, new_n10262);
nand_5 g09877(new_n10262, new_n679, new_n10263);
nand_5 g09878(new_n10263, new_n685, new_n10264);
nand_5 g09879(new_n10264, new_n691, new_n10265);
nand_5 g09880(new_n10265, new_n508, new_n10266);
nand_5 g09881(new_n10266, new_n698, new_n10267);
nand_5 g09882(new_n10267, n13814, new_n10268);
nor_5  g09883(new_n10268, new_n10183, n11664);
not_4  g09884(new_n1787, new_n10270);
nand_5 g09885(new_n1607, new_n1024, new_n10271);
nand_5 g09886(new_n10271, new_n1021, new_n10272);
nand_5 g09887(new_n10272, new_n1017, new_n10273);
nand_5 g09888(new_n10273, new_n1012, new_n10274);
nand_5 g09889(new_n10274, new_n1009, new_n10275);
nand_5 g09890(new_n10275, new_n1004, new_n10276);
nand_5 g09891(new_n10276, new_n1000, new_n10277);
nand_5 g09892(new_n10277, new_n995, new_n10278_1);
nand_5 g09893(new_n10278_1, new_n990, new_n10279);
nand_5 g09894(new_n10279, new_n985, new_n10280);
nand_5 g09895(new_n10280, new_n981, new_n10281);
nand_5 g09896(new_n10281, new_n1179, new_n10282);
nand_5 g09897(new_n10282, new_n976, new_n10283_1);
nand_5 g09898(new_n10283_1, new_n971, new_n10284);
nand_5 g09899(new_n10284, new_n966, new_n10285);
nand_5 g09900(new_n10285, new_n961, new_n10286);
nand_5 g09901(new_n10286, new_n957, new_n10287);
nand_5 g09902(new_n10287, new_n952, new_n10288);
nand_5 g09903(new_n10288, new_n948_1, new_n10289);
nand_5 g09904(new_n10289, new_n943, new_n10290);
nand_5 g09905(new_n10290, new_n941, new_n10291);
nand_5 g09906(new_n10291, new_n938, new_n10292);
nand_5 g09907(new_n10292, new_n936, new_n10293);
nand_5 g09908(new_n10293, new_n931, new_n10294);
nand_5 g09909(new_n10294, new_n927, new_n10295);
nand_5 g09910(new_n10295, new_n922, new_n10296);
nand_5 g09911(new_n10296, new_n917, new_n10297);
nand_5 g09912(new_n10297, new_n912, new_n10298);
nand_5 g09913(new_n10298, new_n907, new_n10299);
nand_5 g09914(new_n10299, new_n903, new_n10300);
nand_5 g09915(new_n10300, new_n2066, new_n10301);
nand_5 g09916(new_n10301, new_n2063, new_n10302);
nand_5 g09917(new_n10302, new_n2062, new_n10303);
nand_5 g09918(new_n10303, new_n2058, new_n10304);
nand_5 g09919(new_n10304, new_n2055, new_n10305);
nand_5 g09920(new_n10305, new_n2051, new_n10306);
nand_5 g09921(new_n10306, new_n2046, new_n10307);
nand_5 g09922(new_n10307, new_n2042, new_n10308);
nand_5 g09923(new_n10308, new_n2039, new_n10309);
nand_5 g09924(new_n10309, new_n2036, new_n10310);
nand_5 g09925(new_n10310, new_n2033, new_n10311);
nand_5 g09926(new_n10311, new_n2029, new_n10312);
nand_5 g09927(new_n10312, new_n2026, new_n10313);
nand_5 g09928(new_n10313, new_n2022, new_n10314);
nand_5 g09929(new_n10314, new_n2018, new_n10315);
nand_5 g09930(new_n10315, new_n1726, new_n10316);
nand_5 g09931(new_n10316, new_n1722, new_n10317);
nand_5 g09932(new_n10317, new_n1718, new_n10318);
nand_5 g09933(new_n10318, new_n1713, new_n10319);
nand_5 g09934(new_n10319, new_n1737, new_n10320);
nand_5 g09935(new_n10320, new_n1709, new_n10321);
nand_5 g09936(new_n10321, new_n1742, new_n10322);
nand_5 g09937(new_n10322, new_n1704, new_n10323);
nand_5 g09938(new_n10323, new_n1702_1, new_n10324);
nand_5 g09939(new_n10324, new_n1698, new_n10325);
nand_5 g09940(new_n10325, new_n1695, new_n10326);
nand_5 g09941(new_n10326, new_n1692, new_n10327);
nand_5 g09942(new_n10327, new_n1752, new_n10328);
nand_5 g09943(new_n10328, new_n1688, new_n10329);
nand_5 g09944(new_n10329, new_n1685, new_n10330);
nand_5 g09945(new_n10330, new_n1680, new_n10331);
nand_5 g09946(new_n10331, new_n1676, new_n10332);
nand_5 g09947(new_n10332, new_n1672, new_n10333);
nand_5 g09948(new_n10333, new_n1669, new_n10334);
nand_5 g09949(new_n10334, new_n1666, new_n10335);
nand_5 g09950(new_n10335, new_n1663, new_n10336);
nand_5 g09951(new_n10336, new_n1658, new_n10337);
nand_5 g09952(new_n10337, new_n1653, new_n10338);
nand_5 g09953(new_n10338, new_n1651, new_n10339);
nand_5 g09954(new_n10339, new_n1649, new_n10340);
nand_5 g09955(new_n10340, new_n1646, new_n10341);
nand_5 g09956(new_n10341, new_n1643, new_n10342);
nand_5 g09957(new_n10342, new_n1641, new_n10343);
nand_5 g09958(new_n10343, new_n1638, new_n10344);
nand_5 g09959(new_n10344, new_n1635, new_n10345);
nand_5 g09960(new_n10345, new_n1632, new_n10346);
nand_5 g09961(new_n10346, new_n1628, new_n10347);
nand_5 g09962(new_n10347, new_n1625, new_n10348);
nand_5 g09963(new_n10348, new_n1621, new_n10349);
nand_5 g09964(new_n10349, new_n1618, new_n10350);
nand_5 g09965(new_n10350, new_n1778, new_n10351);
nand_5 g09966(new_n10351, new_n1782, new_n10352);
nand_5 g09967(new_n10352, new_n1614, new_n10353);
nand_5 g09968(new_n10353, new_n1611, new_n10354);
nand_5 g09969(new_n10354, n8746, new_n10355);
nor_5  g09970(new_n10355, new_n10270, n11822);
not_4  g09971(new_n696, new_n10357);
nand_5 g09972(new_n1576, new_n10357, new_n10358);
nand_5 g09973(new_n10358, new_n1573, new_n10359);
nand_5 g09974(new_n10359, new_n1570, new_n10360);
nand_5 g09975(new_n10360, new_n1567, new_n10361);
nand_5 g09976(new_n10361, new_n1564, new_n10362);
nand_5 g09977(new_n10362, new_n1561, new_n10363);
nand_5 g09978(new_n10363, new_n1338, new_n10364);
nand_5 g09979(new_n10364, new_n1331, new_n10365);
nand_5 g09980(new_n10365, new_n1326, new_n10366);
nand_5 g09981(new_n10366, new_n1321, new_n10367);
nand_5 g09982(new_n10367, new_n1318, new_n10368);
nand_5 g09983(new_n10368, new_n1315, new_n10369);
nand_5 g09984(new_n10369, new_n1312, new_n10370);
nand_5 g09985(new_n10370, new_n1309, new_n10371);
nand_5 g09986(new_n10371, new_n1307, new_n10372);
nand_5 g09987(new_n10372, new_n1304, new_n10373);
nand_5 g09988(new_n10373, new_n1300, new_n10374);
nand_5 g09989(new_n10374, new_n1297, new_n10375);
nand_5 g09990(new_n10375, new_n1294, new_n10376);
nand_5 g09991(new_n10376, new_n1355, new_n10377);
nand_5 g09992(new_n10377, new_n1291, new_n10378_1);
nand_5 g09993(new_n10378_1, new_n1288, new_n10379);
nand_5 g09994(new_n10379, new_n1283, new_n10380);
nand_5 g09995(new_n10380, new_n1363, new_n10381);
nand_5 g09996(new_n10381, new_n1280, new_n10382);
nand_5 g09997(new_n10382, new_n1370, new_n10383);
nand_5 g09998(new_n10383, new_n1373, new_n10384);
nand_5 g09999(new_n10384, new_n1277, new_n10385);
nand_5 g10000(new_n10385, new_n1272, new_n10386);
nand_5 g10001(new_n10386, new_n1269, new_n10387);
nand_5 g10002(new_n10387, new_n1380, new_n10388);
nand_5 g10003(new_n10388, new_n1264, new_n10389);
nand_5 g10004(new_n10389, new_n1259, new_n10390);
nand_5 g10005(new_n10390, new_n1388, new_n10391);
nand_5 g10006(new_n10391, new_n1392, new_n10392);
nand_5 g10007(new_n10392, new_n1256, new_n10393);
nand_5 g10008(new_n10393, new_n1252, new_n10394);
nand_5 g10009(new_n10394, new_n1249, new_n10395);
nand_5 g10010(new_n10395, new_n1244, new_n10396);
nand_5 g10011(new_n10396, new_n1240, new_n10397);
nand_5 g10012(new_n10397, new_n1234, new_n10398);
nand_5 g10013(new_n10398, new_n1231, new_n10399);
nand_5 g10014(new_n10399, new_n1227, new_n10400);
nand_5 g10015(new_n10400, new_n1407, new_n10401);
nand_5 g10016(new_n10401, new_n1223, new_n10402);
nand_5 g10017(new_n10402, new_n1218, new_n10403);
nand_5 g10018(new_n10403, new_n1213, new_n10404);
nand_5 g10019(new_n10404, new_n1210, new_n10405);
nand_5 g10020(new_n10405, new_n1206, new_n10406);
nand_5 g10021(new_n10406, new_n1418, new_n10407_1);
nand_5 g10022(new_n10407_1, new_n1422, new_n10408);
nand_5 g10023(new_n10408, new_n1428, new_n10409);
nand_5 g10024(new_n10409, new_n1203, new_n10410);
nand_5 g10025(new_n10410, new_n1433, new_n10411);
nand_5 g10026(new_n10411, new_n581, new_n10412);
nand_5 g10027(new_n10412, new_n574, new_n10413);
nand_5 g10028(new_n10413, new_n568, new_n10414);
nand_5 g10029(new_n10414, new_n589, new_n10415);
nand_5 g10030(new_n10415, new_n595, new_n10416);
nand_5 g10031(new_n10416, new_n601, new_n10417);
nand_5 g10032(new_n10417, new_n563, new_n10418);
nand_5 g10033(new_n10418, new_n608, new_n10419);
nand_5 g10034(new_n10419, new_n558, new_n10420);
nand_5 g10035(new_n10420, new_n615, new_n10421);
nand_5 g10036(new_n10421, new_n553, new_n10422);
nand_5 g10037(new_n10422, new_n622, new_n10423);
nand_5 g10038(new_n10423, new_n628, new_n10424);
nand_5 g10039(new_n10424, new_n548, new_n10425);
nand_5 g10040(new_n10425, new_n543_1, new_n10426_1);
nand_5 g10041(new_n10426_1, new_n636, new_n10427);
nand_5 g10042(new_n10427, new_n642, new_n10428);
nand_5 g10043(new_n10428, new_n538, new_n10429);
nand_5 g10044(new_n10429, new_n533, new_n10430);
nand_5 g10045(new_n10430, new_n650_1, new_n10431);
nand_5 g10046(new_n10431, new_n528, new_n10432);
nand_5 g10047(new_n10432, new_n523, new_n10433);
nand_5 g10048(new_n10433, new_n518, new_n10434);
nand_5 g10049(new_n10434, new_n659, new_n10435);
nand_5 g10050(new_n10435, new_n665, new_n10436);
nand_5 g10051(new_n10436, new_n672, new_n10437);
nand_5 g10052(new_n10437, new_n513, new_n10438);
nand_5 g10053(new_n10438, new_n679, new_n10439);
nand_5 g10054(new_n10439, new_n685, new_n10440);
nand_5 g10055(new_n10440, new_n691, new_n10441);
nand_5 g10056(new_n10441, n203, new_n10442);
nor_5  g10057(new_n10442, new_n505, n11847);
nand_5 g10058(new_n1603, new_n649, new_n10444);
nand_5 g10059(new_n10444, new_n1795, new_n10445);
nand_5 g10060(new_n10445, new_n1799, new_n10446_1);
nand_5 g10061(new_n10446_1, new_n1602, new_n10447);
nand_5 g10062(new_n10447, new_n1599, new_n10448);
nand_5 g10063(new_n10448, new_n1596, new_n10449);
nand_5 g10064(new_n10449, new_n1593, new_n10450);
nand_5 g10065(new_n10450, new_n1806, new_n10451);
nand_5 g10066(new_n10451, new_n1589, new_n10452);
nand_5 g10067(new_n10452, new_n1586, new_n10453);
nand_5 g10068(new_n10453, new_n1583, new_n10454);
nand_5 g10069(new_n10454, new_n1580, new_n10455);
nand_5 g10070(new_n10455, new_n1576, new_n10456);
nand_5 g10071(new_n10456, new_n1573, new_n10457);
nand_5 g10072(new_n10457, new_n1570, new_n10458);
nand_5 g10073(new_n10458, new_n1567, new_n10459);
nand_5 g10074(new_n10459, new_n1564, new_n10460);
nand_5 g10075(new_n10460, new_n1561, new_n10461);
nand_5 g10076(new_n10461, new_n1338, new_n10462);
nand_5 g10077(new_n10462, new_n1331, new_n10463);
nand_5 g10078(new_n10463, new_n1326, new_n10464);
nand_5 g10079(new_n10464, new_n1321, new_n10465);
nand_5 g10080(new_n10465, new_n1318, new_n10466_1);
nand_5 g10081(new_n10466_1, new_n1315, new_n10467);
nand_5 g10082(new_n10467, new_n1312, new_n10468);
nand_5 g10083(new_n10468, new_n1309, new_n10469);
nand_5 g10084(new_n10469, new_n1307, new_n10470_1);
nand_5 g10085(new_n10470_1, new_n1304, new_n10471);
nand_5 g10086(new_n10471, new_n1300, new_n10472);
nand_5 g10087(new_n10472, new_n1297, new_n10473);
nand_5 g10088(new_n10473, new_n1294, new_n10474);
nand_5 g10089(new_n10474, new_n1355, new_n10475);
nand_5 g10090(new_n10475, new_n1291, new_n10476);
nand_5 g10091(new_n10476, new_n1288, new_n10477);
nand_5 g10092(new_n10477, new_n1283, new_n10478);
nand_5 g10093(new_n10478, new_n1363, new_n10479);
nand_5 g10094(new_n10479, new_n1280, new_n10480);
nand_5 g10095(new_n10480, new_n1370, new_n10481);
nand_5 g10096(new_n10481, new_n1373, new_n10482);
nand_5 g10097(new_n10482, new_n1277, new_n10483);
nand_5 g10098(new_n10483, new_n1272, new_n10484);
nand_5 g10099(new_n10484, new_n1269, new_n10485);
nand_5 g10100(new_n10485, new_n1380, new_n10486);
nand_5 g10101(new_n10486, new_n1264, new_n10487);
nand_5 g10102(new_n10487, new_n1259, new_n10488);
nand_5 g10103(new_n10488, new_n1388, new_n10489);
nand_5 g10104(new_n10489, new_n1392, new_n10490);
nand_5 g10105(new_n10490, new_n1256, new_n10491);
nand_5 g10106(new_n10491, new_n1252, new_n10492);
nand_5 g10107(new_n10492, new_n1249, new_n10493);
nand_5 g10108(new_n10493, new_n1244, new_n10494);
nand_5 g10109(new_n10494, new_n1240, new_n10495);
nand_5 g10110(new_n10495, new_n1234, new_n10496);
nand_5 g10111(new_n10496, new_n1231, new_n10497);
nand_5 g10112(new_n10497, new_n1227, new_n10498);
nand_5 g10113(new_n10498, new_n1407, new_n10499);
nand_5 g10114(new_n10499, new_n1223, new_n10500);
nand_5 g10115(new_n10500, new_n1218, new_n10501);
nand_5 g10116(new_n10501, new_n1213, new_n10502);
nand_5 g10117(new_n10502, new_n1210, new_n10503);
nand_5 g10118(new_n10503, new_n1206, new_n10504);
nand_5 g10119(new_n10504, new_n1418, new_n10505);
nand_5 g10120(new_n10505, new_n1422, new_n10506);
nand_5 g10121(new_n10506, new_n1428, new_n10507);
nand_5 g10122(new_n10507, new_n1203, new_n10508);
nand_5 g10123(new_n10508, new_n1433, new_n10509);
nand_5 g10124(new_n10509, new_n581, new_n10510);
nand_5 g10125(new_n10510, new_n574, new_n10511);
nand_5 g10126(new_n10511, new_n568, new_n10512);
nand_5 g10127(new_n10512, new_n589, new_n10513);
nand_5 g10128(new_n10513, new_n595, new_n10514);
nand_5 g10129(new_n10514, new_n601, new_n10515_1);
nand_5 g10130(new_n10515_1, new_n563, new_n10516);
nand_5 g10131(new_n10516, new_n608, new_n10517);
nand_5 g10132(new_n10517, new_n558, new_n10518);
nand_5 g10133(new_n10518, new_n615, new_n10519);
nand_5 g10134(new_n10519, new_n553, new_n10520);
nand_5 g10135(new_n10520, new_n622, new_n10521);
nand_5 g10136(new_n10521, new_n628, new_n10522);
nand_5 g10137(new_n10522, new_n548, new_n10523);
nand_5 g10138(new_n10523, new_n543_1, new_n10524);
nand_5 g10139(new_n10524, new_n636, new_n10525);
nand_5 g10140(new_n10525, new_n642, new_n10526);
nand_5 g10141(new_n10526, new_n538, new_n10527);
nand_5 g10142(new_n10527, n8550, new_n10528);
nor_5  g10143(new_n10528, new_n530, n12032);
nand_5 g10144(new_n1639, new_n600, new_n10530);
nand_5 g10145(new_n10530, new_n1638, new_n10531);
nand_5 g10146(new_n10531, new_n1635, new_n10532);
nand_5 g10147(new_n10532, new_n1632, new_n10533);
nand_5 g10148(new_n10533, new_n1628, new_n10534);
nand_5 g10149(new_n10534, new_n1625, new_n10535);
nand_5 g10150(new_n10535, new_n1621, new_n10536);
nand_5 g10151(new_n10536, new_n1618, new_n10537);
nand_5 g10152(new_n10537, new_n1778, new_n10538);
nand_5 g10153(new_n10538, new_n1782, new_n10539);
nand_5 g10154(new_n10539, new_n1614, new_n10540);
nand_5 g10155(new_n10540, new_n1611, new_n10541);
nand_5 g10156(new_n10541, new_n1789, new_n10542);
nand_5 g10157(new_n10542, new_n1608, new_n10543);
nand_5 g10158(new_n10543, new_n1605, new_n10544);
nand_5 g10159(new_n10544, new_n1795, new_n10545);
nand_5 g10160(new_n10545, new_n1799, new_n10546);
nand_5 g10161(new_n10546, new_n1602, new_n10547);
nand_5 g10162(new_n10547, new_n1599, new_n10548);
nand_5 g10163(new_n10548, new_n1596, new_n10549);
nand_5 g10164(new_n10549, new_n1593, new_n10550);
nand_5 g10165(new_n10550, new_n1806, new_n10551);
nand_5 g10166(new_n10551, new_n1589, new_n10552);
nand_5 g10167(new_n10552, new_n1586, new_n10553);
nand_5 g10168(new_n10553, new_n1583, new_n10554);
nand_5 g10169(new_n10554, new_n1580, new_n10555);
nand_5 g10170(new_n10555, new_n1576, new_n10556);
nand_5 g10171(new_n10556, new_n1573, new_n10557);
nand_5 g10172(new_n10557, new_n1570, new_n10558);
nand_5 g10173(new_n10558, new_n1567, new_n10559);
nand_5 g10174(new_n10559, new_n1564, new_n10560);
nand_5 g10175(new_n10560, new_n1561, new_n10561);
nand_5 g10176(new_n10561, new_n1338, new_n10562);
nand_5 g10177(new_n10562, new_n1331, new_n10563);
nand_5 g10178(new_n10563, new_n1326, new_n10564);
nand_5 g10179(new_n10564, new_n1321, new_n10565);
nand_5 g10180(new_n10565, new_n1318, new_n10566);
nand_5 g10181(new_n10566, new_n1315, new_n10567);
nand_5 g10182(new_n10567, new_n1312, new_n10568);
nand_5 g10183(new_n10568, new_n1309, new_n10569);
nand_5 g10184(new_n10569, new_n1307, new_n10570);
nand_5 g10185(new_n10570, new_n1304, new_n10571);
nand_5 g10186(new_n10571, new_n1300, new_n10572);
nand_5 g10187(new_n10572, new_n1297, new_n10573_1);
nand_5 g10188(new_n10573_1, new_n1294, new_n10574);
nand_5 g10189(new_n10574, new_n1355, new_n10575);
nand_5 g10190(new_n10575, new_n1291, new_n10576);
nand_5 g10191(new_n10576, new_n1288, new_n10577);
nand_5 g10192(new_n10577, new_n1283, new_n10578);
nand_5 g10193(new_n10578, new_n1363, new_n10579);
nand_5 g10194(new_n10579, new_n1280, new_n10580);
nand_5 g10195(new_n10580, new_n1370, new_n10581);
nand_5 g10196(new_n10581, new_n1373, new_n10582);
nand_5 g10197(new_n10582, new_n1277, new_n10583);
nand_5 g10198(new_n10583, new_n1272, new_n10584);
nand_5 g10199(new_n10584, new_n1269, new_n10585);
nand_5 g10200(new_n10585, new_n1380, new_n10586);
nand_5 g10201(new_n10586, new_n1264, new_n10587);
nand_5 g10202(new_n10587, new_n1259, new_n10588);
nand_5 g10203(new_n10588, new_n1388, new_n10589);
nand_5 g10204(new_n10589, new_n1392, new_n10590);
nand_5 g10205(new_n10590, new_n1256, new_n10591_1);
nand_5 g10206(new_n10591_1, new_n1252, new_n10592);
nand_5 g10207(new_n10592, new_n1249, new_n10593);
nand_5 g10208(new_n10593, new_n1244, new_n10594);
nand_5 g10209(new_n10594, new_n1240, new_n10595);
nand_5 g10210(new_n10595, new_n1234, new_n10596);
nand_5 g10211(new_n10596, new_n1231, new_n10597);
nand_5 g10212(new_n10597, new_n1227, new_n10598);
nand_5 g10213(new_n10598, new_n1407, new_n10599);
nand_5 g10214(new_n10599, new_n1223, new_n10600);
nand_5 g10215(new_n10600, new_n1218, new_n10601);
nand_5 g10216(new_n10601, new_n1213, new_n10602);
nand_5 g10217(new_n10602, new_n1210, new_n10603);
nand_5 g10218(new_n10603, new_n1206, new_n10604);
nand_5 g10219(new_n10604, new_n1418, new_n10605);
nand_5 g10220(new_n10605, new_n1422, new_n10606);
nand_5 g10221(new_n10606, new_n1428, new_n10607);
nand_5 g10222(new_n10607, new_n1203, new_n10608);
nand_5 g10223(new_n10608, new_n1433, new_n10609);
nand_5 g10224(new_n10609, new_n581, new_n10610);
nand_5 g10225(new_n10610, new_n574, new_n10611);
nand_5 g10226(new_n10611, new_n568, new_n10612);
nand_5 g10227(new_n10612, new_n589, new_n10613);
nand_5 g10228(new_n10613, n7354, new_n10614);
nor_5  g10229(new_n10614, new_n592, n12166);
nand_5 g10230(new_n1072, new_n1070, new_n10616);
nand_5 g10231(new_n10616, new_n1143, new_n10617);
nand_5 g10232(new_n10617, new_n1148, new_n10618);
nand_5 g10233(new_n10618, new_n1065, new_n10619);
nand_5 g10234(new_n10619, new_n1062, new_n10620);
nand_5 g10235(new_n10620, new_n1156, new_n10621);
nand_5 g10236(new_n10621, new_n1057, new_n10622);
nand_5 g10237(new_n10622, new_n1053, new_n10623);
nand_5 g10238(new_n10623, new_n1050, new_n10624);
nand_5 g10239(new_n10624, new_n1045, new_n10625);
nand_5 g10240(new_n10625, new_n1040, new_n10626);
nand_5 g10241(new_n10626, new_n1036, new_n10627);
nand_5 g10242(new_n10627, new_n1033, new_n10628);
nand_5 g10243(new_n10628, new_n1028, new_n10629);
nand_5 g10244(new_n10629, new_n1026, new_n10630_1);
nand_5 g10245(new_n10630_1, new_n1021, new_n10631);
nand_5 g10246(new_n10631, new_n1017, new_n10632);
nand_5 g10247(new_n10632, new_n1012, new_n10633);
nand_5 g10248(new_n10633, new_n1009, new_n10634);
nand_5 g10249(new_n10634, new_n1004, new_n10635);
nand_5 g10250(new_n10635, new_n1000, new_n10636);
nand_5 g10251(new_n10636, new_n995, new_n10637);
nand_5 g10252(new_n10637, new_n990, new_n10638);
nand_5 g10253(new_n10638, new_n985, new_n10639);
nand_5 g10254(new_n10639, new_n981, new_n10640);
nand_5 g10255(new_n10640, new_n1179, new_n10641);
nand_5 g10256(new_n10641, new_n976, new_n10642);
nand_5 g10257(new_n10642, new_n971, new_n10643);
nand_5 g10258(new_n10643, new_n966, new_n10644);
nand_5 g10259(new_n10644, new_n961, new_n10645);
nand_5 g10260(new_n10645, new_n957, new_n10646);
nand_5 g10261(new_n10646, new_n952, new_n10647);
nand_5 g10262(new_n10647, new_n948_1, new_n10648);
nand_5 g10263(new_n10648, new_n943, new_n10649);
nand_5 g10264(new_n10649, new_n941, new_n10650);
nand_5 g10265(new_n10650, new_n938, new_n10651);
nand_5 g10266(new_n10651, new_n936, new_n10652);
nand_5 g10267(new_n10652, new_n931, new_n10653);
nand_5 g10268(new_n10653, new_n927, new_n10654);
nand_5 g10269(new_n10654, new_n922, new_n10655);
nand_5 g10270(new_n10655, new_n917, new_n10656);
nand_5 g10271(new_n10656, new_n912, new_n10657);
nand_5 g10272(new_n10657, new_n907, new_n10658);
nand_5 g10273(new_n10658, new_n903, new_n10659);
nand_5 g10274(new_n10659, new_n2066, new_n10660);
nand_5 g10275(new_n10660, new_n2063, new_n10661);
nand_5 g10276(new_n10661, new_n2062, new_n10662);
nand_5 g10277(new_n10662, new_n2058, new_n10663);
nand_5 g10278(new_n10663, new_n2055, new_n10664);
nand_5 g10279(new_n10664, new_n2051, new_n10665);
nand_5 g10280(new_n10665, new_n2046, new_n10666);
nand_5 g10281(new_n10666, new_n2042, new_n10667);
nand_5 g10282(new_n10667, new_n2039, new_n10668);
nand_5 g10283(new_n10668, new_n2036, new_n10669);
nand_5 g10284(new_n10669, new_n2033, new_n10670);
nand_5 g10285(new_n10670, new_n2029, new_n10671);
nand_5 g10286(new_n10671, new_n2026, new_n10672);
nand_5 g10287(new_n10672, new_n2022, new_n10673);
nand_5 g10288(new_n10673, new_n2018, new_n10674);
nand_5 g10289(new_n10674, new_n1726, new_n10675);
nand_5 g10290(new_n10675, new_n1722, new_n10676);
nand_5 g10291(new_n10676, new_n1718, new_n10677);
nand_5 g10292(new_n10677, new_n1713, new_n10678);
nand_5 g10293(new_n10678, new_n1737, new_n10679);
nand_5 g10294(new_n10679, new_n1709, new_n10680);
nand_5 g10295(new_n10680, new_n1742, new_n10681);
nand_5 g10296(new_n10681, new_n1704, new_n10682);
nand_5 g10297(new_n10682, new_n1702_1, new_n10683);
nand_5 g10298(new_n10683, new_n1698, new_n10684);
nand_5 g10299(new_n10684, new_n1695, new_n10685);
nand_5 g10300(new_n10685, new_n1692, new_n10686);
nand_5 g10301(new_n10686, new_n1752, new_n10687);
nand_5 g10302(new_n10687, new_n1688, new_n10688);
nand_5 g10303(new_n10688, new_n1685, new_n10689);
nand_5 g10304(new_n10689, new_n1680, new_n10690);
nand_5 g10305(new_n10690, new_n1676, new_n10691);
nand_5 g10306(new_n10691, new_n1672, new_n10692);
nand_5 g10307(new_n10692, new_n1669, new_n10693);
nand_5 g10308(new_n10693, new_n1666, new_n10694);
nand_5 g10309(new_n10694, new_n1663, new_n10695);
nand_5 g10310(new_n10695, new_n1658, new_n10696);
nand_5 g10311(new_n10696, new_n1653, new_n10697);
nand_5 g10312(new_n10697, new_n1651, new_n10698);
nand_5 g10313(new_n10698, new_n1649, new_n10699);
nand_5 g10314(new_n10699, n13102, new_n10700);
nor_5  g10315(new_n10700, new_n586, n12232);
nand_5 g10316(new_n1250, new_n827, new_n10702);
nand_5 g10317(new_n10702, new_n1249, new_n10703);
nand_5 g10318(new_n10703, new_n1244, new_n10704);
nand_5 g10319(new_n10704, new_n1240, new_n10705);
nand_5 g10320(new_n10705, new_n1234, new_n10706);
nand_5 g10321(new_n10706, new_n1231, new_n10707);
nand_5 g10322(new_n10707, new_n1227, new_n10708);
nand_5 g10323(new_n10708, new_n1407, new_n10709);
nand_5 g10324(new_n10709, new_n1223, new_n10710);
nand_5 g10325(new_n10710, new_n1218, new_n10711);
nand_5 g10326(new_n10711, new_n1213, new_n10712);
nand_5 g10327(new_n10712, new_n1210, new_n10713);
nand_5 g10328(new_n10713, new_n1206, new_n10714);
nand_5 g10329(new_n10714, new_n1418, new_n10715);
nand_5 g10330(new_n10715, new_n1422, new_n10716);
nand_5 g10331(new_n10716, new_n1428, new_n10717);
nand_5 g10332(new_n10717, new_n1203, new_n10718);
nand_5 g10333(new_n10718, new_n1433, new_n10719);
nand_5 g10334(new_n10719, new_n581, new_n10720);
nand_5 g10335(new_n10720, new_n574, new_n10721);
nand_5 g10336(new_n10721, new_n568, new_n10722);
nand_5 g10337(new_n10722, new_n589, new_n10723);
nand_5 g10338(new_n10723, new_n595, new_n10724);
nand_5 g10339(new_n10724, new_n601, new_n10725);
nand_5 g10340(new_n10725, new_n563, new_n10726);
nand_5 g10341(new_n10726, new_n608, new_n10727);
nand_5 g10342(new_n10727, new_n558, new_n10728);
nand_5 g10343(new_n10728, new_n615, new_n10729);
nand_5 g10344(new_n10729, new_n553, new_n10730);
nand_5 g10345(new_n10730, new_n622, new_n10731);
nand_5 g10346(new_n10731, new_n628, new_n10732);
nand_5 g10347(new_n10732, new_n548, new_n10733);
nand_5 g10348(new_n10733, new_n543_1, new_n10734);
nand_5 g10349(new_n10734, new_n636, new_n10735);
nand_5 g10350(new_n10735, new_n642, new_n10736_1);
nand_5 g10351(new_n10736_1, new_n538, new_n10737);
nand_5 g10352(new_n10737, new_n533, new_n10738);
nand_5 g10353(new_n10738, new_n650_1, new_n10739);
nand_5 g10354(new_n10739, new_n528, new_n10740);
nand_5 g10355(new_n10740, new_n523, new_n10741);
nand_5 g10356(new_n10741, new_n518, new_n10742);
nand_5 g10357(new_n10742, new_n659, new_n10743);
nand_5 g10358(new_n10743, new_n665, new_n10744);
nand_5 g10359(new_n10744, new_n672, new_n10745);
nand_5 g10360(new_n10745, new_n513, new_n10746);
nand_5 g10361(new_n10746, new_n679, new_n10747);
nand_5 g10362(new_n10747, new_n685, new_n10748);
nand_5 g10363(new_n10748, new_n691, new_n10749);
nand_5 g10364(new_n10749, new_n508, new_n10750_1);
nand_5 g10365(new_n10750_1, new_n698, new_n10751);
nand_5 g10366(new_n10751, new_n503, new_n10752);
nand_5 g10367(new_n10752, new_n704, new_n10753);
nand_5 g10368(new_n10753, new_n498_1, new_n10754);
nand_5 g10369(new_n10754, new_n711, new_n10755);
nand_5 g10370(new_n10755, new_n493, new_n10756);
nand_5 g10371(new_n10756, new_n718, new_n10757);
nand_5 g10372(new_n10757, new_n488, new_n10758);
nand_5 g10373(new_n10758, new_n725, new_n10759);
nand_5 g10374(new_n10759, new_n483, new_n10760);
nand_5 g10375(new_n10760, new_n732, new_n10761);
nand_5 g10376(new_n10761, new_n478, new_n10762);
nand_5 g10377(new_n10762, new_n739, new_n10763);
nand_5 g10378(new_n10763, new_n745, new_n10764);
nand_5 g10379(new_n10764, new_n751, new_n10765_1);
nand_5 g10380(new_n10765_1, new_n473, new_n10766);
nand_5 g10381(new_n10766, new_n758, new_n10767);
nand_5 g10382(new_n10767, new_n764, new_n10768);
nand_5 g10383(new_n10768, new_n770, new_n10769);
nand_5 g10384(new_n10769, new_n468, new_n10770);
nand_5 g10385(new_n10770, new_n777, new_n10771);
nand_5 g10386(new_n10771, new_n783, new_n10772);
nand_5 g10387(new_n10772, new_n789, new_n10773);
nand_5 g10388(new_n10773, new_n463, new_n10774);
nand_5 g10389(new_n10774, new_n796, new_n10775);
nand_5 g10390(new_n10775, new_n458, new_n10776);
nand_5 g10391(new_n10776, new_n453, new_n10777);
nand_5 g10392(new_n10777, new_n447, new_n10778);
nand_5 g10393(new_n10778, new_n805, new_n10779);
nand_5 g10394(new_n10779, new_n811, new_n10780);
nand_5 g10395(new_n10780, new_n442, new_n10781);
nand_5 g10396(new_n10781, new_n437, new_n10782);
nand_5 g10397(new_n10782, new_n819, new_n10783);
nand_5 g10398(new_n10783, new_n432, new_n10784);
nand_5 g10399(new_n10784, new_n427_1, new_n10785);
nand_5 g10400(new_n10785, n14464, new_n10786);
nor_5  g10401(new_n10786, new_n419, n12355);
nand_5 g10402(new_n1652, new_n1082, new_n10788);
nand_5 g10403(new_n10788, new_n1134, new_n10789);
nand_5 g10404(new_n10789, new_n1080, new_n10790);
nand_5 g10405(new_n10790, new_n1075, new_n10791_1);
nand_5 g10406(new_n10791_1, new_n1070, new_n10792);
nand_5 g10407(new_n10792, new_n1143, new_n10793);
nand_5 g10408(new_n10793, new_n1148, new_n10794);
nand_5 g10409(new_n10794, new_n1065, new_n10795);
nand_5 g10410(new_n10795, new_n1062, new_n10796);
nand_5 g10411(new_n10796, new_n1156, new_n10797);
nand_5 g10412(new_n10797, new_n1057, new_n10798);
nand_5 g10413(new_n10798, new_n1053, new_n10799);
nand_5 g10414(new_n10799, new_n1050, new_n10800);
nand_5 g10415(new_n10800, new_n1045, new_n10801);
nand_5 g10416(new_n10801, new_n1040, new_n10802_1);
nand_5 g10417(new_n10802_1, new_n1036, new_n10803);
nand_5 g10418(new_n10803, new_n1033, new_n10804);
nand_5 g10419(new_n10804, new_n1028, new_n10805);
nand_5 g10420(new_n10805, new_n1026, new_n10806);
nand_5 g10421(new_n10806, new_n1021, new_n10807);
nand_5 g10422(new_n10807, new_n1017, new_n10808);
nand_5 g10423(new_n10808, new_n1012, new_n10809);
nand_5 g10424(new_n10809, new_n1009, new_n10810);
nand_5 g10425(new_n10810, new_n1004, new_n10811);
nand_5 g10426(new_n10811, new_n1000, new_n10812);
nand_5 g10427(new_n10812, new_n995, new_n10813);
nand_5 g10428(new_n10813, new_n990, new_n10814);
nand_5 g10429(new_n10814, new_n985, new_n10815);
nand_5 g10430(new_n10815, new_n981, new_n10816);
nand_5 g10431(new_n10816, new_n1179, new_n10817);
nand_5 g10432(new_n10817, new_n976, new_n10818);
nand_5 g10433(new_n10818, new_n971, new_n10819);
nand_5 g10434(new_n10819, new_n966, new_n10820);
nand_5 g10435(new_n10820, new_n961, new_n10821);
nand_5 g10436(new_n10821, new_n957, new_n10822);
nand_5 g10437(new_n10822, new_n952, new_n10823);
nand_5 g10438(new_n10823, new_n948_1, new_n10824);
nand_5 g10439(new_n10824, new_n943, new_n10825);
nand_5 g10440(new_n10825, new_n941, new_n10826);
nand_5 g10441(new_n10826, new_n938, new_n10827);
nand_5 g10442(new_n10827, new_n936, new_n10828);
nand_5 g10443(new_n10828, new_n931, new_n10829);
nand_5 g10444(new_n10829, new_n927, new_n10830);
nand_5 g10445(new_n10830, new_n922, new_n10831);
nand_5 g10446(new_n10831, new_n917, new_n10832);
nand_5 g10447(new_n10832, new_n912, new_n10833);
nand_5 g10448(new_n10833, new_n907, new_n10834);
nand_5 g10449(new_n10834, new_n903, new_n10835);
nand_5 g10450(new_n10835, new_n2066, new_n10836);
nand_5 g10451(new_n10836, new_n2063, new_n10837);
nand_5 g10452(new_n10837, new_n2062, new_n10838);
nand_5 g10453(new_n10838, new_n2058, new_n10839);
nand_5 g10454(new_n10839, new_n2055, new_n10840);
nand_5 g10455(new_n10840, new_n2051, new_n10841);
nand_5 g10456(new_n10841, new_n2046, new_n10842);
nand_5 g10457(new_n10842, new_n2042, new_n10843);
nand_5 g10458(new_n10843, new_n2039, new_n10844);
nand_5 g10459(new_n10844, new_n2036, new_n10845);
nand_5 g10460(new_n10845, new_n2033, new_n10846);
nand_5 g10461(new_n10846, new_n2029, new_n10847);
nand_5 g10462(new_n10847, new_n2026, new_n10848);
nand_5 g10463(new_n10848, new_n2022, new_n10849);
nand_5 g10464(new_n10849, new_n2018, new_n10850);
nand_5 g10465(new_n10850, new_n1726, new_n10851);
nand_5 g10466(new_n10851, new_n1722, new_n10852);
nand_5 g10467(new_n10852, new_n1718, new_n10853);
nand_5 g10468(new_n10853, new_n1713, new_n10854);
nand_5 g10469(new_n10854, new_n1737, new_n10855);
nand_5 g10470(new_n10855, new_n1709, new_n10856);
nand_5 g10471(new_n10856, new_n1742, new_n10857);
nand_5 g10472(new_n10857, new_n1704, new_n10858);
nand_5 g10473(new_n10858, new_n1702_1, new_n10859);
nand_5 g10474(new_n10859, new_n1698, new_n10860);
nand_5 g10475(new_n10860, new_n1695, new_n10861);
nand_5 g10476(new_n10861, new_n1692, new_n10862_1);
nand_5 g10477(new_n10862_1, new_n1752, new_n10863);
nand_5 g10478(new_n10863, new_n1688, new_n10864);
nand_5 g10479(new_n10864, new_n1685, new_n10865);
nand_5 g10480(new_n10865, new_n1680, new_n10866);
nand_5 g10481(new_n10866, new_n1676, new_n10867);
nand_5 g10482(new_n10867, new_n1672, new_n10868);
nand_5 g10483(new_n10868, new_n1669, new_n10869);
nand_5 g10484(new_n10869, new_n1666, new_n10870);
nand_5 g10485(new_n10870, new_n1663, new_n10871);
nand_5 g10486(new_n10871, n2201, new_n10872);
nor_5  g10487(new_n10872, new_n1655, n12535);
not_4  g10488(new_n1584, new_n10874);
nand_5 g10489(new_n10874, new_n981, new_n10875);
nand_5 g10490(new_n10875, new_n1179, new_n10876);
nand_5 g10491(new_n10876, new_n976, new_n10877);
nand_5 g10492(new_n10877, new_n971, new_n10878);
nand_5 g10493(new_n10878, new_n966, new_n10879);
nand_5 g10494(new_n10879, new_n961, new_n10880);
nand_5 g10495(new_n10880, new_n957, new_n10881);
nand_5 g10496(new_n10881, new_n952, new_n10882);
nand_5 g10497(new_n10882, new_n948_1, new_n10883);
nand_5 g10498(new_n10883, new_n943, new_n10884);
nand_5 g10499(new_n10884, new_n941, new_n10885);
nand_5 g10500(new_n10885, new_n938, new_n10886);
nand_5 g10501(new_n10886, new_n936, new_n10887);
nand_5 g10502(new_n10887, new_n931, new_n10888);
nand_5 g10503(new_n10888, new_n927, new_n10889);
nand_5 g10504(new_n10889, new_n922, new_n10890);
nand_5 g10505(new_n10890, new_n917, new_n10891);
nand_5 g10506(new_n10891, new_n912, new_n10892);
nand_5 g10507(new_n10892, new_n907, new_n10893);
nand_5 g10508(new_n10893, new_n903, new_n10894);
nand_5 g10509(new_n10894, new_n2066, new_n10895);
nand_5 g10510(new_n10895, new_n2063, new_n10896);
nand_5 g10511(new_n10896, new_n2062, new_n10897);
nand_5 g10512(new_n10897, new_n2058, new_n10898);
nand_5 g10513(new_n10898, new_n2055, new_n10899);
nand_5 g10514(new_n10899, new_n2051, new_n10900);
nand_5 g10515(new_n10900, new_n2046, new_n10901);
nand_5 g10516(new_n10901, new_n2042, new_n10902);
nand_5 g10517(new_n10902, new_n2039, new_n10903);
nand_5 g10518(new_n10903, new_n2036, new_n10904);
nand_5 g10519(new_n10904, new_n2033, new_n10905);
nand_5 g10520(new_n10905, new_n2029, new_n10906);
nand_5 g10521(new_n10906, new_n2026, new_n10907);
nand_5 g10522(new_n10907, new_n2022, new_n10908);
nand_5 g10523(new_n10908, new_n2018, new_n10909);
nand_5 g10524(new_n10909, new_n1726, new_n10910);
nand_5 g10525(new_n10910, new_n1722, new_n10911);
nand_5 g10526(new_n10911, new_n1718, new_n10912_1);
nand_5 g10527(new_n10912_1, new_n1713, new_n10913);
nand_5 g10528(new_n10913, new_n1737, new_n10914);
nand_5 g10529(new_n10914, new_n1709, new_n10915_1);
nand_5 g10530(new_n10915_1, new_n1742, new_n10916);
nand_5 g10531(new_n10916, new_n1704, new_n10917);
nand_5 g10532(new_n10917, new_n1702_1, new_n10918);
nand_5 g10533(new_n10918, new_n1698, new_n10919);
nand_5 g10534(new_n10919, new_n1695, new_n10920);
nand_5 g10535(new_n10920, new_n1692, new_n10921);
nand_5 g10536(new_n10921, new_n1752, new_n10922);
nand_5 g10537(new_n10922, new_n1688, new_n10923);
nand_5 g10538(new_n10923, new_n1685, new_n10924);
nand_5 g10539(new_n10924, new_n1680, new_n10925);
nand_5 g10540(new_n10925, new_n1676, new_n10926);
nand_5 g10541(new_n10926, new_n1672, new_n10927);
nand_5 g10542(new_n10927, new_n1669, new_n10928);
nand_5 g10543(new_n10928, new_n1666, new_n10929);
nand_5 g10544(new_n10929, new_n1663, new_n10930);
nand_5 g10545(new_n10930, new_n1658, new_n10931);
nand_5 g10546(new_n10931, new_n1653, new_n10932);
nand_5 g10547(new_n10932, new_n1651, new_n10933);
nand_5 g10548(new_n10933, new_n1649, new_n10934);
nand_5 g10549(new_n10934, new_n1646, new_n10935);
nand_5 g10550(new_n10935, new_n1643, new_n10936);
nand_5 g10551(new_n10936, new_n1641, new_n10937);
nand_5 g10552(new_n10937, new_n1638, new_n10938);
nand_5 g10553(new_n10938, new_n1635, new_n10939);
nand_5 g10554(new_n10939, new_n1632, new_n10940);
nand_5 g10555(new_n10940, new_n1628, new_n10941);
nand_5 g10556(new_n10941, new_n1625, new_n10942);
nand_5 g10557(new_n10942, new_n1621, new_n10943);
nand_5 g10558(new_n10943, new_n1618, new_n10944);
nand_5 g10559(new_n10944, new_n1778, new_n10945_1);
nand_5 g10560(new_n10945_1, new_n1782, new_n10946);
nand_5 g10561(new_n10946, new_n1614, new_n10947);
nand_5 g10562(new_n10947, new_n1611, new_n10948);
nand_5 g10563(new_n10948, new_n1789, new_n10949);
nand_5 g10564(new_n10949, new_n1608, new_n10950);
nand_5 g10565(new_n10950, new_n1605, new_n10951);
nand_5 g10566(new_n10951, new_n1795, new_n10952);
nand_5 g10567(new_n10952, new_n1799, new_n10953);
nand_5 g10568(new_n10953, new_n1602, new_n10954);
nand_5 g10569(new_n10954, new_n1599, new_n10955);
nand_5 g10570(new_n10955, new_n1596, new_n10956);
nand_5 g10571(new_n10956, new_n1593, new_n10957);
nand_5 g10572(new_n10957, new_n1806, new_n10958);
nand_5 g10573(new_n10958, n3893, new_n10959);
nor_5  g10574(new_n10959, new_n676, n12989);
nand_5 g10575(new_n951, new_n491, new_n10961);
nand_5 g10576(new_n10961, new_n718, new_n10962);
nand_5 g10577(new_n10962, new_n488, new_n10963);
nand_5 g10578(new_n10963, new_n725, new_n10964);
nand_5 g10579(new_n10964, new_n483, new_n10965);
nand_5 g10580(new_n10965, new_n732, new_n10966);
nand_5 g10581(new_n10966, new_n478, new_n10967);
nand_5 g10582(new_n10967, new_n739, new_n10968);
nand_5 g10583(new_n10968, new_n745, new_n10969);
nand_5 g10584(new_n10969, new_n751, new_n10970);
nand_5 g10585(new_n10970, new_n473, new_n10971);
nand_5 g10586(new_n10971, new_n758, new_n10972);
nand_5 g10587(new_n10972, new_n764, new_n10973);
nand_5 g10588(new_n10973, new_n770, new_n10974);
nand_5 g10589(new_n10974, new_n468, new_n10975);
nand_5 g10590(new_n10975, new_n777, new_n10976);
nand_5 g10591(new_n10976, new_n783, new_n10977);
nand_5 g10592(new_n10977, new_n789, new_n10978);
nand_5 g10593(new_n10978, new_n463, new_n10979);
nand_5 g10594(new_n10979, new_n796, new_n10980);
nand_5 g10595(new_n10980, new_n458, new_n10981);
nand_5 g10596(new_n10981, new_n453, new_n10982);
nand_5 g10597(new_n10982, new_n447, new_n10983);
nand_5 g10598(new_n10983, new_n805, new_n10984);
nand_5 g10599(new_n10984, new_n811, new_n10985);
nand_5 g10600(new_n10985, new_n442, new_n10986);
nand_5 g10601(new_n10986, new_n437, new_n10987);
nand_5 g10602(new_n10987, new_n819, new_n10988);
nand_5 g10603(new_n10988, new_n432, new_n10989);
nand_5 g10604(new_n10989, new_n427_1, new_n10990);
nand_5 g10605(new_n10990, new_n422, new_n10991);
nand_5 g10606(new_n10991, new_n828, new_n10992);
nand_5 g10607(new_n10992, new_n834, new_n10993);
nand_5 g10608(new_n10993, new_n840, new_n10994);
nand_5 g10609(new_n10994, new_n417, new_n10995);
nand_5 g10610(new_n10995, new_n847, new_n10996);
nand_5 g10611(new_n10996, new_n853, new_n10997);
nand_5 g10612(new_n10997, new_n859, new_n10998);
nand_5 g10613(new_n10998, new_n412, new_n10999);
nand_5 g10614(new_n10999, new_n866, new_n11000);
nand_5 g10615(new_n11000, new_n872, new_n11001);
nand_5 g10616(new_n11001, new_n878, new_n11002);
nand_5 g10617(new_n11002, new_n407, new_n11003);
nand_5 g10618(new_n11003, new_n885, new_n11004);
nand_5 g10619(new_n11004, new_n402, new_n11005);
nand_5 g10620(new_n11005, new_n397, new_n11006);
nand_5 g10621(new_n11006, new_n392, new_n11007);
nand_5 g10622(new_n11007, new_n894, new_n11008);
nand_5 g10623(new_n11008, new_n1087, new_n11009);
nand_5 g10624(new_n11009, new_n1129, new_n11010);
nand_5 g10625(new_n11010, new_n1084, new_n11011);
nand_5 g10626(new_n11011, new_n1134, new_n11012);
nand_5 g10627(new_n11012, new_n1080, new_n11013);
nand_5 g10628(new_n11013, new_n1075, new_n11014);
nand_5 g10629(new_n11014, new_n1070, new_n11015);
nand_5 g10630(new_n11015, new_n1143, new_n11016);
nand_5 g10631(new_n11016, new_n1148, new_n11017);
nand_5 g10632(new_n11017, new_n1065, new_n11018);
nand_5 g10633(new_n11018, new_n1062, new_n11019);
nand_5 g10634(new_n11019, new_n1156, new_n11020);
nand_5 g10635(new_n11020, new_n1057, new_n11021);
nand_5 g10636(new_n11021, new_n1053, new_n11022);
nand_5 g10637(new_n11022, new_n1050, new_n11023);
nand_5 g10638(new_n11023, new_n1045, new_n11024);
nand_5 g10639(new_n11024, new_n1040, new_n11025);
nand_5 g10640(new_n11025, new_n1036, new_n11026);
nand_5 g10641(new_n11026, new_n1033, new_n11027);
nand_5 g10642(new_n11027, new_n1028, new_n11028);
nand_5 g10643(new_n11028, new_n1026, new_n11029);
nand_5 g10644(new_n11029, new_n1021, new_n11030);
nand_5 g10645(new_n11030, new_n1017, new_n11031);
nand_5 g10646(new_n11031, new_n1012, new_n11032);
nand_5 g10647(new_n11032, new_n1009, new_n11033);
nand_5 g10648(new_n11033, new_n1004, new_n11034);
nand_5 g10649(new_n11034, new_n1000, new_n11035);
nand_5 g10650(new_n11035, new_n995, new_n11036);
nand_5 g10651(new_n11036, new_n990, new_n11037);
nand_5 g10652(new_n11037, new_n985, new_n11038);
nand_5 g10653(new_n11038, new_n981, new_n11039);
nand_5 g10654(new_n11039, new_n1179, new_n11040);
nand_5 g10655(new_n11040, new_n976, new_n11041);
nand_5 g10656(new_n11041, new_n971, new_n11042);
nand_5 g10657(new_n11042, new_n966, new_n11043);
nand_5 g10658(new_n11043, new_n961, new_n11044);
nand_5 g10659(new_n11044, n10061, new_n11045);
nor_5  g10660(new_n11045, new_n954, n13010);
nand_5 g10661(new_n909, new_n907, new_n11047);
nand_5 g10662(new_n11047, new_n903, new_n11048);
nand_5 g10663(new_n11048, new_n2066, new_n11049);
nand_5 g10664(new_n11049, new_n2063, new_n11050);
nand_5 g10665(new_n11050, new_n2062, new_n11051);
nand_5 g10666(new_n11051, new_n2058, new_n11052);
nand_5 g10667(new_n11052, new_n2055, new_n11053);
nand_5 g10668(new_n11053, new_n2051, new_n11054);
nand_5 g10669(new_n11054, new_n2046, new_n11055);
nand_5 g10670(new_n11055, new_n2042, new_n11056);
nand_5 g10671(new_n11056, new_n2039, new_n11057);
nand_5 g10672(new_n11057, new_n2036, new_n11058);
nand_5 g10673(new_n11058, new_n2033, new_n11059);
nand_5 g10674(new_n11059, new_n2029, new_n11060);
nand_5 g10675(new_n11060, new_n2026, new_n11061);
nand_5 g10676(new_n11061, new_n2022, new_n11062);
nand_5 g10677(new_n11062, new_n2018, new_n11063);
nand_5 g10678(new_n11063, new_n1726, new_n11064);
nand_5 g10679(new_n11064, new_n1722, new_n11065);
nand_5 g10680(new_n11065, new_n1718, new_n11066);
nand_5 g10681(new_n11066, new_n1713, new_n11067);
nand_5 g10682(new_n11067, new_n1737, new_n11068);
nand_5 g10683(new_n11068, new_n1709, new_n11069);
nand_5 g10684(new_n11069, new_n1742, new_n11070);
nand_5 g10685(new_n11070, new_n1704, new_n11071);
nand_5 g10686(new_n11071, new_n1702_1, new_n11072);
nand_5 g10687(new_n11072, new_n1698, new_n11073);
nand_5 g10688(new_n11073, new_n1695, new_n11074);
nand_5 g10689(new_n11074, new_n1692, new_n11075);
nand_5 g10690(new_n11075, new_n1752, new_n11076);
nand_5 g10691(new_n11076, new_n1688, new_n11077);
nand_5 g10692(new_n11077, new_n1685, new_n11078);
nand_5 g10693(new_n11078, new_n1680, new_n11079);
nand_5 g10694(new_n11079, new_n1676, new_n11080);
nand_5 g10695(new_n11080, new_n1672, new_n11081);
nand_5 g10696(new_n11081, new_n1669, new_n11082);
nand_5 g10697(new_n11082, new_n1666, new_n11083);
nand_5 g10698(new_n11083, new_n1663, new_n11084);
nand_5 g10699(new_n11084, new_n1658, new_n11085);
nand_5 g10700(new_n11085, new_n1653, new_n11086);
nand_5 g10701(new_n11086, new_n1651, new_n11087);
nand_5 g10702(new_n11087, new_n1649, new_n11088);
nand_5 g10703(new_n11088, new_n1646, new_n11089);
nand_5 g10704(new_n11089, new_n1643, new_n11090);
nand_5 g10705(new_n11090, new_n1641, new_n11091);
nand_5 g10706(new_n11091, new_n1638, new_n11092);
nand_5 g10707(new_n11092, new_n1635, new_n11093);
nand_5 g10708(new_n11093, new_n1632, new_n11094);
nand_5 g10709(new_n11094, new_n1628, new_n11095);
nand_5 g10710(new_n11095, new_n1625, new_n11096);
nand_5 g10711(new_n11096, new_n1621, new_n11097);
nand_5 g10712(new_n11097, new_n1618, new_n11098);
nand_5 g10713(new_n11098, new_n1778, new_n11099);
nand_5 g10714(new_n11099, new_n1782, new_n11100);
nand_5 g10715(new_n11100, new_n1614, new_n11101);
nand_5 g10716(new_n11101, new_n1611, new_n11102);
nand_5 g10717(new_n11102, new_n1789, new_n11103);
nand_5 g10718(new_n11103, new_n1608, new_n11104);
nand_5 g10719(new_n11104, new_n1605, new_n11105);
nand_5 g10720(new_n11105, new_n1795, new_n11106);
nand_5 g10721(new_n11106, new_n1799, new_n11107);
nand_5 g10722(new_n11107, new_n1602, new_n11108);
nand_5 g10723(new_n11108, new_n1599, new_n11109);
nand_5 g10724(new_n11109, new_n1596, new_n11110);
nand_5 g10725(new_n11110, new_n1593, new_n11111);
nand_5 g10726(new_n11111, new_n1806, new_n11112);
nand_5 g10727(new_n11112, new_n1589, new_n11113);
nand_5 g10728(new_n11113, new_n1586, new_n11114);
nand_5 g10729(new_n11114, new_n1583, new_n11115);
nand_5 g10730(new_n11115, new_n1580, new_n11116);
nand_5 g10731(new_n11116, new_n1576, new_n11117);
nand_5 g10732(new_n11117, new_n1573, new_n11118);
nand_5 g10733(new_n11118, new_n1570, new_n11119);
nand_5 g10734(new_n11119, new_n1567, new_n11120);
nand_5 g10735(new_n11120, new_n1564, new_n11121);
nand_5 g10736(new_n11121, new_n1561, new_n11122_1);
nand_5 g10737(new_n11122_1, new_n1338, new_n11123);
nand_5 g10738(new_n11123, new_n1331, new_n11124);
nand_5 g10739(new_n11124, new_n1326, new_n11125);
nand_5 g10740(new_n11125, new_n1321, new_n11126);
nand_5 g10741(new_n11126, new_n1318, new_n11127);
nand_5 g10742(new_n11127, new_n1315, new_n11128);
nand_5 g10743(new_n11128, new_n1312, new_n11129);
nand_5 g10744(new_n11129, new_n1309, new_n11130);
nand_5 g10745(new_n11130, n12321, new_n11131);
nor_5  g10746(new_n11131, new_n748, n13045);
nand_5 g10747(new_n930, new_n476, new_n11133);
nand_5 g10748(new_n11133, new_n739, new_n11134);
nand_5 g10749(new_n11134, new_n745, new_n11135);
nand_5 g10750(new_n11135, new_n751, new_n11136);
nand_5 g10751(new_n11136, new_n473, new_n11137);
nand_5 g10752(new_n11137, new_n758, new_n11138);
nand_5 g10753(new_n11138, new_n764, new_n11139);
nand_5 g10754(new_n11139, new_n770, new_n11140);
nand_5 g10755(new_n11140, new_n468, new_n11141);
nand_5 g10756(new_n11141, new_n777, new_n11142);
nand_5 g10757(new_n11142, new_n783, new_n11143_1);
nand_5 g10758(new_n11143_1, new_n789, new_n11144);
nand_5 g10759(new_n11144, new_n463, new_n11145);
nand_5 g10760(new_n11145, new_n796, new_n11146);
nand_5 g10761(new_n11146, new_n458, new_n11147);
nand_5 g10762(new_n11147, new_n453, new_n11148);
nand_5 g10763(new_n11148, new_n447, new_n11149);
nand_5 g10764(new_n11149, new_n805, new_n11150);
nand_5 g10765(new_n11150, new_n811, new_n11151);
nand_5 g10766(new_n11151, new_n442, new_n11152);
nand_5 g10767(new_n11152, new_n437, new_n11153);
nand_5 g10768(new_n11153, new_n819, new_n11154);
nand_5 g10769(new_n11154, new_n432, new_n11155);
nand_5 g10770(new_n11155, new_n427_1, new_n11156);
nand_5 g10771(new_n11156, new_n422, new_n11157);
nand_5 g10772(new_n11157, new_n828, new_n11158_1);
nand_5 g10773(new_n11158_1, new_n834, new_n11159);
nand_5 g10774(new_n11159, new_n840, new_n11160);
nand_5 g10775(new_n11160, new_n417, new_n11161);
nand_5 g10776(new_n11161, new_n847, new_n11162);
nand_5 g10777(new_n11162, new_n853, new_n11163);
nand_5 g10778(new_n11163, new_n859, new_n11164);
nand_5 g10779(new_n11164, new_n412, new_n11165);
nand_5 g10780(new_n11165, new_n866, new_n11166);
nand_5 g10781(new_n11166, new_n872, new_n11167);
nand_5 g10782(new_n11167, new_n878, new_n11168);
nand_5 g10783(new_n11168, new_n407, new_n11169);
nand_5 g10784(new_n11169, new_n885, new_n11170);
nand_5 g10785(new_n11170, new_n402, new_n11171);
nand_5 g10786(new_n11171, new_n397, new_n11172);
nand_5 g10787(new_n11172, new_n392, new_n11173);
nand_5 g10788(new_n11173, new_n894, new_n11174);
nand_5 g10789(new_n11174, new_n1087, new_n11175);
nand_5 g10790(new_n11175, new_n1129, new_n11176);
nand_5 g10791(new_n11176, new_n1084, new_n11177);
nand_5 g10792(new_n11177, new_n1134, new_n11178);
nand_5 g10793(new_n11178, new_n1080, new_n11179);
nand_5 g10794(new_n11179, new_n1075, new_n11180);
nand_5 g10795(new_n11180, new_n1070, new_n11181);
nand_5 g10796(new_n11181, new_n1143, new_n11182);
nand_5 g10797(new_n11182, new_n1148, new_n11183);
nand_5 g10798(new_n11183, new_n1065, new_n11184);
nand_5 g10799(new_n11184, new_n1062, new_n11185);
nand_5 g10800(new_n11185, new_n1156, new_n11186);
nand_5 g10801(new_n11186, new_n1057, new_n11187);
nand_5 g10802(new_n11187, new_n1053, new_n11188);
nand_5 g10803(new_n11188, new_n1050, new_n11189);
nand_5 g10804(new_n11189, new_n1045, new_n11190);
nand_5 g10805(new_n11190, new_n1040, new_n11191);
nand_5 g10806(new_n11191, new_n1036, new_n11192);
nand_5 g10807(new_n11192, new_n1033, new_n11193);
nand_5 g10808(new_n11193, new_n1028, new_n11194);
nand_5 g10809(new_n11194, new_n1026, new_n11195);
nand_5 g10810(new_n11195, new_n1021, new_n11196);
nand_5 g10811(new_n11196, new_n1017, new_n11197);
nand_5 g10812(new_n11197, new_n1012, new_n11198);
nand_5 g10813(new_n11198, new_n1009, new_n11199);
nand_5 g10814(new_n11199, new_n1004, new_n11200);
nand_5 g10815(new_n11200, new_n1000, new_n11201);
nand_5 g10816(new_n11201, new_n995, new_n11202);
nand_5 g10817(new_n11202, new_n990, new_n11203);
nand_5 g10818(new_n11203, new_n985, new_n11204);
nand_5 g10819(new_n11204, new_n981, new_n11205);
nand_5 g10820(new_n11205, new_n1179, new_n11206);
nand_5 g10821(new_n11206, new_n976, new_n11207);
nand_5 g10822(new_n11207, new_n971, new_n11208);
nand_5 g10823(new_n11208, new_n966, new_n11209);
nand_5 g10824(new_n11209, new_n961, new_n11210);
nand_5 g10825(new_n11210, new_n957, new_n11211);
nand_5 g10826(new_n11211, new_n952, new_n11212);
nand_5 g10827(new_n11212, new_n948_1, new_n11213);
nand_5 g10828(new_n11213, new_n943, new_n11214);
nand_5 g10829(new_n11214, new_n941, new_n11215);
nand_5 g10830(new_n11215, new_n938, new_n11216);
nand_5 g10831(new_n11216, n10470, new_n11217);
nor_5  g10832(new_n11217, new_n933, n13114);
nand_5 g10833(new_n2064, new_n1296, new_n11219);
nand_5 g10834(new_n11219, new_n2063, new_n11220);
nand_5 g10835(new_n11220, new_n2062, new_n11221);
nand_5 g10836(new_n11221, new_n2058, new_n11222);
nand_5 g10837(new_n11222, new_n2055, new_n11223);
nand_5 g10838(new_n11223, new_n2051, new_n11224);
nand_5 g10839(new_n11224, new_n2046, new_n11225);
nand_5 g10840(new_n11225, new_n2042, new_n11226);
nand_5 g10841(new_n11226, new_n2039, new_n11227);
nand_5 g10842(new_n11227, new_n2036, new_n11228);
nand_5 g10843(new_n11228, new_n2033, new_n11229);
nand_5 g10844(new_n11229, new_n2029, new_n11230);
nand_5 g10845(new_n11230, new_n2026, new_n11231);
nand_5 g10846(new_n11231, new_n2022, new_n11232);
nand_5 g10847(new_n11232, new_n2018, new_n11233);
nand_5 g10848(new_n11233, new_n1726, new_n11234);
nand_5 g10849(new_n11234, new_n1722, new_n11235);
nand_5 g10850(new_n11235, new_n1718, new_n11236);
nand_5 g10851(new_n11236, new_n1713, new_n11237);
nand_5 g10852(new_n11237, new_n1737, new_n11238);
nand_5 g10853(new_n11238, new_n1709, new_n11239);
nand_5 g10854(new_n11239, new_n1742, new_n11240);
nand_5 g10855(new_n11240, new_n1704, new_n11241);
nand_5 g10856(new_n11241, new_n1702_1, new_n11242);
nand_5 g10857(new_n11242, new_n1698, new_n11243);
nand_5 g10858(new_n11243, new_n1695, new_n11244);
nand_5 g10859(new_n11244, new_n1692, new_n11245);
nand_5 g10860(new_n11245, new_n1752, new_n11246);
nand_5 g10861(new_n11246, new_n1688, new_n11247);
nand_5 g10862(new_n11247, new_n1685, new_n11248);
nand_5 g10863(new_n11248, new_n1680, new_n11249);
nand_5 g10864(new_n11249, new_n1676, new_n11250);
nand_5 g10865(new_n11250, new_n1672, new_n11251);
nand_5 g10866(new_n11251, new_n1669, new_n11252);
nand_5 g10867(new_n11252, new_n1666, new_n11253);
nand_5 g10868(new_n11253, new_n1663, new_n11254);
nand_5 g10869(new_n11254, new_n1658, new_n11255);
nand_5 g10870(new_n11255, new_n1653, new_n11256);
nand_5 g10871(new_n11256, new_n1651, new_n11257);
nand_5 g10872(new_n11257, new_n1649, new_n11258);
nand_5 g10873(new_n11258, new_n1646, new_n11259);
nand_5 g10874(new_n11259, new_n1643, new_n11260);
nand_5 g10875(new_n11260, new_n1641, new_n11261);
nand_5 g10876(new_n11261, new_n1638, new_n11262);
nand_5 g10877(new_n11262, new_n1635, new_n11263);
nand_5 g10878(new_n11263, new_n1632, new_n11264);
nand_5 g10879(new_n11264, new_n1628, new_n11265);
nand_5 g10880(new_n11265, new_n1625, new_n11266);
nand_5 g10881(new_n11266, new_n1621, new_n11267);
nand_5 g10882(new_n11267, new_n1618, new_n11268);
nand_5 g10883(new_n11268, new_n1778, new_n11269_1);
nand_5 g10884(new_n11269_1, new_n1782, new_n11270);
nand_5 g10885(new_n11270, new_n1614, new_n11271);
nand_5 g10886(new_n11271, new_n1611, new_n11272);
nand_5 g10887(new_n11272, new_n1789, new_n11273);
nand_5 g10888(new_n11273, new_n1608, new_n11274);
nand_5 g10889(new_n11274, new_n1605, new_n11275);
nand_5 g10890(new_n11275, new_n1795, new_n11276);
nand_5 g10891(new_n11276, new_n1799, new_n11277);
nand_5 g10892(new_n11277, new_n1602, new_n11278);
nand_5 g10893(new_n11278, new_n1599, new_n11279);
nand_5 g10894(new_n11279, new_n1596, new_n11280);
nand_5 g10895(new_n11280, new_n1593, new_n11281);
nand_5 g10896(new_n11281, new_n1806, new_n11282);
nand_5 g10897(new_n11282, new_n1589, new_n11283);
nand_5 g10898(new_n11283, new_n1586, new_n11284);
nand_5 g10899(new_n11284, new_n1583, new_n11285);
nand_5 g10900(new_n11285, new_n1580, new_n11286);
nand_5 g10901(new_n11286, new_n1576, new_n11287);
nand_5 g10902(new_n11287, new_n1573, new_n11288);
nand_5 g10903(new_n11288, new_n1570, new_n11289);
nand_5 g10904(new_n11289, new_n1567, new_n11290);
nand_5 g10905(new_n11290, new_n1564, new_n11291);
nand_5 g10906(new_n11291, new_n1561, new_n11292);
nand_5 g10907(new_n11292, new_n1338, new_n11293);
nand_5 g10908(new_n11293, new_n1331, new_n11294);
nand_5 g10909(new_n11294, new_n1326, new_n11295);
nand_5 g10910(new_n11295, new_n1321, new_n11296);
nand_5 g10911(new_n11296, new_n1318, new_n11297);
nand_5 g10912(new_n11297, new_n1315, new_n11298);
nand_5 g10913(new_n11298, new_n1312, new_n11299);
nand_5 g10914(new_n11299, new_n1309, new_n11300);
nand_5 g10915(new_n11300, new_n1307, new_n11301);
nand_5 g10916(new_n11301, new_n1304, new_n11302);
nand_5 g10917(new_n11302, n4147, new_n11303);
nor_5  g10918(new_n11303, new_n755, n13141);
nand_5 g10919(new_n1686, new_n1217, new_n11305);
nand_5 g10920(new_n11305, new_n1685, new_n11306);
nand_5 g10921(new_n11306, new_n1680, new_n11307);
nand_5 g10922(new_n11307, new_n1676, new_n11308);
nand_5 g10923(new_n11308, new_n1672, new_n11309);
nand_5 g10924(new_n11309, new_n1669, new_n11310);
nand_5 g10925(new_n11310, new_n1666, new_n11311);
nand_5 g10926(new_n11311, new_n1663, new_n11312);
nand_5 g10927(new_n11312, new_n1658, new_n11313);
nand_5 g10928(new_n11313, new_n1653, new_n11314);
nand_5 g10929(new_n11314, new_n1651, new_n11315);
nand_5 g10930(new_n11315, new_n1649, new_n11316);
nand_5 g10931(new_n11316, new_n1646, new_n11317);
nand_5 g10932(new_n11317, new_n1643, new_n11318);
nand_5 g10933(new_n11318, new_n1641, new_n11319);
nand_5 g10934(new_n11319, new_n1638, new_n11320);
nand_5 g10935(new_n11320, new_n1635, new_n11321);
nand_5 g10936(new_n11321, new_n1632, new_n11322);
nand_5 g10937(new_n11322, new_n1628, new_n11323);
nand_5 g10938(new_n11323, new_n1625, new_n11324);
nand_5 g10939(new_n11324, new_n1621, new_n11325);
nand_5 g10940(new_n11325, new_n1618, new_n11326);
nand_5 g10941(new_n11326, new_n1778, new_n11327);
nand_5 g10942(new_n11327, new_n1782, new_n11328);
nand_5 g10943(new_n11328, new_n1614, new_n11329);
nand_5 g10944(new_n11329, new_n1611, new_n11330);
nand_5 g10945(new_n11330, new_n1789, new_n11331);
nand_5 g10946(new_n11331, new_n1608, new_n11332);
nand_5 g10947(new_n11332, new_n1605, new_n11333);
nand_5 g10948(new_n11333, new_n1795, new_n11334);
nand_5 g10949(new_n11334, new_n1799, new_n11335);
nand_5 g10950(new_n11335, new_n1602, new_n11336);
nand_5 g10951(new_n11336, new_n1599, new_n11337);
nand_5 g10952(new_n11337, new_n1596, new_n11338);
nand_5 g10953(new_n11338, new_n1593, new_n11339);
nand_5 g10954(new_n11339, new_n1806, new_n11340);
nand_5 g10955(new_n11340, new_n1589, new_n11341);
nand_5 g10956(new_n11341, new_n1586, new_n11342);
nand_5 g10957(new_n11342, new_n1583, new_n11343);
nand_5 g10958(new_n11343, new_n1580, new_n11344);
nand_5 g10959(new_n11344, new_n1576, new_n11345_1);
nand_5 g10960(new_n11345_1, new_n1573, new_n11346);
nand_5 g10961(new_n11346, new_n1570, new_n11347);
nand_5 g10962(new_n11347, new_n1567, new_n11348);
nand_5 g10963(new_n11348, new_n1564, new_n11349);
nand_5 g10964(new_n11349, new_n1561, new_n11350);
nand_5 g10965(new_n11350, new_n1338, new_n11351);
nand_5 g10966(new_n11351, new_n1331, new_n11352);
nand_5 g10967(new_n11352, new_n1326, new_n11353);
nand_5 g10968(new_n11353, new_n1321, new_n11354);
nand_5 g10969(new_n11354, new_n1318, new_n11355);
nand_5 g10970(new_n11355, new_n1315, new_n11356);
nand_5 g10971(new_n11356, new_n1312, new_n11357);
nand_5 g10972(new_n11357, new_n1309, new_n11358);
nand_5 g10973(new_n11358, new_n1307, new_n11359);
nand_5 g10974(new_n11359, new_n1304, new_n11360);
nand_5 g10975(new_n11360, new_n1300, new_n11361);
nand_5 g10976(new_n11361, new_n1297, new_n11362);
nand_5 g10977(new_n11362, new_n1294, new_n11363);
nand_5 g10978(new_n11363, new_n1355, new_n11364);
nand_5 g10979(new_n11364, new_n1291, new_n11365);
nand_5 g10980(new_n11365, new_n1288, new_n11366);
nand_5 g10981(new_n11366, new_n1283, new_n11367);
nand_5 g10982(new_n11367, new_n1363, new_n11368);
nand_5 g10983(new_n11368, new_n1280, new_n11369);
nand_5 g10984(new_n11369, new_n1370, new_n11370);
nand_5 g10985(new_n11370, new_n1373, new_n11371);
nand_5 g10986(new_n11371, new_n1277, new_n11372);
nand_5 g10987(new_n11372, new_n1272, new_n11373);
nand_5 g10988(new_n11373, new_n1269, new_n11374);
nand_5 g10989(new_n11374, new_n1380, new_n11375);
nand_5 g10990(new_n11375, new_n1264, new_n11376);
nand_5 g10991(new_n11376, new_n1259, new_n11377);
nand_5 g10992(new_n11377, new_n1388, new_n11378);
nand_5 g10993(new_n11378, new_n1392, new_n11379);
nand_5 g10994(new_n11379, new_n1256, new_n11380);
nand_5 g10995(new_n11380, new_n1252, new_n11381);
nand_5 g10996(new_n11381, new_n1249, new_n11382);
nand_5 g10997(new_n11382, new_n1244, new_n11383);
nand_5 g10998(new_n11383, new_n1240, new_n11384);
nand_5 g10999(new_n11384, new_n1234, new_n11385);
nand_5 g11000(new_n11385, new_n1231, new_n11386);
nand_5 g11001(new_n11386, new_n1227, new_n11387);
nand_5 g11002(new_n11387, new_n1407, new_n11388);
nand_5 g11003(new_n11388, n5467, new_n11389);
nor_5  g11004(new_n11389, new_n1220, n13316);
nand_5 g11005(new_n1154, new_n1623, new_n11391);
nand_5 g11006(new_n11391, new_n551, new_n11392);
nand_5 g11007(new_n11392, new_n622, new_n11393_1);
nand_5 g11008(new_n11393_1, new_n628, new_n11394);
nand_5 g11009(new_n11394, new_n548, new_n11395);
nand_5 g11010(new_n11395, new_n543_1, new_n11396);
nand_5 g11011(new_n11396, new_n636, new_n11397);
nand_5 g11012(new_n11397, new_n642, new_n11398);
nand_5 g11013(new_n11398, new_n538, new_n11399);
nand_5 g11014(new_n11399, new_n533, new_n11400);
nand_5 g11015(new_n11400, new_n650_1, new_n11401);
nand_5 g11016(new_n11401, new_n528, new_n11402);
nand_5 g11017(new_n11402, new_n523, new_n11403);
nand_5 g11018(new_n11403, new_n518, new_n11404_1);
nand_5 g11019(new_n11404_1, new_n659, new_n11405);
nand_5 g11020(new_n11405, new_n665, new_n11406);
nand_5 g11021(new_n11406, new_n672, new_n11407);
nand_5 g11022(new_n11407, new_n513, new_n11408);
nand_5 g11023(new_n11408, new_n679, new_n11409);
nand_5 g11024(new_n11409, new_n685, new_n11410);
nand_5 g11025(new_n11410, new_n691, new_n11411);
nand_5 g11026(new_n11411, new_n508, new_n11412);
nand_5 g11027(new_n11412, new_n698, new_n11413);
nand_5 g11028(new_n11413, new_n503, new_n11414);
nand_5 g11029(new_n11414, new_n704, new_n11415);
nand_5 g11030(new_n11415, new_n498_1, new_n11416);
nand_5 g11031(new_n11416, new_n711, new_n11417);
nand_5 g11032(new_n11417, new_n493, new_n11418);
nand_5 g11033(new_n11418, new_n718, new_n11419);
nand_5 g11034(new_n11419, new_n488, new_n11420);
nand_5 g11035(new_n11420, new_n725, new_n11421);
nand_5 g11036(new_n11421, new_n483, new_n11422);
nand_5 g11037(new_n11422, new_n732, new_n11423);
nand_5 g11038(new_n11423, new_n478, new_n11424);
nand_5 g11039(new_n11424, new_n739, new_n11425);
nand_5 g11040(new_n11425, new_n745, new_n11426);
nand_5 g11041(new_n11426, new_n751, new_n11427);
nand_5 g11042(new_n11427, new_n473, new_n11428);
nand_5 g11043(new_n11428, new_n758, new_n11429);
nand_5 g11044(new_n11429, new_n764, new_n11430);
nand_5 g11045(new_n11430, new_n770, new_n11431);
nand_5 g11046(new_n11431, new_n468, new_n11432);
nand_5 g11047(new_n11432, new_n777, new_n11433);
nand_5 g11048(new_n11433, new_n783, new_n11434);
nand_5 g11049(new_n11434, new_n789, new_n11435);
nand_5 g11050(new_n11435, new_n463, new_n11436);
nand_5 g11051(new_n11436, new_n796, new_n11437);
nand_5 g11052(new_n11437, new_n458, new_n11438);
nand_5 g11053(new_n11438, new_n453, new_n11439);
nand_5 g11054(new_n11439, new_n447, new_n11440);
nand_5 g11055(new_n11440, new_n805, new_n11441);
nand_5 g11056(new_n11441, new_n811, new_n11442);
nand_5 g11057(new_n11442, new_n442, new_n11443);
nand_5 g11058(new_n11443, new_n437, new_n11444);
nand_5 g11059(new_n11444, new_n819, new_n11445);
nand_5 g11060(new_n11445, new_n432, new_n11446);
nand_5 g11061(new_n11446, new_n427_1, new_n11447);
nand_5 g11062(new_n11447, new_n422, new_n11448);
nand_5 g11063(new_n11448, new_n828, new_n11449);
nand_5 g11064(new_n11449, new_n834, new_n11450);
nand_5 g11065(new_n11450, new_n840, new_n11451);
nand_5 g11066(new_n11451, new_n417, new_n11452);
nand_5 g11067(new_n11452, new_n847, new_n11453);
nand_5 g11068(new_n11453, new_n853, new_n11454);
nand_5 g11069(new_n11454, new_n859, new_n11455);
nand_5 g11070(new_n11455, new_n412, new_n11456);
nand_5 g11071(new_n11456, new_n866, new_n11457);
nand_5 g11072(new_n11457, new_n872, new_n11458);
nand_5 g11073(new_n11458, new_n878, new_n11459);
nand_5 g11074(new_n11459, new_n407, new_n11460);
nand_5 g11075(new_n11460, new_n885, new_n11461);
nand_5 g11076(new_n11461, new_n402, new_n11462);
nand_5 g11077(new_n11462, new_n397, new_n11463_1);
nand_5 g11078(new_n11463_1, new_n392, new_n11464);
nand_5 g11079(new_n11464, new_n894, new_n11465);
nand_5 g11080(new_n11465, new_n1087, new_n11466);
nand_5 g11081(new_n11466, new_n1129, new_n11467);
nand_5 g11082(new_n11467, new_n1084, new_n11468);
nand_5 g11083(new_n11468, new_n1134, new_n11469);
nand_5 g11084(new_n11469, new_n1080, new_n11470);
nand_5 g11085(new_n11470, new_n1075, new_n11471);
nand_5 g11086(new_n11471, new_n1070, new_n11472);
nand_5 g11087(new_n11472, new_n1143, new_n11473);
nand_5 g11088(new_n11473, new_n1148, new_n11474);
nand_5 g11089(new_n11474, new_n1065, new_n11475);
nand_5 g11090(new_n11475, n9110, new_n11476);
nor_5  g11091(new_n11476, new_n1059, n13577);
nand_5 g11092(new_n1204, new_n884_1, new_n11478);
nand_5 g11093(new_n11478, new_n1418, new_n11479);
nand_5 g11094(new_n11479, new_n1422, new_n11480);
nand_5 g11095(new_n11480, new_n1428, new_n11481);
nand_5 g11096(new_n11481, new_n1203, new_n11482);
nand_5 g11097(new_n11482, new_n1433, new_n11483);
nand_5 g11098(new_n11483, new_n581, new_n11484);
nand_5 g11099(new_n11484, new_n574, new_n11485);
nand_5 g11100(new_n11485, new_n568, new_n11486);
nand_5 g11101(new_n11486, new_n589, new_n11487);
nand_5 g11102(new_n11487, new_n595, new_n11488);
nand_5 g11103(new_n11488, new_n601, new_n11489);
nand_5 g11104(new_n11489, new_n563, new_n11490);
nand_5 g11105(new_n11490, new_n608, new_n11491);
nand_5 g11106(new_n11491, new_n558, new_n11492);
nand_5 g11107(new_n11492, new_n615, new_n11493);
nand_5 g11108(new_n11493, new_n553, new_n11494);
nand_5 g11109(new_n11494, new_n622, new_n11495);
nand_5 g11110(new_n11495, new_n628, new_n11496);
nand_5 g11111(new_n11496, new_n548, new_n11497);
nand_5 g11112(new_n11497, new_n543_1, new_n11498);
nand_5 g11113(new_n11498, new_n636, new_n11499);
nand_5 g11114(new_n11499, new_n642, new_n11500);
nand_5 g11115(new_n11500, new_n538, new_n11501);
nand_5 g11116(new_n11501, new_n533, new_n11502);
nand_5 g11117(new_n11502, new_n650_1, new_n11503);
nand_5 g11118(new_n11503, new_n528, new_n11504);
nand_5 g11119(new_n11504, new_n523, new_n11505);
nand_5 g11120(new_n11505, new_n518, new_n11506);
nand_5 g11121(new_n11506, new_n659, new_n11507);
nand_5 g11122(new_n11507, new_n665, new_n11508);
nand_5 g11123(new_n11508, new_n672, new_n11509);
nand_5 g11124(new_n11509, new_n513, new_n11510);
nand_5 g11125(new_n11510, new_n679, new_n11511);
nand_5 g11126(new_n11511, new_n685, new_n11512);
nand_5 g11127(new_n11512, new_n691, new_n11513);
nand_5 g11128(new_n11513, new_n508, new_n11514);
nand_5 g11129(new_n11514, new_n698, new_n11515);
nand_5 g11130(new_n11515, new_n503, new_n11516);
nand_5 g11131(new_n11516, new_n704, new_n11517);
nand_5 g11132(new_n11517, new_n498_1, new_n11518);
nand_5 g11133(new_n11518, new_n711, new_n11519);
nand_5 g11134(new_n11519, new_n493, new_n11520);
nand_5 g11135(new_n11520, new_n718, new_n11521);
nand_5 g11136(new_n11521, new_n488, new_n11522);
nand_5 g11137(new_n11522, new_n725, new_n11523);
nand_5 g11138(new_n11523, new_n483, new_n11524);
nand_5 g11139(new_n11524, new_n732, new_n11525);
nand_5 g11140(new_n11525, new_n478, new_n11526);
nand_5 g11141(new_n11526, new_n739, new_n11527);
nand_5 g11142(new_n11527, new_n745, new_n11528);
nand_5 g11143(new_n11528, new_n751, new_n11529_1);
nand_5 g11144(new_n11529_1, new_n473, new_n11530);
nand_5 g11145(new_n11530, new_n758, new_n11531);
nand_5 g11146(new_n11531, new_n764, new_n11532);
nand_5 g11147(new_n11532, new_n770, new_n11533);
nand_5 g11148(new_n11533, new_n468, new_n11534_1);
nand_5 g11149(new_n11534_1, new_n777, new_n11535);
nand_5 g11150(new_n11535, new_n783, new_n11536);
nand_5 g11151(new_n11536, new_n789, new_n11537);
nand_5 g11152(new_n11537, new_n463, new_n11538);
nand_5 g11153(new_n11538, new_n796, new_n11539);
nand_5 g11154(new_n11539, new_n458, new_n11540);
nand_5 g11155(new_n11540, new_n453, new_n11541);
nand_5 g11156(new_n11541, new_n447, new_n11542);
nand_5 g11157(new_n11542, new_n805, new_n11543);
nand_5 g11158(new_n11543, new_n811, new_n11544);
nand_5 g11159(new_n11544, new_n442, new_n11545);
nand_5 g11160(new_n11545, new_n437, new_n11546);
nand_5 g11161(new_n11546, new_n819, new_n11547);
nand_5 g11162(new_n11547, new_n432, new_n11548);
nand_5 g11163(new_n11548, new_n427_1, new_n11549);
nand_5 g11164(new_n11549, new_n422, new_n11550);
nand_5 g11165(new_n11550, new_n828, new_n11551);
nand_5 g11166(new_n11551, new_n834, new_n11552);
nand_5 g11167(new_n11552, new_n840, new_n11553);
nand_5 g11168(new_n11553, new_n417, new_n11554);
nand_5 g11169(new_n11554, new_n847, new_n11555);
nand_5 g11170(new_n11555, new_n853, new_n11556);
nand_5 g11171(new_n11556, new_n859, new_n11557);
nand_5 g11172(new_n11557, new_n412, new_n11558);
nand_5 g11173(new_n11558, new_n866, new_n11559);
nand_5 g11174(new_n11559, new_n872, new_n11560);
nand_5 g11175(new_n11560, new_n878, new_n11561);
nand_5 g11176(new_n11561, n12927, new_n11562);
nor_5  g11177(new_n11562, new_n404, n13639);
nand_5 g11178(new_n1211, new_n877, new_n11564);
nand_5 g11179(new_n11564, new_n1210, new_n11565);
nand_5 g11180(new_n11565, new_n1206, new_n11566);
nand_5 g11181(new_n11566, new_n1418, new_n11567);
nand_5 g11182(new_n11567, new_n1422, new_n11568);
nand_5 g11183(new_n11568, new_n1428, new_n11569);
nand_5 g11184(new_n11569, new_n1203, new_n11570);
nand_5 g11185(new_n11570, new_n1433, new_n11571);
nand_5 g11186(new_n11571, new_n581, new_n11572);
nand_5 g11187(new_n11572, new_n574, new_n11573);
nand_5 g11188(new_n11573, new_n568, new_n11574);
nand_5 g11189(new_n11574, new_n589, new_n11575);
nand_5 g11190(new_n11575, new_n595, new_n11576);
nand_5 g11191(new_n11576, new_n601, new_n11577);
nand_5 g11192(new_n11577, new_n563, new_n11578);
nand_5 g11193(new_n11578, new_n608, new_n11579);
nand_5 g11194(new_n11579, new_n558, new_n11580);
nand_5 g11195(new_n11580, new_n615, new_n11581);
nand_5 g11196(new_n11581, new_n553, new_n11582);
nand_5 g11197(new_n11582, new_n622, new_n11583);
nand_5 g11198(new_n11583, new_n628, new_n11584);
nand_5 g11199(new_n11584, new_n548, new_n11585);
nand_5 g11200(new_n11585, new_n543_1, new_n11586);
nand_5 g11201(new_n11586, new_n636, new_n11587);
nand_5 g11202(new_n11587, new_n642, new_n11588);
nand_5 g11203(new_n11588, new_n538, new_n11589);
nand_5 g11204(new_n11589, new_n533, new_n11590_1);
nand_5 g11205(new_n11590_1, new_n650_1, new_n11591);
nand_5 g11206(new_n11591, new_n528, new_n11592);
nand_5 g11207(new_n11592, new_n523, new_n11593);
nand_5 g11208(new_n11593, new_n518, new_n11594);
nand_5 g11209(new_n11594, new_n659, new_n11595);
nand_5 g11210(new_n11595, new_n665, new_n11596);
nand_5 g11211(new_n11596, new_n672, new_n11597);
nand_5 g11212(new_n11597, new_n513, new_n11598);
nand_5 g11213(new_n11598, new_n679, new_n11599);
nand_5 g11214(new_n11599, new_n685, new_n11600);
nand_5 g11215(new_n11600, new_n691, new_n11601);
nand_5 g11216(new_n11601, new_n508, new_n11602);
nand_5 g11217(new_n11602, new_n698, new_n11603);
nand_5 g11218(new_n11603, new_n503, new_n11604);
nand_5 g11219(new_n11604, new_n704, new_n11605_1);
nand_5 g11220(new_n11605_1, new_n498_1, new_n11606);
nand_5 g11221(new_n11606, new_n711, new_n11607);
nand_5 g11222(new_n11607, new_n493, new_n11608);
nand_5 g11223(new_n11608, new_n718, new_n11609);
nand_5 g11224(new_n11609, new_n488, new_n11610);
nand_5 g11225(new_n11610, new_n725, new_n11611);
nand_5 g11226(new_n11611, new_n483, new_n11612);
nand_5 g11227(new_n11612, new_n732, new_n11613);
nand_5 g11228(new_n11613, new_n478, new_n11614);
nand_5 g11229(new_n11614, new_n739, new_n11615);
nand_5 g11230(new_n11615, new_n745, new_n11616);
nand_5 g11231(new_n11616, new_n751, new_n11617);
nand_5 g11232(new_n11617, new_n473, new_n11618);
nand_5 g11233(new_n11618, new_n758, new_n11619);
nand_5 g11234(new_n11619, new_n764, new_n11620);
nand_5 g11235(new_n11620, new_n770, new_n11621);
nand_5 g11236(new_n11621, new_n468, new_n11622);
nand_5 g11237(new_n11622, new_n777, new_n11623);
nand_5 g11238(new_n11623, new_n783, new_n11624);
nand_5 g11239(new_n11624, new_n789, new_n11625);
nand_5 g11240(new_n11625, new_n463, new_n11626);
nand_5 g11241(new_n11626, new_n796, new_n11627_1);
nand_5 g11242(new_n11627_1, new_n458, new_n11628);
nand_5 g11243(new_n11628, new_n453, new_n11629);
nand_5 g11244(new_n11629, new_n447, new_n11630);
nand_5 g11245(new_n11630, new_n805, new_n11631);
nand_5 g11246(new_n11631, new_n811, new_n11632);
nand_5 g11247(new_n11632, new_n442, new_n11633);
nand_5 g11248(new_n11633, new_n437, new_n11634);
nand_5 g11249(new_n11634, new_n819, new_n11635);
nand_5 g11250(new_n11635, new_n432, new_n11636);
nand_5 g11251(new_n11636, new_n427_1, new_n11637);
nand_5 g11252(new_n11637, new_n422, new_n11638);
nand_5 g11253(new_n11638, new_n828, new_n11639);
nand_5 g11254(new_n11639, new_n834, new_n11640);
nand_5 g11255(new_n11640, new_n840, new_n11641);
nand_5 g11256(new_n11641, new_n417, new_n11642);
nand_5 g11257(new_n11642, new_n847, new_n11643);
nand_5 g11258(new_n11643, new_n853, new_n11644);
nand_5 g11259(new_n11644, new_n859, new_n11645);
nand_5 g11260(new_n11645, new_n412, new_n11646);
nand_5 g11261(new_n11646, new_n866, new_n11647);
nand_5 g11262(new_n11647, n7282, new_n11648);
nor_5  g11263(new_n11648, new_n869, n13658);
not_4  g11264(n13231, new_n11650);
nand_5 g11265(new_n1630, new_n11650, new_n11651);
nand_5 g11266(new_n11651, new_n1060, new_n11652);
nand_5 g11267(new_n11652, new_n1156, new_n11653);
nand_5 g11268(new_n11653, new_n1057, new_n11654);
nand_5 g11269(new_n11654, new_n1053, new_n11655);
nand_5 g11270(new_n11655, new_n1050, new_n11656);
nand_5 g11271(new_n11656, new_n1045, new_n11657);
nand_5 g11272(new_n11657, new_n1040, new_n11658);
nand_5 g11273(new_n11658, new_n1036, new_n11659);
nand_5 g11274(new_n11659, new_n1033, new_n11660);
nand_5 g11275(new_n11660, new_n1028, new_n11661);
nand_5 g11276(new_n11661, new_n1026, new_n11662);
nand_5 g11277(new_n11662, new_n1021, new_n11663);
nand_5 g11278(new_n11663, new_n1017, new_n11664_1);
nand_5 g11279(new_n11664_1, new_n1012, new_n11665);
nand_5 g11280(new_n11665, new_n1009, new_n11666_1);
nand_5 g11281(new_n11666_1, new_n1004, new_n11667);
nand_5 g11282(new_n11667, new_n1000, new_n11668);
nand_5 g11283(new_n11668, new_n995, new_n11669);
nand_5 g11284(new_n11669, new_n990, new_n11670);
nand_5 g11285(new_n11670, new_n985, new_n11671);
nand_5 g11286(new_n11671, new_n981, new_n11672);
nand_5 g11287(new_n11672, new_n1179, new_n11673);
nand_5 g11288(new_n11673, new_n976, new_n11674);
nand_5 g11289(new_n11674, new_n971, new_n11675);
nand_5 g11290(new_n11675, new_n966, new_n11676);
nand_5 g11291(new_n11676, new_n961, new_n11677);
nand_5 g11292(new_n11677, new_n957, new_n11678);
nand_5 g11293(new_n11678, new_n952, new_n11679);
nand_5 g11294(new_n11679, new_n948_1, new_n11680);
nand_5 g11295(new_n11680, new_n943, new_n11681);
nand_5 g11296(new_n11681, new_n941, new_n11682);
nand_5 g11297(new_n11682, new_n938, new_n11683);
nand_5 g11298(new_n11683, new_n936, new_n11684);
nand_5 g11299(new_n11684, new_n931, new_n11685);
nand_5 g11300(new_n11685, new_n927, new_n11686);
nand_5 g11301(new_n11686, new_n922, new_n11687);
nand_5 g11302(new_n11687, new_n917, new_n11688);
nand_5 g11303(new_n11688, new_n912, new_n11689);
nand_5 g11304(new_n11689, new_n907, new_n11690);
nand_5 g11305(new_n11690, new_n903, new_n11691);
nand_5 g11306(new_n11691, new_n2066, new_n11692);
nand_5 g11307(new_n11692, new_n2063, new_n11693);
nand_5 g11308(new_n11693, new_n2062, new_n11694);
nand_5 g11309(new_n11694, new_n2058, new_n11695);
nand_5 g11310(new_n11695, new_n2055, new_n11696);
nand_5 g11311(new_n11696, new_n2051, new_n11697);
nand_5 g11312(new_n11697, new_n2046, new_n11698);
nand_5 g11313(new_n11698, new_n2042, new_n11699);
nand_5 g11314(new_n11699, new_n2039, new_n11700);
nand_5 g11315(new_n11700, new_n2036, new_n11701);
nand_5 g11316(new_n11701, new_n2033, new_n11702);
nand_5 g11317(new_n11702, new_n2029, new_n11703);
nand_5 g11318(new_n11703, new_n2026, new_n11704);
nand_5 g11319(new_n11704, new_n2022, new_n11705);
nand_5 g11320(new_n11705, new_n2018, new_n11706);
nand_5 g11321(new_n11706, new_n1726, new_n11707);
nand_5 g11322(new_n11707, new_n1722, new_n11708);
nand_5 g11323(new_n11708, new_n1718, new_n11709);
nand_5 g11324(new_n11709, new_n1713, new_n11710);
nand_5 g11325(new_n11710, new_n1737, new_n11711);
nand_5 g11326(new_n11711, new_n1709, new_n11712);
nand_5 g11327(new_n11712, new_n1742, new_n11713);
nand_5 g11328(new_n11713, new_n1704, new_n11714);
nand_5 g11329(new_n11714, new_n1702_1, new_n11715);
nand_5 g11330(new_n11715, new_n1698, new_n11716);
nand_5 g11331(new_n11716, new_n1695, new_n11717);
nand_5 g11332(new_n11717, new_n1692, new_n11718);
nand_5 g11333(new_n11718, new_n1752, new_n11719);
nand_5 g11334(new_n11719, new_n1688, new_n11720);
nand_5 g11335(new_n11720, new_n1685, new_n11721);
nand_5 g11336(new_n11721, new_n1680, new_n11722);
nand_5 g11337(new_n11722, new_n1676, new_n11723);
nand_5 g11338(new_n11723, new_n1672, new_n11724);
nand_5 g11339(new_n11724, new_n1669, new_n11725);
nand_5 g11340(new_n11725, new_n1666, new_n11726);
nand_5 g11341(new_n11726, new_n1663, new_n11727);
nand_5 g11342(new_n11727, new_n1658, new_n11728);
nand_5 g11343(new_n11728, new_n1653, new_n11729);
nand_5 g11344(new_n11729, new_n1651, new_n11730);
nand_5 g11345(new_n11730, new_n1649, new_n11731);
nand_5 g11346(new_n11731, new_n1646, new_n11732);
nand_5 g11347(new_n11732, new_n1643, new_n11733);
nand_5 g11348(new_n11733, new_n1641, new_n11734);
nand_5 g11349(new_n11734, new_n1638, new_n11735);
nand_5 g11350(new_n11735, n74, new_n11736);
nor_5  g11351(new_n11736, new_n605, n13693);
not_4  g11352(new_n2044, new_n11738);
nand_5 g11353(new_n2041, new_n456, new_n11739);
nand_5 g11354(new_n11739, new_n453, new_n11740);
nand_5 g11355(new_n11740, new_n447, new_n11741);
nand_5 g11356(new_n11741, new_n805, new_n11742);
nand_5 g11357(new_n11742, new_n811, new_n11743);
nand_5 g11358(new_n11743, new_n442, new_n11744);
nand_5 g11359(new_n11744, new_n437, new_n11745);
nand_5 g11360(new_n11745, new_n819, new_n11746);
nand_5 g11361(new_n11746, new_n432, new_n11747);
nand_5 g11362(new_n11747, new_n427_1, new_n11748);
nand_5 g11363(new_n11748, new_n422, new_n11749);
nand_5 g11364(new_n11749, new_n828, new_n11750);
nand_5 g11365(new_n11750, new_n834, new_n11751);
nand_5 g11366(new_n11751, new_n840, new_n11752);
nand_5 g11367(new_n11752, new_n417, new_n11753);
nand_5 g11368(new_n11753, new_n847, new_n11754);
nand_5 g11369(new_n11754, new_n853, new_n11755);
nand_5 g11370(new_n11755, new_n859, new_n11756_1);
nand_5 g11371(new_n11756_1, new_n412, new_n11757);
nand_5 g11372(new_n11757, new_n866, new_n11758);
nand_5 g11373(new_n11758, new_n872, new_n11759);
nand_5 g11374(new_n11759, new_n878, new_n11760);
nand_5 g11375(new_n11760, new_n407, new_n11761);
nand_5 g11376(new_n11761, new_n885, new_n11762);
nand_5 g11377(new_n11762, new_n402, new_n11763);
nand_5 g11378(new_n11763, new_n397, new_n11764);
nand_5 g11379(new_n11764, new_n392, new_n11765);
nand_5 g11380(new_n11765, new_n894, new_n11766);
nand_5 g11381(new_n11766, new_n1087, new_n11767);
nand_5 g11382(new_n11767, new_n1129, new_n11768);
nand_5 g11383(new_n11768, new_n1084, new_n11769);
nand_5 g11384(new_n11769, new_n1134, new_n11770);
nand_5 g11385(new_n11770, new_n1080, new_n11771);
nand_5 g11386(new_n11771, new_n1075, new_n11772);
nand_5 g11387(new_n11772, new_n1070, new_n11773);
nand_5 g11388(new_n11773, new_n1143, new_n11774);
nand_5 g11389(new_n11774, new_n1148, new_n11775);
nand_5 g11390(new_n11775, new_n1065, new_n11776_1);
nand_5 g11391(new_n11776_1, new_n1062, new_n11777);
nand_5 g11392(new_n11777, new_n1156, new_n11778);
nand_5 g11393(new_n11778, new_n1057, new_n11779);
nand_5 g11394(new_n11779, new_n1053, new_n11780);
nand_5 g11395(new_n11780, new_n1050, new_n11781);
nand_5 g11396(new_n11781, new_n1045, new_n11782);
nand_5 g11397(new_n11782, new_n1040, new_n11783);
nand_5 g11398(new_n11783, new_n1036, new_n11784);
nand_5 g11399(new_n11784, new_n1033, new_n11785);
nand_5 g11400(new_n11785, new_n1028, new_n11786);
nand_5 g11401(new_n11786, new_n1026, new_n11787);
nand_5 g11402(new_n11787, new_n1021, new_n11788);
nand_5 g11403(new_n11788, new_n1017, new_n11789);
nand_5 g11404(new_n11789, new_n1012, new_n11790);
nand_5 g11405(new_n11790, new_n1009, new_n11791);
nand_5 g11406(new_n11791, new_n1004, new_n11792);
nand_5 g11407(new_n11792, new_n1000, new_n11793);
nand_5 g11408(new_n11793, new_n995, new_n11794);
nand_5 g11409(new_n11794, new_n990, new_n11795);
nand_5 g11410(new_n11795, new_n985, new_n11796);
nand_5 g11411(new_n11796, new_n981, new_n11797);
nand_5 g11412(new_n11797, new_n1179, new_n11798);
nand_5 g11413(new_n11798, new_n976, new_n11799);
nand_5 g11414(new_n11799, new_n971, new_n11800);
nand_5 g11415(new_n11800, new_n966, new_n11801);
nand_5 g11416(new_n11801, new_n961, new_n11802);
nand_5 g11417(new_n11802, new_n957, new_n11803);
nand_5 g11418(new_n11803, new_n952, new_n11804);
nand_5 g11419(new_n11804, new_n948_1, new_n11805);
nand_5 g11420(new_n11805, new_n943, new_n11806);
nand_5 g11421(new_n11806, new_n941, new_n11807);
nand_5 g11422(new_n11807, new_n938, new_n11808);
nand_5 g11423(new_n11808, new_n936, new_n11809);
nand_5 g11424(new_n11809, new_n931, new_n11810);
nand_5 g11425(new_n11810, new_n927, new_n11811);
nand_5 g11426(new_n11811, new_n922, new_n11812);
nand_5 g11427(new_n11812, new_n917, new_n11813);
nand_5 g11428(new_n11813, new_n912, new_n11814);
nand_5 g11429(new_n11814, new_n907, new_n11815);
nand_5 g11430(new_n11815, new_n903, new_n11816);
nand_5 g11431(new_n11816, new_n2066, new_n11817);
nand_5 g11432(new_n11817, new_n2063, new_n11818);
nand_5 g11433(new_n11818, new_n2062, new_n11819);
nand_5 g11434(new_n11819, new_n2058, new_n11820);
nand_5 g11435(new_n11820, new_n2055, new_n11821);
nand_5 g11436(new_n11821, new_n2051, new_n11822_1);
nand_5 g11437(new_n11822_1, n9921, new_n11823);
nor_5  g11438(new_n11823, new_n11738, n13760);
nand_5 g11439(new_n1042, new_n1040, new_n11825);
nand_5 g11440(new_n11825, new_n1036, new_n11826);
nand_5 g11441(new_n11826, new_n1033, new_n11827);
nand_5 g11442(new_n11827, new_n1028, new_n11828);
nand_5 g11443(new_n11828, new_n1026, new_n11829);
nand_5 g11444(new_n11829, new_n1021, new_n11830);
nand_5 g11445(new_n11830, new_n1017, new_n11831);
nand_5 g11446(new_n11831, new_n1012, new_n11832);
nand_5 g11447(new_n11832, new_n1009, new_n11833);
nand_5 g11448(new_n11833, new_n1004, new_n11834);
nand_5 g11449(new_n11834, new_n1000, new_n11835);
nand_5 g11450(new_n11835, new_n995, new_n11836);
nand_5 g11451(new_n11836, new_n990, new_n11837);
nand_5 g11452(new_n11837, new_n985, new_n11838);
nand_5 g11453(new_n11838, new_n981, new_n11839);
nand_5 g11454(new_n11839, new_n1179, new_n11840);
nand_5 g11455(new_n11840, new_n976, new_n11841);
nand_5 g11456(new_n11841, new_n971, new_n11842_1);
nand_5 g11457(new_n11842_1, new_n966, new_n11843);
nand_5 g11458(new_n11843, new_n961, new_n11844);
nand_5 g11459(new_n11844, new_n957, new_n11845);
nand_5 g11460(new_n11845, new_n952, new_n11846);
nand_5 g11461(new_n11846, new_n948_1, new_n11847_1);
nand_5 g11462(new_n11847_1, new_n943, new_n11848);
nand_5 g11463(new_n11848, new_n941, new_n11849);
nand_5 g11464(new_n11849, new_n938, new_n11850);
nand_5 g11465(new_n11850, new_n936, new_n11851);
nand_5 g11466(new_n11851, new_n931, new_n11852);
nand_5 g11467(new_n11852, new_n927, new_n11853);
nand_5 g11468(new_n11853, new_n922, new_n11854_1);
nand_5 g11469(new_n11854_1, new_n917, new_n11855);
nand_5 g11470(new_n11855, new_n912, new_n11856);
nand_5 g11471(new_n11856, new_n907, new_n11857);
nand_5 g11472(new_n11857, new_n903, new_n11858);
nand_5 g11473(new_n11858, new_n2066, new_n11859);
nand_5 g11474(new_n11859, new_n2063, new_n11860);
nand_5 g11475(new_n11860, new_n2062, new_n11861);
nand_5 g11476(new_n11861, new_n2058, new_n11862);
nand_5 g11477(new_n11862, new_n2055, new_n11863);
nand_5 g11478(new_n11863, new_n2051, new_n11864);
nand_5 g11479(new_n11864, new_n2046, new_n11865);
nand_5 g11480(new_n11865, new_n2042, new_n11866);
nand_5 g11481(new_n11866, new_n2039, new_n11867);
nand_5 g11482(new_n11867, new_n2036, new_n11868);
nand_5 g11483(new_n11868, new_n2033, new_n11869);
nand_5 g11484(new_n11869, new_n2029, new_n11870);
nand_5 g11485(new_n11870, new_n2026, new_n11871);
nand_5 g11486(new_n11871, new_n2022, new_n11872);
nand_5 g11487(new_n11872, new_n2018, new_n11873);
nand_5 g11488(new_n11873, new_n1726, new_n11874);
nand_5 g11489(new_n11874, new_n1722, new_n11875_1);
nand_5 g11490(new_n11875_1, new_n1718, new_n11876);
nand_5 g11491(new_n11876, new_n1713, new_n11877);
nand_5 g11492(new_n11877, new_n1737, new_n11878);
nand_5 g11493(new_n11878, new_n1709, new_n11879);
nand_5 g11494(new_n11879, new_n1742, new_n11880);
nand_5 g11495(new_n11880, new_n1704, new_n11881);
nand_5 g11496(new_n11881, new_n1702_1, new_n11882);
nand_5 g11497(new_n11882, new_n1698, new_n11883);
nand_5 g11498(new_n11883, new_n1695, new_n11884);
nand_5 g11499(new_n11884, new_n1692, new_n11885);
nand_5 g11500(new_n11885, new_n1752, new_n11886);
nand_5 g11501(new_n11886, new_n1688, new_n11887);
nand_5 g11502(new_n11887, new_n1685, new_n11888);
nand_5 g11503(new_n11888, new_n1680, new_n11889);
nand_5 g11504(new_n11889, new_n1676, new_n11890);
nand_5 g11505(new_n11890, new_n1672, new_n11891);
nand_5 g11506(new_n11891, new_n1669, new_n11892);
nand_5 g11507(new_n11892, new_n1666, new_n11893);
nand_5 g11508(new_n11893, new_n1663, new_n11894);
nand_5 g11509(new_n11894, new_n1658, new_n11895);
nand_5 g11510(new_n11895, new_n1653, new_n11896);
nand_5 g11511(new_n11896, new_n1651, new_n11897);
nand_5 g11512(new_n11897, new_n1649, new_n11898);
nand_5 g11513(new_n11898, new_n1646, new_n11899);
nand_5 g11514(new_n11899, new_n1643, new_n11900);
nand_5 g11515(new_n11900, new_n1641, new_n11901);
nand_5 g11516(new_n11901, new_n1638, new_n11902_1);
nand_5 g11517(new_n11902_1, new_n1635, new_n11903);
nand_5 g11518(new_n11903, new_n1632, new_n11904);
nand_5 g11519(new_n11904, new_n1628, new_n11905);
nand_5 g11520(new_n11905, new_n1625, new_n11906);
nand_5 g11521(new_n11906, new_n1621, new_n11907);
nand_5 g11522(new_n11907, new_n1618, new_n11908);
nand_5 g11523(new_n11908, n3367, new_n11909);
nor_5  g11524(new_n11909, new_n545, n13853);
not_4  g11525(n7450, new_n11911);
nand_5 g11526(new_n920, new_n11911, new_n11912);
nand_5 g11527(new_n11912, new_n743, new_n11913);
nand_5 g11528(new_n11913, new_n751, new_n11914);
nand_5 g11529(new_n11914, new_n473, new_n11915);
nand_5 g11530(new_n11915, new_n758, new_n11916);
nand_5 g11531(new_n11916, new_n764, new_n11917);
nand_5 g11532(new_n11917, new_n770, new_n11918);
nand_5 g11533(new_n11918, new_n468, new_n11919);
nand_5 g11534(new_n11919, new_n777, new_n11920);
nand_5 g11535(new_n11920, new_n783, new_n11921);
nand_5 g11536(new_n11921, new_n789, new_n11922);
nand_5 g11537(new_n11922, new_n463, new_n11923);
nand_5 g11538(new_n11923, new_n796, new_n11924);
nand_5 g11539(new_n11924, new_n458, new_n11925);
nand_5 g11540(new_n11925, new_n453, new_n11926);
nand_5 g11541(new_n11926, new_n447, new_n11927);
nand_5 g11542(new_n11927, new_n805, new_n11928);
nand_5 g11543(new_n11928, new_n811, new_n11929);
nand_5 g11544(new_n11929, new_n442, new_n11930_1);
nand_5 g11545(new_n11930_1, new_n437, new_n11931);
nand_5 g11546(new_n11931, new_n819, new_n11932);
nand_5 g11547(new_n11932, new_n432, new_n11933_1);
nand_5 g11548(new_n11933_1, new_n427_1, new_n11934);
nand_5 g11549(new_n11934, new_n422, new_n11935);
nand_5 g11550(new_n11935, new_n828, new_n11936);
nand_5 g11551(new_n11936, new_n834, new_n11937);
nand_5 g11552(new_n11937, new_n840, new_n11938);
nand_5 g11553(new_n11938, new_n417, new_n11939);
nand_5 g11554(new_n11939, new_n847, new_n11940);
nand_5 g11555(new_n11940, new_n853, new_n11941);
nand_5 g11556(new_n11941, new_n859, new_n11942);
nand_5 g11557(new_n11942, new_n412, new_n11943);
nand_5 g11558(new_n11943, new_n866, new_n11944);
nand_5 g11559(new_n11944, new_n872, new_n11945);
nand_5 g11560(new_n11945, new_n878, new_n11946);
nand_5 g11561(new_n11946, new_n407, new_n11947);
nand_5 g11562(new_n11947, new_n885, new_n11948);
nand_5 g11563(new_n11948, new_n402, new_n11949);
nand_5 g11564(new_n11949, new_n397, new_n11950);
nand_5 g11565(new_n11950, new_n392, new_n11951);
nand_5 g11566(new_n11951, new_n894, new_n11952);
nand_5 g11567(new_n11952, new_n1087, new_n11953);
nand_5 g11568(new_n11953, new_n1129, new_n11954);
nand_5 g11569(new_n11954, new_n1084, new_n11955);
nand_5 g11570(new_n11955, new_n1134, new_n11956);
nand_5 g11571(new_n11956, new_n1080, new_n11957);
nand_5 g11572(new_n11957, new_n1075, new_n11958);
nand_5 g11573(new_n11958, new_n1070, new_n11959);
nand_5 g11574(new_n11959, new_n1143, new_n11960);
nand_5 g11575(new_n11960, new_n1148, new_n11961_1);
nand_5 g11576(new_n11961_1, new_n1065, new_n11962);
nand_5 g11577(new_n11962, new_n1062, new_n11963);
nand_5 g11578(new_n11963, new_n1156, new_n11964);
nand_5 g11579(new_n11964, new_n1057, new_n11965);
nand_5 g11580(new_n11965, new_n1053, new_n11966);
nand_5 g11581(new_n11966, new_n1050, new_n11967);
nand_5 g11582(new_n11967, new_n1045, new_n11968);
nand_5 g11583(new_n11968, new_n1040, new_n11969);
nand_5 g11584(new_n11969, new_n1036, new_n11970);
nand_5 g11585(new_n11970, new_n1033, new_n11971);
nand_5 g11586(new_n11971, new_n1028, new_n11972);
nand_5 g11587(new_n11972, new_n1026, new_n11973);
nand_5 g11588(new_n11973, new_n1021, new_n11974);
nand_5 g11589(new_n11974, new_n1017, new_n11975);
nand_5 g11590(new_n11975, new_n1012, new_n11976);
nand_5 g11591(new_n11976, new_n1009, new_n11977);
nand_5 g11592(new_n11977, new_n1004, new_n11978);
nand_5 g11593(new_n11978, new_n1000, new_n11979);
nand_5 g11594(new_n11979, new_n995, new_n11980);
nand_5 g11595(new_n11980, new_n990, new_n11981);
nand_5 g11596(new_n11981, new_n985, new_n11982);
nand_5 g11597(new_n11982, new_n981, new_n11983);
nand_5 g11598(new_n11983, new_n1179, new_n11984);
nand_5 g11599(new_n11984, new_n976, new_n11985);
nand_5 g11600(new_n11985, new_n971, new_n11986);
nand_5 g11601(new_n11986, new_n966, new_n11987);
nand_5 g11602(new_n11987, new_n961, new_n11988);
nand_5 g11603(new_n11988, new_n957, new_n11989);
nand_5 g11604(new_n11989, new_n952, new_n11990);
nand_5 g11605(new_n11990, new_n948_1, new_n11991);
nand_5 g11606(new_n11991, new_n943, new_n11992);
nand_5 g11607(new_n11992, new_n941, new_n11993);
nand_5 g11608(new_n11993, new_n938, new_n11994);
nand_5 g11609(new_n11994, new_n936, new_n11995);
nand_5 g11610(new_n11995, new_n931, new_n11996);
nand_5 g11611(new_n11996, n7972, new_n11997);
nor_5  g11612(new_n11997, new_n924, n13870);
nand_5 g11613(new_n1328, new_n1326, new_n11999);
nand_5 g11614(new_n11999, new_n1321, new_n12000);
nand_5 g11615(new_n12000, new_n1318, new_n12001);
nand_5 g11616(new_n12001, new_n1315, new_n12002);
nand_5 g11617(new_n12002, new_n1312, new_n12003);
nand_5 g11618(new_n12003, new_n1309, new_n12004);
nand_5 g11619(new_n12004, new_n1307, new_n12005);
nand_5 g11620(new_n12005, new_n1304, new_n12006);
nand_5 g11621(new_n12006, new_n1300, new_n12007);
nand_5 g11622(new_n12007, new_n1297, new_n12008);
nand_5 g11623(new_n12008, new_n1294, new_n12009_1);
nand_5 g11624(new_n12009_1, new_n1355, new_n12010);
nand_5 g11625(new_n12010, new_n1291, new_n12011);
nand_5 g11626(new_n12011, new_n1288, new_n12012_1);
nand_5 g11627(new_n12012_1, new_n1283, new_n12013);
nand_5 g11628(new_n12013, new_n1363, new_n12014);
nand_5 g11629(new_n12014, new_n1280, new_n12015);
nand_5 g11630(new_n12015, new_n1370, new_n12016);
nand_5 g11631(new_n12016, new_n1373, new_n12017);
nand_5 g11632(new_n12017, new_n1277, new_n12018);
nand_5 g11633(new_n12018, new_n1272, new_n12019);
nand_5 g11634(new_n12019, new_n1269, new_n12020);
nand_5 g11635(new_n12020, new_n1380, new_n12021);
nand_5 g11636(new_n12021, new_n1264, new_n12022);
nand_5 g11637(new_n12022, new_n1259, new_n12023);
nand_5 g11638(new_n12023, new_n1388, new_n12024);
nand_5 g11639(new_n12024, new_n1392, new_n12025_1);
nand_5 g11640(new_n12025_1, new_n1256, new_n12026);
nand_5 g11641(new_n12026, new_n1252, new_n12027);
nand_5 g11642(new_n12027, new_n1249, new_n12028);
nand_5 g11643(new_n12028, new_n1244, new_n12029);
nand_5 g11644(new_n12029, new_n1240, new_n12030);
nand_5 g11645(new_n12030, new_n1234, new_n12031);
nand_5 g11646(new_n12031, new_n1231, new_n12032_1);
nand_5 g11647(new_n12032_1, new_n1227, new_n12033);
nand_5 g11648(new_n12033, new_n1407, new_n12034);
nand_5 g11649(new_n12034, new_n1223, new_n12035);
nand_5 g11650(new_n12035, new_n1218, new_n12036);
nand_5 g11651(new_n12036, new_n1213, new_n12037);
nand_5 g11652(new_n12037, new_n1210, new_n12038);
nand_5 g11653(new_n12038, new_n1206, new_n12039);
nand_5 g11654(new_n12039, new_n1418, new_n12040);
nand_5 g11655(new_n12040, new_n1422, new_n12041);
nand_5 g11656(new_n12041, new_n1428, new_n12042);
nand_5 g11657(new_n12042, new_n1203, new_n12043);
nand_5 g11658(new_n12043, new_n1433, new_n12044);
nand_5 g11659(new_n12044, new_n581, new_n12045);
nand_5 g11660(new_n12045, new_n574, new_n12046);
nand_5 g11661(new_n12046, new_n568, new_n12047);
nand_5 g11662(new_n12047, new_n589, new_n12048);
nand_5 g11663(new_n12048, new_n595, new_n12049);
nand_5 g11664(new_n12049, new_n601, new_n12050);
nand_5 g11665(new_n12050, new_n563, new_n12051);
nand_5 g11666(new_n12051, new_n608, new_n12052);
nand_5 g11667(new_n12052, new_n558, new_n12053);
nand_5 g11668(new_n12053, new_n615, new_n12054);
nand_5 g11669(new_n12054, new_n553, new_n12055);
nand_5 g11670(new_n12055, new_n622, new_n12056);
nand_5 g11671(new_n12056, new_n628, new_n12057);
nand_5 g11672(new_n12057, new_n548, new_n12058);
nand_5 g11673(new_n12058, new_n543_1, new_n12059);
nand_5 g11674(new_n12059, new_n636, new_n12060);
nand_5 g11675(new_n12060, new_n642, new_n12061);
nand_5 g11676(new_n12061, new_n538, new_n12062);
nand_5 g11677(new_n12062, new_n533, new_n12063);
nand_5 g11678(new_n12063, new_n650_1, new_n12064);
nand_5 g11679(new_n12064, new_n528, new_n12065);
nand_5 g11680(new_n12065, new_n523, new_n12066);
nand_5 g11681(new_n12066, new_n518, new_n12067);
nand_5 g11682(new_n12067, new_n659, new_n12068);
nand_5 g11683(new_n12068, new_n665, new_n12069);
nand_5 g11684(new_n12069, new_n672, new_n12070);
nand_5 g11685(new_n12070, new_n513, new_n12071);
nand_5 g11686(new_n12071, new_n679, new_n12072);
nand_5 g11687(new_n12072, new_n685, new_n12073);
nand_5 g11688(new_n12073, new_n691, new_n12074);
nand_5 g11689(new_n12074, new_n508, new_n12075);
nand_5 g11690(new_n12075, new_n698, new_n12076);
nand_5 g11691(new_n12076, new_n503, new_n12077);
nand_5 g11692(new_n12077, new_n704, new_n12078);
nand_5 g11693(new_n12078, new_n498_1, new_n12079);
nand_5 g11694(new_n12079, new_n711, new_n12080);
nand_5 g11695(new_n12080, new_n493, new_n12081);
nand_5 g11696(new_n12081, new_n718, new_n12082);
nand_5 g11697(new_n12082, n11158, new_n12083);
nor_5  g11698(new_n12083, new_n485, n13953);
nand_5 g11699(new_n1776_1, new_n547, new_n12085);
nand_5 g11700(new_n12085, new_n1782, new_n12086);
nand_5 g11701(new_n12086, new_n1614, new_n12087);
nand_5 g11702(new_n12087, new_n1611, new_n12088);
nand_5 g11703(new_n12088, new_n1789, new_n12089);
nand_5 g11704(new_n12089, new_n1608, new_n12090);
nand_5 g11705(new_n12090, new_n1605, new_n12091);
nand_5 g11706(new_n12091, new_n1795, new_n12092);
nand_5 g11707(new_n12092, new_n1799, new_n12093);
nand_5 g11708(new_n12093, new_n1602, new_n12094);
nand_5 g11709(new_n12094, new_n1599, new_n12095);
nand_5 g11710(new_n12095, new_n1596, new_n12096);
nand_5 g11711(new_n12096, new_n1593, new_n12097);
nand_5 g11712(new_n12097, new_n1806, new_n12098);
nand_5 g11713(new_n12098, new_n1589, new_n12099);
nand_5 g11714(new_n12099, new_n1586, new_n12100);
nand_5 g11715(new_n12100, new_n1583, new_n12101);
nand_5 g11716(new_n12101, new_n1580, new_n12102);
nand_5 g11717(new_n12102, new_n1576, new_n12103);
nand_5 g11718(new_n12103, new_n1573, new_n12104);
nand_5 g11719(new_n12104, new_n1570, new_n12105);
nand_5 g11720(new_n12105, new_n1567, new_n12106);
nand_5 g11721(new_n12106, new_n1564, new_n12107);
nand_5 g11722(new_n12107, new_n1561, new_n12108);
nand_5 g11723(new_n12108, new_n1338, new_n12109);
nand_5 g11724(new_n12109, new_n1331, new_n12110);
nand_5 g11725(new_n12110, new_n1326, new_n12111);
nand_5 g11726(new_n12111, new_n1321, new_n12112);
nand_5 g11727(new_n12112, new_n1318, new_n12113);
nand_5 g11728(new_n12113, new_n1315, new_n12114);
nand_5 g11729(new_n12114, new_n1312, new_n12115);
nand_5 g11730(new_n12115, new_n1309, new_n12116);
nand_5 g11731(new_n12116, new_n1307, new_n12117);
nand_5 g11732(new_n12117, new_n1304, new_n12118);
nand_5 g11733(new_n12118, new_n1300, new_n12119);
nand_5 g11734(new_n12119, new_n1297, new_n12120);
nand_5 g11735(new_n12120, new_n1294, new_n12121);
nand_5 g11736(new_n12121, new_n1355, new_n12122);
nand_5 g11737(new_n12122, new_n1291, new_n12123);
nand_5 g11738(new_n12123, new_n1288, new_n12124);
nand_5 g11739(new_n12124, new_n1283, new_n12125);
nand_5 g11740(new_n12125, new_n1363, new_n12126);
nand_5 g11741(new_n12126, new_n1280, new_n12127);
nand_5 g11742(new_n12127, new_n1370, new_n12128);
nand_5 g11743(new_n12128, new_n1373, new_n12129);
nand_5 g11744(new_n12129, new_n1277, new_n12130);
nand_5 g11745(new_n12130, new_n1272, new_n12131);
nand_5 g11746(new_n12131, new_n1269, new_n12132);
nand_5 g11747(new_n12132, new_n1380, new_n12133);
nand_5 g11748(new_n12133, new_n1264, new_n12134);
nand_5 g11749(new_n12134, new_n1259, new_n12135);
nand_5 g11750(new_n12135, new_n1388, new_n12136);
nand_5 g11751(new_n12136, new_n1392, new_n12137);
nand_5 g11752(new_n12137, new_n1256, new_n12138);
nand_5 g11753(new_n12138, new_n1252, new_n12139);
nand_5 g11754(new_n12139, new_n1249, new_n12140);
nand_5 g11755(new_n12140, new_n1244, new_n12141);
nand_5 g11756(new_n12141, new_n1240, new_n12142_1);
nand_5 g11757(new_n12142_1, new_n1234, new_n12143);
nand_5 g11758(new_n12143, new_n1231, new_n12144);
nand_5 g11759(new_n12144, new_n1227, new_n12145);
nand_5 g11760(new_n12145, new_n1407, new_n12146);
nand_5 g11761(new_n12146, new_n1223, new_n12147);
nand_5 g11762(new_n12147, new_n1218, new_n12148);
nand_5 g11763(new_n12148, new_n1213, new_n12149);
nand_5 g11764(new_n12149, new_n1210, new_n12150);
nand_5 g11765(new_n12150, new_n1206, new_n12151);
nand_5 g11766(new_n12151, new_n1418, new_n12152);
nand_5 g11767(new_n12152, new_n1422, new_n12153);
nand_5 g11768(new_n12153, new_n1428, new_n12154);
nand_5 g11769(new_n12154, new_n1203, new_n12155);
nand_5 g11770(new_n12155, new_n1433, new_n12156);
nand_5 g11771(new_n12156, new_n581, new_n12157);
nand_5 g11772(new_n12157, new_n574, new_n12158);
nand_5 g11773(new_n12158, new_n568, new_n12159);
nand_5 g11774(new_n12159, new_n589, new_n12160);
nand_5 g11775(new_n12160, new_n595, new_n12161);
nand_5 g11776(new_n12161, new_n601, new_n12162);
nand_5 g11777(new_n12162, new_n563, new_n12163);
nand_5 g11778(new_n12163, new_n608, new_n12164);
nand_5 g11779(new_n12164, new_n558, new_n12165);
nand_5 g11780(new_n12165, new_n615, new_n12166_1);
nand_5 g11781(new_n12166_1, new_n553, new_n12167);
nand_5 g11782(new_n12167, new_n622, new_n12168);
nand_5 g11783(new_n12168, n2334, new_n12169);
nor_5  g11784(new_n12169, new_n625, n13959);
not_4  g11785(new_n425, new_n12171);
nand_5 g11786(new_n1392, new_n12171, new_n12172);
nand_5 g11787(new_n12172, new_n1256, new_n12173);
nand_5 g11788(new_n12173, new_n1252, new_n12174);
nand_5 g11789(new_n12174, new_n1249, new_n12175);
nand_5 g11790(new_n12175, new_n1244, new_n12176);
nand_5 g11791(new_n12176, new_n1240, new_n12177);
nand_5 g11792(new_n12177, new_n1234, new_n12178);
nand_5 g11793(new_n12178, new_n1231, new_n12179);
nand_5 g11794(new_n12179, new_n1227, new_n12180);
nand_5 g11795(new_n12180, new_n1407, new_n12181);
nand_5 g11796(new_n12181, new_n1223, new_n12182);
nand_5 g11797(new_n12182, new_n1218, new_n12183);
nand_5 g11798(new_n12183, new_n1213, new_n12184);
nand_5 g11799(new_n12184, new_n1210, new_n12185);
nand_5 g11800(new_n12185, new_n1206, new_n12186);
nand_5 g11801(new_n12186, new_n1418, new_n12187);
nand_5 g11802(new_n12187, new_n1422, new_n12188);
nand_5 g11803(new_n12188, new_n1428, new_n12189);
nand_5 g11804(new_n12189, new_n1203, new_n12190);
nand_5 g11805(new_n12190, new_n1433, new_n12191);
nand_5 g11806(new_n12191, new_n581, new_n12192);
nand_5 g11807(new_n12192, new_n574, new_n12193);
nand_5 g11808(new_n12193, new_n568, new_n12194);
nand_5 g11809(new_n12194, new_n589, new_n12195);
nand_5 g11810(new_n12195, new_n595, new_n12196);
nand_5 g11811(new_n12196, new_n601, new_n12197);
nand_5 g11812(new_n12197, new_n563, new_n12198);
nand_5 g11813(new_n12198, new_n608, new_n12199);
nand_5 g11814(new_n12199, new_n558, new_n12200);
nand_5 g11815(new_n12200, new_n615, new_n12201);
nand_5 g11816(new_n12201, new_n553, new_n12202);
nand_5 g11817(new_n12202, new_n622, new_n12203);
nand_5 g11818(new_n12203, new_n628, new_n12204);
nand_5 g11819(new_n12204, new_n548, new_n12205);
nand_5 g11820(new_n12205, new_n543_1, new_n12206);
nand_5 g11821(new_n12206, new_n636, new_n12207);
nand_5 g11822(new_n12207, new_n642, new_n12208);
nand_5 g11823(new_n12208, new_n538, new_n12209);
nand_5 g11824(new_n12209, new_n533, new_n12210);
nand_5 g11825(new_n12210, new_n650_1, new_n12211);
nand_5 g11826(new_n12211, new_n528, new_n12212);
nand_5 g11827(new_n12212, new_n523, new_n12213);
nand_5 g11828(new_n12213, new_n518, new_n12214);
nand_5 g11829(new_n12214, new_n659, new_n12215);
nand_5 g11830(new_n12215, new_n665, new_n12216);
nand_5 g11831(new_n12216, new_n672, new_n12217);
nand_5 g11832(new_n12217, new_n513, new_n12218_1);
nand_5 g11833(new_n12218_1, new_n679, new_n12219);
nand_5 g11834(new_n12219, new_n685, new_n12220);
nand_5 g11835(new_n12220, new_n691, new_n12221);
nand_5 g11836(new_n12221, new_n508, new_n12222);
nand_5 g11837(new_n12222, new_n698, new_n12223);
nand_5 g11838(new_n12223, new_n503, new_n12224);
nand_5 g11839(new_n12224, new_n704, new_n12225);
nand_5 g11840(new_n12225, new_n498_1, new_n12226);
nand_5 g11841(new_n12226, new_n711, new_n12227);
nand_5 g11842(new_n12227, new_n493, new_n12228);
nand_5 g11843(new_n12228, new_n718, new_n12229);
nand_5 g11844(new_n12229, new_n488, new_n12230);
nand_5 g11845(new_n12230, new_n725, new_n12231);
nand_5 g11846(new_n12231, new_n483, new_n12232_1);
nand_5 g11847(new_n12232_1, new_n732, new_n12233);
nand_5 g11848(new_n12233, new_n478, new_n12234);
nand_5 g11849(new_n12234, new_n739, new_n12235);
nand_5 g11850(new_n12235, new_n745, new_n12236);
nand_5 g11851(new_n12236, new_n751, new_n12237);
nand_5 g11852(new_n12237, new_n473, new_n12238);
nand_5 g11853(new_n12238, new_n758, new_n12239);
nand_5 g11854(new_n12239, new_n764, new_n12240);
nand_5 g11855(new_n12240, new_n770, new_n12241);
nand_5 g11856(new_n12241, new_n468, new_n12242);
nand_5 g11857(new_n12242, new_n777, new_n12243);
nand_5 g11858(new_n12243, new_n783, new_n12244);
nand_5 g11859(new_n12244, new_n789, new_n12245);
nand_5 g11860(new_n12245, new_n463, new_n12246);
nand_5 g11861(new_n12246, new_n796, new_n12247);
nand_5 g11862(new_n12247, new_n458, new_n12248);
nand_5 g11863(new_n12248, new_n453, new_n12249);
nand_5 g11864(new_n12249, new_n447, new_n12250);
nand_5 g11865(new_n12250, new_n805, new_n12251);
nand_5 g11866(new_n12251, new_n811, new_n12252);
nand_5 g11867(new_n12252, new_n442, new_n12253);
nand_5 g11868(new_n12253, new_n437, new_n12254);
nand_5 g11869(new_n12254, new_n819, new_n12255);
nand_5 g11870(new_n12255, n14303, new_n12256);
nor_5  g11871(new_n12256, new_n429, n14289);
nand_5 g11872(new_n2037, new_n1369, new_n12258);
nand_5 g11873(new_n12258, new_n2036, new_n12259);
nand_5 g11874(new_n12259, new_n2033, new_n12260);
nand_5 g11875(new_n12260, new_n2029, new_n12261);
nand_5 g11876(new_n12261, new_n2026, new_n12262);
nand_5 g11877(new_n12262, new_n2022, new_n12263);
nand_5 g11878(new_n12263, new_n2018, new_n12264);
nand_5 g11879(new_n12264, new_n1726, new_n12265);
nand_5 g11880(new_n12265, new_n1722, new_n12266);
nand_5 g11881(new_n12266, new_n1718, new_n12267);
nand_5 g11882(new_n12267, new_n1713, new_n12268);
nand_5 g11883(new_n12268, new_n1737, new_n12269);
nand_5 g11884(new_n12269, new_n1709, new_n12270_1);
nand_5 g11885(new_n12270_1, new_n1742, new_n12271);
nand_5 g11886(new_n12271, new_n1704, new_n12272);
nand_5 g11887(new_n12272, new_n1702_1, new_n12273);
nand_5 g11888(new_n12273, new_n1698, new_n12274);
nand_5 g11889(new_n12274, new_n1695, new_n12275);
nand_5 g11890(new_n12275, new_n1692, new_n12276);
nand_5 g11891(new_n12276, new_n1752, new_n12277);
nand_5 g11892(new_n12277, new_n1688, new_n12278);
nand_5 g11893(new_n12278, new_n1685, new_n12279);
nand_5 g11894(new_n12279, new_n1680, new_n12280);
nand_5 g11895(new_n12280, new_n1676, new_n12281);
nand_5 g11896(new_n12281, new_n1672, new_n12282);
nand_5 g11897(new_n12282, new_n1669, new_n12283);
nand_5 g11898(new_n12283, new_n1666, new_n12284);
nand_5 g11899(new_n12284, new_n1663, new_n12285);
nand_5 g11900(new_n12285, new_n1658, new_n12286);
nand_5 g11901(new_n12286, new_n1653, new_n12287);
nand_5 g11902(new_n12287, new_n1651, new_n12288);
nand_5 g11903(new_n12288, new_n1649, new_n12289);
nand_5 g11904(new_n12289, new_n1646, new_n12290);
nand_5 g11905(new_n12290, new_n1643, new_n12291);
nand_5 g11906(new_n12291, new_n1641, new_n12292);
nand_5 g11907(new_n12292, new_n1638, new_n12293);
nand_5 g11908(new_n12293, new_n1635, new_n12294);
nand_5 g11909(new_n12294, new_n1632, new_n12295);
nand_5 g11910(new_n12295, new_n1628, new_n12296);
nand_5 g11911(new_n12296, new_n1625, new_n12297);
nand_5 g11912(new_n12297, new_n1621, new_n12298);
nand_5 g11913(new_n12298, new_n1618, new_n12299);
nand_5 g11914(new_n12299, new_n1778, new_n12300);
nand_5 g11915(new_n12300, new_n1782, new_n12301);
nand_5 g11916(new_n12301, new_n1614, new_n12302);
nand_5 g11917(new_n12302, new_n1611, new_n12303);
nand_5 g11918(new_n12303, new_n1789, new_n12304);
nand_5 g11919(new_n12304, new_n1608, new_n12305);
nand_5 g11920(new_n12305, new_n1605, new_n12306);
nand_5 g11921(new_n12306, new_n1795, new_n12307);
nand_5 g11922(new_n12307, new_n1799, new_n12308);
nand_5 g11923(new_n12308, new_n1602, new_n12309);
nand_5 g11924(new_n12309, new_n1599, new_n12310);
nand_5 g11925(new_n12310, new_n1596, new_n12311);
nand_5 g11926(new_n12311, new_n1593, new_n12312);
nand_5 g11927(new_n12312, new_n1806, new_n12313);
nand_5 g11928(new_n12313, new_n1589, new_n12314);
nand_5 g11929(new_n12314, new_n1586, new_n12315);
nand_5 g11930(new_n12315, new_n1583, new_n12316);
nand_5 g11931(new_n12316, new_n1580, new_n12317);
nand_5 g11932(new_n12317, new_n1576, new_n12318);
nand_5 g11933(new_n12318, new_n1573, new_n12319);
nand_5 g11934(new_n12319, new_n1570, new_n12320);
nand_5 g11935(new_n12320, new_n1567, new_n12321_1);
nand_5 g11936(new_n12321_1, new_n1564, new_n12322);
nand_5 g11937(new_n12322, new_n1561, new_n12323);
nand_5 g11938(new_n12323, new_n1338, new_n12324);
nand_5 g11939(new_n12324, new_n1331, new_n12325);
nand_5 g11940(new_n12325, new_n1326, new_n12326);
nand_5 g11941(new_n12326, new_n1321, new_n12327);
nand_5 g11942(new_n12327, new_n1318, new_n12328);
nand_5 g11943(new_n12328, new_n1315, new_n12329);
nand_5 g11944(new_n12329, new_n1312, new_n12330);
nand_5 g11945(new_n12330, new_n1309, new_n12331);
nand_5 g11946(new_n12331, new_n1307, new_n12332);
nand_5 g11947(new_n12332, new_n1304, new_n12333);
nand_5 g11948(new_n12333, new_n1300, new_n12334);
nand_5 g11949(new_n12334, new_n1297, new_n12335);
nand_5 g11950(new_n12335, new_n1294, new_n12336_1);
nand_5 g11951(new_n12336_1, new_n1355, new_n12337);
nand_5 g11952(new_n12337, new_n1291, new_n12338);
nand_5 g11953(new_n12338, new_n1288, new_n12339);
nand_5 g11954(new_n12339, new_n1283, new_n12340);
nand_5 g11955(new_n12340, new_n1363, new_n12341);
nand_5 g11956(new_n12341, n6480, new_n12342);
nor_5  g11957(new_n12342, new_n793, n14307);
nand_5 g11958(new_n1020, new_n526, new_n12344);
nand_5 g11959(new_n12344, new_n523, new_n12345);
nand_5 g11960(new_n12345, new_n518, new_n12346);
nand_5 g11961(new_n12346, new_n659, new_n12347);
nand_5 g11962(new_n12347, new_n665, new_n12348);
nand_5 g11963(new_n12348, new_n672, new_n12349);
nand_5 g11964(new_n12349, new_n513, new_n12350);
nand_5 g11965(new_n12350, new_n679, new_n12351);
nand_5 g11966(new_n12351, new_n685, new_n12352);
nand_5 g11967(new_n12352, new_n691, new_n12353);
nand_5 g11968(new_n12353, new_n508, new_n12354);
nand_5 g11969(new_n12354, new_n698, new_n12355_1);
nand_5 g11970(new_n12355_1, new_n503, new_n12356);
nand_5 g11971(new_n12356, new_n704, new_n12357);
nand_5 g11972(new_n12357, new_n498_1, new_n12358);
nand_5 g11973(new_n12358, new_n711, new_n12359);
nand_5 g11974(new_n12359, new_n493, new_n12360);
nand_5 g11975(new_n12360, new_n718, new_n12361);
nand_5 g11976(new_n12361, new_n488, new_n12362);
nand_5 g11977(new_n12362, new_n725, new_n12363);
nand_5 g11978(new_n12363, new_n483, new_n12364);
nand_5 g11979(new_n12364, new_n732, new_n12365);
nand_5 g11980(new_n12365, new_n478, new_n12366);
nand_5 g11981(new_n12366, new_n739, new_n12367);
nand_5 g11982(new_n12367, new_n745, new_n12368);
nand_5 g11983(new_n12368, new_n751, new_n12369);
nand_5 g11984(new_n12369, new_n473, new_n12370);
nand_5 g11985(new_n12370, new_n758, new_n12371);
nand_5 g11986(new_n12371, new_n764, new_n12372);
nand_5 g11987(new_n12372, new_n770, new_n12373);
nand_5 g11988(new_n12373, new_n468, new_n12374);
nand_5 g11989(new_n12374, new_n777, new_n12375);
nand_5 g11990(new_n12375, new_n783, new_n12376);
nand_5 g11991(new_n12376, new_n789, new_n12377);
nand_5 g11992(new_n12377, new_n463, new_n12378);
nand_5 g11993(new_n12378, new_n796, new_n12379);
nand_5 g11994(new_n12379, new_n458, new_n12380);
nand_5 g11995(new_n12380, new_n453, new_n12381);
nand_5 g11996(new_n12381, new_n447, new_n12382);
nand_5 g11997(new_n12382, new_n805, new_n12383);
nand_5 g11998(new_n12383, new_n811, new_n12384);
nand_5 g11999(new_n12384, new_n442, new_n12385);
nand_5 g12000(new_n12385, new_n437, new_n12386);
nand_5 g12001(new_n12386, new_n819, new_n12387);
nand_5 g12002(new_n12387, new_n432, new_n12388);
nand_5 g12003(new_n12388, new_n427_1, new_n12389);
nand_5 g12004(new_n12389, new_n422, new_n12390);
nand_5 g12005(new_n12390, new_n828, new_n12391);
nand_5 g12006(new_n12391, new_n834, new_n12392);
nand_5 g12007(new_n12392, new_n840, new_n12393);
nand_5 g12008(new_n12393, new_n417, new_n12394);
nand_5 g12009(new_n12394, new_n847, new_n12395);
nand_5 g12010(new_n12395, new_n853, new_n12396);
nand_5 g12011(new_n12396, new_n859, new_n12397);
nand_5 g12012(new_n12397, new_n412, new_n12398);
nand_5 g12013(new_n12398, new_n866, new_n12399);
nand_5 g12014(new_n12399, new_n872, new_n12400);
nand_5 g12015(new_n12400, new_n878, new_n12401);
nand_5 g12016(new_n12401, new_n407, new_n12402);
nand_5 g12017(new_n12402, new_n885, new_n12403);
nand_5 g12018(new_n12403, new_n402, new_n12404);
nand_5 g12019(new_n12404, new_n397, new_n12405);
nand_5 g12020(new_n12405, new_n392, new_n12406);
nand_5 g12021(new_n12406, new_n894, new_n12407);
nand_5 g12022(new_n12407, new_n1087, new_n12408);
nand_5 g12023(new_n12408, new_n1129, new_n12409);
nand_5 g12024(new_n12409, new_n1084, new_n12410);
nand_5 g12025(new_n12410, new_n1134, new_n12411);
nand_5 g12026(new_n12411, new_n1080, new_n12412);
nand_5 g12027(new_n12412, new_n1075, new_n12413);
nand_5 g12028(new_n12413, new_n1070, new_n12414);
nand_5 g12029(new_n12414, new_n1143, new_n12415);
nand_5 g12030(new_n12415, new_n1148, new_n12416);
nand_5 g12031(new_n12416, new_n1065, new_n12417);
nand_5 g12032(new_n12417, new_n1062, new_n12418);
nand_5 g12033(new_n12418, new_n1156, new_n12419);
nand_5 g12034(new_n12419, new_n1057, new_n12420);
nand_5 g12035(new_n12420, new_n1053, new_n12421);
nand_5 g12036(new_n12421, new_n1050, new_n12422);
nand_5 g12037(new_n12422, new_n1045, new_n12423);
nand_5 g12038(new_n12423, new_n1040, new_n12424);
nand_5 g12039(new_n12424, new_n1036, new_n12425);
nand_5 g12040(new_n12425, new_n1033, new_n12426);
nand_5 g12041(new_n12426, new_n1028, new_n12427);
nand_5 g12042(new_n12427, n5725, new_n12428);
nor_5  g12043(new_n12428, new_n1023, n14330);
nand_5 g12044(new_n668, new_n513, new_n12430);
nand_5 g12045(new_n12430, new_n679, new_n12431);
nand_5 g12046(new_n12431, new_n685, new_n12432);
nand_5 g12047(new_n12432, new_n691, new_n12433);
nand_5 g12048(new_n12433, new_n508, new_n12434);
nand_5 g12049(new_n12434, new_n698, new_n12435);
nand_5 g12050(new_n12435, new_n503, new_n12436);
nand_5 g12051(new_n12436, new_n704, new_n12437);
nand_5 g12052(new_n12437, new_n498_1, new_n12438);
nand_5 g12053(new_n12438, new_n711, new_n12439);
nand_5 g12054(new_n12439, new_n493, new_n12440);
nand_5 g12055(new_n12440, new_n718, new_n12441);
nand_5 g12056(new_n12441, new_n488, new_n12442);
nand_5 g12057(new_n12442, new_n725, new_n12443);
nand_5 g12058(new_n12443, new_n483, new_n12444);
nand_5 g12059(new_n12444, new_n732, new_n12445);
nand_5 g12060(new_n12445, new_n478, new_n12446);
nand_5 g12061(new_n12446, new_n739, new_n12447);
nand_5 g12062(new_n12447, new_n745, new_n12448);
nand_5 g12063(new_n12448, new_n751, new_n12449);
nand_5 g12064(new_n12449, new_n473, new_n12450);
nand_5 g12065(new_n12450, new_n758, new_n12451);
nand_5 g12066(new_n12451, new_n764, new_n12452);
nand_5 g12067(new_n12452, new_n770, new_n12453);
nand_5 g12068(new_n12453, new_n468, new_n12454);
nand_5 g12069(new_n12454, new_n777, new_n12455);
nand_5 g12070(new_n12455, new_n783, new_n12456);
nand_5 g12071(new_n12456, new_n789, new_n12457);
nand_5 g12072(new_n12457, new_n463, new_n12458);
nand_5 g12073(new_n12458, new_n796, new_n12459);
nand_5 g12074(new_n12459, new_n458, new_n12460);
nand_5 g12075(new_n12460, new_n453, new_n12461);
nand_5 g12076(new_n12461, new_n447, new_n12462);
nand_5 g12077(new_n12462, new_n805, new_n12463);
nand_5 g12078(new_n12463, new_n811, new_n12464);
nand_5 g12079(new_n12464, new_n442, new_n12465);
nand_5 g12080(new_n12465, new_n437, new_n12466);
nand_5 g12081(new_n12466, new_n819, new_n12467);
nand_5 g12082(new_n12467, new_n432, new_n12468);
nand_5 g12083(new_n12468, new_n427_1, new_n12469);
nand_5 g12084(new_n12469, new_n422, new_n12470);
nand_5 g12085(new_n12470, new_n828, new_n12471);
nand_5 g12086(new_n12471, new_n834, new_n12472);
nand_5 g12087(new_n12472, new_n840, new_n12473);
nand_5 g12088(new_n12473, new_n417, new_n12474);
nand_5 g12089(new_n12474, new_n847, new_n12475);
nand_5 g12090(new_n12475, new_n853, new_n12476);
nand_5 g12091(new_n12476, new_n859, new_n12477);
nand_5 g12092(new_n12477, new_n412, new_n12478);
nand_5 g12093(new_n12478, new_n866, new_n12479);
nand_5 g12094(new_n12479, new_n872, new_n12480);
nand_5 g12095(new_n12480, new_n878, new_n12481);
nand_5 g12096(new_n12481, new_n407, new_n12482);
nand_5 g12097(new_n12482, new_n885, new_n12483);
nand_5 g12098(new_n12483, new_n402, new_n12484);
nand_5 g12099(new_n12484, new_n397, new_n12485);
nand_5 g12100(new_n12485, new_n392, new_n12486);
nand_5 g12101(new_n12486, new_n894, new_n12487);
nand_5 g12102(new_n12487, new_n1087, new_n12488);
nand_5 g12103(new_n12488, new_n1129, new_n12489);
nand_5 g12104(new_n12489, new_n1084, new_n12490);
nand_5 g12105(new_n12490, new_n1134, new_n12491);
nand_5 g12106(new_n12491, new_n1080, new_n12492);
nand_5 g12107(new_n12492, new_n1075, new_n12493);
nand_5 g12108(new_n12493, new_n1070, new_n12494);
nand_5 g12109(new_n12494, new_n1143, new_n12495);
nand_5 g12110(new_n12495, new_n1148, new_n12496);
nand_5 g12111(new_n12496, new_n1065, new_n12497);
nand_5 g12112(new_n12497, new_n1062, new_n12498);
nand_5 g12113(new_n12498, new_n1156, new_n12499);
nand_5 g12114(new_n12499, new_n1057, new_n12500);
nand_5 g12115(new_n12500, new_n1053, new_n12501);
nand_5 g12116(new_n12501, new_n1050, new_n12502);
nand_5 g12117(new_n12502, new_n1045, new_n12503);
nand_5 g12118(new_n12503, new_n1040, new_n12504);
nand_5 g12119(new_n12504, new_n1036, new_n12505);
nand_5 g12120(new_n12505, new_n1033, new_n12506);
nand_5 g12121(new_n12506, new_n1028, new_n12507);
nand_5 g12122(new_n12507, new_n1026, new_n12508);
nand_5 g12123(new_n12508, new_n1021, new_n12509);
nand_5 g12124(new_n12509, new_n1017, new_n12510);
nand_5 g12125(new_n12510, new_n1012, new_n12511);
nand_5 g12126(new_n12511, new_n1009, new_n12512);
nand_5 g12127(new_n12512, new_n1004, new_n12513);
nand_5 g12128(new_n12513, n10765, new_n12514);
nor_5  g12129(new_n12514, new_n997, n14399);
not_4  g12130(new_n634, new_n12516);
nand_5 g12131(new_n1614, new_n12516, new_n12517);
nand_5 g12132(new_n12517, new_n1611, new_n12518);
nand_5 g12133(new_n12518, new_n1789, new_n12519);
nand_5 g12134(new_n12519, new_n1608, new_n12520);
nand_5 g12135(new_n12520, new_n1605, new_n12521);
nand_5 g12136(new_n12521, new_n1795, new_n12522);
nand_5 g12137(new_n12522, new_n1799, new_n12523);
nand_5 g12138(new_n12523, new_n1602, new_n12524);
nand_5 g12139(new_n12524, new_n1599, new_n12525);
nand_5 g12140(new_n12525, new_n1596, new_n12526);
nand_5 g12141(new_n12526, new_n1593, new_n12527);
nand_5 g12142(new_n12527, new_n1806, new_n12528);
nand_5 g12143(new_n12528, new_n1589, new_n12529);
nand_5 g12144(new_n12529, new_n1586, new_n12530);
nand_5 g12145(new_n12530, new_n1583, new_n12531);
nand_5 g12146(new_n12531, new_n1580, new_n12532);
nand_5 g12147(new_n12532, new_n1576, new_n12533);
nand_5 g12148(new_n12533, new_n1573, new_n12534);
nand_5 g12149(new_n12534, new_n1570, new_n12535_1);
nand_5 g12150(new_n12535_1, new_n1567, new_n12536);
nand_5 g12151(new_n12536, new_n1564, new_n12537);
nand_5 g12152(new_n12537, new_n1561, new_n12538);
nand_5 g12153(new_n12538, new_n1338, new_n12539);
nand_5 g12154(new_n12539, new_n1331, new_n12540);
nand_5 g12155(new_n12540, new_n1326, new_n12541);
nand_5 g12156(new_n12541, new_n1321, new_n12542);
nand_5 g12157(new_n12542, new_n1318, new_n12543);
nand_5 g12158(new_n12543, new_n1315, new_n12544);
nand_5 g12159(new_n12544, new_n1312, new_n12545);
nand_5 g12160(new_n12545, new_n1309, new_n12546);
nand_5 g12161(new_n12546, new_n1307, new_n12547);
nand_5 g12162(new_n12547, new_n1304, new_n12548);
nand_5 g12163(new_n12548, new_n1300, new_n12549);
nand_5 g12164(new_n12549, new_n1297, new_n12550);
nand_5 g12165(new_n12550, new_n1294, new_n12551);
nand_5 g12166(new_n12551, new_n1355, new_n12552);
nand_5 g12167(new_n12552, new_n1291, new_n12553);
nand_5 g12168(new_n12553, new_n1288, new_n12554);
nand_5 g12169(new_n12554, new_n1283, new_n12555);
nand_5 g12170(new_n12555, new_n1363, new_n12556);
nand_5 g12171(new_n12556, new_n1280, new_n12557);
nand_5 g12172(new_n12557, new_n1370, new_n12558);
nand_5 g12173(new_n12558, new_n1373, new_n12559);
nand_5 g12174(new_n12559, new_n1277, new_n12560);
nand_5 g12175(new_n12560, new_n1272, new_n12561);
nand_5 g12176(new_n12561, new_n1269, new_n12562);
nand_5 g12177(new_n12562, new_n1380, new_n12563);
nand_5 g12178(new_n12563, new_n1264, new_n12564);
nand_5 g12179(new_n12564, new_n1259, new_n12565);
nand_5 g12180(new_n12565, new_n1388, new_n12566);
nand_5 g12181(new_n12566, new_n1392, new_n12567);
nand_5 g12182(new_n12567, new_n1256, new_n12568);
nand_5 g12183(new_n12568, new_n1252, new_n12569);
nand_5 g12184(new_n12569, new_n1249, new_n12570);
nand_5 g12185(new_n12570, new_n1244, new_n12571);
nand_5 g12186(new_n12571, new_n1240, new_n12572);
nand_5 g12187(new_n12572, new_n1234, new_n12573_1);
nand_5 g12188(new_n12573_1, new_n1231, new_n12574);
nand_5 g12189(new_n12574, new_n1227, new_n12575);
nand_5 g12190(new_n12575, new_n1407, new_n12576);
nand_5 g12191(new_n12576, new_n1223, new_n12577);
nand_5 g12192(new_n12577, new_n1218, new_n12578);
nand_5 g12193(new_n12578, new_n1213, new_n12579);
nand_5 g12194(new_n12579, new_n1210, new_n12580);
nand_5 g12195(new_n12580, new_n1206, new_n12581);
nand_5 g12196(new_n12581, new_n1418, new_n12582);
nand_5 g12197(new_n12582, new_n1422, new_n12583);
nand_5 g12198(new_n12583, new_n1428, new_n12584);
nand_5 g12199(new_n12584, new_n1203, new_n12585);
nand_5 g12200(new_n12585, new_n1433, new_n12586);
nand_5 g12201(new_n12586, new_n581, new_n12587);
nand_5 g12202(new_n12587, new_n574, new_n12588);
nand_5 g12203(new_n12588, new_n568, new_n12589);
nand_5 g12204(new_n12589, new_n589, new_n12590);
nand_5 g12205(new_n12590, new_n595, new_n12591);
nand_5 g12206(new_n12591, new_n601, new_n12592);
nand_5 g12207(new_n12592, new_n563, new_n12593);
nand_5 g12208(new_n12593, new_n608, new_n12594);
nand_5 g12209(new_n12594, new_n558, new_n12595);
nand_5 g12210(new_n12595, new_n615, new_n12596);
nand_5 g12211(new_n12596, new_n553, new_n12597);
nand_5 g12212(new_n12597, new_n622, new_n12598);
nand_5 g12213(new_n12598, new_n628, new_n12599);
nand_5 g12214(new_n12599, new_n548, new_n12600);
nand_5 g12215(new_n12600, n11776, new_n12601);
nor_5  g12216(new_n12601, new_n540, n14463);
endmodule


