// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Thu Jun 27 14:29:42 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2528, new_n2529, new_n2530,
    new_n2531, new_n2533_1, new_n2534, new_n2535_1, new_n2536, new_n2537_1,
    new_n2538, new_n2539, new_n2540, new_n2541, new_n2542, new_n2543,
    new_n2544, new_n2545, new_n2546, new_n2547_1, new_n2548, new_n2549,
    new_n2550, new_n2551, new_n2552, new_n2553_1, new_n2554, new_n2555_1,
    new_n2556, new_n2557, new_n2558, new_n2559, new_n2560_1, new_n2561_1,
    new_n2562, new_n2563, new_n2564, new_n2565, new_n2566, new_n2567,
    new_n2568, new_n2569, new_n2570_1, new_n2571, new_n2572, new_n2573_1,
    new_n2574, new_n2575, new_n2576, new_n2577, new_n2578_1, new_n2579,
    new_n2580, new_n2581, new_n2582_1, new_n2583, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602_1, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619_1, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772,
    new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777, new_n2778,
    new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1, new_n2784,
    new_n2785, new_n2786, new_n2787, new_n2788, new_n2789, new_n2790,
    new_n2791, new_n2792, new_n2793, new_n2794, new_n2795, new_n2796,
    new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802,
    new_n2803, new_n2804, new_n2805, new_n2806, new_n2807, new_n2808,
    new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813, new_n2814,
    new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819, new_n2820,
    new_n2821, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826_1,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886_1,
    new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945, new_n2946,
    new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2967, new_n2968, new_n2969, new_n2970, new_n2971_1,
    new_n2972, new_n2973, new_n2974, new_n2975, new_n2976, new_n2977,
    new_n2978_1, new_n2979_1, new_n2980, new_n2981, new_n2982, new_n2983,
    new_n2984, new_n2985_1, new_n2986, new_n2987, new_n2988, new_n2989,
    new_n2990, new_n2991, new_n2992, new_n2993, new_n2994, new_n2995,
    new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000, new_n3001,
    new_n3002, new_n3003, new_n3004, new_n3005, new_n3006, new_n3007,
    new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012, new_n3013,
    new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1, new_n3019,
    new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024, new_n3025,
    new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1, new_n3031,
    new_n3032, new_n3033, new_n3034, new_n3035, new_n3036, new_n3037,
    new_n3038, new_n3039, new_n3040, new_n3041, new_n3042, new_n3043,
    new_n3044, new_n3045, new_n3046, new_n3047, new_n3048, new_n3049,
    new_n3050, new_n3051, new_n3052, new_n3053, new_n3054, new_n3055,
    new_n3056, new_n3057, new_n3058, new_n3059, new_n3060, new_n3061,
    new_n3062, new_n3063, new_n3064, new_n3065, new_n3066, new_n3067_1,
    new_n3068, new_n3069, new_n3070, new_n3071, new_n3072, new_n3073,
    new_n3074, new_n3075, new_n3076_1, new_n3077, new_n3078, new_n3079,
    new_n3080, new_n3081, new_n3082, new_n3083, new_n3084, new_n3085,
    new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090, new_n3091,
    new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097,
    new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3162, new_n3163,
    new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235_1,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3252, new_n3253_1, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260_1,
    new_n3261, new_n3262, new_n3263_1, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279_1, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287, new_n3288, new_n3289_1, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301_1, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306_1, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319, new_n3320_1,
    new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332_1,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505, new_n3506_1,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528_1, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541_1, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555_1,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561_1,
    new_n3562, new_n3563_1, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570_1, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582_1, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616, new_n3617_1, new_n3618_1, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642_1, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649_1, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661, new_n3662, new_n3663,
    new_n3664, new_n3665_1, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677, new_n3678, new_n3679_1, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710_1, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725_1, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733_1, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740_1, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755_1, new_n3756, new_n3757, new_n3758_1, new_n3759, new_n3760_1,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781_1, new_n3782, new_n3783, new_n3784,
    new_n3785_1, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794_1, new_n3795_1, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828_1, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3842_1, new_n3843, new_n3844, new_n3845,
    new_n3846, new_n3847, new_n3848, new_n3849, new_n3850_1, new_n3851,
    new_n3852, new_n3853, new_n3854, new_n3855, new_n3856, new_n3857,
    new_n3858, new_n3859, new_n3860, new_n3861, new_n3862, new_n3863,
    new_n3864, new_n3865, new_n3866, new_n3867, new_n3868, new_n3869_1,
    new_n3870, new_n3871_1, new_n3872, new_n3873, new_n3874, new_n3875,
    new_n3876, new_n3877, new_n3878, new_n3879, new_n3880, new_n3881,
    new_n3882, new_n3883, new_n3884, new_n3885, new_n3886, new_n3887,
    new_n3888, new_n3890, new_n3891_1, new_n3892, new_n3893, new_n3894,
    new_n3895, new_n3896, new_n3897, new_n3898, new_n3899, new_n3900,
    new_n3901, new_n3902, new_n3903, new_n3904, new_n3905, new_n3906,
    new_n3907, new_n3908, new_n3909_1, new_n3910, new_n3911, new_n3912,
    new_n3913, new_n3914, new_n3915, new_n3916, new_n3917, new_n3918_1,
    new_n3919, new_n3920, new_n3921, new_n3922, new_n3923, new_n3924,
    new_n3925_1, new_n3926, new_n3927, new_n3928, new_n3929, new_n3930,
    new_n3931, new_n3932_1, new_n3933, new_n3934_1, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945_1, new_n3946, new_n3947, new_n3948,
    new_n3949, new_n3950, new_n3951, new_n3952_1, new_n3953, new_n3954,
    new_n3955, new_n3956, new_n3957, new_n3958, new_n3959_1, new_n3960,
    new_n3961, new_n3962_1, new_n3963, new_n3964, new_n3965, new_n3966,
    new_n3967, new_n3968, new_n3969, new_n3970, new_n3971_1, new_n3972,
    new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978,
    new_n3979, new_n3980, new_n3981, new_n3982, new_n3983_1, new_n3984_1,
    new_n3985, new_n3986, new_n3987, new_n3988, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000_1, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4006, new_n4007, new_n4008, new_n4009,
    new_n4010_1, new_n4011, new_n4012, new_n4013, new_n4014_1, new_n4015,
    new_n4016, new_n4017, new_n4018, new_n4019, new_n4020, new_n4021,
    new_n4022, new_n4023, new_n4024, new_n4025, new_n4026, new_n4027,
    new_n4028, new_n4029, new_n4030, new_n4031, new_n4032, new_n4033,
    new_n4034, new_n4035, new_n4036, new_n4037, new_n4038, new_n4039,
    new_n4040, new_n4041, new_n4042, new_n4043, new_n4044, new_n4045,
    new_n4046, new_n4047, new_n4048, new_n4049, new_n4050, new_n4051,
    new_n4052, new_n4053, new_n4054, new_n4055, new_n4056, new_n4057,
    new_n4058, new_n4059, new_n4060, new_n4061, new_n4062, new_n4063,
    new_n4064, new_n4065, new_n4066, new_n4067, new_n4068, new_n4069,
    new_n4070, new_n4071_1, new_n4072, new_n4073, new_n4074, new_n4075,
    new_n4076, new_n4077, new_n4078, new_n4079, new_n4080, new_n4081,
    new_n4082, new_n4083, new_n4084, new_n4085_1, new_n4086, new_n4087,
    new_n4088_1, new_n4089_1, new_n4090, new_n4091, new_n4092, new_n4093,
    new_n4094, new_n4095, new_n4096, new_n4097, new_n4098, new_n4099,
    new_n4100_1, new_n4101, new_n4102, new_n4103_1, new_n4104, new_n4105,
    new_n4106, new_n4107, new_n4108, new_n4109, new_n4110, new_n4111,
    new_n4112, new_n4113, new_n4114, new_n4115, new_n4116, new_n4117,
    new_n4118, new_n4119_1, new_n4120, new_n4121, new_n4122, new_n4123_1,
    new_n4124, new_n4125, new_n4126, new_n4127, new_n4128, new_n4129,
    new_n4130, new_n4131, new_n4132, new_n4133, new_n4134_1, new_n4135,
    new_n4136, new_n4137, new_n4138, new_n4139, new_n4140, new_n4141,
    new_n4142, new_n4143, new_n4144, new_n4145, new_n4146_1, new_n4147,
    new_n4148, new_n4149, new_n4150_1, new_n4151_1, new_n4152_1,
    new_n4153_1, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165_1, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172_1, new_n4173_1, new_n4174, new_n4175, new_n4176_1,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186_1, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204_1, new_n4205_1, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215_1, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221_1, new_n4222, new_n4223, new_n4224_1,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231_1, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256_1, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266_1,
    new_n4268, new_n4269, new_n4270, new_n4271, new_n4272_1, new_n4273,
    new_n4274, new_n4275, new_n4276, new_n4277, new_n4278, new_n4279,
    new_n4280, new_n4281, new_n4282, new_n4283, new_n4284, new_n4285,
    new_n4286, new_n4287, new_n4288, new_n4289, new_n4290, new_n4291,
    new_n4292, new_n4293, new_n4294, new_n4295, new_n4296, new_n4297,
    new_n4298, new_n4299, new_n4300, new_n4301, new_n4302, new_n4303,
    new_n4304, new_n4305, new_n4306_1, new_n4307, new_n4308, new_n4309,
    new_n4310, new_n4311, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319_1, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325_1, new_n4326_1, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340_1, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374_1, new_n4375,
    new_n4376_1, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401_1, new_n4402, new_n4404, new_n4405, new_n4406,
    new_n4407, new_n4408, new_n4409_1, new_n4410, new_n4411, new_n4412,
    new_n4413, new_n4414, new_n4415, new_n4416, new_n4417, new_n4418,
    new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424_1,
    new_n4425, new_n4426_1, new_n4427, new_n4428, new_n4429, new_n4430,
    new_n4431, new_n4432_1, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437, new_n4438, new_n4439, new_n4440, new_n4441_1, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451_1, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476_1, new_n4477, new_n4478_1,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514_1,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529_1, new_n4530, new_n4531, new_n4532,
    new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538,
    new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544,
    new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550,
    new_n4551, new_n4552_1, new_n4553, new_n4554, new_n4555, new_n4556,
    new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562,
    new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568,
    new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574,
    new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4587, new_n4588_1, new_n4589, new_n4590_1, new_n4591, new_n4592,
    new_n4593, new_n4594, new_n4595_1, new_n4596, new_n4597, new_n4598,
    new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604,
    new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610,
    new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624_1, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646_1,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665_1,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674_1, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689,
    new_n4690, new_n4691, new_n4692, new_n4693_1, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4703, new_n4704, new_n4705, new_n4706, new_n4707, new_n4708,
    new_n4709, new_n4710, new_n4711, new_n4712, new_n4713, new_n4714,
    new_n4715, new_n4716, new_n4717, new_n4718, new_n4719, new_n4720,
    new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725, new_n4726,
    new_n4727, new_n4728, new_n4729, new_n4730, new_n4731_1, new_n4732,
    new_n4733, new_n4734, new_n4735, new_n4736, new_n4737, new_n4738,
    new_n4739, new_n4740, new_n4741, new_n4742, new_n4743, new_n4744,
    new_n4745_1, new_n4746, new_n4747_1, new_n4748, new_n4749, new_n4750,
    new_n4751, new_n4752, new_n4753, new_n4754, new_n4755, new_n4756,
    new_n4757, new_n4758, new_n4759, new_n4760, new_n4761, new_n4762,
    new_n4763, new_n4764, new_n4765, new_n4766_1, new_n4767, new_n4768,
    new_n4769, new_n4770_1, new_n4771, new_n4772, new_n4773, new_n4774,
    new_n4775, new_n4776, new_n4777_1, new_n4778, new_n4779, new_n4780,
    new_n4781, new_n4782, new_n4783, new_n4784, new_n4785_1, new_n4786,
    new_n4787, new_n4788, new_n4789, new_n4790, new_n4791, new_n4792,
    new_n4793, new_n4794, new_n4795, new_n4796, new_n4797, new_n4798,
    new_n4799, new_n4800, new_n4801, new_n4802, new_n4803, new_n4804_1,
    new_n4805, new_n4806, new_n4807, new_n4808, new_n4809, new_n4810_1,
    new_n4811, new_n4812_1, new_n4813, new_n4814_1, new_n4815, new_n4816,
    new_n4817, new_n4819, new_n4820, new_n4821, new_n4822, new_n4823,
    new_n4824, new_n4825, new_n4826, new_n4827, new_n4828, new_n4829,
    new_n4830, new_n4831, new_n4832, new_n4833, new_n4834, new_n4835,
    new_n4836, new_n4837, new_n4838, new_n4839, new_n4840, new_n4841,
    new_n4842, new_n4843, new_n4844, new_n4845, new_n4846, new_n4847,
    new_n4848, new_n4849, new_n4850_1, new_n4851, new_n4852, new_n4853,
    new_n4854, new_n4855, new_n4856, new_n4857, new_n4858_1, new_n4859,
    new_n4860, new_n4861, new_n4862, new_n4863, new_n4864, new_n4865,
    new_n4866, new_n4867, new_n4868, new_n4869, new_n4870, new_n4871,
    new_n4872, new_n4873, new_n4874, new_n4875, new_n4876, new_n4877,
    new_n4878, new_n4879, new_n4880, new_n4881, new_n4882, new_n4883,
    new_n4884, new_n4885, new_n4886, new_n4887, new_n4888, new_n4889,
    new_n4890, new_n4891_1, new_n4892, new_n4893, new_n4894, new_n4895,
    new_n4896, new_n4897, new_n4898, new_n4899, new_n4900, new_n4901,
    new_n4902, new_n4903, new_n4904, new_n4905, new_n4906, new_n4907,
    new_n4908, new_n4909, new_n4910, new_n4911, new_n4912, new_n4913_1,
    new_n4914, new_n4915, new_n4916, new_n4917, new_n4918, new_n4919,
    new_n4920, new_n4921, new_n4922, new_n4923, new_n4924, new_n4925_1,
    new_n4926, new_n4927, new_n4928, new_n4929, new_n4930, new_n4931,
    new_n4932, new_n4933, new_n4934, new_n4935, new_n4936, new_n4937,
    new_n4938, new_n4939_1, new_n4940, new_n4941, new_n4942, new_n4943,
    new_n4944, new_n4945, new_n4946, new_n4947_1, new_n4948, new_n4949,
    new_n4950, new_n4951, new_n4952_1, new_n4953, new_n4954, new_n4955,
    new_n4956, new_n4957_1, new_n4958, new_n4959, new_n4960, new_n4961,
    new_n4962, new_n4963, new_n4964_1, new_n4965, new_n4966_1, new_n4967_1,
    new_n4968, new_n4969, new_n4970, new_n4971, new_n4972_1, new_n4973,
    new_n4974, new_n4975, new_n4976, new_n4977, new_n4978, new_n4979,
    new_n4980, new_n4981, new_n4982, new_n4983, new_n4984, new_n4985,
    new_n4986, new_n4987, new_n4988, new_n4989, new_n4990, new_n4991,
    new_n4992, new_n4993, new_n4994, new_n4995, new_n4996, new_n4997,
    new_n4998, new_n4999, new_n5000, new_n5001, new_n5002, new_n5003,
    new_n5004, new_n5005, new_n5006, new_n5007, new_n5008, new_n5009,
    new_n5010, new_n5011_1, new_n5012, new_n5013, new_n5014, new_n5015,
    new_n5016, new_n5017, new_n5018, new_n5019, new_n5020_1, new_n5021,
    new_n5022, new_n5024_1, new_n5025_1, new_n5026_1, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031_1, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046_1,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060_1, new_n5061, new_n5062_1, new_n5063, new_n5064_1,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077_1, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082_1,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098_1, new_n5099, new_n5100,
    new_n5101_1, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115_1, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120_1, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128_1, new_n5129, new_n5130,
    new_n5131_1, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140_1, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158_1, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168_1, new_n5169, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178,
    new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184_1,
    new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190,
    new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196,
    new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5202,
    new_n5203, new_n5204, new_n5205, new_n5206, new_n5207, new_n5208,
    new_n5209, new_n5210, new_n5211_1, new_n5212, new_n5213_1, new_n5214,
    new_n5215, new_n5216, new_n5217, new_n5218, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226_1,
    new_n5227, new_n5228_1, new_n5229, new_n5230, new_n5231, new_n5232,
    new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238,
    new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255_1, new_n5256_1,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265_1, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273_1, new_n5274_1,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300_1, new_n5301, new_n5302_1, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5310, new_n5311,
    new_n5312, new_n5313, new_n5314, new_n5315, new_n5316, new_n5317,
    new_n5318, new_n5319, new_n5320, new_n5321, new_n5322, new_n5323,
    new_n5324, new_n5325_1, new_n5326, new_n5327, new_n5329, new_n5330_1,
    new_n5331, new_n5334, new_n5335, new_n5336, new_n5337_1, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351_1, new_n5352, new_n5353_1, new_n5354, new_n5356, new_n5357,
    new_n5358, new_n5359, new_n5360, new_n5361, new_n5362, new_n5363,
    new_n5364, new_n5365, new_n5366, new_n5367, new_n5368, new_n5369,
    new_n5370, new_n5371, new_n5372, new_n5373, new_n5374, new_n5375,
    new_n5376_1, new_n5377, new_n5378, new_n5379, new_n5380, new_n5384,
    new_n5385, new_n5386_1, new_n5387, new_n5388, new_n5389, new_n5390,
    new_n5391, new_n5392, new_n5393, new_n5394, new_n5395, new_n5396,
    new_n5397, new_n5398, new_n5399_1, new_n5400_1, new_n5401, new_n5402,
    new_n5403_1, new_n5404, new_n5405, new_n5406, new_n5407, new_n5408,
    new_n5409, new_n5410, new_n5411, new_n5412, new_n5413, new_n5414,
    new_n5415, new_n5416, new_n5417, new_n5418, new_n5419, new_n5420,
    new_n5421, new_n5422, new_n5423, new_n5424, new_n5425, new_n5426,
    new_n5427, new_n5428, new_n5429, new_n5430_1, new_n5431, new_n5432,
    new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438_1,
    new_n5439_1, new_n5440, new_n5441, new_n5442, new_n5443_1, new_n5444,
    new_n5445, new_n5446, new_n5447, new_n5448, new_n5449, new_n5450,
    new_n5451_1, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472_1, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485_1, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516,
    new_n5517_1, new_n5518, new_n5519, new_n5520, new_n5521_1, new_n5522,
    new_n5523, new_n5524_1, new_n5525, new_n5526, new_n5527, new_n5528,
    new_n5529, new_n5530, new_n5531, new_n5532_1, new_n5533, new_n5534,
    new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540,
    new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546,
    new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552,
    new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564_1,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579_1, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593_1, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603_1, new_n5604, new_n5605_1, new_n5606,
    new_n5607, new_n5608, new_n5609_1, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5624, new_n5625,
    new_n5626, new_n5627, new_n5628, new_n5629, new_n5630, new_n5631,
    new_n5632, new_n5633, new_n5634_1, new_n5635, new_n5636, new_n5637,
    new_n5638, new_n5639, new_n5640, new_n5641, new_n5642, new_n5643_1,
    new_n5644, new_n5645, new_n5646, new_n5647, new_n5648, new_n5649,
    new_n5650, new_n5651, new_n5652, new_n5653, new_n5654, new_n5655,
    new_n5656, new_n5657, new_n5658, new_n5659, new_n5660, new_n5661,
    new_n5662, new_n5663, new_n5664, new_n5665, new_n5666, new_n5667,
    new_n5668, new_n5669, new_n5670, new_n5671, new_n5672, new_n5673,
    new_n5674, new_n5675, new_n5676, new_n5677, new_n5678, new_n5679,
    new_n5680_1, new_n5681, new_n5682, new_n5683, new_n5684, new_n5685,
    new_n5686, new_n5687_1, new_n5688, new_n5689, new_n5690, new_n5691,
    new_n5692, new_n5693, new_n5694, new_n5695, new_n5696_1, new_n5697,
    new_n5698, new_n5699, new_n5700_1, new_n5701, new_n5702, new_n5703,
    new_n5704_1, new_n5705, new_n5706, new_n5707, new_n5708, new_n5709,
    new_n5710, new_n5711, new_n5712, new_n5713, new_n5714, new_n5715,
    new_n5716, new_n5717, new_n5718, new_n5719, new_n5720, new_n5721,
    new_n5722, new_n5723, new_n5724, new_n5725, new_n5726, new_n5727,
    new_n5728, new_n5729, new_n5730, new_n5731, new_n5732_1, new_n5733,
    new_n5734, new_n5735, new_n5736, new_n5737, new_n5738, new_n5739,
    new_n5740, new_n5741, new_n5742_1, new_n5743, new_n5744, new_n5745,
    new_n5746, new_n5747, new_n5748, new_n5749, new_n5750, new_n5751,
    new_n5752_1, new_n5753, new_n5754, new_n5755, new_n5756, new_n5757,
    new_n5758, new_n5759, new_n5760, new_n5761, new_n5762, new_n5763,
    new_n5764, new_n5765_1, new_n5766, new_n5767, new_n5768, new_n5769,
    new_n5770, new_n5771, new_n5772, new_n5773, new_n5774, new_n5775,
    new_n5776_1, new_n5777, new_n5778, new_n5779, new_n5780, new_n5781,
    new_n5782_1, new_n5783, new_n5784, new_n5785, new_n5786, new_n5787,
    new_n5788, new_n5789, new_n5790, new_n5791, new_n5792, new_n5793,
    new_n5794, new_n5795, new_n5796, new_n5797, new_n5798, new_n5799,
    new_n5800, new_n5801, new_n5802, new_n5803, new_n5804, new_n5805,
    new_n5806, new_n5807, new_n5808, new_n5809, new_n5810, new_n5811,
    new_n5812, new_n5813, new_n5814, new_n5815, new_n5816, new_n5817,
    new_n5818, new_n5819, new_n5820, new_n5821, new_n5822_1, new_n5823,
    new_n5824, new_n5825, new_n5826, new_n5827, new_n5828, new_n5829,
    new_n5830, new_n5831, new_n5832, new_n5833_1, new_n5834_1, new_n5835,
    new_n5836, new_n5837, new_n5838, new_n5840_1, new_n5841_1, new_n5842_1,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850_1, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882_1, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903_1, new_n5904_1, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911_1, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934, new_n5935, new_n5936_1, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943_1, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980_1,
    new_n5981, new_n5983, new_n5984, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012_1,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022_1, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031_1, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044_1, new_n6045, new_n6046_1, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6055,
    new_n6056, new_n6057, new_n6058, new_n6059, new_n6060, new_n6061,
    new_n6062, new_n6063, new_n6064, new_n6065, new_n6066, new_n6067,
    new_n6068, new_n6069, new_n6070, new_n6071, new_n6072, new_n6073,
    new_n6074, new_n6075, new_n6076, new_n6077, new_n6078, new_n6079,
    new_n6080, new_n6081, new_n6082, new_n6083, new_n6084_1, new_n6085,
    new_n6086, new_n6087, new_n6088, new_n6089, new_n6090, new_n6091,
    new_n6092, new_n6093, new_n6094, new_n6095, new_n6096, new_n6097,
    new_n6098, new_n6099, new_n6100, new_n6101, new_n6102, new_n6103,
    new_n6104_1, new_n6105_1, new_n6106, new_n6107, new_n6108, new_n6109,
    new_n6110, new_n6111, new_n6112, new_n6113, new_n6114, new_n6115,
    new_n6116, new_n6117, new_n6118, new_n6119, new_n6120, new_n6121,
    new_n6122, new_n6123, new_n6124, new_n6126, new_n6127, new_n6128,
    new_n6129, new_n6130, new_n6131, new_n6132, new_n6133, new_n6134,
    new_n6135, new_n6136, new_n6137, new_n6138, new_n6139, new_n6140,
    new_n6141, new_n6142, new_n6143, new_n6144, new_n6145, new_n6146,
    new_n6147, new_n6148, new_n6149, new_n6150, new_n6151, new_n6152,
    new_n6153, new_n6154, new_n6155, new_n6156, new_n6157, new_n6158,
    new_n6159, new_n6160_1, new_n6161, new_n6162, new_n6163, new_n6164,
    new_n6165, new_n6166, new_n6167, new_n6168, new_n6169, new_n6170,
    new_n6171_1, new_n6172, new_n6173, new_n6174, new_n6175, new_n6176,
    new_n6177, new_n6178, new_n6179, new_n6180, new_n6181, new_n6182,
    new_n6183_1, new_n6184, new_n6185, new_n6186, new_n6187, new_n6188,
    new_n6189_1, new_n6190, new_n6191, new_n6192, new_n6193, new_n6194,
    new_n6195, new_n6196, new_n6197, new_n6198, new_n6199, new_n6200,
    new_n6201, new_n6202, new_n6203, new_n6204_1, new_n6205, new_n6206,
    new_n6207, new_n6208, new_n6209, new_n6210, new_n6211, new_n6212,
    new_n6213, new_n6214, new_n6215, new_n6216, new_n6217, new_n6218_1,
    new_n6219, new_n6220, new_n6221, new_n6222, new_n6223_1, new_n6224,
    new_n6225, new_n6226, new_n6227, new_n6228, new_n6229, new_n6230,
    new_n6231, new_n6232, new_n6233_1, new_n6234, new_n6235, new_n6236,
    new_n6237, new_n6238, new_n6239, new_n6240, new_n6241, new_n6242,
    new_n6243, new_n6244, new_n6245_1, new_n6246, new_n6247, new_n6248_1,
    new_n6249, new_n6250, new_n6251, new_n6252, new_n6253, new_n6254,
    new_n6255, new_n6256_1, new_n6257, new_n6258, new_n6259, new_n6260,
    new_n6261, new_n6262, new_n6263, new_n6264, new_n6265, new_n6266,
    new_n6267, new_n6268, new_n6269, new_n6270, new_n6271_1, new_n6272,
    new_n6273, new_n6274, new_n6275, new_n6276_1, new_n6277, new_n6278,
    new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6284,
    new_n6285, new_n6286, new_n6287, new_n6288, new_n6289, new_n6290,
    new_n6291, new_n6292, new_n6293, new_n6294, new_n6295, new_n6296,
    new_n6297, new_n6298, new_n6299, new_n6300, new_n6301, new_n6302,
    new_n6303, new_n6304, new_n6305, new_n6306, new_n6308_1, new_n6309,
    new_n6310, new_n6311_1, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323_1, new_n6324, new_n6325, new_n6326, new_n6327,
    new_n6328, new_n6329, new_n6330_1, new_n6331, new_n6332, new_n6333,
    new_n6334, new_n6335, new_n6336, new_n6337, new_n6338, new_n6339_1,
    new_n6340, new_n6341, new_n6342, new_n6343, new_n6344, new_n6345,
    new_n6346, new_n6347, new_n6348, new_n6349, new_n6350, new_n6351,
    new_n6352, new_n6353, new_n6354_1, new_n6355, new_n6356_1, new_n6357,
    new_n6358, new_n6359, new_n6360, new_n6361, new_n6362, new_n6363,
    new_n6364, new_n6365, new_n6366, new_n6367, new_n6368, new_n6369_1,
    new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375_1,
    new_n6376, new_n6377, new_n6378, new_n6379_1, new_n6380, new_n6381_1,
    new_n6382, new_n6383_1, new_n6384, new_n6385_1, new_n6386, new_n6387,
    new_n6388, new_n6389, new_n6390, new_n6391, new_n6392, new_n6393,
    new_n6394, new_n6395, new_n6396, new_n6397_1, new_n6398, new_n6399,
    new_n6400, new_n6401, new_n6402, new_n6403, new_n6404, new_n6405,
    new_n6406, new_n6407_1, new_n6408, new_n6409, new_n6410, new_n6411,
    new_n6412, new_n6413, new_n6414, new_n6415, new_n6416, new_n6417,
    new_n6418, new_n6419, new_n6420, new_n6421, new_n6422, new_n6423,
    new_n6424, new_n6425, new_n6426, new_n6427_1, new_n6428, new_n6429,
    new_n6430, new_n6431_1, new_n6432, new_n6433, new_n6434, new_n6435,
    new_n6436, new_n6437_1, new_n6438, new_n6439, new_n6440, new_n6441,
    new_n6442, new_n6443, new_n6444, new_n6445, new_n6446, new_n6447,
    new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453,
    new_n6454, new_n6455, new_n6456_1, new_n6457_1, new_n6458, new_n6459,
    new_n6460, new_n6461, new_n6462, new_n6463, new_n6464, new_n6465_1,
    new_n6466, new_n6467, new_n6468, new_n6469, new_n6470_1, new_n6471,
    new_n6472, new_n6473, new_n6474, new_n6475, new_n6476_1, new_n6477,
    new_n6478, new_n6479, new_n6480, new_n6481, new_n6482, new_n6483,
    new_n6484, new_n6485_1, new_n6486, new_n6487, new_n6488, new_n6489,
    new_n6490, new_n6491, new_n6492, new_n6493, new_n6494, new_n6495,
    new_n6496, new_n6497, new_n6498, new_n6499, new_n6500, new_n6501,
    new_n6502_1, new_n6503, new_n6504, new_n6505, new_n6506_1, new_n6507,
    new_n6508, new_n6509, new_n6510, new_n6511, new_n6512, new_n6513_1,
    new_n6514_1, new_n6515, new_n6516, new_n6517, new_n6518, new_n6519,
    new_n6520, new_n6522, new_n6523, new_n6524, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542_1, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556_1, new_n6557,
    new_n6558_1, new_n6559, new_n6560_1, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567_1, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576_1, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587_1,
    new_n6588, new_n6589, new_n6590_1, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596_1, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611_1,
    new_n6612_1, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628_1, new_n6629,
    new_n6630_1, new_n6631_1, new_n6632, new_n6633, new_n6634_1, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6645, new_n6646, new_n6647,
    new_n6648, new_n6649, new_n6650, new_n6651, new_n6652_1, new_n6653,
    new_n6654, new_n6655_1, new_n6656, new_n6657, new_n6658, new_n6659_1,
    new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665,
    new_n6666, new_n6667, new_n6668, new_n6669_1, new_n6670, new_n6671_1,
    new_n6672, new_n6673_1, new_n6674_1, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684_1, new_n6685, new_n6686, new_n6687, new_n6688, new_n6689,
    new_n6690, new_n6691_1, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703, new_n6704, new_n6705, new_n6706_1, new_n6707_1,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729_1, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736_1, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6744,
    new_n6745, new_n6746, new_n6747, new_n6748, new_n6749, new_n6750,
    new_n6751, new_n6752, new_n6753, new_n6754, new_n6755, new_n6756,
    new_n6757, new_n6758, new_n6759, new_n6760, new_n6761, new_n6762,
    new_n6763, new_n6764, new_n6765, new_n6766, new_n6767, new_n6768,
    new_n6769, new_n6770, new_n6771, new_n6772, new_n6773_1, new_n6774,
    new_n6775_1, new_n6776, new_n6777, new_n6778, new_n6779, new_n6780,
    new_n6781, new_n6782, new_n6783, new_n6784, new_n6785_1, new_n6786,
    new_n6787, new_n6788, new_n6789, new_n6790_1, new_n6791_1, new_n6792,
    new_n6793, new_n6794_1, new_n6795, new_n6796, new_n6797, new_n6798,
    new_n6799, new_n6800, new_n6801, new_n6802_1, new_n6803, new_n6804,
    new_n6805, new_n6806, new_n6807, new_n6808, new_n6809, new_n6810,
    new_n6811, new_n6812, new_n6813, new_n6814_1, new_n6815, new_n6816,
    new_n6817, new_n6818, new_n6819, new_n6820, new_n6821, new_n6822,
    new_n6823, new_n6824, new_n6825, new_n6826_1, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835_1, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853_1, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860, new_n6861_1, new_n6862_1, new_n6863_1, new_n6864,
    new_n6865, new_n6866, new_n6867_1, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6924, new_n6925,
    new_n6926, new_n6927, new_n6928, new_n6929, new_n6930, new_n6931,
    new_n6932, new_n6933, new_n6934, new_n6935, new_n6936, new_n6937,
    new_n6938, new_n6939, new_n6940, new_n6941, new_n6942, new_n6943,
    new_n6944, new_n6945, new_n6946, new_n6947, new_n6948, new_n6949,
    new_n6950, new_n6951, new_n6952, new_n6953, new_n6954, new_n6955,
    new_n6956, new_n6957, new_n6958, new_n6959, new_n6960, new_n6961,
    new_n6962, new_n6963, new_n6964, new_n6965_1, new_n6966, new_n6967_1,
    new_n6968, new_n6969, new_n6970, new_n6971_1, new_n6972, new_n6973,
    new_n6974, new_n6975_1, new_n6976, new_n6977, new_n6978, new_n6979,
    new_n6980, new_n6981, new_n6982, new_n6983_1, new_n6984, new_n6985_1,
    new_n6986, new_n6987, new_n6988, new_n6989, new_n6990, new_n6991,
    new_n6992, new_n6993, new_n6994, new_n6995, new_n6996, new_n6997,
    new_n6998_1, new_n6999, new_n7000, new_n7001, new_n7002, new_n7003,
    new_n7004, new_n7005, new_n7006, new_n7007, new_n7008, new_n7009,
    new_n7010, new_n7011, new_n7012, new_n7013, new_n7014, new_n7015,
    new_n7016, new_n7017, new_n7018, new_n7019, new_n7020, new_n7021,
    new_n7022, new_n7023, new_n7024, new_n7025, new_n7026_1, new_n7027,
    new_n7028, new_n7029, new_n7030, new_n7031, new_n7032_1, new_n7033,
    new_n7034, new_n7035, new_n7036, new_n7037, new_n7038_1, new_n7039,
    new_n7040, new_n7041, new_n7042, new_n7043, new_n7044, new_n7045,
    new_n7046, new_n7047, new_n7048, new_n7049, new_n7050, new_n7051,
    new_n7052, new_n7053, new_n7054, new_n7055, new_n7056, new_n7057_1,
    new_n7058, new_n7059, new_n7060, new_n7061, new_n7062, new_n7063,
    new_n7064, new_n7065, new_n7066, new_n7067, new_n7068, new_n7069,
    new_n7070, new_n7071, new_n7072, new_n7073, new_n7074, new_n7075,
    new_n7076, new_n7077, new_n7078, new_n7079_1, new_n7080, new_n7081,
    new_n7082, new_n7083, new_n7084, new_n7085, new_n7086, new_n7087,
    new_n7088, new_n7089, new_n7090, new_n7091, new_n7092, new_n7093,
    new_n7094, new_n7095, new_n7096, new_n7097, new_n7098, new_n7099_1,
    new_n7100, new_n7101, new_n7102, new_n7103, new_n7104, new_n7105,
    new_n7106, new_n7107, new_n7108, new_n7109, new_n7110, new_n7111,
    new_n7112, new_n7113, new_n7114, new_n7115, new_n7116, new_n7117,
    new_n7118, new_n7119, new_n7120, new_n7121, new_n7122, new_n7123,
    new_n7124, new_n7125, new_n7126, new_n7127, new_n7128, new_n7129,
    new_n7130, new_n7131, new_n7132, new_n7133, new_n7134, new_n7135,
    new_n7136, new_n7137, new_n7138, new_n7139_1, new_n7140, new_n7141,
    new_n7142, new_n7143, new_n7144, new_n7145, new_n7146, new_n7147,
    new_n7148, new_n7149_1, new_n7150, new_n7151, new_n7152, new_n7153,
    new_n7154, new_n7155, new_n7156, new_n7157, new_n7158, new_n7159,
    new_n7160, new_n7161, new_n7162, new_n7163, new_n7164, new_n7165,
    new_n7166, new_n7167, new_n7168, new_n7169, new_n7170, new_n7171,
    new_n7172, new_n7173, new_n7174, new_n7175, new_n7176, new_n7177,
    new_n7178, new_n7179, new_n7180, new_n7181, new_n7182, new_n7183,
    new_n7184, new_n7185, new_n7186, new_n7187, new_n7188, new_n7189,
    new_n7190_1, new_n7191, new_n7192, new_n7193, new_n7194, new_n7195,
    new_n7196, new_n7197, new_n7198, new_n7199, new_n7200, new_n7201,
    new_n7202, new_n7204, new_n7205, new_n7206, new_n7207, new_n7208,
    new_n7209, new_n7210, new_n7211, new_n7212, new_n7213, new_n7214,
    new_n7215, new_n7216, new_n7217, new_n7218, new_n7219, new_n7220,
    new_n7221, new_n7222, new_n7223, new_n7224, new_n7225, new_n7226,
    new_n7227, new_n7228, new_n7229_1, new_n7230_1, new_n7231, new_n7232,
    new_n7233_1, new_n7234, new_n7235, new_n7236_1, new_n7237, new_n7238,
    new_n7239, new_n7240, new_n7241, new_n7242, new_n7243, new_n7244,
    new_n7245, new_n7246, new_n7247, new_n7248, new_n7249, new_n7250,
    new_n7251, new_n7252, new_n7253_1, new_n7254, new_n7255, new_n7256_1,
    new_n7257, new_n7258, new_n7259, new_n7260, new_n7261, new_n7262,
    new_n7263, new_n7264, new_n7265, new_n7266, new_n7267, new_n7268_1,
    new_n7269, new_n7270, new_n7271, new_n7272, new_n7273, new_n7274,
    new_n7275, new_n7276, new_n7277_1, new_n7278, new_n7279, new_n7280_1,
    new_n7281, new_n7282, new_n7283, new_n7284, new_n7285, new_n7286,
    new_n7287, new_n7288, new_n7289, new_n7290, new_n7291, new_n7292,
    new_n7293, new_n7294, new_n7295, new_n7296, new_n7297, new_n7298_1,
    new_n7299, new_n7300, new_n7301, new_n7302, new_n7303, new_n7304,
    new_n7305_1, new_n7306, new_n7307, new_n7308_1, new_n7309, new_n7310,
    new_n7311, new_n7312, new_n7313_1, new_n7314, new_n7315, new_n7316,
    new_n7317, new_n7318, new_n7319, new_n7320, new_n7321, new_n7322,
    new_n7323, new_n7324, new_n7325, new_n7326, new_n7327, new_n7328,
    new_n7329, new_n7330_1, new_n7331, new_n7332, new_n7333, new_n7334,
    new_n7335_1, new_n7336, new_n7337, new_n7338, new_n7339_1, new_n7340,
    new_n7341, new_n7342, new_n7343, new_n7344, new_n7345, new_n7346_1,
    new_n7347, new_n7348, new_n7349_1, new_n7350, new_n7351, new_n7352,
    new_n7353, new_n7354, new_n7355, new_n7356, new_n7357, new_n7358,
    new_n7359, new_n7360, new_n7361, new_n7362, new_n7363_1, new_n7364,
    new_n7365, new_n7366, new_n7367, new_n7368, new_n7369, new_n7370,
    new_n7371, new_n7372, new_n7373, new_n7374, new_n7375, new_n7376,
    new_n7377_1, new_n7378, new_n7379, new_n7380, new_n7381, new_n7382,
    new_n7383, new_n7384, new_n7385, new_n7386, new_n7387, new_n7388,
    new_n7389, new_n7390_1, new_n7391, new_n7392, new_n7393, new_n7394,
    new_n7395, new_n7396, new_n7397, new_n7398, new_n7399, new_n7400,
    new_n7401, new_n7402, new_n7403_1, new_n7404, new_n7405, new_n7406,
    new_n7407, new_n7408_1, new_n7409, new_n7410, new_n7411, new_n7412,
    new_n7413, new_n7414, new_n7415, new_n7416, new_n7417, new_n7418,
    new_n7419, new_n7420, new_n7421_1, new_n7422, new_n7423, new_n7424,
    new_n7425, new_n7426, new_n7427, new_n7428_1, new_n7429, new_n7430,
    new_n7431, new_n7432_1, new_n7433, new_n7434, new_n7435, new_n7436,
    new_n7437_1, new_n7438, new_n7439, new_n7440, new_n7441, new_n7442,
    new_n7443, new_n7444, new_n7445, new_n7446, new_n7447, new_n7448,
    new_n7449, new_n7450, new_n7451, new_n7452, new_n7453, new_n7454,
    new_n7455, new_n7456, new_n7457, new_n7458, new_n7459, new_n7460_1,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475_1, new_n7476, new_n7477_1, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507_1, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514_1, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524_1, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558_1,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566_1, new_n7567, new_n7568, new_n7569_1, new_n7570,
    new_n7571, new_n7572_1, new_n7573, new_n7574, new_n7575_1, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585_1, new_n7586, new_n7587, new_n7588_1,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593_1, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598_1, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607_1, new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616_1, new_n7617, new_n7618,
    new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624,
    new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630_1,
    new_n7631, new_n7632, new_n7633, new_n7634, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643_1,
    new_n7644, new_n7645, new_n7646, new_n7647_1, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657_1, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670_1, new_n7671, new_n7672, new_n7674_1,
    new_n7675, new_n7676, new_n7677, new_n7678_1, new_n7679_1, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686_1,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692_1,
    new_n7693_1, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698_1,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708_1, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7714, new_n7715, new_n7716, new_n7717,
    new_n7718, new_n7719, new_n7720, new_n7721_1, new_n7722, new_n7723,
    new_n7724, new_n7725, new_n7726, new_n7727, new_n7728, new_n7729,
    new_n7730, new_n7731_1, new_n7732, new_n7733, new_n7734, new_n7735,
    new_n7736, new_n7737, new_n7738, new_n7739, new_n7740, new_n7741,
    new_n7742, new_n7743, new_n7744, new_n7745, new_n7746, new_n7747,
    new_n7748, new_n7749, new_n7750, new_n7751_1, new_n7752, new_n7753,
    new_n7754, new_n7755, new_n7756, new_n7757, new_n7758, new_n7759_1,
    new_n7760, new_n7761, new_n7762, new_n7763, new_n7764, new_n7765,
    new_n7766, new_n7767, new_n7768, new_n7769_1, new_n7770, new_n7771,
    new_n7772, new_n7773_1, new_n7774, new_n7775, new_n7776, new_n7777,
    new_n7778, new_n7779, new_n7780_1, new_n7781, new_n7782, new_n7783,
    new_n7784, new_n7785, new_n7786, new_n7787, new_n7788_1, new_n7789,
    new_n7790, new_n7791, new_n7792, new_n7793, new_n7794_1, new_n7795,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811_1, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820,
    new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826,
    new_n7827, new_n7828, new_n7829, new_n7830_1, new_n7831, new_n7832,
    new_n7833, new_n7834_1, new_n7835, new_n7836, new_n7837, new_n7838,
    new_n7839, new_n7840, new_n7841_1, new_n7842, new_n7843, new_n7844,
    new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850,
    new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856,
    new_n7857, new_n7859, new_n7860, new_n7861, new_n7862, new_n7863,
    new_n7864, new_n7865, new_n7866, new_n7867, new_n7868, new_n7869,
    new_n7870, new_n7871, new_n7872, new_n7873, new_n7874, new_n7875,
    new_n7876_1, new_n7877, new_n7878, new_n7879, new_n7880, new_n7881,
    new_n7882, new_n7883, new_n7884_1, new_n7885, new_n7886, new_n7887,
    new_n7888, new_n7889, new_n7890, new_n7891, new_n7892, new_n7893,
    new_n7894, new_n7895, new_n7896, new_n7897, new_n7898, new_n7899,
    new_n7900, new_n7901, new_n7902, new_n7903, new_n7904, new_n7905,
    new_n7906, new_n7907, new_n7908, new_n7909, new_n7910, new_n7911,
    new_n7912, new_n7913, new_n7914, new_n7915, new_n7916, new_n7917_1,
    new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923,
    new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929,
    new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935,
    new_n7936, new_n7937_1, new_n7938, new_n7939, new_n7940, new_n7941,
    new_n7942, new_n7943_1, new_n7944, new_n7945, new_n7946, new_n7947,
    new_n7948, new_n7949_1, new_n7950_1, new_n7951, new_n7952, new_n7953,
    new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959_1,
    new_n7960, new_n7961, new_n7962, new_n7963_1, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968_1, new_n7969, new_n7970, new_n7971,
    new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989,
    new_n7990, new_n7991, new_n7992_1, new_n7993, new_n7994, new_n7995,
    new_n7996, new_n7997, new_n7998, new_n7999_1, new_n8000, new_n8001,
    new_n8002, new_n8003, new_n8004, new_n8005, new_n8006_1, new_n8007,
    new_n8008, new_n8009, new_n8010, new_n8011, new_n8012, new_n8013,
    new_n8014, new_n8015, new_n8016, new_n8017, new_n8018, new_n8019,
    new_n8020, new_n8021, new_n8022, new_n8023, new_n8024, new_n8025,
    new_n8026, new_n8027_1, new_n8028, new_n8029, new_n8030, new_n8031_1,
    new_n8032, new_n8033, new_n8034, new_n8035, new_n8036, new_n8037,
    new_n8038, new_n8039, new_n8040, new_n8041, new_n8042_1, new_n8043,
    new_n8044, new_n8045, new_n8046, new_n8047, new_n8048, new_n8049,
    new_n8050, new_n8051, new_n8052_1, new_n8053, new_n8054, new_n8055,
    new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061,
    new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067_1,
    new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073,
    new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079,
    new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085,
    new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091,
    new_n8092, new_n8093, new_n8094, new_n8095_1, new_n8096, new_n8097,
    new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8104,
    new_n8105, new_n8106, new_n8108, new_n8109_1, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127_1, new_n8128, new_n8129,
    new_n8130_1, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135_1,
    new_n8136, new_n8137, new_n8138, new_n8139_1, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148_1, new_n8149_1, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159_1,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179_1, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194_1, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215_1, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244_1, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8256_1,
    new_n8257, new_n8258, new_n8259_1, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267_1, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285_1, new_n8286,
    new_n8287, new_n8288_1, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304,
    new_n8305_1, new_n8306_1, new_n8307, new_n8308, new_n8309_1, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320_1, new_n8321_1, new_n8322,
    new_n8323, new_n8324_1, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336, new_n8337, new_n8338, new_n8339_1, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363_1, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376_1,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381_1, new_n8382,
    new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399_1, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405_1, new_n8406,
    new_n8407, new_n8408_1, new_n8409, new_n8410, new_n8415, new_n8416,
    new_n8417_1, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422,
    new_n8423, new_n8424, new_n8425, new_n8426, new_n8427, new_n8428,
    new_n8429, new_n8430, new_n8431, new_n8432_1, new_n8433, new_n8434,
    new_n8435, new_n8436, new_n8437, new_n8438, new_n8439_1, new_n8440,
    new_n8441, new_n8442, new_n8443, new_n8444, new_n8445, new_n8446,
    new_n8447, new_n8448, new_n8449, new_n8450, new_n8451, new_n8452,
    new_n8453_1, new_n8454, new_n8455, new_n8456, new_n8457, new_n8458,
    new_n8459, new_n8460, new_n8461, new_n8462, new_n8463, new_n8464,
    new_n8465, new_n8466, new_n8467, new_n8468, new_n8469, new_n8470,
    new_n8471, new_n8472, new_n8473, new_n8474, new_n8475, new_n8476,
    new_n8477, new_n8478, new_n8479, new_n8480_1, new_n8481, new_n8482,
    new_n8483, new_n8484, new_n8485, new_n8486, new_n8487, new_n8488,
    new_n8489_1, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494,
    new_n8495, new_n8496, new_n8497, new_n8498, new_n8499, new_n8500,
    new_n8501, new_n8502, new_n8503, new_n8504, new_n8505_1, new_n8506,
    new_n8507, new_n8508, new_n8509, new_n8510_1, new_n8511, new_n8512,
    new_n8513, new_n8514, new_n8515, new_n8516, new_n8517, new_n8518,
    new_n8519_1, new_n8520, new_n8521, new_n8522, new_n8523, new_n8524,
    new_n8525, new_n8526_1, new_n8527, new_n8528, new_n8529, new_n8530,
    new_n8531, new_n8532, new_n8533, new_n8534, new_n8535_1, new_n8536,
    new_n8537, new_n8538, new_n8539, new_n8540, new_n8541, new_n8542,
    new_n8543, new_n8544, new_n8545, new_n8546, new_n8547, new_n8548,
    new_n8549, new_n8550_1, new_n8551, new_n8552, new_n8553, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563_1, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581_1, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594_1, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608_1, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614_1, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620_1, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8633, new_n8634, new_n8635,
    new_n8636, new_n8637_1, new_n8638_1, new_n8639, new_n8640, new_n8641,
    new_n8642, new_n8643, new_n8644, new_n8645, new_n8646, new_n8647,
    new_n8648, new_n8649, new_n8650, new_n8651, new_n8652, new_n8653,
    new_n8654, new_n8655, new_n8656_1, new_n8657, new_n8658, new_n8659,
    new_n8660, new_n8661, new_n8662_1, new_n8663, new_n8664, new_n8665,
    new_n8666, new_n8667, new_n8668, new_n8669, new_n8670, new_n8671,
    new_n8672, new_n8673, new_n8674, new_n8675, new_n8676, new_n8677,
    new_n8678_1, new_n8679, new_n8680, new_n8681, new_n8682, new_n8683,
    new_n8684, new_n8685, new_n8686, new_n8687_1, new_n8688, new_n8689,
    new_n8690, new_n8691, new_n8692, new_n8693, new_n8694_1, new_n8695,
    new_n8696, new_n8697, new_n8698, new_n8699, new_n8700, new_n8701,
    new_n8702, new_n8703, new_n8704, new_n8705, new_n8706, new_n8707,
    new_n8708, new_n8709, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716_1, new_n8717, new_n8718, new_n8719, new_n8720,
    new_n8721_1, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744_1,
    new_n8745_1, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782_1, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803_1, new_n8804,
    new_n8805, new_n8806_1, new_n8807, new_n8808, new_n8809_1, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819, new_n8820, new_n8821_1, new_n8822,
    new_n8823, new_n8824_1, new_n8825, new_n8826, new_n8827_1, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8834, new_n8836,
    new_n8837, new_n8838, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849_1,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8857, new_n8859, new_n8860, new_n8861_1, new_n8862_1, new_n8863,
    new_n8864, new_n8865, new_n8866, new_n8867, new_n8868, new_n8869_1,
    new_n8870, new_n8871, new_n8872, new_n8873, new_n8874, new_n8875,
    new_n8876, new_n8877, new_n8878, new_n8879, new_n8880, new_n8881,
    new_n8882, new_n8883, new_n8884_1, new_n8885, new_n8886, new_n8887,
    new_n8888, new_n8889, new_n8890, new_n8891, new_n8892, new_n8893,
    new_n8894, new_n8895, new_n8896, new_n8897, new_n8898, new_n8899,
    new_n8900, new_n8901, new_n8902, new_n8903, new_n8904, new_n8905,
    new_n8906, new_n8907, new_n8908, new_n8909_1, new_n8910, new_n8911_1,
    new_n8912, new_n8913, new_n8914, new_n8915, new_n8916, new_n8917,
    new_n8918, new_n8919, new_n8920_1, new_n8921, new_n8922, new_n8923,
    new_n8924, new_n8925, new_n8926, new_n8927, new_n8928, new_n8929,
    new_n8930, new_n8931, new_n8932, new_n8933, new_n8934, new_n8935,
    new_n8936, new_n8937, new_n8938, new_n8939, new_n8940, new_n8941,
    new_n8942, new_n8943_1, new_n8944, new_n8945, new_n8946, new_n8947,
    new_n8948, new_n8949, new_n8950, new_n8951, new_n8952, new_n8953,
    new_n8954, new_n8955, new_n8956, new_n8957, new_n8958, new_n8959,
    new_n8960, new_n8961, new_n8962, new_n8963, new_n8964_1, new_n8965,
    new_n8966, new_n8967, new_n8968, new_n8969, new_n8970, new_n8971_1,
    new_n8972, new_n8973, new_n8974, new_n8975, new_n8976, new_n8977,
    new_n8978, new_n8979, new_n8980, new_n8981, new_n8982_1, new_n8983,
    new_n8984, new_n8985, new_n8986, new_n8987, new_n8988, new_n8989,
    new_n8990, new_n8991, new_n8992, new_n8993_1, new_n8994, new_n8995,
    new_n8996, new_n8997, new_n8998, new_n8999, new_n9000, new_n9001,
    new_n9002, new_n9003_1, new_n9004, new_n9005, new_n9006, new_n9007,
    new_n9008, new_n9009, new_n9010, new_n9011, new_n9012_1, new_n9013,
    new_n9014, new_n9015, new_n9016, new_n9017, new_n9018, new_n9019,
    new_n9020, new_n9021, new_n9022, new_n9023, new_n9024, new_n9025,
    new_n9026, new_n9027, new_n9028, new_n9029, new_n9030, new_n9031,
    new_n9032_1, new_n9033, new_n9034, new_n9035, new_n9036, new_n9037,
    new_n9038, new_n9039, new_n9040, new_n9041, new_n9042_1, new_n9043,
    new_n9044, new_n9045, new_n9046_1, new_n9047_1, new_n9048, new_n9049,
    new_n9050, new_n9051, new_n9052, new_n9053, new_n9054, new_n9055,
    new_n9056, new_n9057, new_n9058, new_n9059, new_n9060, new_n9061,
    new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067,
    new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073,
    new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079,
    new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085,
    new_n9086, new_n9087, new_n9088, new_n9089, new_n9090_1, new_n9091,
    new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104_1,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129_1, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146_1,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164_1,
    new_n9165, new_n9166_1, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172_1, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182_1,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189, new_n9190, new_n9191_1, new_n9192, new_n9193, new_n9194,
    new_n9195, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217_1, new_n9218,
    new_n9219, new_n9220_1, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246_1, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251_1, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259_1, new_n9260,
    new_n9261_1, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9270, new_n9271, new_n9272, new_n9273,
    new_n9274, new_n9275, new_n9276, new_n9277, new_n9278, new_n9279,
    new_n9280, new_n9281, new_n9282, new_n9283, new_n9284, new_n9285,
    new_n9286, new_n9287_1, new_n9288, new_n9289, new_n9290, new_n9291,
    new_n9292, new_n9293, new_n9294, new_n9295, new_n9296, new_n9297,
    new_n9298, new_n9299, new_n9300, new_n9301, new_n9302, new_n9303,
    new_n9304, new_n9305, new_n9306, new_n9307, new_n9308_1, new_n9309,
    new_n9310, new_n9311, new_n9312, new_n9313, new_n9314, new_n9315,
    new_n9316, new_n9317, new_n9318_1, new_n9319, new_n9320, new_n9321,
    new_n9322, new_n9323_1, new_n9324, new_n9325, new_n9326, new_n9327,
    new_n9328, new_n9329, new_n9330, new_n9331, new_n9332, new_n9333,
    new_n9334, new_n9335, new_n9336, new_n9337, new_n9338, new_n9339,
    new_n9340, new_n9341, new_n9342, new_n9343, new_n9344_1, new_n9345,
    new_n9346, new_n9347, new_n9348, new_n9349, new_n9350, new_n9351,
    new_n9352, new_n9353, new_n9354, new_n9355, new_n9356, new_n9357,
    new_n9358, new_n9359, new_n9360, new_n9361, new_n9362, new_n9363,
    new_n9364_1, new_n9365, new_n9366, new_n9367, new_n9368, new_n9369,
    new_n9370, new_n9371_1, new_n9372_1, new_n9373, new_n9374, new_n9375,
    new_n9376, new_n9377, new_n9378, new_n9379, new_n9380_1, new_n9381,
    new_n9382_1, new_n9383, new_n9384, new_n9385, new_n9386, new_n9387,
    new_n9388, new_n9389, new_n9390, new_n9391, new_n9392, new_n9393,
    new_n9394, new_n9395, new_n9396_1, new_n9397, new_n9398, new_n9399_1,
    new_n9400, new_n9401, new_n9402, new_n9403_1, new_n9404, new_n9405,
    new_n9406, new_n9407, new_n9408, new_n9409, new_n9410, new_n9411,
    new_n9412, new_n9413, new_n9414, new_n9415, new_n9416, new_n9417,
    new_n9418, new_n9419_1, new_n9420, new_n9421, new_n9422, new_n9423_1,
    new_n9424, new_n9425, new_n9426, new_n9427, new_n9428, new_n9429,
    new_n9430_1, new_n9431, new_n9432, new_n9433, new_n9434, new_n9435_1,
    new_n9436, new_n9437, new_n9438, new_n9439, new_n9440, new_n9441,
    new_n9442, new_n9443, new_n9444, new_n9445_1, new_n9446, new_n9447,
    new_n9448, new_n9449, new_n9450, new_n9451_1, new_n9452, new_n9453,
    new_n9454, new_n9455, new_n9456, new_n9457, new_n9458_1, new_n9459_1,
    new_n9460_1, new_n9461, new_n9462, new_n9463, new_n9464, new_n9465,
    new_n9466, new_n9467, new_n9468, new_n9469, new_n9470, new_n9471,
    new_n9472, new_n9473, new_n9474, new_n9475, new_n9476, new_n9477,
    new_n9478, new_n9479, new_n9480, new_n9481, new_n9482, new_n9483,
    new_n9484, new_n9485, new_n9486, new_n9487, new_n9488, new_n9489,
    new_n9490, new_n9491, new_n9493_1, new_n9494, new_n9495, new_n9496,
    new_n9497, new_n9498, new_n9499, new_n9500, new_n9501, new_n9502,
    new_n9503, new_n9504, new_n9505, new_n9506, new_n9507_1, new_n9508_1,
    new_n9509, new_n9510, new_n9511, new_n9512_1, new_n9513, new_n9514,
    new_n9515, new_n9516, new_n9517, new_n9518, new_n9519, new_n9520,
    new_n9521, new_n9522, new_n9523, new_n9524, new_n9525, new_n9526,
    new_n9527, new_n9528, new_n9529, new_n9530, new_n9531, new_n9532,
    new_n9533, new_n9534, new_n9535, new_n9536, new_n9537, new_n9538,
    new_n9539, new_n9540, new_n9541, new_n9542, new_n9543, new_n9544,
    new_n9545, new_n9546, new_n9547, new_n9548, new_n9549, new_n9550,
    new_n9551, new_n9552_1, new_n9553, new_n9554_1, new_n9555, new_n9556_1,
    new_n9557_1, new_n9558_1, new_n9559, new_n9560, new_n9561, new_n9562,
    new_n9563, new_n9564, new_n9565, new_n9566, new_n9567, new_n9568,
    new_n9569, new_n9570, new_n9571, new_n9572, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598_1, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616_1, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622_1, new_n9623,
    new_n9624, new_n9625, new_n9626_1, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633_1, new_n9634, new_n9635_1,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646_1, new_n9647,
    new_n9648_1, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655_1, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689_1, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695_1, new_n9696,
    new_n9697, new_n9698, new_n9699_1, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726_1,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753_1, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761_1, new_n9762,
    new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1, new_n9768,
    new_n9769, new_n9770, new_n9771_1, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778_1, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783_1, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803_1, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9814, new_n9815, new_n9817, new_n9818,
    new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832_1, new_n9833_1, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838_1, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848,
    new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867_1, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872_1,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890_1,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9897,
    new_n9898, new_n9899, new_n9900, new_n9901, new_n9902, new_n9903,
    new_n9904, new_n9905, new_n9906, new_n9907, new_n9908, new_n9909,
    new_n9910, new_n9911, new_n9912, new_n9913, new_n9914, new_n9915,
    new_n9916, new_n9917_1, new_n9918, new_n9919_1, new_n9920, new_n9921,
    new_n9922, new_n9923, new_n9924, new_n9925, new_n9926_1, new_n9927,
    new_n9928, new_n9929, new_n9930, new_n9931, new_n9932, new_n9933,
    new_n9934_1, new_n9935, new_n9936, new_n9937, new_n9938_1, new_n9939,
    new_n9940, new_n9941, new_n9942_1, new_n9943, new_n9944, new_n9945,
    new_n9946_1, new_n9947, new_n9948, new_n9949, new_n9950, new_n9951,
    new_n9952, new_n9953, new_n9954, new_n9955, new_n9956, new_n9957,
    new_n9958, new_n9959, new_n9960, new_n9961, new_n9962, new_n9963,
    new_n9964, new_n9965, new_n9966, new_n9967_1, new_n9968_1, new_n9969,
    new_n9970, new_n9971, new_n9972, new_n9973, new_n9974, new_n9975,
    new_n9976, new_n9977, new_n9978, new_n9979, new_n9980, new_n9981,
    new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009_1, new_n10010_1,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017_1, new_n10018_1, new_n10019_1, new_n10020, new_n10021_1,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051,
    new_n10052, new_n10053_1, new_n10054, new_n10055_1, new_n10056,
    new_n10057_1, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10094, new_n10095, new_n10096_1, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101_1, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111_1, new_n10112, new_n10113,
    new_n10114, new_n10115, new_n10116, new_n10117_1, new_n10118,
    new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125_1, new_n10126, new_n10127, new_n10128, new_n10129,
    new_n10130, new_n10131, new_n10132, new_n10133, new_n10134, new_n10135,
    new_n10136, new_n10137, new_n10138, new_n10139, new_n10140, new_n10141,
    new_n10142, new_n10143, new_n10144, new_n10145, new_n10146, new_n10147,
    new_n10148, new_n10149, new_n10151, new_n10152, new_n10153, new_n10154,
    new_n10155, new_n10156, new_n10158_1, new_n10159, new_n10160,
    new_n10161, new_n10162, new_n10163, new_n10164, new_n10165_1,
    new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177,
    new_n10178, new_n10179, new_n10180, new_n10181, new_n10182, new_n10183,
    new_n10184, new_n10185, new_n10186, new_n10187, new_n10188, new_n10189,
    new_n10190, new_n10191, new_n10192, new_n10193, new_n10194, new_n10195,
    new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201_1, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229,
    new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236_1, new_n10237, new_n10238, new_n10239_1, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244_1, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250_1,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261_1,
    new_n10262_1, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10279, new_n10280, new_n10281, new_n10282,
    new_n10283, new_n10284, new_n10285, new_n10286, new_n10287_1,
    new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293,
    new_n10294, new_n10295_1, new_n10296, new_n10297, new_n10298,
    new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304,
    new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310,
    new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316,
    new_n10317, new_n10318, new_n10319, new_n10320, new_n10321_1,
    new_n10322, new_n10323, new_n10324, new_n10325, new_n10326_1,
    new_n10327_1, new_n10328, new_n10329, new_n10330_1, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340_1, new_n10341, new_n10342,
    new_n10343, new_n10344, new_n10345_1, new_n10346, new_n10347,
    new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356_1, new_n10357, new_n10358,
    new_n10359, new_n10360, new_n10361, new_n10362, new_n10363, new_n10364,
    new_n10365, new_n10366, new_n10367, new_n10368, new_n10369, new_n10370,
    new_n10371, new_n10372_1, new_n10373, new_n10374, new_n10375,
    new_n10376, new_n10377, new_n10378, new_n10379, new_n10380, new_n10381,
    new_n10382, new_n10383, new_n10384, new_n10385_1, new_n10386,
    new_n10387_1, new_n10388_1, new_n10389, new_n10390_1, new_n10391,
    new_n10392, new_n10393, new_n10394, new_n10395, new_n10396, new_n10397,
    new_n10398, new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404_1, new_n10405_1, new_n10406, new_n10408, new_n10409_1,
    new_n10410, new_n10411_1, new_n10412, new_n10413, new_n10414,
    new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420_1, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432_1, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476, new_n10477,
    new_n10478, new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484_1, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489_1, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505,
    new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514_1, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525_1, new_n10526, new_n10527,
    new_n10528, new_n10529, new_n10530, new_n10531, new_n10532, new_n10533,
    new_n10534, new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540_1, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561_1,
    new_n10562, new_n10563, new_n10564_1, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588_1, new_n10589, new_n10593_1, new_n10594, new_n10595_1,
    new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601,
    new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607,
    new_n10608, new_n10609, new_n10610, new_n10611_1, new_n10612,
    new_n10613, new_n10614_1, new_n10615, new_n10616, new_n10617_1,
    new_n10618, new_n10619, new_n10620, new_n10623, new_n10624, new_n10625,
    new_n10626, new_n10627, new_n10628_1, new_n10629, new_n10630,
    new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636,
    new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642,
    new_n10643, new_n10644, new_n10645, new_n10646, new_n10647_1,
    new_n10648, new_n10649, new_n10650_1, new_n10651, new_n10652,
    new_n10653_1, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692_1,
    new_n10693, new_n10694_1, new_n10695, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10701_1, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710_1, new_n10711, new_n10712_1, new_n10713,
    new_n10714, new_n10715, new_n10716, new_n10717, new_n10718, new_n10719,
    new_n10720, new_n10721, new_n10722, new_n10723, new_n10724, new_n10725,
    new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731,
    new_n10732, new_n10733, new_n10734, new_n10735, new_n10736, new_n10737,
    new_n10738, new_n10739_1, new_n10740, new_n10741, new_n10742,
    new_n10743, new_n10744, new_n10745, new_n10746, new_n10747, new_n10748,
    new_n10749, new_n10750, new_n10751, new_n10752, new_n10753, new_n10754,
    new_n10755, new_n10756_1, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763_1, new_n10764,
    new_n10765, new_n10768, new_n10769, new_n10770, new_n10771, new_n10772,
    new_n10773, new_n10774, new_n10775_1, new_n10776, new_n10777,
    new_n10778, new_n10779, new_n10780_1, new_n10781, new_n10782,
    new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788,
    new_n10789, new_n10790, new_n10791, new_n10792_1, new_n10793,
    new_n10794, new_n10795, new_n10796, new_n10797, new_n10798, new_n10799,
    new_n10800, new_n10801, new_n10802, new_n10803, new_n10804, new_n10805,
    new_n10806, new_n10807, new_n10808, new_n10809, new_n10810, new_n10811,
    new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817_1, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834_1, new_n10835, new_n10836, new_n10837, new_n10838,
    new_n10839, new_n10840, new_n10841, new_n10842, new_n10843, new_n10844,
    new_n10845, new_n10846, new_n10847, new_n10848, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874_1, new_n10875, new_n10876, new_n10877, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903,
    new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909,
    new_n10910, new_n10911, new_n10912, new_n10913, new_n10914, new_n10915,
    new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921,
    new_n10922, new_n10923, new_n10924_1, new_n10925, new_n10926,
    new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943_1,
    new_n10944, new_n10945, new_n10946, new_n10947, new_n10948, new_n10949,
    new_n10950, new_n10951, new_n10952, new_n10953, new_n10954, new_n10955,
    new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961_1, new_n10962, new_n10963, new_n10964, new_n10965,
    new_n10966, new_n10967, new_n10968, new_n10969, new_n10970, new_n10971,
    new_n10972, new_n10973, new_n10974, new_n10975, new_n10976, new_n10977,
    new_n10978, new_n10979, new_n10980, new_n10981, new_n10982, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005_1, new_n11006, new_n11007,
    new_n11008, new_n11009, new_n11010, new_n11011_1, new_n11012,
    new_n11013, new_n11017, new_n11018, new_n11019, new_n11020, new_n11021,
    new_n11022, new_n11023_1, new_n11024, new_n11025_1, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043,
    new_n11044_1, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056_1, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063_1, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078_1, new_n11079, new_n11080_1, new_n11081,
    new_n11082, new_n11085, new_n11086, new_n11087, new_n11088, new_n11089,
    new_n11090, new_n11091, new_n11092, new_n11093, new_n11094_1,
    new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101_1, new_n11102, new_n11103_1, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120_1, new_n11121_1, new_n11122,
    new_n11123, new_n11124, new_n11125, new_n11126, new_n11127_1,
    new_n11128, new_n11129, new_n11130, new_n11131, new_n11132_1,
    new_n11133, new_n11134_1, new_n11135, new_n11136, new_n11137,
    new_n11138_1, new_n11139, new_n11140, new_n11141, new_n11142,
    new_n11143, new_n11144, new_n11145, new_n11146, new_n11147, new_n11148,
    new_n11149, new_n11150, new_n11151, new_n11152, new_n11153, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182_1, new_n11183,
    new_n11184_1, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192_1, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201_1, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220_1, new_n11221,
    new_n11222, new_n11223_1, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234_1, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245_1, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254,
    new_n11255, new_n11256, new_n11257, new_n11258, new_n11259, new_n11260,
    new_n11261_1, new_n11262, new_n11263, new_n11264, new_n11265,
    new_n11266_1, new_n11267, new_n11268, new_n11269, new_n11270,
    new_n11271, new_n11272, new_n11273_1, new_n11274, new_n11275_1,
    new_n11276, new_n11277, new_n11278, new_n11279, new_n11280, new_n11281,
    new_n11282, new_n11283, new_n11284, new_n11285, new_n11286, new_n11287,
    new_n11288, new_n11289, new_n11290_1, new_n11291, new_n11292,
    new_n11293, new_n11294, new_n11295, new_n11296, new_n11297, new_n11298,
    new_n11299, new_n11300, new_n11301, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313_1, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325_1, new_n11326_1, new_n11327, new_n11328,
    new_n11329, new_n11330_1, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11339, new_n11340,
    new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346,
    new_n11347_1, new_n11348_1, new_n11349, new_n11350, new_n11351,
    new_n11352_1, new_n11353, new_n11354, new_n11355, new_n11356_1,
    new_n11357, new_n11358, new_n11359, new_n11360, new_n11361, new_n11362,
    new_n11363, new_n11364, new_n11365, new_n11366, new_n11367, new_n11368,
    new_n11369, new_n11370, new_n11371, new_n11372, new_n11373, new_n11374,
    new_n11375_1, new_n11376, new_n11377, new_n11378, new_n11379_1,
    new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385,
    new_n11386_1, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391_1, new_n11392, new_n11393, new_n11394, new_n11395,
    new_n11396, new_n11397, new_n11398_1, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403_1, new_n11404, new_n11405,
    new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11411,
    new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11417,
    new_n11418, new_n11419_1, new_n11420, new_n11421, new_n11422,
    new_n11423, new_n11424_1, new_n11425, new_n11426, new_n11427,
    new_n11428, new_n11429, new_n11430, new_n11431, new_n11432, new_n11433,
    new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439_1, new_n11440, new_n11441, new_n11442, new_n11443,
    new_n11444, new_n11445, new_n11446, new_n11447, new_n11448, new_n11449,
    new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455_1, new_n11456, new_n11457, new_n11458, new_n11459,
    new_n11460, new_n11461, new_n11462_1, new_n11463, new_n11464,
    new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470_1, new_n11471, new_n11472_1, new_n11473_1, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479_1,
    new_n11480, new_n11481_1, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486_1, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496_1, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503_1, new_n11504, new_n11505,
    new_n11506_1, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515_1,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537, new_n11538_1,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548_1, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564_1, new_n11565, new_n11566_1,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579_1, new_n11580_1, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589,
    new_n11590, new_n11591_1, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607_1, new_n11608, new_n11609, new_n11610, new_n11611,
    new_n11612, new_n11613, new_n11614, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627, new_n11628, new_n11629, new_n11630_1,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647_1,
    new_n11648, new_n11649, new_n11650, new_n11651, new_n11652, new_n11653,
    new_n11654, new_n11655, new_n11656, new_n11657, new_n11658, new_n11659,
    new_n11660, new_n11661, new_n11662, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667_1, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674_1, new_n11679,
    new_n11680, new_n11681, new_n11682_1, new_n11683, new_n11684,
    new_n11685, new_n11686, new_n11687, new_n11688, new_n11689, new_n11690,
    new_n11691, new_n11692, new_n11693, new_n11694, new_n11698, new_n11699,
    new_n11700, new_n11701, new_n11702, new_n11703, new_n11704, new_n11705,
    new_n11706, new_n11707, new_n11708, new_n11709, new_n11710_1,
    new_n11711, new_n11712_1, new_n11713, new_n11714, new_n11715,
    new_n11716, new_n11717, new_n11721, new_n11722, new_n11723,
    new_n11724_1, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736_1, new_n11737, new_n11738, new_n11739,
    new_n11740, new_n11741_1, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11750, new_n11751,
    new_n11752, new_n11753, new_n11754, new_n11755, new_n11756, new_n11757,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770_1, new_n11771_1, new_n11772, new_n11773, new_n11774,
    new_n11775_1, new_n11779, new_n11780, new_n11781, new_n11782,
    new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788,
    new_n11789, new_n11790, new_n11791, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837_1,
    new_n11838, new_n11839, new_n11840, new_n11841_1, new_n11842_1,
    new_n11843_1, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898_1, new_n11899, new_n11900,
    new_n11901, new_n11902, new_n11903, new_n11904, new_n11905_1,
    new_n11906, new_n11907, new_n11908, new_n11909, new_n11910, new_n11911,
    new_n11912, new_n11913, new_n11914, new_n11915, new_n11916, new_n11917,
    new_n11918, new_n11919, new_n11920, new_n11921, new_n11922, new_n11923,
    new_n11925, new_n11926_1, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964,
    new_n11965_1, new_n11966, new_n11967, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980_1,
    new_n11981, new_n11982, new_n11983, new_n11984, new_n11985, new_n11986,
    new_n11987, new_n11988, new_n11989, new_n11990, new_n11991, new_n11992,
    new_n11993, new_n11994, new_n11995, new_n11996, new_n11997, new_n11998,
    new_n11999, new_n12000_1, new_n12001, new_n12002, new_n12003_1,
    new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011_1, new_n12012, new_n12013, new_n12014,
    new_n12015, new_n12016, new_n12017, new_n12018, new_n12019, new_n12020,
    new_n12021, new_n12022, new_n12023, new_n12024, new_n12025, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12042, new_n12043, new_n12044, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068, new_n12071,
    new_n12072_1, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12078, new_n12079, new_n12080, new_n12081, new_n12082, new_n12083,
    new_n12084, new_n12085, new_n12086, new_n12087, new_n12088, new_n12089,
    new_n12090, new_n12091, new_n12092, new_n12093, new_n12094, new_n12095,
    new_n12096, new_n12097, new_n12098, new_n12099, new_n12100, new_n12101,
    new_n12102, new_n12103, new_n12104, new_n12105, new_n12106, new_n12107,
    new_n12108, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113_1, new_n12114, new_n12115, new_n12116, new_n12117,
    new_n12118, new_n12119, new_n12120, new_n12121_1, new_n12122,
    new_n12123, new_n12124, new_n12125, new_n12126, new_n12127, new_n12128,
    new_n12129, new_n12130, new_n12131_1, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145,
    new_n12146_1, new_n12147, new_n12148, new_n12149, new_n12150,
    new_n12151, new_n12152_1, new_n12153_1, new_n12154, new_n12155,
    new_n12156, new_n12157_1, new_n12158_1, new_n12159, new_n12160,
    new_n12161_1, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166, new_n12167, new_n12168, new_n12169, new_n12170, new_n12171,
    new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177,
    new_n12178, new_n12179_1, new_n12180, new_n12181, new_n12182,
    new_n12183, new_n12184, new_n12185, new_n12186, new_n12187, new_n12188,
    new_n12189, new_n12190, new_n12191, new_n12192_1, new_n12193,
    new_n12194, new_n12195, new_n12196, new_n12197, new_n12198, new_n12199,
    new_n12200, new_n12201, new_n12202, new_n12203, new_n12204, new_n12205,
    new_n12206, new_n12207, new_n12208, new_n12209_1, new_n12210,
    new_n12211, new_n12212, new_n12213, new_n12214, new_n12215, new_n12216,
    new_n12217, new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223_1, new_n12224, new_n12225_1, new_n12226, new_n12227,
    new_n12228_1, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235_1, new_n12238, new_n12239,
    new_n12240, new_n12241, new_n12242, new_n12243, new_n12244, new_n12245,
    new_n12246, new_n12247, new_n12248, new_n12249, new_n12250, new_n12251,
    new_n12252, new_n12253, new_n12254, new_n12255, new_n12256, new_n12257,
    new_n12258, new_n12259, new_n12260, new_n12261, new_n12262, new_n12263,
    new_n12264, new_n12265, new_n12266, new_n12267, new_n12268, new_n12269,
    new_n12270, new_n12271, new_n12272, new_n12273, new_n12274, new_n12275,
    new_n12276, new_n12277, new_n12278, new_n12279, new_n12280, new_n12281,
    new_n12282, new_n12283, new_n12284, new_n12285, new_n12286, new_n12287,
    new_n12288, new_n12289, new_n12290, new_n12291, new_n12292, new_n12293,
    new_n12294, new_n12295, new_n12296, new_n12297, new_n12298, new_n12299,
    new_n12300, new_n12301, new_n12302_1, new_n12303, new_n12304_1,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12311,
    new_n12312, new_n12313, new_n12314, new_n12315_1, new_n12316,
    new_n12317, new_n12320, new_n12321, new_n12322, new_n12323,
    new_n12324_1, new_n12325_1, new_n12326, new_n12327, new_n12328,
    new_n12329_1, new_n12330_1, new_n12331, new_n12332, new_n12333,
    new_n12334, new_n12335, new_n12336, new_n12337, new_n12338, new_n12339,
    new_n12340, new_n12341_1, new_n12342, new_n12343, new_n12344,
    new_n12345, new_n12346_1, new_n12347, new_n12348, new_n12349_1,
    new_n12350, new_n12351, new_n12352, new_n12353, new_n12354, new_n12355,
    new_n12356, new_n12357, new_n12358, new_n12359, new_n12360, new_n12361,
    new_n12362, new_n12363, new_n12364_1, new_n12365, new_n12366,
    new_n12367, new_n12368, new_n12369, new_n12370, new_n12371, new_n12372,
    new_n12373, new_n12374, new_n12375, new_n12376, new_n12377, new_n12378,
    new_n12379, new_n12380_1, new_n12381, new_n12382, new_n12383_1,
    new_n12384_1, new_n12385, new_n12386, new_n12387, new_n12388,
    new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394,
    new_n12395, new_n12396, new_n12397_1, new_n12398_1, new_n12399,
    new_n12401, new_n12402, new_n12403, new_n12404, new_n12405, new_n12406,
    new_n12407, new_n12408_1, new_n12409, new_n12410, new_n12411,
    new_n12412, new_n12413, new_n12414, new_n12415, new_n12416, new_n12417,
    new_n12418, new_n12419, new_n12420, new_n12421, new_n12422, new_n12423,
    new_n12424, new_n12425, new_n12426, new_n12427, new_n12428, new_n12429,
    new_n12430, new_n12431, new_n12432, new_n12433, new_n12434, new_n12435,
    new_n12436, new_n12437, new_n12438, new_n12439, new_n12440, new_n12441,
    new_n12442, new_n12443, new_n12444, new_n12445, new_n12446_1,
    new_n12447, new_n12448, new_n12449_1, new_n12450, new_n12451,
    new_n12452, new_n12453, new_n12454, new_n12455, new_n12456, new_n12457,
    new_n12458, new_n12459, new_n12460, new_n12461_1, new_n12462_1,
    new_n12463, new_n12464, new_n12465, new_n12466, new_n12467_1,
    new_n12468, new_n12469_1, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490,
    new_n12491, new_n12492, new_n12493, new_n12494, new_n12495_1,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506,
    new_n12507_1, new_n12508, new_n12509, new_n12510, new_n12511,
    new_n12512, new_n12515_1, new_n12516_1, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540_1, new_n12541,
    new_n12542, new_n12543, new_n12544, new_n12545_1, new_n12546_1,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552_1, new_n12553, new_n12554, new_n12555, new_n12558,
    new_n12559, new_n12560, new_n12561, new_n12562_1, new_n12563,
    new_n12564, new_n12565, new_n12566_1, new_n12567, new_n12568,
    new_n12569_1, new_n12570, new_n12571, new_n12572, new_n12573,
    new_n12574, new_n12575, new_n12576, new_n12577, new_n12578, new_n12579,
    new_n12580, new_n12581, new_n12582, new_n12583, new_n12584, new_n12585,
    new_n12586, new_n12587_1, new_n12588, new_n12589, new_n12590,
    new_n12591, new_n12592, new_n12593_1, new_n12594, new_n12595,
    new_n12596, new_n12597, new_n12598, new_n12599, new_n12600, new_n12601,
    new_n12602, new_n12603, new_n12604, new_n12605, new_n12606,
    new_n12607_1, new_n12608, new_n12609, new_n12610, new_n12611,
    new_n12612, new_n12613, new_n12614, new_n12615, new_n12616, new_n12617,
    new_n12618, new_n12619, new_n12620_1, new_n12621_1, new_n12622,
    new_n12623, new_n12624, new_n12625, new_n12626_1, new_n12627,
    new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648, new_n12649, new_n12650_1,
    new_n12651, new_n12652, new_n12653, new_n12654_1, new_n12655,
    new_n12656, new_n12657_1, new_n12658, new_n12659, new_n12660,
    new_n12661, new_n12662, new_n12663, new_n12664, new_n12665_1,
    new_n12666, new_n12667, new_n12668, new_n12669, new_n12670_1,
    new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676,
    new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682,
    new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688,
    new_n12689, new_n12690, new_n12691, new_n12693, new_n12694, new_n12695,
    new_n12696, new_n12697, new_n12698, new_n12699, new_n12700, new_n12701,
    new_n12702_1, new_n12703, new_n12704, new_n12705, new_n12706,
    new_n12707_1, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12720, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725_1, new_n12726, new_n12727_1, new_n12728, new_n12729,
    new_n12730, new_n12731, new_n12732, new_n12733, new_n12734, new_n12735,
    new_n12736, new_n12737, new_n12738, new_n12739, new_n12740_1,
    new_n12741, new_n12742_1, new_n12743, new_n12744, new_n12745,
    new_n12746_1, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753, new_n12754, new_n12755,
    new_n12756_1, new_n12757, new_n12758, new_n12759, new_n12760,
    new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766,
    new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772,
    new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783_1,
    new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789,
    new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795,
    new_n12796, new_n12797, new_n12798, new_n12799, new_n12800,
    new_n12801_1, new_n12802, new_n12803, new_n12804, new_n12805,
    new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811_1, new_n12812_1, new_n12813, new_n12814, new_n12815,
    new_n12816_1, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821_1, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837,
    new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843_1, new_n12844, new_n12845, new_n12846, new_n12847,
    new_n12848, new_n12849, new_n12850, new_n12851, new_n12852, new_n12853,
    new_n12854, new_n12855, new_n12856, new_n12857, new_n12858, new_n12859,
    new_n12860, new_n12861_1, new_n12862, new_n12863, new_n12864_1,
    new_n12865_1, new_n12866, new_n12867, new_n12868, new_n12869,
    new_n12870_1, new_n12871_1, new_n12872, new_n12873_1, new_n12874,
    new_n12875_1, new_n12876, new_n12877, new_n12878, new_n12879,
    new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892_1, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12898, new_n12899, new_n12900_1, new_n12901, new_n12902,
    new_n12903, new_n12904_1, new_n12905, new_n12906, new_n12907,
    new_n12908, new_n12909, new_n12910, new_n12911, new_n12912, new_n12913,
    new_n12914, new_n12915, new_n12916, new_n12917_1, new_n12918,
    new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924,
    new_n12925, new_n12926, new_n12927, new_n12928, new_n12929, new_n12930,
    new_n12931, new_n12932, new_n12933, new_n12934, new_n12935, new_n12936,
    new_n12937, new_n12938, new_n12939, new_n12940, new_n12941_1,
    new_n12942_1, new_n12943, new_n12944, new_n12945, new_n12946,
    new_n12947, new_n12948, new_n12949, new_n12950, new_n12951, new_n12952,
    new_n12953, new_n12954, new_n12955, new_n12956_1, new_n12957,
    new_n12958, new_n12959, new_n12960, new_n12961, new_n12962, new_n12963,
    new_n12964, new_n12965, new_n12966, new_n12967, new_n12968, new_n12969,
    new_n12970, new_n12971, new_n12972, new_n12973, new_n12974, new_n12975,
    new_n12976, new_n12977, new_n12978_1, new_n12979, new_n12980_1,
    new_n12981, new_n12982, new_n12983, new_n12984, new_n12985_1,
    new_n12986, new_n12987_1, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992_1, new_n12993, new_n12994, new_n12995,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002, new_n13003, new_n13004, new_n13005_1, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026_1, new_n13027, new_n13028, new_n13029,
    new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043_1, new_n13044_1, new_n13045, new_n13047,
    new_n13048_1, new_n13049, new_n13050, new_n13051, new_n13052,
    new_n13053, new_n13054_1, new_n13055, new_n13056, new_n13057,
    new_n13058, new_n13059, new_n13060, new_n13061, new_n13062, new_n13063,
    new_n13064, new_n13065, new_n13066, new_n13067, new_n13068, new_n13069,
    new_n13070, new_n13071, new_n13072, new_n13073, new_n13074_1,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082_1, new_n13083, new_n13084, new_n13085,
    new_n13086, new_n13087, new_n13088, new_n13089, new_n13090, new_n13091,
    new_n13092, new_n13093, new_n13094, new_n13095, new_n13096_1,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110_1, new_n13111, new_n13112, new_n13113,
    new_n13114, new_n13115, new_n13116_1, new_n13117, new_n13118,
    new_n13119, new_n13120, new_n13121, new_n13122_1, new_n13123,
    new_n13124, new_n13125, new_n13126, new_n13127, new_n13128, new_n13129,
    new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135,
    new_n13136, new_n13137_1, new_n13138, new_n13139, new_n13140,
    new_n13141_1, new_n13142, new_n13143, new_n13144_1, new_n13145,
    new_n13146, new_n13147, new_n13148, new_n13149, new_n13150, new_n13151,
    new_n13152, new_n13153, new_n13154, new_n13155, new_n13156, new_n13157,
    new_n13158, new_n13159, new_n13160, new_n13161, new_n13162, new_n13163,
    new_n13164, new_n13165, new_n13166, new_n13167, new_n13168_1,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13187,
    new_n13188, new_n13189, new_n13190_1, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197,
    new_n13198_1, new_n13199_1, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13204_1, new_n13205, new_n13206, new_n13207,
    new_n13208, new_n13209_1, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263_1, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270_1,
    new_n13271, new_n13272, new_n13273_1, new_n13274, new_n13275,
    new_n13276, new_n13277, new_n13278, new_n13279, new_n13280, new_n13281,
    new_n13282, new_n13283, new_n13284, new_n13285_1, new_n13286,
    new_n13287, new_n13288, new_n13289, new_n13291, new_n13292, new_n13293,
    new_n13294, new_n13295, new_n13296, new_n13297, new_n13298, new_n13299,
    new_n13300, new_n13301, new_n13302, new_n13303, new_n13304, new_n13305,
    new_n13306, new_n13307, new_n13308, new_n13309, new_n13310, new_n13311,
    new_n13312, new_n13313, new_n13314, new_n13315, new_n13316, new_n13317,
    new_n13318, new_n13319_1, new_n13320, new_n13321, new_n13322,
    new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328,
    new_n13329, new_n13330, new_n13331, new_n13332, new_n13333_1,
    new_n13334, new_n13335, new_n13336, new_n13337, new_n13338_1,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367_1, new_n13368, new_n13369,
    new_n13370, new_n13371, new_n13372, new_n13373, new_n13374, new_n13375,
    new_n13376, new_n13377, new_n13378, new_n13379, new_n13380, new_n13381,
    new_n13382, new_n13383, new_n13384, new_n13385, new_n13386, new_n13387,
    new_n13388, new_n13389, new_n13390, new_n13391, new_n13392, new_n13393,
    new_n13394, new_n13395, new_n13396, new_n13397, new_n13398, new_n13399,
    new_n13400, new_n13401, new_n13402, new_n13403, new_n13404, new_n13405,
    new_n13406, new_n13407_1, new_n13408, new_n13409_1, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419_1, new_n13420, new_n13421,
    new_n13422, new_n13423, new_n13424_1, new_n13425, new_n13426,
    new_n13427, new_n13428, new_n13429, new_n13430, new_n13431, new_n13432,
    new_n13433, new_n13434, new_n13435, new_n13436, new_n13437, new_n13438,
    new_n13439, new_n13440, new_n13441, new_n13442, new_n13443, new_n13444,
    new_n13445, new_n13446, new_n13447, new_n13448, new_n13449, new_n13450,
    new_n13451, new_n13452, new_n13453_1, new_n13454, new_n13455,
    new_n13456_1, new_n13457_1, new_n13458, new_n13459, new_n13460_1,
    new_n13461, new_n13462, new_n13463, new_n13464, new_n13465, new_n13466,
    new_n13467, new_n13468, new_n13469, new_n13470, new_n13471, new_n13472,
    new_n13473, new_n13474, new_n13475, new_n13476, new_n13477_1,
    new_n13478, new_n13479, new_n13480, new_n13481, new_n13482, new_n13483,
    new_n13484_1, new_n13485, new_n13487_1, new_n13488, new_n13489,
    new_n13490_1, new_n13491, new_n13492, new_n13493, new_n13494_1,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499,
    new_n13500_1, new_n13501_1, new_n13502, new_n13503, new_n13504,
    new_n13505, new_n13506_1, new_n13507, new_n13508, new_n13509,
    new_n13510, new_n13511, new_n13512, new_n13513, new_n13514, new_n13515,
    new_n13516, new_n13517, new_n13518, new_n13519, new_n13520, new_n13521,
    new_n13522, new_n13523, new_n13524, new_n13525, new_n13526, new_n13527,
    new_n13528, new_n13529, new_n13530, new_n13531, new_n13532, new_n13533,
    new_n13534, new_n13535, new_n13536, new_n13537, new_n13538, new_n13539,
    new_n13540, new_n13541, new_n13542, new_n13543, new_n13544, new_n13545,
    new_n13546, new_n13547, new_n13548_1, new_n13549_1, new_n13550,
    new_n13551_1, new_n13552, new_n13553, new_n13554, new_n13555,
    new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561,
    new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13596,
    new_n13599, new_n13600, new_n13601, new_n13603, new_n13604, new_n13605,
    new_n13606, new_n13607, new_n13608, new_n13609, new_n13610, new_n13611,
    new_n13612, new_n13613, new_n13614, new_n13615, new_n13616, new_n13617,
    new_n13618, new_n13619, new_n13620, new_n13621, new_n13622, new_n13623,
    new_n13624, new_n13625, new_n13626_1, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13634, new_n13635, new_n13636,
    new_n13637, new_n13638, new_n13639, new_n13640, new_n13641, new_n13642,
    new_n13643, new_n13644, new_n13645, new_n13646, new_n13647, new_n13648,
    new_n13649, new_n13650, new_n13651, new_n13652, new_n13653, new_n13654,
    new_n13655, new_n13656, new_n13657, new_n13658, new_n13659, new_n13660,
    new_n13661, new_n13662, new_n13663, new_n13664, new_n13665, new_n13666,
    new_n13667, new_n13668_1, new_n13669, new_n13670, new_n13671,
    new_n13672, new_n13673, new_n13674, new_n13675, new_n13676,
    new_n13677_1, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683_1, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13704, new_n13705, new_n13706, new_n13707, new_n13708_1,
    new_n13709, new_n13710_1, new_n13711, new_n13712, new_n13713,
    new_n13714_1, new_n13715, new_n13716, new_n13717, new_n13718,
    new_n13719_1, new_n13720, new_n13721, new_n13722_1, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13727, new_n13728, new_n13729,
    new_n13730, new_n13731, new_n13732, new_n13733, new_n13734, new_n13735,
    new_n13736, new_n13737, new_n13738, new_n13739, new_n13740, new_n13741,
    new_n13742, new_n13743, new_n13744, new_n13745, new_n13746, new_n13747,
    new_n13748, new_n13749, new_n13750, new_n13751, new_n13752, new_n13753,
    new_n13754_1, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763,
    new_n13764_1, new_n13765, new_n13766, new_n13767, new_n13768,
    new_n13769, new_n13770, new_n13771, new_n13772, new_n13773, new_n13774,
    new_n13775_1, new_n13776, new_n13777, new_n13778, new_n13779,
    new_n13780, new_n13781_1, new_n13782, new_n13783_1, new_n13784,
    new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790,
    new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798_1, new_n13799, new_n13800, new_n13801,
    new_n13802, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807,
    new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813,
    new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819,
    new_n13820, new_n13821, new_n13822, new_n13825, new_n13826, new_n13827,
    new_n13828, new_n13829, new_n13830, new_n13831, new_n13832, new_n13833,
    new_n13834, new_n13835_1, new_n13836, new_n13837, new_n13838,
    new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844,
    new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850_1, new_n13851_1, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872,
    new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878,
    new_n13879, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13913, new_n13914_1, new_n13915, new_n13916,
    new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922_1, new_n13923_1, new_n13924, new_n13925, new_n13926,
    new_n13927, new_n13928, new_n13929, new_n13930, new_n13931, new_n13932,
    new_n13933, new_n13934, new_n13935, new_n13936, new_n13937, new_n13938,
    new_n13939, new_n13940, new_n13941, new_n13942, new_n13943, new_n13944,
    new_n13945, new_n13946, new_n13947, new_n13948, new_n13949, new_n13950,
    new_n13951_1, new_n13953, new_n13954, new_n13955, new_n13956,
    new_n13957, new_n13958, new_n13959, new_n13960, new_n13961, new_n13962,
    new_n13963, new_n13964, new_n13965, new_n13966, new_n13967, new_n13968,
    new_n13969, new_n13970, new_n13971, new_n13972, new_n13973, new_n13974,
    new_n13975, new_n13976, new_n13977, new_n13978, new_n13979, new_n13980,
    new_n13981, new_n13982, new_n13983, new_n13984, new_n13985, new_n13986,
    new_n13987, new_n13988, new_n13989, new_n13990, new_n13991, new_n13992,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004_1,
    new_n14005, new_n14006, new_n14007, new_n14008, new_n14009, new_n14010,
    new_n14011, new_n14012, new_n14013, new_n14014, new_n14015, new_n14016,
    new_n14017, new_n14018, new_n14019, new_n14020, new_n14021, new_n14022,
    new_n14023, new_n14024, new_n14025, new_n14026, new_n14027, new_n14028,
    new_n14029, new_n14030, new_n14031, new_n14032, new_n14033, new_n14034,
    new_n14035, new_n14036_1, new_n14037, new_n14038, new_n14039,
    new_n14040, new_n14041, new_n14042, new_n14043, new_n14044, new_n14045,
    new_n14046, new_n14047, new_n14048, new_n14049, new_n14050, new_n14051,
    new_n14052, new_n14053, new_n14054, new_n14055, new_n14056, new_n14057,
    new_n14058, new_n14059_1, new_n14060, new_n14061, new_n14062,
    new_n14063, new_n14064, new_n14065, new_n14066, new_n14067, new_n14068,
    new_n14069, new_n14070, new_n14071_1, new_n14072, new_n14073,
    new_n14074, new_n14075, new_n14076, new_n14077, new_n14078, new_n14079,
    new_n14080, new_n14081_1, new_n14082, new_n14083, new_n14084,
    new_n14085, new_n14086, new_n14087, new_n14088, new_n14089,
    new_n14090_1, new_n14091, new_n14092, new_n14093, new_n14094,
    new_n14095_1, new_n14096, new_n14097, new_n14098, new_n14099,
    new_n14100, new_n14101, new_n14102, new_n14103, new_n14104, new_n14105,
    new_n14106, new_n14107_1, new_n14108, new_n14109, new_n14110,
    new_n14111, new_n14112, new_n14113, new_n14114, new_n14115, new_n14116,
    new_n14117, new_n14118, new_n14119, new_n14120, new_n14121_1,
    new_n14122, new_n14123, new_n14124, new_n14125, new_n14126_1,
    new_n14127, new_n14128, new_n14129, new_n14130_1, new_n14131,
    new_n14132, new_n14133, new_n14134, new_n14135, new_n14136_1,
    new_n14137, new_n14138, new_n14139, new_n14140, new_n14141, new_n14142,
    new_n14143, new_n14144, new_n14145, new_n14146, new_n14147_1,
    new_n14148_1, new_n14149, new_n14150, new_n14151, new_n14152,
    new_n14153, new_n14154, new_n14155, new_n14156, new_n14157, new_n14158,
    new_n14159, new_n14160, new_n14165, new_n14166, new_n14167, new_n14168,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173,
    new_n14174_1, new_n14175, new_n14176, new_n14177, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190_1, new_n14191,
    new_n14192, new_n14193, new_n14194, new_n14195, new_n14196, new_n14197,
    new_n14198, new_n14199, new_n14200, new_n14201, new_n14202, new_n14203,
    new_n14204, new_n14205, new_n14206, new_n14207, new_n14208, new_n14209,
    new_n14210, new_n14211_1, new_n14212, new_n14213, new_n14214,
    new_n14215, new_n14216, new_n14217, new_n14218, new_n14219, new_n14220,
    new_n14221, new_n14222_1, new_n14223, new_n14224, new_n14225,
    new_n14226, new_n14227, new_n14228, new_n14229, new_n14230_1,
    new_n14231, new_n14232, new_n14233, new_n14234, new_n14235, new_n14236,
    new_n14237, new_n14238, new_n14239, new_n14240, new_n14241, new_n14242,
    new_n14243, new_n14244, new_n14245, new_n14246, new_n14247, new_n14248,
    new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254,
    new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260,
    new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267_1, new_n14268, new_n14269, new_n14270, new_n14271_1,
    new_n14272, new_n14273, new_n14276, new_n14277_1, new_n14278,
    new_n14279, new_n14280, new_n14281, new_n14282, new_n14283, new_n14284,
    new_n14285, new_n14286, new_n14287, new_n14288, new_n14289, new_n14290,
    new_n14291, new_n14292, new_n14293, new_n14294_1, new_n14295,
    new_n14296, new_n14297, new_n14298, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310_1, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14322, new_n14323_1, new_n14324, new_n14325, new_n14326_1,
    new_n14327, new_n14328, new_n14329, new_n14330, new_n14331, new_n14332,
    new_n14333, new_n14334, new_n14335, new_n14336, new_n14337, new_n14338,
    new_n14339, new_n14340, new_n14341, new_n14342_1, new_n14343,
    new_n14344, new_n14345_1, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353_1,
    new_n14354, new_n14355, new_n14356, new_n14357, new_n14358, new_n14359,
    new_n14360, new_n14361, new_n14362, new_n14364_1, new_n14365,
    new_n14366, new_n14367, new_n14368, new_n14369, new_n14370, new_n14371,
    new_n14372, new_n14373, new_n14374, new_n14375_1, new_n14376,
    new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382,
    new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388,
    new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394,
    new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400,
    new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406,
    new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412_1, new_n14413, new_n14414_1, new_n14415, new_n14416,
    new_n14417, new_n14418, new_n14419, new_n14420, new_n14421, new_n14422,
    new_n14423, new_n14424, new_n14425, new_n14426, new_n14427, new_n14428,
    new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440_1, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457_1, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464_1, new_n14465, new_n14466,
    new_n14467, new_n14468, new_n14469, new_n14470, new_n14471_1,
    new_n14472, new_n14473, new_n14474, new_n14475_1, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510_1, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14532, new_n14533, new_n14534, new_n14535, new_n14536,
    new_n14537, new_n14538, new_n14539, new_n14540, new_n14541_1,
    new_n14542, new_n14543, new_n14544, new_n14545, new_n14546_1,
    new_n14547_1, new_n14548, new_n14549, new_n14550, new_n14551,
    new_n14552, new_n14553, new_n14554, new_n14555, new_n14556, new_n14557,
    new_n14558, new_n14559, new_n14560, new_n14561, new_n14562, new_n14563,
    new_n14564, new_n14565, new_n14566, new_n14567, new_n14568, new_n14569,
    new_n14570_1, new_n14571, new_n14572, new_n14573, new_n14574,
    new_n14575_1, new_n14576_1, new_n14577, new_n14578, new_n14579,
    new_n14580, new_n14581, new_n14582, new_n14583, new_n14584, new_n14585,
    new_n14586, new_n14587, new_n14588, new_n14589, new_n14590, new_n14591,
    new_n14592, new_n14593_1, new_n14594, new_n14595, new_n14596,
    new_n14597, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602,
    new_n14603_1, new_n14604, new_n14605, new_n14606, new_n14607,
    new_n14608, new_n14609, new_n14610, new_n14611, new_n14612, new_n14613,
    new_n14614, new_n14615, new_n14616, new_n14617, new_n14618, new_n14619,
    new_n14620, new_n14621, new_n14622, new_n14623, new_n14624, new_n14625,
    new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631,
    new_n14632, new_n14633_1, new_n14636_1, new_n14637, new_n14638,
    new_n14639, new_n14640, new_n14641, new_n14642, new_n14643, new_n14644,
    new_n14645, new_n14646, new_n14647, new_n14648, new_n14649, new_n14650,
    new_n14651, new_n14652, new_n14653, new_n14654, new_n14655, new_n14656,
    new_n14657, new_n14658, new_n14659, new_n14660, new_n14661, new_n14662,
    new_n14663, new_n14664, new_n14665, new_n14666, new_n14667, new_n14668,
    new_n14669, new_n14670, new_n14671, new_n14672, new_n14673, new_n14674,
    new_n14675, new_n14676, new_n14677, new_n14678, new_n14679,
    new_n14680_1, new_n14681, new_n14682, new_n14683, new_n14684_1,
    new_n14685, new_n14686, new_n14687, new_n14688, new_n14689, new_n14690,
    new_n14691, new_n14692_1, new_n14693, new_n14694, new_n14695,
    new_n14696, new_n14697, new_n14698, new_n14699, new_n14700,
    new_n14701_1, new_n14702_1, new_n14703, new_n14704_1, new_n14705,
    new_n14706, new_n14707, new_n14708, new_n14709, new_n14710, new_n14711,
    new_n14712, new_n14713, new_n14714, new_n14715, new_n14716, new_n14717,
    new_n14718, new_n14719, new_n14720, new_n14721, new_n14722, new_n14723,
    new_n14724, new_n14725, new_n14726, new_n14727, new_n14728, new_n14729,
    new_n14730, new_n14731, new_n14733, new_n14734_1, new_n14735,
    new_n14736, new_n14737, new_n14738, new_n14739, new_n14740, new_n14741,
    new_n14742, new_n14743, new_n14744, new_n14745, new_n14746_1,
    new_n14747, new_n14748, new_n14749, new_n14750, new_n14751, new_n14752,
    new_n14753, new_n14754, new_n14755, new_n14756, new_n14757, new_n14758,
    new_n14759, new_n14760, new_n14761, new_n14762, new_n14763_1,
    new_n14764, new_n14765, new_n14766, new_n14767, new_n14768, new_n14769,
    new_n14770, new_n14771, new_n14772_1, new_n14773, new_n14774,
    new_n14775, new_n14776, new_n14777, new_n14778, new_n14779, new_n14780,
    new_n14781, new_n14782, new_n14783, new_n14784, new_n14785, new_n14787,
    new_n14788, new_n14789, new_n14790_1, new_n14791, new_n14792,
    new_n14793, new_n14794, new_n14795, new_n14796, new_n14797, new_n14798,
    new_n14799, new_n14800, new_n14801_1, new_n14802, new_n14803,
    new_n14804, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819_1, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826_1, new_n14827_1,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839_1, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14848,
    new_n14849_1, new_n14850, new_n14851, new_n14852, new_n14853,
    new_n14854, new_n14855, new_n14856, new_n14857, new_n14858, new_n14859,
    new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865,
    new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871,
    new_n14872, new_n14873, new_n14874, new_n14875, new_n14876, new_n14877,
    new_n14878, new_n14879, new_n14883, new_n14884, new_n14885, new_n14886,
    new_n14887, new_n14888, new_n14889, new_n14890, new_n14891_1,
    new_n14892, new_n14896, new_n14897, new_n14898, new_n14899_1,
    new_n14900, new_n14901, new_n14902, new_n14903, new_n14904, new_n14905,
    new_n14906, new_n14907, new_n14908, new_n14909, new_n14910, new_n14911,
    new_n14912, new_n14913, new_n14914, new_n14915, new_n14916, new_n14917,
    new_n14918, new_n14919, new_n14922, new_n14923, new_n14924, new_n14925,
    new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931_1, new_n14932, new_n14933, new_n14934, new_n14935,
    new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941,
    new_n14942, new_n14943, new_n14944_1, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954_1, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977_1, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986,
    new_n14987, new_n14988, new_n14989_1, new_n14990, new_n14991,
    new_n14992, new_n14993, new_n14994, new_n14995, new_n14996, new_n14997,
    new_n14998, new_n14999, new_n15000, new_n15001, new_n15002_1,
    new_n15003, new_n15004_1, new_n15005, new_n15006, new_n15007,
    new_n15008, new_n15009, new_n15010, new_n15011_1, new_n15012,
    new_n15013, new_n15014, new_n15015, new_n15016, new_n15017, new_n15018,
    new_n15019_1, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031_1, new_n15035, new_n15036, new_n15037,
    new_n15038, new_n15039, new_n15040, new_n15041, new_n15042, new_n15043,
    new_n15044, new_n15045, new_n15046, new_n15047, new_n15048, new_n15049,
    new_n15050, new_n15051, new_n15052_1, new_n15053_1, new_n15054,
    new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060,
    new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066,
    new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072,
    new_n15073, new_n15074, new_n15075, new_n15076, new_n15077_1,
    new_n15078, new_n15079, new_n15080, new_n15081, new_n15082_1,
    new_n15083, new_n15084, new_n15085, new_n15086, new_n15087, new_n15088,
    new_n15089, new_n15090, new_n15091, new_n15092, new_n15093,
    new_n15094_1, new_n15095, new_n15096, new_n15097, new_n15098,
    new_n15099, new_n15100, new_n15101, new_n15102, new_n15103, new_n15104,
    new_n15105, new_n15106, new_n15107, new_n15108, new_n15109, new_n15110,
    new_n15111, new_n15112, new_n15113, new_n15114, new_n15115, new_n15116,
    new_n15117, new_n15118_1, new_n15119, new_n15120, new_n15121,
    new_n15122, new_n15123, new_n15124, new_n15125, new_n15126, new_n15127,
    new_n15128_1, new_n15129, new_n15130, new_n15131, new_n15132,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139_1, new_n15140, new_n15141, new_n15142, new_n15143,
    new_n15144, new_n15145_1, new_n15146_1, new_n15147, new_n15148,
    new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154,
    new_n15155, new_n15156, new_n15157, new_n15158, new_n15159, new_n15160,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165_1,
    new_n15166, new_n15167_1, new_n15169, new_n15170, new_n15171,
    new_n15172, new_n15173, new_n15174, new_n15175, new_n15176_1,
    new_n15177, new_n15178, new_n15180_1, new_n15181, new_n15182_1,
    new_n15183, new_n15184, new_n15185, new_n15186, new_n15187, new_n15188,
    new_n15189, new_n15190, new_n15191, new_n15192, new_n15193, new_n15194,
    new_n15195, new_n15196, new_n15197, new_n15198, new_n15199, new_n15200,
    new_n15201, new_n15202, new_n15203, new_n15204, new_n15205_1,
    new_n15206, new_n15207, new_n15208, new_n15209, new_n15210, new_n15211,
    new_n15212, new_n15213, new_n15214, new_n15215, new_n15216, new_n15217,
    new_n15218, new_n15220, new_n15221, new_n15222, new_n15223, new_n15224,
    new_n15225, new_n15226, new_n15227, new_n15228, new_n15229,
    new_n15230_1, new_n15231, new_n15232, new_n15233, new_n15234,
    new_n15235, new_n15236, new_n15237, new_n15238, new_n15239, new_n15240,
    new_n15241_1, new_n15242, new_n15243, new_n15244, new_n15245,
    new_n15246, new_n15247, new_n15248, new_n15249, new_n15250, new_n15251,
    new_n15252, new_n15253, new_n15254, new_n15255_1, new_n15256,
    new_n15257, new_n15258_1, new_n15259, new_n15261, new_n15262,
    new_n15263, new_n15264, new_n15265, new_n15266, new_n15267, new_n15268,
    new_n15269, new_n15270, new_n15271_1, new_n15272, new_n15273,
    new_n15274, new_n15275_1, new_n15276, new_n15277, new_n15278,
    new_n15279, new_n15280, new_n15281, new_n15282, new_n15283, new_n15284,
    new_n15285, new_n15286, new_n15287, new_n15288, new_n15289_1,
    new_n15292, new_n15293, new_n15294, new_n15295, new_n15296, new_n15297,
    new_n15298, new_n15299, new_n15300_1, new_n15301, new_n15302,
    new_n15303, new_n15304, new_n15305, new_n15306, new_n15307_1,
    new_n15308, new_n15309, new_n15310, new_n15311, new_n15312, new_n15313,
    new_n15314, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327_1, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332_1, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342,
    new_n15343, new_n15344, new_n15345_1, new_n15346, new_n15347,
    new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353_1, new_n15354, new_n15355, new_n15356, new_n15357,
    new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363,
    new_n15364, new_n15365, new_n15366_1, new_n15367, new_n15368,
    new_n15369, new_n15370, new_n15371, new_n15372, new_n15373, new_n15374,
    new_n15375, new_n15377, new_n15378_1, new_n15379, new_n15380,
    new_n15381, new_n15382_1, new_n15383, new_n15384, new_n15385,
    new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391,
    new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397,
    new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403,
    new_n15404, new_n15405, new_n15406, new_n15407_1, new_n15408,
    new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414,
    new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420,
    new_n15421, new_n15422, new_n15423, new_n15424_1, new_n15425,
    new_n15426, new_n15427, new_n15428_1, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435_1,
    new_n15436, new_n15437, new_n15438_1, new_n15439, new_n15440,
    new_n15441, new_n15442, new_n15443, new_n15444, new_n15445, new_n15446,
    new_n15447, new_n15448, new_n15449, new_n15450, new_n15451, new_n15452,
    new_n15453, new_n15454, new_n15455, new_n15456, new_n15457, new_n15458,
    new_n15459, new_n15460, new_n15461, new_n15462, new_n15463, new_n15464,
    new_n15465_1, new_n15466, new_n15467_1, new_n15468, new_n15469,
    new_n15470_1, new_n15471, new_n15472, new_n15473, new_n15474,
    new_n15475, new_n15476, new_n15477_1, new_n15478, new_n15479,
    new_n15480, new_n15481_1, new_n15482, new_n15483, new_n15484,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489,
    new_n15490_1, new_n15491, new_n15492, new_n15493, new_n15494,
    new_n15495, new_n15496_1, new_n15497, new_n15498, new_n15499,
    new_n15500, new_n15501_1, new_n15502, new_n15503, new_n15504,
    new_n15505, new_n15506_1, new_n15507, new_n15508_1, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527,
    new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534,
    new_n15535, new_n15536, new_n15537, new_n15538, new_n15539_1,
    new_n15540, new_n15541, new_n15542, new_n15545, new_n15546_1,
    new_n15547, new_n15548, new_n15549, new_n15550, new_n15551, new_n15552,
    new_n15553, new_n15554, new_n15555_1, new_n15560, new_n15561,
    new_n15562, new_n15563, new_n15564, new_n15565, new_n15566, new_n15567,
    new_n15568, new_n15569, new_n15570_1, new_n15571, new_n15572,
    new_n15573_1, new_n15580, new_n15581, new_n15582, new_n15583,
    new_n15584, new_n15585, new_n15586, new_n15587, new_n15588_1,
    new_n15589, new_n15590_1, new_n15591, new_n15592, new_n15593,
    new_n15594, new_n15595, new_n15596, new_n15597, new_n15598_1,
    new_n15599, new_n15600, new_n15601, new_n15602_1, new_n15603,
    new_n15604, new_n15605, new_n15606, new_n15607, new_n15608, new_n15609,
    new_n15610, new_n15611, new_n15612, new_n15613, new_n15614_1,
    new_n15615, new_n15616, new_n15617, new_n15618, new_n15619, new_n15620,
    new_n15621, new_n15622, new_n15623, new_n15624, new_n15625, new_n15626,
    new_n15627, new_n15628, new_n15629, new_n15630, new_n15631, new_n15632,
    new_n15633, new_n15634, new_n15635, new_n15636_1, new_n15637,
    new_n15638, new_n15639, new_n15640, new_n15641, new_n15642, new_n15643,
    new_n15644, new_n15645, new_n15646, new_n15647, new_n15648, new_n15649,
    new_n15650, new_n15651, new_n15652_1, new_n15653, new_n15654,
    new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660,
    new_n15661, new_n15662_1, new_n15663, new_n15664, new_n15665,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15714, new_n15715,
    new_n15716_1, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743_1,
    new_n15744, new_n15745, new_n15746, new_n15747, new_n15748,
    new_n15749_1, new_n15750, new_n15751, new_n15752, new_n15753,
    new_n15754, new_n15755, new_n15756, new_n15757, new_n15758, new_n15759,
    new_n15760, new_n15761_1, new_n15762_1, new_n15763, new_n15764,
    new_n15765, new_n15766_1, new_n15767, new_n15768, new_n15769,
    new_n15770, new_n15771, new_n15772, new_n15773, new_n15774, new_n15775,
    new_n15776, new_n15777, new_n15778, new_n15779, new_n15780_1,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793_1, new_n15794, new_n15795, new_n15796, new_n15797,
    new_n15798, new_n15799, new_n15800, new_n15801, new_n15802, new_n15803,
    new_n15804, new_n15805, new_n15806, new_n15807, new_n15808, new_n15809,
    new_n15810, new_n15811, new_n15812_1, new_n15813, new_n15814,
    new_n15815_1, new_n15816_1, new_n15817, new_n15818, new_n15819,
    new_n15820, new_n15821, new_n15822, new_n15823, new_n15824, new_n15825,
    new_n15826, new_n15827, new_n15828, new_n15829, new_n15830,
    new_n15831_1, new_n15832, new_n15833, new_n15834, new_n15835,
    new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841,
    new_n15842, new_n15843, new_n15845, new_n15846_1, new_n15847,
    new_n15848, new_n15849, new_n15850, new_n15851, new_n15852, new_n15853,
    new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859_1, new_n15860, new_n15861, new_n15862, new_n15863,
    new_n15864, new_n15865, new_n15866, new_n15867, new_n15868,
    new_n15869_1, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884_1,
    new_n15885_1, new_n15886, new_n15889_1, new_n15890, new_n15891,
    new_n15892, new_n15893, new_n15894, new_n15895, new_n15896, new_n15897,
    new_n15898, new_n15899, new_n15900, new_n15901, new_n15902, new_n15903,
    new_n15906, new_n15907, new_n15908, new_n15909, new_n15910, new_n15911,
    new_n15912, new_n15913, new_n15914, new_n15918_1, new_n15919,
    new_n15920, new_n15921, new_n15922_1, new_n15923, new_n15924,
    new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930,
    new_n15931, new_n15932, new_n15933, new_n15934, new_n15935,
    new_n15936_1, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947_1, new_n15948, new_n15949, new_n15950, new_n15951,
    new_n15952, new_n15953, new_n15954, new_n15955, new_n15956_1,
    new_n15957, new_n15958_1, new_n15961, new_n15962, new_n15963,
    new_n15964, new_n15965, new_n15966, new_n15967_1, new_n15968,
    new_n15969, new_n15970, new_n15971, new_n15972, new_n15973, new_n15974,
    new_n15975, new_n15976, new_n15977, new_n15978, new_n15979_1,
    new_n15980, new_n15981, new_n15982, new_n15983, new_n15984, new_n15985,
    new_n15986_1, new_n15987, new_n15988, new_n15989, new_n15990,
    new_n15991, new_n15992, new_n15993, new_n15994, new_n15995, new_n15996,
    new_n15997, new_n15998, new_n15999, new_n16000, new_n16001, new_n16002,
    new_n16003, new_n16004, new_n16005, new_n16006, new_n16007, new_n16008,
    new_n16009, new_n16010, new_n16011, new_n16012, new_n16013_1,
    new_n16014, new_n16015, new_n16016, new_n16017, new_n16018, new_n16019,
    new_n16020, new_n16021, new_n16022, new_n16023, new_n16024, new_n16025,
    new_n16026, new_n16027, new_n16028, new_n16029_1, new_n16030,
    new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036,
    new_n16037, new_n16038, new_n16039, new_n16040, new_n16042, new_n16043,
    new_n16044, new_n16045, new_n16046, new_n16047, new_n16048, new_n16049,
    new_n16050, new_n16051, new_n16052, new_n16053, new_n16054, new_n16055,
    new_n16056, new_n16057, new_n16058, new_n16059, new_n16060_1,
    new_n16061, new_n16062_1, new_n16063, new_n16064, new_n16065,
    new_n16066, new_n16067, new_n16068_1, new_n16069, new_n16070,
    new_n16071, new_n16072, new_n16073, new_n16074, new_n16075, new_n16076,
    new_n16077, new_n16078, new_n16079, new_n16080_1, new_n16082,
    new_n16083, new_n16084, new_n16085, new_n16086, new_n16087, new_n16088,
    new_n16089, new_n16090, new_n16091, new_n16092, new_n16093, new_n16094,
    new_n16095, new_n16096, new_n16097, new_n16098_1, new_n16099,
    new_n16100, new_n16101, new_n16102, new_n16103, new_n16104, new_n16105,
    new_n16106, new_n16107, new_n16108, new_n16109, new_n16110_1,
    new_n16111, new_n16112, new_n16113, new_n16114, new_n16115, new_n16116,
    new_n16117, new_n16118, new_n16119, new_n16120, new_n16121, new_n16122,
    new_n16123, new_n16124, new_n16125, new_n16126, new_n16127, new_n16128,
    new_n16129, new_n16130, new_n16131, new_n16132, new_n16133, new_n16134,
    new_n16135, new_n16141, new_n16142_1, new_n16143, new_n16144,
    new_n16145, new_n16146, new_n16147, new_n16148, new_n16149, new_n16150,
    new_n16151, new_n16152, new_n16153, new_n16154, new_n16155, new_n16156,
    new_n16157, new_n16158_1, new_n16159, new_n16160, new_n16161,
    new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167_1, new_n16168, new_n16169, new_n16170, new_n16171,
    new_n16172, new_n16173, new_n16174, new_n16175, new_n16176, new_n16177,
    new_n16178, new_n16179, new_n16180, new_n16181, new_n16182, new_n16183,
    new_n16184, new_n16185_1, new_n16186, new_n16187, new_n16188,
    new_n16189, new_n16190, new_n16191, new_n16192, new_n16193, new_n16194,
    new_n16195, new_n16196_1, new_n16197, new_n16198, new_n16199,
    new_n16200, new_n16201, new_n16202, new_n16205, new_n16206_1,
    new_n16207, new_n16208, new_n16209, new_n16210, new_n16211, new_n16212,
    new_n16213, new_n16214, new_n16215_1, new_n16216, new_n16217_1,
    new_n16218_1, new_n16219_1, new_n16220, new_n16221, new_n16222,
    new_n16223_1, new_n16224, new_n16225, new_n16226, new_n16227,
    new_n16228, new_n16229, new_n16230_1, new_n16233, new_n16234,
    new_n16235, new_n16236, new_n16237, new_n16238, new_n16239, new_n16240,
    new_n16241, new_n16242, new_n16243_1, new_n16244, new_n16245,
    new_n16246, new_n16247_1, new_n16248, new_n16249, new_n16251,
    new_n16256, new_n16257, new_n16258, new_n16259, new_n16260, new_n16261,
    new_n16262, new_n16263, new_n16264, new_n16265, new_n16266, new_n16267,
    new_n16268, new_n16269, new_n16270, new_n16271, new_n16272, new_n16273,
    new_n16274, new_n16275_1, new_n16276, new_n16277, new_n16278,
    new_n16279_1, new_n16280, new_n16281, new_n16282, new_n16283,
    new_n16284, new_n16285, new_n16286, new_n16287, new_n16288, new_n16289,
    new_n16290, new_n16291, new_n16292, new_n16293, new_n16294, new_n16295,
    new_n16296, new_n16297, new_n16298, new_n16299, new_n16300, new_n16301,
    new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307,
    new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313,
    new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319,
    new_n16320, new_n16321, new_n16322_1, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327_1, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350_1, new_n16351, new_n16352,
    new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358,
    new_n16359, new_n16360, new_n16361, new_n16365, new_n16366,
    new_n16367_1, new_n16368, new_n16369, new_n16370, new_n16371,
    new_n16372, new_n16373, new_n16374, new_n16375, new_n16376_1,
    new_n16377, new_n16378, new_n16379_1, new_n16380, new_n16381,
    new_n16382, new_n16383, new_n16384, new_n16385, new_n16386, new_n16387,
    new_n16388, new_n16389, new_n16396_1, new_n16397, new_n16398_1,
    new_n16399, new_n16400, new_n16401, new_n16402, new_n16403, new_n16404,
    new_n16405, new_n16406_1, new_n16407_1, new_n16408, new_n16409,
    new_n16410, new_n16411, new_n16412, new_n16413, new_n16414, new_n16415,
    new_n16416, new_n16417, new_n16418, new_n16419_1, new_n16420,
    new_n16421, new_n16422, new_n16423, new_n16424_1, new_n16425,
    new_n16426, new_n16427, new_n16428_1, new_n16429, new_n16430,
    new_n16431, new_n16432, new_n16433_1, new_n16434, new_n16435,
    new_n16436, new_n16437, new_n16438, new_n16439_1, new_n16440_1,
    new_n16441, new_n16442, new_n16443, new_n16444, new_n16445_1,
    new_n16446, new_n16447, new_n16448, new_n16449, new_n16450, new_n16451,
    new_n16452, new_n16453, new_n16454, new_n16455, new_n16456, new_n16457,
    new_n16458, new_n16459, new_n16460_1, new_n16461, new_n16462,
    new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470,
    new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476_1, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481_1, new_n16482_1, new_n16483, new_n16484, new_n16485,
    new_n16486, new_n16487, new_n16488, new_n16489, new_n16490, new_n16491,
    new_n16492, new_n16493_1, new_n16494, new_n16495, new_n16496,
    new_n16497, new_n16498, new_n16499, new_n16500, new_n16501,
    new_n16502_1, new_n16503, new_n16504, new_n16505, new_n16506_1,
    new_n16507_1, new_n16508, new_n16509, new_n16510, new_n16511,
    new_n16512, new_n16513, new_n16514, new_n16515, new_n16516_1,
    new_n16517_1, new_n16518, new_n16519, new_n16520, new_n16521_1,
    new_n16522, new_n16523, new_n16524_1, new_n16525, new_n16526,
    new_n16527_1, new_n16528, new_n16529, new_n16530, new_n16531,
    new_n16532, new_n16533, new_n16534, new_n16535, new_n16537, new_n16538,
    new_n16539, new_n16540, new_n16541, new_n16542, new_n16543,
    new_n16544_1, new_n16545, new_n16546, new_n16547, new_n16548,
    new_n16549, new_n16550, new_n16551, new_n16552, new_n16553,
    new_n16554_1, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583_1, new_n16584_1, new_n16586, new_n16587, new_n16588,
    new_n16589_1, new_n16590, new_n16591, new_n16592, new_n16593,
    new_n16594, new_n16595, new_n16596_1, new_n16597, new_n16598,
    new_n16599, new_n16600, new_n16601, new_n16602, new_n16603, new_n16604,
    new_n16605, new_n16606, new_n16607, new_n16608_1, new_n16609,
    new_n16610, new_n16611, new_n16612, new_n16613, new_n16614, new_n16615,
    new_n16616, new_n16617_1, new_n16618, new_n16619, new_n16620,
    new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16630_1, new_n16631, new_n16632, new_n16633, new_n16634,
    new_n16635, new_n16636, new_n16637, new_n16638, new_n16639,
    new_n16640_1, new_n16641, new_n16642, new_n16643, new_n16648,
    new_n16649, new_n16650, new_n16651, new_n16652, new_n16653, new_n16654,
    new_n16655, new_n16656_1, new_n16657, new_n16658, new_n16659,
    new_n16660, new_n16661, new_n16662, new_n16663, new_n16664, new_n16665,
    new_n16666, new_n16667, new_n16668, new_n16669, new_n16670, new_n16671,
    new_n16672, new_n16673, new_n16674_1, new_n16675, new_n16676,
    new_n16677, new_n16678, new_n16679, new_n16680, new_n16681,
    new_n16682_1, new_n16683, new_n16684_1, new_n16685, new_n16686,
    new_n16687, new_n16688_1, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16696, new_n16697, new_n16698,
    new_n16699, new_n16700, new_n16702, new_n16703, new_n16704, new_n16705,
    new_n16706, new_n16707, new_n16708, new_n16709, new_n16710, new_n16711,
    new_n16712, new_n16713, new_n16714, new_n16718, new_n16719, new_n16720,
    new_n16721, new_n16722_1, new_n16723, new_n16724, new_n16725,
    new_n16726, new_n16727, new_n16728, new_n16729, new_n16730, new_n16731,
    new_n16732, new_n16733_1, new_n16734, new_n16735, new_n16736,
    new_n16737, new_n16739, new_n16740, new_n16741, new_n16742,
    new_n16743_1, new_n16744, new_n16745, new_n16746, new_n16747,
    new_n16748, new_n16749, new_n16750, new_n16751, new_n16752, new_n16753,
    new_n16754, new_n16755, new_n16756, new_n16757, new_n16758, new_n16759,
    new_n16760, new_n16761, new_n16762, new_n16763, new_n16764, new_n16765,
    new_n16766, new_n16767, new_n16768, new_n16769, new_n16770, new_n16771,
    new_n16772, new_n16773, new_n16774, new_n16775, new_n16776, new_n16777,
    new_n16778, new_n16779, new_n16780, new_n16781, new_n16782, new_n16783,
    new_n16784, new_n16785, new_n16786, new_n16787, new_n16788, new_n16789,
    new_n16790, new_n16791, new_n16792, new_n16793, new_n16794, new_n16795,
    new_n16796, new_n16798_1, new_n16799, new_n16800, new_n16801,
    new_n16802, new_n16803, new_n16804, new_n16805, new_n16806, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812_1, new_n16813,
    new_n16814, new_n16815, new_n16816, new_n16817, new_n16818_1,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823,
    new_n16824_1, new_n16825, new_n16826, new_n16827, new_n16828,
    new_n16829, new_n16830, new_n16831, new_n16832, new_n16833,
    new_n16834_1, new_n16835, new_n16836, new_n16837_1, new_n16838,
    new_n16839, new_n16840, new_n16841_1, new_n16842, new_n16843,
    new_n16844, new_n16845, new_n16846, new_n16847, new_n16848, new_n16849,
    new_n16850, new_n16851, new_n16852, new_n16853, new_n16854, new_n16855,
    new_n16856, new_n16857, new_n16858, new_n16859, new_n16860, new_n16861,
    new_n16862, new_n16863, new_n16864, new_n16865, new_n16866, new_n16867,
    new_n16868, new_n16869, new_n16870, new_n16871, new_n16872, new_n16873,
    new_n16874, new_n16875, new_n16876, new_n16877, new_n16878, new_n16879,
    new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885_1, new_n16886, new_n16887, new_n16888, new_n16889,
    new_n16890, new_n16891, new_n16892, new_n16893, new_n16894, new_n16895,
    new_n16896, new_n16897, new_n16898, new_n16899, new_n16900, new_n16901,
    new_n16902, new_n16903, new_n16904, new_n16905_1, new_n16906,
    new_n16907, new_n16908, new_n16909, new_n16910, new_n16911_1,
    new_n16912, new_n16913, new_n16914, new_n16915, new_n16916, new_n16917,
    new_n16918, new_n16919, new_n16920, new_n16921, new_n16922, new_n16923,
    new_n16924, new_n16925, new_n16926, new_n16927, new_n16928, new_n16929,
    new_n16930, new_n16931, new_n16932, new_n16933, new_n16934, new_n16935,
    new_n16936, new_n16937, new_n16938, new_n16939, new_n16940, new_n16941,
    new_n16942, new_n16943, new_n16944, new_n16945, new_n16946, new_n16947,
    new_n16948, new_n16949, new_n16950, new_n16951_1, new_n16952,
    new_n16953, new_n16954_1, new_n16955, new_n16956, new_n16957,
    new_n16958, new_n16959, new_n16960, new_n16961, new_n16962, new_n16963,
    new_n16964, new_n16965, new_n16966, new_n16967, new_n16968_1,
    new_n16969, new_n16970, new_n16971_1, new_n16972, new_n16973,
    new_n16974, new_n16975, new_n16976, new_n16977, new_n16978, new_n16979,
    new_n16980, new_n16981, new_n16982, new_n16983, new_n16984, new_n16985,
    new_n16986, new_n16987, new_n16988_1, new_n16989_1, new_n16990,
    new_n16991, new_n16992, new_n16993, new_n16994_1, new_n16995,
    new_n16996, new_n16997, new_n16998, new_n17001, new_n17002, new_n17003,
    new_n17004, new_n17005, new_n17006_1, new_n17007, new_n17008,
    new_n17009, new_n17010, new_n17011, new_n17012, new_n17013, new_n17014,
    new_n17015, new_n17016, new_n17017, new_n17018, new_n17019, new_n17020,
    new_n17021, new_n17022, new_n17023, new_n17024, new_n17026, new_n17027,
    new_n17028, new_n17029, new_n17030, new_n17031, new_n17032, new_n17033,
    new_n17034, new_n17035_1, new_n17036, new_n17037_1, new_n17038,
    new_n17039, new_n17040, new_n17041, new_n17042, new_n17043, new_n17044,
    new_n17045, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052,
    new_n17053, new_n17058, new_n17059, new_n17060, new_n17061, new_n17062,
    new_n17063, new_n17064, new_n17065, new_n17066, new_n17067,
    new_n17068_1, new_n17069_1, new_n17070_1, new_n17071, new_n17072,
    new_n17073, new_n17074, new_n17075_1, new_n17076, new_n17077_1,
    new_n17078, new_n17079, new_n17080, new_n17081, new_n17082, new_n17083,
    new_n17084_1, new_n17085, new_n17086, new_n17087, new_n17088,
    new_n17089, new_n17090_1, new_n17091, new_n17092, new_n17093,
    new_n17094, new_n17095_1, new_n17096, new_n17097, new_n17098,
    new_n17099, new_n17100, new_n17101, new_n17102, new_n17103,
    new_n17104_1, new_n17105, new_n17106_1, new_n17107, new_n17108,
    new_n17109, new_n17110, new_n17111, new_n17112, new_n17113, new_n17114,
    new_n17115, new_n17116, new_n17117, new_n17118, new_n17119_1,
    new_n17120, new_n17121, new_n17122, new_n17123, new_n17124, new_n17125,
    new_n17126, new_n17127, new_n17128, new_n17129, new_n17130_1,
    new_n17131, new_n17132, new_n17133, new_n17134, new_n17135, new_n17136,
    new_n17137, new_n17138_1, new_n17139, new_n17140, new_n17141,
    new_n17142, new_n17143, new_n17144, new_n17145, new_n17146, new_n17147,
    new_n17148, new_n17149, new_n17150, new_n17151, new_n17152, new_n17153,
    new_n17154, new_n17155, new_n17156, new_n17159, new_n17160, new_n17161,
    new_n17162, new_n17163_1, new_n17164, new_n17165, new_n17166,
    new_n17167, new_n17168_1, new_n17169, new_n17170, new_n17171,
    new_n17172, new_n17173, new_n17174, new_n17175, new_n17176, new_n17177,
    new_n17178, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201,
    new_n17202_1, new_n17203, new_n17204, new_n17205, new_n17206,
    new_n17207, new_n17208, new_n17209, new_n17210, new_n17211, new_n17212,
    new_n17213, new_n17214, new_n17215, new_n17216, new_n17217, new_n17218,
    new_n17219_1, new_n17220, new_n17221, new_n17222, new_n17223,
    new_n17224, new_n17225, new_n17226, new_n17227, new_n17228, new_n17229,
    new_n17230, new_n17231, new_n17232_1, new_n17233, new_n17236_1,
    new_n17237, new_n17238, new_n17239, new_n17240, new_n17241, new_n17242,
    new_n17243_1, new_n17244, new_n17245, new_n17246, new_n17247,
    new_n17248, new_n17249, new_n17250_1, new_n17251_1, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263_1,
    new_n17264, new_n17265, new_n17266, new_n17267, new_n17268, new_n17269,
    new_n17270, new_n17271, new_n17273, new_n17274, new_n17275, new_n17276,
    new_n17277, new_n17278, new_n17279, new_n17280, new_n17281, new_n17282,
    new_n17283, new_n17284, new_n17285_1, new_n17286, new_n17287,
    new_n17288, new_n17289, new_n17290, new_n17291, new_n17292, new_n17293,
    new_n17294, new_n17295, new_n17296, new_n17297, new_n17298, new_n17299,
    new_n17300, new_n17301, new_n17302_1, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17315, new_n17316, new_n17317, new_n17318, new_n17319,
    new_n17320_1, new_n17321, new_n17322, new_n17323, new_n17324,
    new_n17325, new_n17326, new_n17327, new_n17328, new_n17329, new_n17330,
    new_n17331, new_n17332, new_n17333, new_n17334, new_n17339, new_n17340,
    new_n17341, new_n17342, new_n17343, new_n17344_1, new_n17345,
    new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351_1, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359_1, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387_1, new_n17388, new_n17389,
    new_n17390, new_n17391_1, new_n17392_1, new_n17393, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17419, new_n17420, new_n17421_1, new_n17422,
    new_n17423, new_n17424, new_n17425, new_n17426, new_n17427, new_n17428,
    new_n17429, new_n17430, new_n17431, new_n17432_1, new_n17433,
    new_n17434, new_n17436_1, new_n17437, new_n17438, new_n17439,
    new_n17440_1, new_n17441, new_n17442, new_n17443, new_n17444,
    new_n17445, new_n17446, new_n17447, new_n17448, new_n17449,
    new_n17450_1, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17458_1, new_n17459,
    new_n17460, new_n17461_1, new_n17462, new_n17463, new_n17464,
    new_n17465, new_n17466_1, new_n17467, new_n17468, new_n17469,
    new_n17470, new_n17471, new_n17472, new_n17473, new_n17474, new_n17475,
    new_n17476, new_n17477, new_n17478, new_n17479, new_n17480, new_n17481,
    new_n17482, new_n17483, new_n17484, new_n17485, new_n17486, new_n17487,
    new_n17488, new_n17489, new_n17490, new_n17491, new_n17492,
    new_n17493_1, new_n17494, new_n17495, new_n17496, new_n17497,
    new_n17498, new_n17499, new_n17500_1, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17508,
    new_n17509, new_n17510, new_n17515, new_n17516, new_n17517, new_n17518,
    new_n17519, new_n17520, new_n17521, new_n17522, new_n17523,
    new_n17524_1, new_n17525, new_n17526, new_n17527, new_n17528,
    new_n17529_1, new_n17530, new_n17531, new_n17532, new_n17533,
    new_n17534, new_n17535, new_n17536, new_n17537, new_n17538, new_n17539,
    new_n17540, new_n17541, new_n17542, new_n17543, new_n17544, new_n17545,
    new_n17546, new_n17547, new_n17548, new_n17549, new_n17550, new_n17551,
    new_n17552, new_n17553, new_n17554, new_n17555, new_n17556,
    new_n17557_1, new_n17558, new_n17559, new_n17560, new_n17561,
    new_n17562, new_n17563, new_n17564, new_n17565, new_n17566, new_n17567,
    new_n17568, new_n17569, new_n17570, new_n17571, new_n17572, new_n17573,
    new_n17574, new_n17575, new_n17576, new_n17577, new_n17578, new_n17579,
    new_n17580, new_n17581, new_n17582, new_n17583_1, new_n17584,
    new_n17585, new_n17586, new_n17587, new_n17590, new_n17591,
    new_n17592_1, new_n17593, new_n17594, new_n17595, new_n17596,
    new_n17597, new_n17598, new_n17599, new_n17600, new_n17601, new_n17602,
    new_n17603, new_n17604, new_n17605, new_n17606, new_n17607, new_n17608,
    new_n17609, new_n17610, new_n17611, new_n17612, new_n17613, new_n17614,
    new_n17615, new_n17616, new_n17617, new_n17618, new_n17619, new_n17620,
    new_n17621, new_n17622, new_n17623, new_n17624, new_n17625, new_n17626,
    new_n17627, new_n17628, new_n17629, new_n17630, new_n17631, new_n17632,
    new_n17633, new_n17634, new_n17635, new_n17636, new_n17637,
    new_n17638_1, new_n17639, new_n17640, new_n17641, new_n17642,
    new_n17643, new_n17644, new_n17645, new_n17646, new_n17647, new_n17648,
    new_n17649, new_n17652, new_n17653, new_n17654, new_n17655, new_n17656,
    new_n17657, new_n17658, new_n17659, new_n17660, new_n17661, new_n17662,
    new_n17663, new_n17664_1, new_n17665, new_n17666, new_n17667,
    new_n17668, new_n17670, new_n17671, new_n17672, new_n17673, new_n17674,
    new_n17675, new_n17676, new_n17677, new_n17678, new_n17679, new_n17680,
    new_n17681, new_n17682, new_n17683, new_n17684, new_n17685, new_n17686,
    new_n17687_1, new_n17688, new_n17689, new_n17691, new_n17692,
    new_n17693, new_n17694, new_n17695, new_n17696, new_n17697, new_n17698,
    new_n17699, new_n17700, new_n17701, new_n17702, new_n17703, new_n17704,
    new_n17705, new_n17706, new_n17707, new_n17708, new_n17709, new_n17710,
    new_n17711, new_n17712, new_n17713, new_n17714, new_n17715, new_n17716,
    new_n17717, new_n17718, new_n17719, new_n17720, new_n17721_1,
    new_n17722, new_n17723, new_n17724, new_n17725, new_n17726, new_n17727,
    new_n17728, new_n17729, new_n17730, new_n17734, new_n17735_1,
    new_n17736, new_n17737, new_n17738_1, new_n17739, new_n17740,
    new_n17741, new_n17742, new_n17743, new_n17744, new_n17745,
    new_n17746_1, new_n17747, new_n17748, new_n17749_1, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17783, new_n17784_1, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17807, new_n17808, new_n17809, new_n17810,
    new_n17811, new_n17812, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820_1, new_n17821, new_n17822,
    new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828,
    new_n17829, new_n17830, new_n17835, new_n17836, new_n17837, new_n17838,
    new_n17839, new_n17840, new_n17841, new_n17842, new_n17843, new_n17846,
    new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852,
    new_n17853, new_n17854, new_n17855_1, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17860, new_n17861, new_n17862, new_n17863,
    new_n17864, new_n17865, new_n17866, new_n17867, new_n17868, new_n17869,
    new_n17870, new_n17871, new_n17872, new_n17873, new_n17874, new_n17875,
    new_n17876, new_n17877_1, new_n17878, new_n17879, new_n17880,
    new_n17881, new_n17882, new_n17883, new_n17884, new_n17885, new_n17886,
    new_n17887, new_n17888, new_n17889_1, new_n17890, new_n17891,
    new_n17892, new_n17893, new_n17894, new_n17895, new_n17896, new_n17897,
    new_n17898, new_n17899, new_n17900, new_n17901, new_n17902, new_n17903,
    new_n17904, new_n17905, new_n17906, new_n17907, new_n17908, new_n17909,
    new_n17910, new_n17915, new_n17916, new_n17917, new_n17918, new_n17919,
    new_n17920, new_n17921, new_n17922, new_n17923, new_n17924, new_n17925,
    new_n17926, new_n17927_1, new_n17928, new_n17929, new_n17930,
    new_n17931_1, new_n17932, new_n17933, new_n17934, new_n17935,
    new_n17939, new_n17940, new_n17941, new_n17942, new_n17943, new_n17944,
    new_n17945, new_n17946, new_n17947, new_n17948_1, new_n17949,
    new_n17950, new_n17951, new_n17952, new_n17953, new_n17954_1,
    new_n17955, new_n17956_1, new_n17957, new_n17958, new_n17959_1,
    new_n17960, new_n17961, new_n17962, new_n17963_1, new_n17964,
    new_n17965, new_n17966, new_n17967, new_n17968_1, new_n17969,
    new_n17970, new_n17971, new_n17972, new_n17973, new_n17974, new_n17975,
    new_n17976_1, new_n17977, new_n17978, new_n17979, new_n17980,
    new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986,
    new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992,
    new_n17993, new_n17994, new_n17995, new_n17996, new_n17997,
    new_n17998_1, new_n17999, new_n18000, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020,
    new_n18021, new_n18022, new_n18023, new_n18024, new_n18025_1,
    new_n18026, new_n18027, new_n18028, new_n18029, new_n18030, new_n18031,
    new_n18032, new_n18040, new_n18041, new_n18042, new_n18043_1,
    new_n18044, new_n18045_1, new_n18046, new_n18047, new_n18048,
    new_n18049, new_n18050, new_n18051, new_n18052, new_n18053, new_n18054,
    new_n18055, new_n18056, new_n18057, new_n18058, new_n18059_1,
    new_n18060, new_n18061_1, new_n18062, new_n18063, new_n18064,
    new_n18065, new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071_1, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18081, new_n18082, new_n18083, new_n18084,
    new_n18085, new_n18086, new_n18087, new_n18088, new_n18089, new_n18090,
    new_n18091, new_n18092, new_n18093, new_n18094, new_n18095, new_n18096,
    new_n18097, new_n18098, new_n18099, new_n18100, new_n18101, new_n18102,
    new_n18103, new_n18104, new_n18105_1, new_n18106, new_n18107,
    new_n18108, new_n18109, new_n18110, new_n18111, new_n18112, new_n18113,
    new_n18114, new_n18115, new_n18116, new_n18117, new_n18118, new_n18119,
    new_n18120, new_n18121, new_n18122, new_n18123, new_n18124, new_n18125,
    new_n18126, new_n18127, new_n18128, new_n18129, new_n18130, new_n18131,
    new_n18132, new_n18133, new_n18134, new_n18135, new_n18136, new_n18137,
    new_n18138, new_n18139, new_n18140, new_n18141, new_n18142,
    new_n18143_1, new_n18144, new_n18145_1, new_n18146, new_n18147,
    new_n18148, new_n18149, new_n18150, new_n18151_1, new_n18152_1,
    new_n18153, new_n18154, new_n18155, new_n18156, new_n18157_1,
    new_n18158, new_n18159, new_n18160, new_n18161, new_n18162, new_n18163,
    new_n18164, new_n18165, new_n18166, new_n18167, new_n18168, new_n18169,
    new_n18170, new_n18171_1, new_n18173, new_n18174, new_n18175,
    new_n18176, new_n18177, new_n18178, new_n18179, new_n18180, new_n18181,
    new_n18185, new_n18186, new_n18187, new_n18188, new_n18189, new_n18190,
    new_n18191, new_n18192, new_n18193_1, new_n18194, new_n18195,
    new_n18196, new_n18197, new_n18198, new_n18199, new_n18200, new_n18201,
    new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207,
    new_n18208, new_n18209, new_n18211, new_n18212, new_n18213, new_n18214,
    new_n18215, new_n18216, new_n18217, new_n18218, new_n18219, new_n18220,
    new_n18221, new_n18222, new_n18223, new_n18224, new_n18225, new_n18226,
    new_n18227_1, new_n18228, new_n18229, new_n18230, new_n18231,
    new_n18232_1, new_n18233, new_n18234, new_n18235, new_n18236,
    new_n18237, new_n18238_1, new_n18239, new_n18240, new_n18241_1,
    new_n18242, new_n18243, new_n18244, new_n18245, new_n18246, new_n18247,
    new_n18248, new_n18249, new_n18250, new_n18251, new_n18252, new_n18253,
    new_n18254_1, new_n18255, new_n18256, new_n18257, new_n18258,
    new_n18259, new_n18260, new_n18261, new_n18262, new_n18263, new_n18264,
    new_n18265, new_n18266, new_n18267, new_n18268, new_n18269, new_n18270,
    new_n18271, new_n18272, new_n18273, new_n18274_1, new_n18275,
    new_n18277, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284,
    new_n18285, new_n18286, new_n18287, new_n18288_1, new_n18289,
    new_n18290_1, new_n18291, new_n18292, new_n18293, new_n18294,
    new_n18295_1, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301_1, new_n18302, new_n18303, new_n18304_1,
    new_n18305, new_n18306, new_n18307, new_n18308, new_n18309,
    new_n18310_1, new_n18311_1, new_n18312, new_n18313, new_n18314,
    new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320,
    new_n18321, new_n18322, new_n18323_1, new_n18324, new_n18325,
    new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332_1, new_n18333, new_n18334, new_n18335, new_n18336,
    new_n18337, new_n18338, new_n18339, new_n18340, new_n18341, new_n18342,
    new_n18343_1, new_n18344, new_n18345_1, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350_1, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362_1, new_n18363,
    new_n18364, new_n18365, new_n18366, new_n18367, new_n18368, new_n18369,
    new_n18370, new_n18371, new_n18372, new_n18373, new_n18374, new_n18375,
    new_n18376, new_n18377_1, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18387, new_n18388,
    new_n18389, new_n18390, new_n18391, new_n18392, new_n18393, new_n18394,
    new_n18395, new_n18396, new_n18397, new_n18398, new_n18399, new_n18400,
    new_n18401, new_n18402, new_n18403, new_n18404, new_n18405_1,
    new_n18406, new_n18407, new_n18408, new_n18409_1, new_n18410,
    new_n18411, new_n18412, new_n18413, new_n18414_1, new_n18415,
    new_n18416, new_n18417, new_n18418_1, new_n18419, new_n18420,
    new_n18421, new_n18422, new_n18423, new_n18424, new_n18425, new_n18426,
    new_n18427, new_n18428, new_n18429, new_n18430, new_n18431, new_n18432,
    new_n18433, new_n18434, new_n18435, new_n18436, new_n18437_1,
    new_n18438, new_n18439_1, new_n18440, new_n18441, new_n18442,
    new_n18443, new_n18444_1, new_n18445_1, new_n18446, new_n18447,
    new_n18448, new_n18449, new_n18450, new_n18451, new_n18452_1,
    new_n18453, new_n18460, new_n18461, new_n18462, new_n18466,
    new_n18467_1, new_n18468, new_n18469, new_n18470, new_n18471,
    new_n18472, new_n18473, new_n18474, new_n18475, new_n18476, new_n18477,
    new_n18478, new_n18479, new_n18480, new_n18481, new_n18482_1,
    new_n18483_1, new_n18484, new_n18485, new_n18486, new_n18487,
    new_n18488, new_n18489, new_n18490, new_n18491, new_n18492, new_n18493,
    new_n18494, new_n18495, new_n18496_1, new_n18497, new_n18498,
    new_n18499, new_n18500, new_n18501, new_n18502, new_n18503, new_n18504,
    new_n18505, new_n18506, new_n18507, new_n18508, new_n18509_1,
    new_n18510, new_n18511, new_n18512, new_n18513_1, new_n18514,
    new_n18515_1, new_n18516, new_n18517, new_n18518, new_n18519,
    new_n18520, new_n18521, new_n18522, new_n18523, new_n18524, new_n18525,
    new_n18526, new_n18527, new_n18528, new_n18529, new_n18530, new_n18531,
    new_n18532, new_n18533, new_n18534, new_n18535, new_n18536,
    new_n18537_1, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18555, new_n18556, new_n18557, new_n18558_1,
    new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564,
    new_n18565, new_n18566, new_n18567, new_n18568, new_n18569, new_n18570,
    new_n18571, new_n18572_1, new_n18573, new_n18574_1, new_n18575,
    new_n18576_1, new_n18577, new_n18578_1, new_n18579, new_n18580,
    new_n18581, new_n18582_1, new_n18583_1, new_n18584_1, new_n18585,
    new_n18586, new_n18587, new_n18588, new_n18589, new_n18590, new_n18591,
    new_n18592, new_n18593, new_n18594, new_n18595, new_n18596, new_n18597,
    new_n18600, new_n18601, new_n18602, new_n18603, new_n18604, new_n18605,
    new_n18606, new_n18607, new_n18608, new_n18609, new_n18610_1,
    new_n18611, new_n18612, new_n18613, new_n18614, new_n18615, new_n18616,
    new_n18617, new_n18618, new_n18619, new_n18620, new_n18621, new_n18622,
    new_n18623, new_n18624, new_n18625, new_n18626, new_n18627, new_n18628,
    new_n18629, new_n18630, new_n18631, new_n18632, new_n18633, new_n18634,
    new_n18635_1, new_n18636, new_n18637, new_n18638, new_n18639,
    new_n18640, new_n18641, new_n18642, new_n18643, new_n18644, new_n18645,
    new_n18646, new_n18647, new_n18648, new_n18649_1, new_n18650,
    new_n18651, new_n18652, new_n18653_1, new_n18654, new_n18655,
    new_n18656, new_n18657, new_n18658, new_n18659, new_n18660, new_n18661,
    new_n18662, new_n18663, new_n18664, new_n18665, new_n18666, new_n18667,
    new_n18668, new_n18669, new_n18670, new_n18671, new_n18672, new_n18673,
    new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679_1, new_n18680, new_n18681, new_n18682, new_n18683,
    new_n18684, new_n18685, new_n18686, new_n18687, new_n18688, new_n18689,
    new_n18694, new_n18695, new_n18696, new_n18697, new_n18698, new_n18699,
    new_n18700, new_n18701, new_n18702, new_n18703, new_n18704, new_n18705,
    new_n18706, new_n18707, new_n18708_1, new_n18709, new_n18710,
    new_n18711, new_n18712, new_n18713, new_n18714, new_n18715, new_n18716,
    new_n18717, new_n18718, new_n18719, new_n18720, new_n18721_1,
    new_n18722, new_n18723, new_n18724, new_n18725_1, new_n18726,
    new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732,
    new_n18733, new_n18734, new_n18735, new_n18736, new_n18737_1,
    new_n18738, new_n18739, new_n18740, new_n18741, new_n18742, new_n18743,
    new_n18744, new_n18745_1, new_n18746, new_n18747, new_n18748,
    new_n18749, new_n18750, new_n18751_1, new_n18752, new_n18753,
    new_n18754, new_n18755, new_n18756, new_n18757, new_n18758, new_n18759,
    new_n18760, new_n18761, new_n18762, new_n18763, new_n18764, new_n18765,
    new_n18766, new_n18767, new_n18768, new_n18769, new_n18770, new_n18771,
    new_n18772, new_n18773, new_n18774, new_n18775, new_n18776, new_n18777,
    new_n18778, new_n18779, new_n18780_1, new_n18781, new_n18782_1,
    new_n18783, new_n18784, new_n18785, new_n18786, new_n18788, new_n18789,
    new_n18790, new_n18791, new_n18792, new_n18793, new_n18794, new_n18795,
    new_n18796, new_n18798, new_n18799, new_n18800, new_n18801,
    new_n18802_1, new_n18803, new_n18804, new_n18805, new_n18806,
    new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812,
    new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818,
    new_n18819, new_n18820, new_n18821, new_n18822, new_n18823, new_n18824,
    new_n18831_1, new_n18832, new_n18833, new_n18834, new_n18835,
    new_n18836, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841,
    new_n18842, new_n18843_1, new_n18844, new_n18845, new_n18846,
    new_n18858_1, new_n18859_1, new_n18860, new_n18861, new_n18862,
    new_n18863, new_n18864_1, new_n18865_1, new_n18866, new_n18867,
    new_n18868, new_n18869, new_n18870, new_n18871, new_n18872, new_n18873,
    new_n18874, new_n18875, new_n18876, new_n18877, new_n18878, new_n18879,
    new_n18880_1, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886_1, new_n18887_1, new_n18888, new_n18889,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18899, new_n18900, new_n18901_1,
    new_n18902, new_n18903, new_n18904, new_n18905, new_n18906,
    new_n18907_1, new_n18908, new_n18909, new_n18910, new_n18911,
    new_n18912, new_n18913, new_n18914, new_n18915, new_n18916, new_n18917,
    new_n18918, new_n18919_1, new_n18920, new_n18921, new_n18922,
    new_n18923, new_n18924, new_n18926_1, new_n18927, new_n18928,
    new_n18929, new_n18930, new_n18931, new_n18932, new_n18933, new_n18934,
    new_n18935, new_n18936, new_n18937, new_n18938, new_n18939,
    new_n18940_1, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945_1, new_n18946, new_n18947, new_n18948, new_n18949,
    new_n18950, new_n18951, new_n18952, new_n18953, new_n18954, new_n18955,
    new_n18956, new_n18957, new_n18958, new_n18959, new_n18960, new_n18961,
    new_n18962_1, new_n18963, new_n18964, new_n18965, new_n18966,
    new_n18967, new_n18968, new_n18969, new_n18970_1, new_n18971,
    new_n18972, new_n18973, new_n18974, new_n18975, new_n18976,
    new_n18977_1, new_n18978, new_n18979, new_n18980, new_n18981,
    new_n18982_1, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999_1, new_n19000, new_n19001, new_n19002, new_n19003,
    new_n19004, new_n19005_1, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033_1, new_n19034, new_n19035, new_n19036, new_n19037,
    new_n19038, new_n19039, new_n19040, new_n19041, new_n19042_1,
    new_n19043, new_n19044_1, new_n19045, new_n19046, new_n19047,
    new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053,
    new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065,
    new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071,
    new_n19072, new_n19073, new_n19074, new_n19075, new_n19076, new_n19077,
    new_n19078, new_n19079, new_n19080, new_n19081_1, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19091, new_n19092,
    new_n19093, new_n19094, new_n19095, new_n19096, new_n19097, new_n19098,
    new_n19099, new_n19100, new_n19101, new_n19102, new_n19103, new_n19104,
    new_n19105, new_n19106, new_n19107_1, new_n19108, new_n19109,
    new_n19112, new_n19113, new_n19114, new_n19115, new_n19116_1,
    new_n19117, new_n19118, new_n19119, new_n19120, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125_1, new_n19126, new_n19127,
    new_n19128, new_n19129, new_n19130, new_n19131, new_n19132, new_n19133,
    new_n19136, new_n19137, new_n19138, new_n19139, new_n19140,
    new_n19141_1, new_n19142, new_n19147, new_n19148, new_n19149,
    new_n19153, new_n19154, new_n19155, new_n19156, new_n19157, new_n19158,
    new_n19159, new_n19160, new_n19161, new_n19162, new_n19163_1,
    new_n19164_1, new_n19165, new_n19166, new_n19167, new_n19168,
    new_n19169, new_n19170, new_n19171, new_n19175, new_n19176_1,
    new_n19177, new_n19178, new_n19179, new_n19180, new_n19181, new_n19182,
    new_n19183, new_n19185, new_n19186, new_n19187, new_n19188, new_n19189,
    new_n19190, new_n19191, new_n19192, new_n19193, new_n19194, new_n19195,
    new_n19196_1, new_n19197, new_n19198, new_n19199, new_n19200,
    new_n19201, new_n19202_1, new_n19203, new_n19205, new_n19206,
    new_n19207, new_n19208, new_n19209, new_n19210, new_n19211, new_n19212,
    new_n19213, new_n19214, new_n19215, new_n19216, new_n19217, new_n19218,
    new_n19219, new_n19220_1, new_n19221_1, new_n19222, new_n19223_1,
    new_n19224_1, new_n19225, new_n19226, new_n19227, new_n19228_1,
    new_n19229, new_n19230, new_n19231, new_n19232, new_n19233_1,
    new_n19234_1, new_n19235, new_n19236, new_n19237, new_n19238,
    new_n19239, new_n19241, new_n19242, new_n19243, new_n19244_1,
    new_n19245, new_n19246, new_n19247, new_n19248, new_n19249, new_n19250,
    new_n19251, new_n19252, new_n19253, new_n19254, new_n19255, new_n19256,
    new_n19257, new_n19258, new_n19259, new_n19260, new_n19261, new_n19262,
    new_n19263, new_n19264, new_n19265, new_n19266, new_n19267, new_n19268,
    new_n19269, new_n19270_1, new_n19271, new_n19272, new_n19273,
    new_n19274, new_n19275, new_n19276, new_n19277, new_n19278, new_n19279,
    new_n19280, new_n19281, new_n19282_1, new_n19283, new_n19284,
    new_n19285, new_n19286, new_n19287, new_n19288, new_n19289, new_n19290,
    new_n19291, new_n19292, new_n19293, new_n19294, new_n19295, new_n19296,
    new_n19297, new_n19298, new_n19299, new_n19300, new_n19301, new_n19302,
    new_n19303, new_n19304, new_n19305, new_n19306, new_n19307, new_n19308,
    new_n19309, new_n19310, new_n19311, new_n19312, new_n19313,
    new_n19314_1, new_n19315_1, new_n19316, new_n19317, new_n19318,
    new_n19323_1, new_n19324, new_n19325, new_n19326, new_n19327_1,
    new_n19328, new_n19329, new_n19330, new_n19331, new_n19332,
    new_n19333_1, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343,
    new_n19344, new_n19345, new_n19346, new_n19347, new_n19348_1,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353,
    new_n19354_1, new_n19355, new_n19356, new_n19357_1, new_n19358,
    new_n19359, new_n19360, new_n19361_1, new_n19362, new_n19363,
    new_n19364, new_n19365, new_n19366, new_n19367_1, new_n19368,
    new_n19369, new_n19370, new_n19371, new_n19372, new_n19373, new_n19374,
    new_n19375, new_n19376, new_n19377, new_n19378, new_n19379, new_n19380,
    new_n19381, new_n19382, new_n19383, new_n19384, new_n19385_1,
    new_n19386, new_n19387, new_n19388, new_n19389_1, new_n19390,
    new_n19391, new_n19392, new_n19393, new_n19394, new_n19395, new_n19396,
    new_n19397, new_n19398, new_n19399, new_n19400, new_n19401_1,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414_1, new_n19415, new_n19416, new_n19417, new_n19418,
    new_n19419, new_n19420, new_n19421, new_n19422, new_n19423,
    new_n19424_1, new_n19425, new_n19426, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19442, new_n19443, new_n19445, new_n19446, new_n19451,
    new_n19454_1, new_n19455, new_n19456, new_n19457, new_n19458_1,
    new_n19459, new_n19460, new_n19461, new_n19462, new_n19463, new_n19464,
    new_n19465, new_n19466, new_n19467_1, new_n19468, new_n19469,
    new_n19470, new_n19471, new_n19472_1, new_n19473, new_n19474,
    new_n19475, new_n19476, new_n19477_1, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19487, new_n19488, new_n19489, new_n19490, new_n19491, new_n19492,
    new_n19493, new_n19494_1, new_n19495, new_n19496_1, new_n19497,
    new_n19498, new_n19499, new_n19500, new_n19501, new_n19502, new_n19503,
    new_n19504, new_n19505, new_n19506, new_n19507, new_n19508, new_n19509,
    new_n19510, new_n19511, new_n19512, new_n19513, new_n19514_1,
    new_n19515_1, new_n19524, new_n19525, new_n19526, new_n19527,
    new_n19528, new_n19529, new_n19530, new_n19531_1, new_n19532,
    new_n19533, new_n19534, new_n19535, new_n19536, new_n19540, new_n19541,
    new_n19542, new_n19543, new_n19544, new_n19545, new_n19546, new_n19547,
    new_n19548, new_n19549, new_n19550, new_n19551, new_n19552, new_n19553,
    new_n19554, new_n19555, new_n19556, new_n19557, new_n19558, new_n19559,
    new_n19560, new_n19561, new_n19562, new_n19563, new_n19564, new_n19565,
    new_n19566, new_n19567, new_n19568, new_n19569, new_n19570_1,
    new_n19571, new_n19574, new_n19575_1, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19639,
    new_n19640, new_n19641_1, new_n19642, new_n19643, new_n19644,
    new_n19645, new_n19646, new_n19647, new_n19648_1, new_n19649,
    new_n19650, new_n19651, new_n19652_1, new_n19653, new_n19654,
    new_n19655, new_n19656, new_n19657, new_n19658, new_n19659, new_n19660,
    new_n19661, new_n19662, new_n19663, new_n19664_1, new_n19665,
    new_n19666, new_n19667, new_n19668, new_n19669, new_n19670, new_n19671,
    new_n19673, new_n19674, new_n19676, new_n19677, new_n19678, new_n19679,
    new_n19680_1, new_n19681, new_n19682, new_n19683, new_n19684,
    new_n19685, new_n19686, new_n19687, new_n19688, new_n19689, new_n19690,
    new_n19691, new_n19692, new_n19693, new_n19694, new_n19695, new_n19696,
    new_n19697, new_n19698, new_n19699, new_n19700, new_n19701_1,
    new_n19702, new_n19703, new_n19704, new_n19705, new_n19706, new_n19707,
    new_n19708, new_n19709, new_n19710, new_n19711, new_n19714, new_n19715,
    new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723,
    new_n19724, new_n19725, new_n19726, new_n19727, new_n19728, new_n19729,
    new_n19730, new_n19731, new_n19732, new_n19733, new_n19734, new_n19735,
    new_n19736_1, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749_1, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756_1,
    new_n19759, new_n19760, new_n19761, new_n19762, new_n19763, new_n19764,
    new_n19765, new_n19766, new_n19767_1, new_n19768, new_n19769,
    new_n19770_1, new_n19771, new_n19772, new_n19773, new_n19774,
    new_n19775, new_n19776, new_n19777, new_n19778, new_n19779,
    new_n19780_1, new_n19781, new_n19789_1, new_n19790, new_n19791,
    new_n19792_1, new_n19793, new_n19794, new_n19795, new_n19796,
    new_n19797, new_n19798_1, new_n19799, new_n19800, new_n19801,
    new_n19802, new_n19803_1, new_n19804, new_n19805, new_n19806,
    new_n19807, new_n19808, new_n19809, new_n19810, new_n19811, new_n19812,
    new_n19813, new_n19814, new_n19815, new_n19816, new_n19817, new_n19818,
    new_n19819, new_n19820, new_n19821, new_n19822, new_n19823, new_n19824,
    new_n19825, new_n19826, new_n19827, new_n19828, new_n19829, new_n19830,
    new_n19831, new_n19832, new_n19833, new_n19834, new_n19835, new_n19836,
    new_n19837, new_n19838, new_n19839, new_n19840, new_n19841, new_n19842,
    new_n19843, new_n19844, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19881, new_n19883, new_n19884, new_n19885,
    new_n19886, new_n19887, new_n19888, new_n19889, new_n19890, new_n19891,
    new_n19892, new_n19893, new_n19894, new_n19895, new_n19896, new_n19897,
    new_n19898, new_n19899, new_n19900, new_n19901, new_n19902, new_n19904,
    new_n19905_1, new_n19906, new_n19907, new_n19908, new_n19909_1,
    new_n19910, new_n19911_1, new_n19912, new_n19913, new_n19914,
    new_n19915, new_n19916_1, new_n19917, new_n19918, new_n19919,
    new_n19920, new_n19922_1, new_n19923_1, new_n19924, new_n19925,
    new_n19926, new_n19927, new_n19928, new_n19929, new_n19930_1,
    new_n19931, new_n19932, new_n19933, new_n19934, new_n19935, new_n19936,
    new_n19941_1, new_n19942, new_n19943, new_n19944, new_n19945,
    new_n19946, new_n19947, new_n19948, new_n19949, new_n19950, new_n19951,
    new_n19952, new_n19953, new_n19954, new_n19955, new_n19956, new_n19957,
    new_n19958, new_n19959, new_n19960, new_n19969, new_n19970, new_n19971,
    new_n19972, new_n19973, new_n19974, new_n19975, new_n19976, new_n19982,
    new_n19983, new_n19984, new_n19985, new_n19986, new_n19987,
    new_n19988_1, new_n19989, new_n19990, new_n19995, new_n20001,
    new_n20002, new_n20003, new_n20004_1, new_n20005, new_n20006,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013_1, new_n20014, new_n20015, new_n20016, new_n20017_1,
    new_n20018, new_n20019, new_n20024, new_n20025, new_n20026, new_n20027,
    new_n20028, new_n20029, new_n20036_1, new_n20037, new_n20038,
    new_n20039, new_n20040_1, new_n20041, new_n20042, new_n20043,
    new_n20044, new_n20045, new_n20046, new_n20047, new_n20048, new_n20049,
    new_n20050, new_n20051, new_n20052, new_n20053, new_n20054, new_n20055,
    new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061_1, new_n20062, new_n20063, new_n20064, new_n20065,
    new_n20066, new_n20067, new_n20068, new_n20069_1, new_n20070,
    new_n20071, new_n20072, new_n20073, new_n20074, new_n20075, new_n20076,
    new_n20077_1, new_n20078, new_n20079, new_n20080, new_n20081,
    new_n20082, new_n20085, new_n20086_1, new_n20087, new_n20088,
    new_n20089, new_n20090, new_n20091, new_n20092, new_n20093, new_n20095,
    new_n20096_1, new_n20097, new_n20098, new_n20099, new_n20100,
    new_n20101, new_n20102, new_n20103_1, new_n20104, new_n20105,
    new_n20106, new_n20107, new_n20108, new_n20109, new_n20110, new_n20111,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125,
    new_n20126_1, new_n20127, new_n20128, new_n20129, new_n20130,
    new_n20131, new_n20132, new_n20133, new_n20134, new_n20135, new_n20136,
    new_n20137, new_n20138_1, new_n20139, new_n20140, new_n20141,
    new_n20142, new_n20143, new_n20144, new_n20145, new_n20146, new_n20147,
    new_n20148, new_n20149_1, new_n20150, new_n20151_1, new_n20157,
    new_n20158, new_n20159, new_n20160, new_n20170, new_n20171, new_n20172,
    new_n20173, new_n20174, new_n20175, new_n20176, new_n20177, new_n20178,
    new_n20179_1, new_n20180, new_n20181, new_n20182, new_n20183,
    new_n20184, new_n20185, new_n20186, new_n20187_1, new_n20188,
    new_n20189, new_n20190, new_n20191, new_n20192, new_n20193, new_n20194,
    new_n20195, new_n20196, new_n20197, new_n20198, new_n20199, new_n20200,
    new_n20201, new_n20202, new_n20203, new_n20204, new_n20205, new_n20206,
    new_n20207, new_n20208, new_n20209, new_n20210, new_n20211, new_n20212,
    new_n20213_1, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229,
    new_n20230, new_n20231, new_n20232, new_n20233, new_n20234,
    new_n20235_1, new_n20236, new_n20237, new_n20238, new_n20239,
    new_n20240, new_n20241, new_n20242, new_n20243, new_n20244, new_n20245,
    new_n20246, new_n20247, new_n20249, new_n20250_1, new_n20251,
    new_n20252, new_n20253, new_n20254, new_n20255, new_n20256, new_n20257,
    new_n20258, new_n20259_1, new_n20260, new_n20261, new_n20262,
    new_n20263, new_n20264, new_n20265, new_n20266, new_n20267, new_n20268,
    new_n20269, new_n20270, new_n20271, new_n20272, new_n20273, new_n20274,
    new_n20275, new_n20276, new_n20277, new_n20278, new_n20279_1,
    new_n20280, new_n20281, new_n20282, new_n20283, new_n20284, new_n20285,
    new_n20286, new_n20287_1, new_n20288, new_n20289, new_n20290,
    new_n20291, new_n20292, new_n20293, new_n20294, new_n20295, new_n20296,
    new_n20297, new_n20298, new_n20299, new_n20300, new_n20301_1,
    new_n20302, new_n20303, new_n20304, new_n20305, new_n20306, new_n20307,
    new_n20308, new_n20309, new_n20310, new_n20311, new_n20312, new_n20315,
    new_n20316, new_n20317, new_n20318, new_n20319, new_n20320, new_n20321,
    new_n20322, new_n20323, new_n20324, new_n20325, new_n20326, new_n20327,
    new_n20333_1, new_n20334, new_n20335, new_n20336, new_n20337,
    new_n20338, new_n20339, new_n20340, new_n20341, new_n20342, new_n20343,
    new_n20344, new_n20345, new_n20346, new_n20347, new_n20348,
    new_n20349_1, new_n20350, new_n20351, new_n20352, new_n20353,
    new_n20354, new_n20355_1, new_n20356, new_n20357, new_n20358,
    new_n20359_1, new_n20360, new_n20361, new_n20362, new_n20363,
    new_n20364, new_n20365, new_n20366_1, new_n20367, new_n20368,
    new_n20369, new_n20370, new_n20371, new_n20372, new_n20373, new_n20374,
    new_n20375, new_n20376, new_n20377, new_n20378, new_n20379, new_n20380,
    new_n20381, new_n20382, new_n20383, new_n20384, new_n20385_1,
    new_n20386, new_n20387, new_n20388_1, new_n20389, new_n20390,
    new_n20391, new_n20392, new_n20393, new_n20394, new_n20395, new_n20396,
    new_n20397, new_n20398, new_n20399, new_n20400, new_n20401,
    new_n20402_1, new_n20403_1, new_n20405, new_n20406, new_n20407,
    new_n20408, new_n20409_1, new_n20410, new_n20411_1, new_n20412,
    new_n20413, new_n20414, new_n20417, new_n20418, new_n20419, new_n20420,
    new_n20421, new_n20422, new_n20423, new_n20424_1, new_n20425,
    new_n20426, new_n20432, new_n20433, new_n20434, new_n20435,
    new_n20436_1, new_n20437, new_n20438, new_n20439, new_n20440,
    new_n20441_1, new_n20442, new_n20443, new_n20444, new_n20445_1,
    new_n20446, new_n20447, new_n20448, new_n20449, new_n20450_1,
    new_n20451, new_n20452, new_n20453, new_n20454, new_n20455_1,
    new_n20456, new_n20457, new_n20458, new_n20459, new_n20460, new_n20461,
    new_n20462, new_n20463, new_n20464, new_n20465, new_n20466, new_n20467,
    new_n20468, new_n20469, new_n20470_1, new_n20471, new_n20472,
    new_n20473, new_n20474, new_n20475, new_n20476, new_n20477,
    new_n20478_1, new_n20479, new_n20480, new_n20481, new_n20482,
    new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489_1, new_n20490_1, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495_1, new_n20496, new_n20497, new_n20498,
    new_n20499, new_n20507, new_n20508, new_n20509, new_n20510, new_n20511,
    new_n20516, new_n20519, new_n20521, new_n20522, new_n20523, new_n20524,
    new_n20525, new_n20526, new_n20527, new_n20528, new_n20529, new_n20530,
    new_n20531, new_n20532, new_n20533_1, new_n20534, new_n20535,
    new_n20536, new_n20537, new_n20538, new_n20539, new_n20540, new_n20541,
    new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547,
    new_n20548, new_n20549, new_n20550, new_n20551, new_n20552, new_n20553,
    new_n20554, new_n20555, new_n20556, new_n20557, new_n20558, new_n20559,
    new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20571, new_n20572, new_n20573,
    new_n20574, new_n20582_1, new_n20583, new_n20584, new_n20585,
    new_n20586, new_n20587, new_n20588, new_n20589, new_n20590_1,
    new_n20594, new_n20602_1, new_n20603, new_n20604_1, new_n20605,
    new_n20606, new_n20607, new_n20608, new_n20609_1, new_n20610,
    new_n20611, new_n20612, new_n20613, new_n20614, new_n20615, new_n20617,
    new_n20618, new_n20619, new_n20620, new_n20621, new_n20622,
    new_n20623_1, new_n20624, new_n20625, new_n20626, new_n20627,
    new_n20628, new_n20629_1, new_n20630, new_n20631, new_n20632,
    new_n20633, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643,
    new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20649,
    new_n20650, new_n20651, new_n20652, new_n20653, new_n20654, new_n20655,
    new_n20656, new_n20657, new_n20658_1, new_n20659, new_n20660,
    new_n20661_1, new_n20662, new_n20663, new_n20664, new_n20665,
    new_n20666, new_n20667, new_n20668, new_n20669, new_n20672,
    new_n20673_1, new_n20674, new_n20675, new_n20676, new_n20677,
    new_n20678_1, new_n20679, new_n20680_1, new_n20681, new_n20682,
    new_n20683, new_n20684, new_n20685_1, new_n20686, new_n20687,
    new_n20688, new_n20689, new_n20690, new_n20691_1, new_n20692,
    new_n20693, new_n20695, new_n20696_1, new_n20697, new_n20698,
    new_n20699, new_n20700_1, new_n20701, new_n20702, new_n20703,
    new_n20704_1, new_n20705_1, new_n20706, new_n20710, new_n20712,
    new_n20713_1, new_n20718, new_n20719, new_n20720, new_n20721,
    new_n20722_1, new_n20723_1, new_n20724, new_n20725, new_n20726,
    new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732,
    new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738,
    new_n20739, new_n20740, new_n20741, new_n20742, new_n20743, new_n20744,
    new_n20745, new_n20746, new_n20747, new_n20748_1, new_n20749,
    new_n20750, new_n20751, new_n20752, new_n20753, new_n20754, new_n20755,
    new_n20756, new_n20757, new_n20758, new_n20759, new_n20760,
    new_n20761_1, new_n20762, new_n20763, new_n20765, new_n20766,
    new_n20767, new_n20768, new_n20769, new_n20770, new_n20771, new_n20772,
    new_n20773, new_n20774_1, new_n20775, new_n20776, new_n20777,
    new_n20778, new_n20779, new_n20780, new_n20781, new_n20782, new_n20783,
    new_n20784, new_n20785, new_n20786, new_n20787, new_n20788_1,
    new_n20789, new_n20790, new_n20791, new_n20792, new_n20793,
    new_n20794_1, new_n20795_1, new_n20796, new_n20797, new_n20798,
    new_n20799, new_n20800, new_n20801, new_n20802, new_n20803_1,
    new_n20804, new_n20805, new_n20806, new_n20807, new_n20808, new_n20809,
    new_n20810, new_n20811, new_n20812, new_n20818, new_n20827, new_n20828,
    new_n20829, new_n20830, new_n20836, new_n20843, new_n20844, new_n20845,
    new_n20846, new_n20847, new_n20848, new_n20849, new_n20850, new_n20851,
    new_n20852, new_n20853, new_n20854, new_n20855, new_n20856, new_n20857,
    new_n20858, new_n20859, new_n20860, new_n20861, new_n20862, new_n20863,
    new_n20864, new_n20865, new_n20866, new_n20867, new_n20868,
    new_n20869_1, new_n20870, new_n20871, new_n20872, new_n20873,
    new_n20874, new_n20875, new_n20876, new_n20877, new_n20880, new_n20881,
    new_n20882, new_n20883, new_n20884, new_n20885, new_n20886, new_n20887,
    new_n20888, new_n20889, new_n20890, new_n20891, new_n20892, new_n20899,
    new_n20900, new_n20901, new_n20902, new_n20903, new_n20904, new_n20905,
    new_n20906, new_n20907, new_n20908, new_n20909, new_n20910, new_n20911,
    new_n20912, new_n20913, new_n20914, new_n20915_1, new_n20916,
    new_n20917, new_n20918, new_n20919, new_n20920, new_n20921, new_n20922,
    new_n20923_1, new_n20924, new_n20925, new_n20926, new_n20927,
    new_n20928, new_n20929_1, new_n20930, new_n20931, new_n20932,
    new_n20933, new_n20934, new_n20935_1, new_n20936_1, new_n20937,
    new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943,
    new_n20944, new_n20945, new_n20946_1, new_n20947, new_n20948,
    new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20954,
    new_n20955, new_n20956, new_n20957, new_n20958, new_n20959, new_n20960,
    new_n20961, new_n20962, new_n20963, new_n20964, new_n20965, new_n20966,
    new_n20967, new_n20968, new_n20969, new_n20970, new_n20971, new_n20972,
    new_n20973, new_n20974, new_n20975, new_n20976, new_n20977, new_n20978,
    new_n20979, new_n20980, new_n20981, new_n20982, new_n20983, new_n20984,
    new_n20985, new_n20986_1, new_n20987, new_n20988, new_n20989,
    new_n20990, new_n20991, new_n20992, new_n20993, new_n20994, new_n20995,
    new_n20996, new_n20997, new_n20998, new_n20999, new_n21000, new_n21001,
    new_n21002, new_n21003, new_n21004, new_n21005, new_n21006, new_n21007,
    new_n21008_1, new_n21009, new_n21010, new_n21011, new_n21012,
    new_n21013, new_n21014, new_n21015, new_n21016, new_n21017_1,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023,
    new_n21027, new_n21030, new_n21031, new_n21032, new_n21033,
    new_n21034_1, new_n21035, new_n21036, new_n21037, new_n21038,
    new_n21039, new_n21040, new_n21041, new_n21042, new_n21043, new_n21044,
    new_n21045, new_n21046_1, new_n21047, new_n21048, new_n21049,
    new_n21050, new_n21055, new_n21056, new_n21057, new_n21058, new_n21059,
    new_n21060, new_n21061, new_n21062_1, new_n21063, new_n21064,
    new_n21065, new_n21066, new_n21067, new_n21068, new_n21069, new_n21070,
    new_n21071, new_n21072, new_n21073, new_n21074, new_n21075, new_n21076,
    new_n21077, new_n21078_1, new_n21080, new_n21081, new_n21082,
    new_n21083, new_n21084, new_n21085, new_n21089, new_n21090, new_n21091,
    new_n21092, new_n21102, new_n21103, new_n21104, new_n21105, new_n21106,
    new_n21107, new_n21108, new_n21109, new_n21110, new_n21111, new_n21112,
    new_n21113, new_n21114, new_n21115, new_n21116, new_n21117, new_n21118,
    new_n21119, new_n21120, new_n21121, new_n21122, new_n21143, new_n21144,
    new_n21145, new_n21146, new_n21147, new_n21148, new_n21149, new_n21150,
    new_n21151, new_n21152, new_n21153, new_n21154_1, new_n21155,
    new_n21156, new_n21157_1, new_n21158, new_n21159, new_n21160,
    new_n21161, new_n21162, new_n21163, new_n21164, new_n21165, new_n21166,
    new_n21167, new_n21168_1, new_n21169, new_n21170, new_n21171,
    new_n21172, new_n21173_1, new_n21174, new_n21175, new_n21176_1,
    new_n21177, new_n21178, new_n21179, new_n21180, new_n21188, new_n21189,
    new_n21190, new_n21191, new_n21192, new_n21193_1, new_n21194,
    new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200,
    new_n21201, new_n21202, new_n21203_1, new_n21207, new_n21208,
    new_n21211, new_n21212, new_n21213, new_n21214, new_n21215, new_n21216,
    new_n21217, new_n21220, new_n21221, new_n21222_1, new_n21223,
    new_n21224, new_n21225_1, new_n21226_1, new_n21227, new_n21228,
    new_n21229, new_n21230, new_n21231, new_n21232, new_n21233, new_n21234,
    new_n21235, new_n21236, new_n21237, new_n21240, new_n21241, new_n21242,
    new_n21243, new_n21244, new_n21245, new_n21246, new_n21247, new_n21248,
    new_n21249, new_n21250, new_n21251, new_n21252, new_n21253,
    new_n21254_1, new_n21255, new_n21256, new_n21257, new_n21258,
    new_n21259, new_n21260, new_n21261, new_n21262, new_n21263, new_n21264,
    new_n21265, new_n21266, new_n21267, new_n21268, new_n21269, new_n21270,
    new_n21271, new_n21272, new_n21273, new_n21274, new_n21275,
    new_n21276_1, new_n21277, new_n21278, new_n21299, new_n21303,
    new_n21304, new_n21305, new_n21306, new_n21307, new_n21308, new_n21309,
    new_n21310, new_n21311, new_n21312, new_n21313, new_n21314, new_n21315,
    new_n21318, new_n21319, new_n21320, new_n21321, new_n21322, new_n21323,
    new_n21324, new_n21325, new_n21326, new_n21327, new_n21328, new_n21329,
    new_n21330, new_n21331, new_n21332, new_n21333, new_n21334, new_n21335,
    new_n21336, new_n21337, new_n21341, new_n21342, new_n21343, new_n21344,
    new_n21345, new_n21346, new_n21350, new_n21355, new_n21356, new_n21357,
    new_n21358, new_n21359, new_n21360, new_n21361, new_n21362, new_n21364,
    new_n21365_1, new_n21366, new_n21367_1, new_n21368, new_n21369,
    new_n21370, new_n21371, new_n21372, new_n21373, new_n21374, new_n21375,
    new_n21376, new_n21377, new_n21378, new_n21379, new_n21380, new_n21381,
    new_n21382, new_n21383, new_n21404_1, new_n21407, new_n21408,
    new_n21409, new_n21410, new_n21411, new_n21412, new_n21413, new_n21414,
    new_n21415, new_n21416, new_n21417, new_n21418, new_n21419, new_n21420,
    new_n21421, new_n21422, new_n21423, new_n21424, new_n21425, new_n21426,
    new_n21427, new_n21432, new_n21433, new_n21434, new_n21435, new_n21447,
    new_n21450, new_n21465, new_n21466, new_n21467, new_n21468, new_n21469,
    new_n21483, new_n21484, new_n21485, new_n21486, new_n21487, new_n21488,
    new_n21489_1, new_n21493, new_n21494, new_n21495, new_n21496,
    new_n21497, new_n21498, new_n21499, new_n21504, new_n21505, new_n21506,
    new_n21507, new_n21508, new_n21509, new_n21510, new_n21511, new_n21514,
    new_n21515, new_n21516, new_n21531, new_n21532, new_n21533, new_n21536,
    new_n21537, new_n21538_1, new_n21539, new_n21547, new_n21548,
    new_n21557, new_n21567, new_n21568, new_n21569, new_n21570, new_n21571,
    new_n21572, new_n21573, new_n21574, new_n21575, new_n21584, new_n21585,
    new_n21586, new_n21587, new_n21588, new_n21589, new_n21590, new_n21591,
    new_n21592, new_n21594, new_n21595, new_n21596, new_n21597, new_n21608,
    new_n21609, new_n21611, new_n21612, new_n21613, new_n21614,
    new_n21615_1, new_n21616, new_n21617, new_n21618, new_n21619,
    new_n21620, new_n21621, new_n21622, new_n21623, new_n21624, new_n21625,
    new_n21643, new_n21644, new_n21645_1, new_n21646, new_n21647,
    new_n21648, new_n21649_1, new_n21650, new_n21651, new_n21652,
    new_n21653, new_n21654_1, new_n21655, new_n21656, new_n21659,
    new_n21660, new_n21661, new_n21666, new_n21667, new_n21668, new_n21669,
    new_n21670, new_n21671, new_n21672, new_n21673, new_n21674_1,
    new_n21677, new_n21678, new_n21679, new_n21680_1, new_n21681,
    new_n21684, new_n21685_1, new_n21686, new_n21687_1, new_n21688,
    new_n21690, new_n21691, new_n21692, new_n21693, new_n21694, new_n21695,
    new_n21696, new_n21697, new_n21698, new_n21699, new_n21700, new_n21701,
    new_n21702, new_n21703, new_n21704, new_n21705, new_n21706, new_n21707,
    new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713,
    new_n21717_1, new_n21718, new_n21719_1, new_n21720, new_n21721,
    new_n21722, new_n21736, new_n21737, new_n21748, new_n21755, new_n21756,
    new_n21757, new_n21758, new_n21759, new_n21760, new_n21768, new_n21787,
    new_n21809, new_n21810, new_n21824, new_n21825, new_n21826, new_n21827,
    new_n21828, new_n21829, new_n21830, new_n21831, new_n21832_1,
    new_n21839_1, new_n21847, new_n21848, new_n21849, new_n21850,
    new_n21851, new_n21852, new_n21853, new_n21854, new_n21855, new_n21856,
    new_n21857, new_n21858, new_n21859, new_n21865, new_n21866, new_n21867,
    new_n21868, new_n21869, new_n21870, new_n21871, new_n21872, new_n21875,
    new_n21876, new_n21877, new_n21878, new_n21884, new_n21885, new_n21886,
    new_n21888, new_n21889, new_n21890, new_n21891, new_n21892, new_n21893,
    new_n21894, new_n21895, new_n21896, new_n21897, new_n21898_1,
    new_n21899, new_n21900, new_n21901, new_n21902, new_n21914, new_n21942,
    new_n21943_1, new_n21944, new_n21945, new_n21956, new_n21962,
    new_n21963, new_n21964, new_n21965, new_n21966, new_n21981_1,
    new_n21988, new_n21989, new_n21990, new_n21991, new_n21992,
    new_n21993_1, new_n21994, new_n21995, new_n22010, new_n22011,
    new_n22012, new_n22013, new_n22014, new_n22015, new_n22016_1,
    new_n22021, new_n22022, new_n22028, new_n22029, new_n22030, new_n22031,
    new_n22032, new_n22033, new_n22034, new_n22035, new_n22036, new_n22037,
    new_n22038, new_n22051, new_n22052, new_n22053, new_n22057, new_n22062,
    new_n22063_1, new_n22064, new_n22065, new_n22072_1, new_n22073,
    new_n22074, new_n22075, new_n22076_1, new_n22077, new_n22078,
    new_n22084, new_n22085, new_n22093, new_n22094, new_n22095, new_n22096,
    new_n22097, new_n22098, new_n22099, new_n22102, new_n22105, new_n22106,
    new_n22107_1, new_n22108, new_n22109, new_n22122, new_n22123,
    new_n22124_1, new_n22125, new_n22127, new_n22138, new_n22139,
    new_n22140, new_n22141, new_n22144_1, new_n22152, new_n22153,
    new_n22154, new_n22155, new_n22156, new_n22157_1, new_n22158,
    new_n22159, new_n22160, new_n22162, new_n22167, new_n22168, new_n22169,
    new_n22170, new_n22172, new_n22173_1, new_n22174, new_n22175,
    new_n22180, new_n22181, new_n22182, new_n22183, new_n22184, new_n22185,
    new_n22186, new_n22187, new_n22188, new_n22189, new_n22190, new_n22191,
    new_n22192, new_n22193, new_n22194, new_n22195, new_n22196, new_n22197,
    new_n22198_1, new_n22199, new_n22200, new_n22201_1, new_n22202,
    new_n22207, new_n22208, new_n22209, new_n22210, new_n22214, new_n22224,
    new_n22225, new_n22226, new_n22227, new_n22228, new_n22229, new_n22230,
    new_n22249, new_n22250, new_n22251, new_n22252, new_n22253_1,
    new_n22254, new_n22256, new_n22257, new_n22258, new_n22259, new_n22260,
    new_n22261, new_n22272, new_n22284, new_n22285, new_n22286,
    new_n22290_1, new_n22291, new_n22292, new_n22293, new_n22295,
    new_n22296, new_n22297, new_n22299, new_n22309_1, new_n22310,
    new_n22311_1, new_n22312, new_n22313, new_n22314, new_n22323,
    new_n22334, new_n22343, new_n22352, new_n22353_1, new_n22363,
    new_n22364, new_n22365, new_n22366, new_n22367, new_n22373, new_n22374,
    new_n22375, new_n22376, new_n22379_1, new_n22380, new_n22381,
    new_n22382, new_n22403, new_n22423, new_n22433_1, new_n22434,
    new_n22435, new_n22436, new_n22450, new_n22451, new_n22466, new_n22482,
    new_n22487, new_n22490, new_n22491, new_n22497, new_n22498, new_n22499,
    new_n22503, new_n22504, new_n22505, new_n22506, new_n22508, new_n22521,
    new_n22524, new_n22525, new_n22526, new_n22527, new_n22530,
    new_n22533_1, new_n22534, new_n22535, new_n22536, new_n22537,
    new_n22551, new_n22552, new_n22555, new_n22567, new_n22569, new_n22570,
    new_n22571, new_n22572, new_n22575, new_n22576, new_n22586,
    new_n22588_1, new_n22593, new_n22594, new_n22595, new_n22596,
    new_n22602, new_n22603, new_n22613, new_n22627, new_n22636, new_n22637,
    new_n22640;
xor_4  g00000(n10739, n9942, new_n2349);
not_10 g00001(n21753, new_n2350);
nor_5  g00002(n25643, new_n2350, new_n2351);
xor_4  g00003(n25643, n21753, new_n2352);
not_10 g00004(n21832, new_n2353);
or_5   g00005(new_n2353, n9557, new_n2354);
xor_4  g00006(n21832, n9557, new_n2355_1);
not_10 g00007(n26913, new_n2356);
or_5   g00008(new_n2356, n3136, new_n2357);
xor_4  g00009(n26913, n3136, new_n2358);
not_10 g00010(n6385, new_n2359);
nor_5  g00011(n16223, new_n2359, new_n2360);
and_5  g00012(n16223, new_n2359, new_n2361_1);
not_10 g00013(n20138, new_n2362);
nor_5  g00014(new_n2362, n19494, new_n2363_1);
not_10 g00015(n19494, new_n2364);
or_5   g00016(n20138, new_n2364, new_n2365);
not_10 g00017(n9251, new_n2366);
nor_5  g00018(new_n2366, n2387, new_n2367);
and_5  g00019(new_n2367, new_n2365, new_n2368);
nor_5  g00020(new_n2368, new_n2363_1, new_n2369);
nor_5  g00021(new_n2369, new_n2361_1, new_n2370);
nor_5  g00022(new_n2370, new_n2360, new_n2371);
not_10 g00023(new_n2371, new_n2372);
or_5   g00024(new_n2372, new_n2358, new_n2373);
and_5  g00025(new_n2373, new_n2357, new_n2374_1);
or_5   g00026(new_n2374_1, new_n2355_1, new_n2375);
and_5  g00027(new_n2375, new_n2354, new_n2376);
nor_5  g00028(new_n2376, new_n2352, new_n2377);
nor_5  g00029(new_n2377, new_n2351, new_n2378);
xnor_4 g00030(new_n2378, new_n2349, new_n2379);
xor_4  g00031(n13781, n5704, new_n2380);
and_5  g00032(n13781, n5704, new_n2381);
xnor_4 g00033(n18409, n11486, new_n2382);
xnor_4 g00034(new_n2382, new_n2381, new_n2383);
nor_5  g00035(new_n2383, new_n2380, new_n2384);
xnor_4 g00036(n16722, n13708, new_n2385);
or_5   g00037(n18409, n11486, new_n2386);
or_5   g00038(new_n2382, new_n2381, new_n2387_1);
and_5  g00039(new_n2387_1, new_n2386, new_n2388_1);
xor_4  g00040(new_n2388_1, new_n2385, new_n2389);
nand_5 g00041(new_n2389, new_n2384, new_n2390);
xnor_4 g00042(n19911, n3480, new_n2391);
nor_5  g00043(n16722, n13708, new_n2392);
nor_5  g00044(new_n2388_1, new_n2385, new_n2393);
nor_5  g00045(new_n2393, new_n2392, new_n2394);
xor_4  g00046(new_n2394, new_n2391, new_n2395);
not_10 g00047(new_n2395, new_n2396);
or_5   g00048(new_n2396, new_n2390, new_n2397);
xnor_4 g00049(n3018, n2731, new_n2398);
nor_5  g00050(n19911, n3480, new_n2399);
nor_5  g00051(new_n2394, new_n2391, new_n2400);
nor_5  g00052(new_n2400, new_n2399, new_n2401);
xor_4  g00053(new_n2401, new_n2398, new_n2402);
not_10 g00054(new_n2402, new_n2403);
or_5   g00055(new_n2403, new_n2397, new_n2404);
xnor_4 g00056(n26660, n18907, new_n2405);
nor_5  g00057(n3018, n2731, new_n2406);
nor_5  g00058(new_n2401, new_n2398, new_n2407);
nor_5  g00059(new_n2407, new_n2406, new_n2408);
xnor_4 g00060(new_n2408, new_n2405, new_n2409_1);
or_5   g00061(new_n2409_1, new_n2404, new_n2410);
xnor_4 g00062(n22332, n13783, new_n2411);
nor_5  g00063(n26660, n18907, new_n2412);
nor_5  g00064(new_n2408, new_n2405, new_n2413);
nor_5  g00065(new_n2413, new_n2412, new_n2414);
xor_4  g00066(new_n2414, new_n2411, new_n2415);
xnor_4 g00067(new_n2415, new_n2410, new_n2416_1);
xnor_4 g00068(n13490, n7751, new_n2417);
nor_5  g00069(n26823, n22660, new_n2418);
xnor_4 g00070(n26823, n22660, new_n2419);
nor_5  g00071(n4812, n1777, new_n2420_1);
xnor_4 g00072(n4812, n1777, new_n2421_1);
nor_5  g00073(n24278, n8745, new_n2422);
xnor_4 g00074(n24278, n8745, new_n2423);
nor_5  g00075(n24618, n15636, new_n2424);
xor_4  g00076(n24618, n15636, new_n2425);
and_5  g00077(n20077, n3952, new_n2426);
or_5   g00078(n20077, n3952, new_n2427);
and_5  g00079(n12315, n6794, new_n2428);
and_5  g00080(new_n2428, new_n2427, new_n2429);
nor_5  g00081(new_n2429, new_n2426, new_n2430);
and_5  g00082(new_n2430, new_n2425, new_n2431);
nor_5  g00083(new_n2431, new_n2424, new_n2432);
nor_5  g00084(new_n2432, new_n2423, new_n2433);
nor_5  g00085(new_n2433, new_n2422, new_n2434);
nor_5  g00086(new_n2434, new_n2421_1, new_n2435);
nor_5  g00087(new_n2435, new_n2420_1, new_n2436);
nor_5  g00088(new_n2436, new_n2419, new_n2437);
nor_5  g00089(new_n2437, new_n2418, new_n2438);
xor_4  g00090(new_n2438, new_n2417, new_n2439);
not_10 g00091(new_n2439, new_n2440_1);
xnor_4 g00092(new_n2440_1, new_n2416_1, new_n2441);
xor_4  g00093(new_n2409_1, new_n2404, new_n2442);
xor_4  g00094(new_n2436, new_n2419, new_n2443);
not_10 g00095(new_n2443, new_n2444_1);
nor_5  g00096(new_n2444_1, new_n2442, new_n2445);
xnor_4 g00097(new_n2402, new_n2397, new_n2446);
xor_4  g00098(new_n2434, new_n2421_1, new_n2447);
not_10 g00099(new_n2447, new_n2448);
nor_5  g00100(new_n2448, new_n2446, new_n2449);
xnor_4 g00101(new_n2448, new_n2446, new_n2450);
xnor_4 g00102(new_n2395, new_n2390, new_n2451);
xor_4  g00103(new_n2432, new_n2423, new_n2452);
not_10 g00104(new_n2452, new_n2453);
nor_5  g00105(new_n2453, new_n2451, new_n2454);
xnor_4 g00106(new_n2388_1, new_n2385, new_n2455);
xnor_4 g00107(new_n2455, new_n2384, new_n2456);
xor_4  g00108(new_n2430, new_n2425, new_n2457);
not_10 g00109(new_n2457, new_n2458);
nor_5  g00110(new_n2458, new_n2456, new_n2459);
xor_4  g00111(new_n2457, new_n2456, new_n2460);
not_10 g00112(new_n2380, new_n2461);
xnor_4 g00113(n12315, n6794, new_n2462);
or_5   g00114(new_n2462, new_n2461, new_n2463);
xnor_4 g00115(n20077, n3952, new_n2464);
xnor_4 g00116(new_n2464, new_n2428, new_n2465);
not_10 g00117(new_n2465, new_n2466);
and_5  g00118(new_n2466, new_n2463, new_n2467);
nor_5  g00119(n13781, n5704, new_n2468);
nor_5  g00120(new_n2387_1, new_n2468, new_n2469);
nor_5  g00121(new_n2469, new_n2384, new_n2470);
nor_5  g00122(new_n2464, new_n2463, new_n2471);
or_5   g00123(new_n2471, new_n2467, new_n2472);
nor_5  g00124(new_n2472, new_n2470, new_n2473);
nor_5  g00125(new_n2473, new_n2467, new_n2474);
nor_5  g00126(new_n2474, new_n2460, new_n2475);
nor_5  g00127(new_n2475, new_n2459, new_n2476);
xor_4  g00128(new_n2452, new_n2451, new_n2477);
nor_5  g00129(new_n2477, new_n2476, new_n2478);
nor_5  g00130(new_n2478, new_n2454, new_n2479_1);
nor_5  g00131(new_n2479_1, new_n2450, new_n2480);
nor_5  g00132(new_n2480, new_n2449, new_n2481);
xnor_4 g00133(new_n2444_1, new_n2442, new_n2482);
nor_5  g00134(new_n2482, new_n2481, new_n2483);
nor_5  g00135(new_n2483, new_n2445, new_n2484);
xor_4  g00136(new_n2484, new_n2441, new_n2485);
xnor_4 g00137(new_n2485, new_n2379, new_n2486);
xnor_4 g00138(new_n2376, new_n2352, new_n2487);
xor_4  g00139(new_n2482, new_n2481, new_n2488);
and_5  g00140(new_n2488, new_n2487, new_n2489);
xnor_4 g00141(new_n2488, new_n2487, new_n2490);
xnor_4 g00142(new_n2374_1, new_n2355_1, new_n2491);
xor_4  g00143(new_n2479_1, new_n2450, new_n2492);
and_5  g00144(new_n2492, new_n2491, new_n2493);
xnor_4 g00145(new_n2492, new_n2491, new_n2494);
xor_4  g00146(new_n2371, new_n2358, new_n2495);
xor_4  g00147(new_n2477, new_n2476, new_n2496);
and_5  g00148(new_n2496, new_n2495, new_n2497);
xnor_4 g00149(new_n2496, new_n2495, new_n2498);
xor_4  g00150(new_n2474, new_n2460, new_n2499);
xnor_4 g00151(n16223, n6385, new_n2500);
xnor_4 g00152(new_n2500, new_n2369, new_n2501);
and_5  g00153(new_n2501, new_n2499, new_n2502);
xnor_4 g00154(new_n2501, new_n2499, new_n2503);
xnor_4 g00155(n9251, n2387, new_n2504);
xor_4  g00156(new_n2462, new_n2380, new_n2505);
or_5   g00157(new_n2505, new_n2504, new_n2506);
xor_4  g00158(n20138, n19494, new_n2507);
xnor_4 g00159(new_n2507, new_n2367, new_n2508);
and_5  g00160(new_n2508, new_n2506, new_n2509);
xor_4  g00161(new_n2472, new_n2470, new_n2510);
xor_4  g00162(new_n2508, new_n2506, new_n2511);
and_5  g00163(new_n2511, new_n2510, new_n2512);
nor_5  g00164(new_n2512, new_n2509, new_n2513_1);
nor_5  g00165(new_n2513_1, new_n2503, new_n2514);
nor_5  g00166(new_n2514, new_n2502, new_n2515_1);
nor_5  g00167(new_n2515_1, new_n2498, new_n2516);
nor_5  g00168(new_n2516, new_n2497, new_n2517);
nor_5  g00169(new_n2517, new_n2494, new_n2518);
nor_5  g00170(new_n2518, new_n2493, new_n2519);
nor_5  g00171(new_n2519, new_n2490, new_n2520);
or_5   g00172(new_n2520, new_n2489, new_n2521);
xor_4  g00173(new_n2521, new_n2486, n7);
xnor_4 g00174(n3618, n1681, new_n2523);
xor_4  g00175(new_n2523, n4588, new_n2524);
xnor_4 g00176(n22843, n583, new_n2525);
xnor_4 g00177(new_n2525, n22201, new_n2526);
xnor_4 g00178(new_n2526, new_n2524, n50);
xor_4  g00179(n19922, n6773, new_n2528);
xnor_4 g00180(new_n2528, n21687, new_n2529);
xor_4  g00181(n21398, n14090, new_n2530);
xnor_4 g00182(new_n2530, n25926, new_n2531);
xor_4  g00183(new_n2531, new_n2529, n55);
xnor_4 g00184(n20040, n9396, new_n2533_1);
nor_5  g00185(n19531, n1999, new_n2534);
xnor_4 g00186(n19531, n1999, new_n2535_1);
nor_5  g00187(n25168, n18345, new_n2536);
xnor_4 g00188(n25168, n18345, new_n2537_1);
nor_5  g00189(n13190, n9318, new_n2538);
xnor_4 g00190(n13190, n9318, new_n2539);
nor_5  g00191(n19477, n3460, new_n2540);
xnor_4 g00192(n19477, n3460, new_n2541);
nor_5  g00193(n11223, n5226, new_n2542);
xnor_4 g00194(n11223, n5226, new_n2543);
nor_5  g00195(n17664, n5115, new_n2544);
xnor_4 g00196(n17664, n5115, new_n2545);
nor_5  g00197(n26572, n23369, new_n2546);
xnor_4 g00198(n26572, n23369, new_n2547_1);
nor_5  g00199(n11667, n1136, new_n2548);
and_5  g00200(n21398, n19234, new_n2549);
xnor_4 g00201(n11667, n1136, new_n2550);
nor_5  g00202(new_n2550, new_n2549, new_n2551);
nor_5  g00203(new_n2551, new_n2548, new_n2552);
nor_5  g00204(new_n2552, new_n2547_1, new_n2553_1);
nor_5  g00205(new_n2553_1, new_n2546, new_n2554);
nor_5  g00206(new_n2554, new_n2545, new_n2555_1);
nor_5  g00207(new_n2555_1, new_n2544, new_n2556);
nor_5  g00208(new_n2556, new_n2543, new_n2557);
nor_5  g00209(new_n2557, new_n2542, new_n2558);
nor_5  g00210(new_n2558, new_n2541, new_n2559);
nor_5  g00211(new_n2559, new_n2540, new_n2560_1);
nor_5  g00212(new_n2560_1, new_n2539, new_n2561_1);
nor_5  g00213(new_n2561_1, new_n2538, new_n2562);
nor_5  g00214(new_n2562, new_n2537_1, new_n2563);
nor_5  g00215(new_n2563, new_n2536, new_n2564);
nor_5  g00216(new_n2564, new_n2535_1, new_n2565);
nor_5  g00217(new_n2565, new_n2534, new_n2566);
xnor_4 g00218(new_n2566, new_n2533_1, new_n2567);
xnor_4 g00219(new_n2567, n25365, new_n2568);
xnor_4 g00220(new_n2564, new_n2535_1, new_n2569);
and_5  g00221(new_n2569, n14704, new_n2570_1);
xnor_4 g00222(new_n2569, n14704, new_n2571);
xnor_4 g00223(new_n2562, new_n2537_1, new_n2572);
and_5  g00224(new_n2572, n19270, new_n2573_1);
xnor_4 g00225(new_n2572, n19270, new_n2574);
xnor_4 g00226(new_n2560_1, new_n2539, new_n2575);
and_5  g00227(new_n2575, n8687, new_n2576);
xnor_4 g00228(new_n2558, new_n2541, new_n2577);
nor_5  g00229(new_n2577, n24768, new_n2578_1);
xnor_4 g00230(new_n2577, n24768, new_n2579);
xnor_4 g00231(new_n2556, new_n2543, new_n2580);
or_5   g00232(new_n2580, n26483, new_n2581);
xnor_4 g00233(new_n2580, n26483, new_n2582_1);
xnor_4 g00234(new_n2554, new_n2545, new_n2583);
and_5  g00235(new_n2583, n15979, new_n2584);
xnor_4 g00236(new_n2583, n15979, new_n2585);
xnor_4 g00237(new_n2552, new_n2547_1, new_n2586);
and_5  g00238(new_n2586, n8638, new_n2587);
xor_4  g00239(new_n2550, new_n2549, new_n2588);
not_10 g00240(new_n2588, new_n2589);
nor_5  g00241(new_n2589, n16247, new_n2590);
xor_4  g00242(n21398, n19234, new_n2591);
nand_5 g00243(new_n2591, n23541, new_n2592);
xnor_4 g00244(new_n2588, n16247, new_n2593);
and_5  g00245(new_n2593, new_n2592, new_n2594);
nor_5  g00246(new_n2594, new_n2590, new_n2595);
xor_4  g00247(new_n2586, n8638, new_n2596);
and_5  g00248(new_n2596, new_n2595, new_n2597);
nor_5  g00249(new_n2597, new_n2587, new_n2598);
nor_5  g00250(new_n2598, new_n2585, new_n2599);
nor_5  g00251(new_n2599, new_n2584, new_n2600);
not_10 g00252(new_n2600, new_n2601);
or_5   g00253(new_n2601, new_n2582_1, new_n2602_1);
and_5  g00254(new_n2602_1, new_n2581, new_n2603);
nor_5  g00255(new_n2603, new_n2579, new_n2604);
or_5   g00256(new_n2604, new_n2578_1, new_n2605);
xnor_4 g00257(new_n2575, n8687, new_n2606);
nor_5  g00258(new_n2606, new_n2605, new_n2607);
nor_5  g00259(new_n2607, new_n2576, new_n2608);
nor_5  g00260(new_n2608, new_n2574, new_n2609);
nor_5  g00261(new_n2609, new_n2573_1, new_n2610);
nor_5  g00262(new_n2610, new_n2571, new_n2611);
nor_5  g00263(new_n2611, new_n2570_1, new_n2612);
xnor_4 g00264(new_n2612, new_n2568, new_n2613);
or_5   g00265(n18151, n11503, new_n2614);
or_5   g00266(new_n2614, n16971, new_n2615);
or_5   g00267(new_n2615, n10411, new_n2616);
or_5   g00268(new_n2616, n23430, new_n2617);
or_5   g00269(new_n2617, n5579, new_n2618);
or_5   g00270(new_n2618, n25523, new_n2619_1);
or_5   g00271(new_n2619_1, n8439, new_n2620);
or_5   g00272(new_n2620, n22793, new_n2621);
xnor_4 g00273(new_n2621, n13951, new_n2622);
xnor_4 g00274(n22270, n2944, new_n2623);
nor_5  g00275(n8806, n767, new_n2624);
xnor_4 g00276(n8806, n767, new_n2625);
nor_5  g00277(n7330, n2479, new_n2626);
xnor_4 g00278(n7330, n2479, new_n2627);
nor_5  g00279(n22492, n9372, new_n2628);
xnor_4 g00280(n22492, n9372, new_n2629);
nor_5  g00281(n12821, n6596, new_n2630);
xnor_4 g00282(n12821, n6596, new_n2631);
nor_5  g00283(n15289, n3468, new_n2632);
xnor_4 g00284(n15289, n3468, new_n2633);
nor_5  g00285(n18558, n6556, new_n2634);
xnor_4 g00286(n18558, n6556, new_n2635);
nor_5  g00287(n22871, n7149, new_n2636);
xnor_4 g00288(n22871, n7149, new_n2637);
nor_5  g00289(n14275, n14148, new_n2638);
and_5  g00290(n25023, n1152, new_n2639);
xnor_4 g00291(n14275, n14148, new_n2640);
nor_5  g00292(new_n2640, new_n2639, new_n2641);
nor_5  g00293(new_n2641, new_n2638, new_n2642);
nor_5  g00294(new_n2642, new_n2637, new_n2643);
nor_5  g00295(new_n2643, new_n2636, new_n2644);
nor_5  g00296(new_n2644, new_n2635, new_n2645);
nor_5  g00297(new_n2645, new_n2634, new_n2646_1);
nor_5  g00298(new_n2646_1, new_n2633, new_n2647);
nor_5  g00299(new_n2647, new_n2632, new_n2648);
nor_5  g00300(new_n2648, new_n2631, new_n2649);
nor_5  g00301(new_n2649, new_n2630, new_n2650);
nor_5  g00302(new_n2650, new_n2629, new_n2651);
nor_5  g00303(new_n2651, new_n2628, new_n2652);
nor_5  g00304(new_n2652, new_n2627, new_n2653);
nor_5  g00305(new_n2653, new_n2626, new_n2654);
nor_5  g00306(new_n2654, new_n2625, new_n2655);
nor_5  g00307(new_n2655, new_n2624, new_n2656);
xor_4  g00308(new_n2656, new_n2623, new_n2657);
xor_4  g00309(new_n2657, new_n2622, new_n2658);
xnor_4 g00310(new_n2620, n22793, new_n2659_1);
xor_4  g00311(new_n2654, new_n2625, new_n2660);
not_10 g00312(new_n2660, new_n2661_1);
nor_5  g00313(new_n2661_1, new_n2659_1, new_n2662);
xnor_4 g00314(new_n2660, new_n2659_1, new_n2663);
xor_4  g00315(new_n2619_1, n8439, new_n2664);
xor_4  g00316(new_n2652, new_n2627, new_n2665);
nor_5  g00317(new_n2665, new_n2664, new_n2666);
xnor_4 g00318(new_n2665, new_n2664, new_n2667);
xor_4  g00319(new_n2618, n25523, new_n2668);
xor_4  g00320(new_n2650, new_n2629, new_n2669);
nor_5  g00321(new_n2669, new_n2668, new_n2670);
xnor_4 g00322(new_n2669, new_n2668, new_n2671);
xor_4  g00323(new_n2617, n5579, new_n2672);
xor_4  g00324(new_n2648, new_n2631, new_n2673);
nor_5  g00325(new_n2673, new_n2672, new_n2674);
xnor_4 g00326(new_n2673, new_n2672, new_n2675);
xor_4  g00327(new_n2616, n23430, new_n2676);
xor_4  g00328(new_n2646_1, new_n2633, new_n2677);
nor_5  g00329(new_n2677, new_n2676, new_n2678);
xor_4  g00330(new_n2615, n10411, new_n2679);
xor_4  g00331(new_n2644, new_n2635, new_n2680_1);
nor_5  g00332(new_n2680_1, new_n2679, new_n2681);
xnor_4 g00333(new_n2680_1, new_n2679, new_n2682);
xor_4  g00334(new_n2614, n16971, new_n2683);
xor_4  g00335(new_n2642, new_n2637, new_n2684);
nor_5  g00336(new_n2684, new_n2683, new_n2685);
xnor_4 g00337(new_n2684, new_n2683, new_n2686);
xor_4  g00338(n18151, n11503, new_n2687);
xor_4  g00339(new_n2640, new_n2639, new_n2688);
nor_5  g00340(new_n2688, new_n2687, new_n2689);
xnor_4 g00341(n25023, n1152, new_n2690);
nor_5  g00342(new_n2690, n18151, new_n2691);
xor_4  g00343(new_n2688, new_n2687, new_n2692);
and_5  g00344(new_n2692, new_n2691, new_n2693_1);
nor_5  g00345(new_n2693_1, new_n2689, new_n2694);
nor_5  g00346(new_n2694, new_n2686, new_n2695);
nor_5  g00347(new_n2695, new_n2685, new_n2696);
nor_5  g00348(new_n2696, new_n2682, new_n2697);
nor_5  g00349(new_n2697, new_n2681, new_n2698);
xnor_4 g00350(new_n2677, new_n2676, new_n2699);
nor_5  g00351(new_n2699, new_n2698, new_n2700);
nor_5  g00352(new_n2700, new_n2678, new_n2701);
nor_5  g00353(new_n2701, new_n2675, new_n2702);
nor_5  g00354(new_n2702, new_n2674, new_n2703_1);
nor_5  g00355(new_n2703_1, new_n2671, new_n2704);
nor_5  g00356(new_n2704, new_n2670, new_n2705);
nor_5  g00357(new_n2705, new_n2667, new_n2706_1);
nor_5  g00358(new_n2706_1, new_n2666, new_n2707);
and_5  g00359(new_n2707, new_n2663, new_n2708);
nor_5  g00360(new_n2708, new_n2662, new_n2709);
xor_4  g00361(new_n2709, new_n2658, new_n2710);
xnor_4 g00362(new_n2710, new_n2613, new_n2711_1);
xor_4  g00363(new_n2610, new_n2571, new_n2712);
xor_4  g00364(new_n2707, new_n2663, new_n2713);
and_5  g00365(new_n2713, new_n2712, new_n2714);
xnor_4 g00366(new_n2713, new_n2712, new_n2715);
xnor_4 g00367(new_n2608, new_n2574, new_n2716);
xor_4  g00368(new_n2705, new_n2667, new_n2717);
and_5  g00369(new_n2717, new_n2716, new_n2718);
xnor_4 g00370(new_n2717, new_n2716, new_n2719);
nor_5  g00371(new_n2604, new_n2578_1, new_n2720);
xor_4  g00372(new_n2606, new_n2720, new_n2721);
xor_4  g00373(new_n2703_1, new_n2671, new_n2722);
and_5  g00374(new_n2722, new_n2721, new_n2723);
xnor_4 g00375(new_n2606, new_n2720, new_n2724);
xnor_4 g00376(new_n2722, new_n2724, new_n2725);
xor_4  g00377(new_n2603, new_n2579, new_n2726);
xor_4  g00378(new_n2701, new_n2675, new_n2727);
nor_5  g00379(new_n2727, new_n2726, new_n2728);
xnor_4 g00380(new_n2727, new_n2726, new_n2729);
xnor_4 g00381(new_n2600, new_n2582_1, new_n2730);
xor_4  g00382(new_n2699, new_n2698, new_n2731_1);
and_5  g00383(new_n2731_1, new_n2730, new_n2732);
xnor_4 g00384(new_n2731_1, new_n2730, new_n2733);
xnor_4 g00385(new_n2696, new_n2682, new_n2734);
xor_4  g00386(new_n2598, new_n2585, new_n2735);
nor_5  g00387(new_n2735, new_n2734, new_n2736);
xor_4  g00388(new_n2735, new_n2734, new_n2737);
xnor_4 g00389(new_n2694, new_n2686, new_n2738);
xor_4  g00390(new_n2596, new_n2595, new_n2739);
and_5  g00391(new_n2739, new_n2738, new_n2740);
xnor_4 g00392(new_n2739, new_n2738, new_n2741);
xnor_4 g00393(new_n2692, new_n2691, new_n2742);
xor_4  g00394(new_n2593, new_n2592, new_n2743_1);
not_10 g00395(new_n2743_1, new_n2744);
nor_5  g00396(new_n2744, new_n2742, new_n2745);
xnor_4 g00397(new_n2591, n23541, new_n2746);
xor_4  g00398(new_n2690, n18151, new_n2747);
or_5   g00399(new_n2747, new_n2746, new_n2748);
xnor_4 g00400(new_n2743_1, new_n2742, new_n2749);
and_5  g00401(new_n2749, new_n2748, new_n2750);
or_5   g00402(new_n2750, new_n2745, new_n2751);
nor_5  g00403(new_n2751, new_n2741, new_n2752);
nor_5  g00404(new_n2752, new_n2740, new_n2753);
and_5  g00405(new_n2753, new_n2737, new_n2754);
nor_5  g00406(new_n2754, new_n2736, new_n2755);
nor_5  g00407(new_n2755, new_n2733, new_n2756);
or_5   g00408(new_n2756, new_n2732, new_n2757);
nor_5  g00409(new_n2757, new_n2729, new_n2758);
nor_5  g00410(new_n2758, new_n2728, new_n2759);
and_5  g00411(new_n2759, new_n2725, new_n2760);
nor_5  g00412(new_n2760, new_n2723, new_n2761_1);
nor_5  g00413(new_n2761_1, new_n2719, new_n2762);
or_5   g00414(new_n2762, new_n2718, new_n2763);
nor_5  g00415(new_n2763, new_n2715, new_n2764);
nor_5  g00416(new_n2764, new_n2714, new_n2765);
xnor_4 g00417(new_n2765, new_n2711_1, n108);
xor_4  g00418(n22379, n767, new_n2767);
not_10 g00419(n1662, new_n2768);
nor_5  g00420(n7330, new_n2768, new_n2769);
xor_4  g00421(n7330, n1662, new_n2770);
not_10 g00422(n12875, new_n2771);
nor_5  g00423(n22492, new_n2771, new_n2772);
xor_4  g00424(n22492, n12875, new_n2773);
not_10 g00425(n2035, new_n2774_1);
nor_5  g00426(n12821, new_n2774_1, new_n2775);
xor_4  g00427(n12821, n2035, new_n2776);
not_10 g00428(n5213, new_n2777);
nor_5  g00429(new_n2777, n3468, new_n2778);
xor_4  g00430(n5213, n3468, new_n2779_1);
not_10 g00431(n4665, new_n2780);
nor_5  g00432(n18558, new_n2780, new_n2781);
xor_4  g00433(n18558, n4665, new_n2782);
not_10 g00434(n7149, new_n2783_1);
nor_5  g00435(n19005, new_n2783_1, new_n2784);
not_10 g00436(n19005, new_n2785);
nor_5  g00437(new_n2785, n7149, new_n2786);
not_10 g00438(n14148, new_n2787);
nor_5  g00439(new_n2787, n4326, new_n2788);
not_10 g00440(n4326, new_n2789);
or_5   g00441(n14148, new_n2789, new_n2790);
not_10 g00442(n5438, new_n2791);
and_5  g00443(new_n2791, n1152, new_n2792);
and_5  g00444(new_n2792, new_n2790, new_n2793);
nor_5  g00445(new_n2793, new_n2788, new_n2794);
nor_5  g00446(new_n2794, new_n2786, new_n2795);
or_5   g00447(new_n2795, new_n2784, new_n2796);
nor_5  g00448(new_n2796, new_n2782, new_n2797);
nor_5  g00449(new_n2797, new_n2781, new_n2798);
nor_5  g00450(new_n2798, new_n2779_1, new_n2799);
nor_5  g00451(new_n2799, new_n2778, new_n2800);
nor_5  g00452(new_n2800, new_n2776, new_n2801);
nor_5  g00453(new_n2801, new_n2775, new_n2802);
nor_5  g00454(new_n2802, new_n2773, new_n2803);
nor_5  g00455(new_n2803, new_n2772, new_n2804);
nor_5  g00456(new_n2804, new_n2770, new_n2805);
nor_5  g00457(new_n2805, new_n2769, new_n2806);
xor_4  g00458(new_n2806, new_n2767, new_n2807);
xnor_4 g00459(n10763, n6814, new_n2808);
nor_5  g00460(n19701, n7437, new_n2809_1);
xnor_4 g00461(n19701, n7437, new_n2810);
nor_5  g00462(n23529, n20700, new_n2811);
xnor_4 g00463(n23529, n20700, new_n2812);
nor_5  g00464(n24620, n7099, new_n2813);
xnor_4 g00465(n24620, n7099, new_n2814);
nor_5  g00466(n12811, n5211, new_n2815);
xnor_4 g00467(n12811, n5211, new_n2816_1);
nor_5  g00468(n12956, n1118, new_n2817);
xnor_4 g00469(n12956, n1118, new_n2818);
nor_5  g00470(n25974, n18295, new_n2819);
xnor_4 g00471(n25974, n18295, new_n2820);
nor_5  g00472(n6502, n1630, new_n2821);
and_5  g00473(n15780, n1451, new_n2822);
xnor_4 g00474(n6502, n1630, new_n2823);
nor_5  g00475(new_n2823, new_n2822, new_n2824);
nor_5  g00476(new_n2824, new_n2821, new_n2825);
nor_5  g00477(new_n2825, new_n2820, new_n2826_1);
nor_5  g00478(new_n2826_1, new_n2819, new_n2827);
nor_5  g00479(new_n2827, new_n2818, new_n2828);
nor_5  g00480(new_n2828, new_n2817, new_n2829);
nor_5  g00481(new_n2829, new_n2816_1, new_n2830);
nor_5  g00482(new_n2830, new_n2815, new_n2831);
nor_5  g00483(new_n2831, new_n2814, new_n2832);
nor_5  g00484(new_n2832, new_n2813, new_n2833);
nor_5  g00485(new_n2833, new_n2812, new_n2834);
nor_5  g00486(new_n2834, new_n2811, new_n2835);
nor_5  g00487(new_n2835, new_n2810, new_n2836);
nor_5  g00488(new_n2836, new_n2809_1, new_n2837);
xnor_4 g00489(new_n2837, new_n2808, new_n2838);
xnor_4 g00490(n27089, n12657, new_n2839);
nor_5  g00491(n17077, n11841, new_n2840);
xnor_4 g00492(n17077, n11841, new_n2841);
nor_5  g00493(n26510, n10710, new_n2842);
xnor_4 g00494(n26510, n10710, new_n2843);
nor_5  g00495(n23068, n20929, new_n2844);
xnor_4 g00496(n23068, n20929, new_n2845);
nor_5  g00497(n19514, n8006, new_n2846);
xnor_4 g00498(n19514, n8006, new_n2847);
nor_5  g00499(n25074, n10053, new_n2848);
xnor_4 g00500(n25074, n10053, new_n2849);
nor_5  g00501(n16396, n8399, new_n2850);
xnor_4 g00502(n16396, n8399, new_n2851);
nor_5  g00503(n9507, n9399, new_n2852);
and_5  g00504(n26979, n2088, new_n2853_1);
xnor_4 g00505(n9507, n9399, new_n2854);
nor_5  g00506(new_n2854, new_n2853_1, new_n2855);
nor_5  g00507(new_n2855, new_n2852, new_n2856);
nor_5  g00508(new_n2856, new_n2851, new_n2857);
nor_5  g00509(new_n2857, new_n2850, new_n2858_1);
nor_5  g00510(new_n2858_1, new_n2849, new_n2859);
nor_5  g00511(new_n2859, new_n2848, new_n2860_1);
nor_5  g00512(new_n2860_1, new_n2847, new_n2861);
nor_5  g00513(new_n2861, new_n2846, new_n2862);
nor_5  g00514(new_n2862, new_n2845, new_n2863);
nor_5  g00515(new_n2863, new_n2844, new_n2864);
nor_5  g00516(new_n2864, new_n2843, new_n2865);
nor_5  g00517(new_n2865, new_n2842, new_n2866);
nor_5  g00518(new_n2866, new_n2841, new_n2867);
nor_5  g00519(new_n2867, new_n2840, new_n2868);
xor_4  g00520(new_n2868, new_n2839, new_n2869);
xnor_4 g00521(new_n2869, new_n2838, new_n2870);
xnor_4 g00522(new_n2835, new_n2810, new_n2871);
xor_4  g00523(new_n2866, new_n2841, new_n2872);
and_5  g00524(new_n2872, new_n2871, new_n2873);
xnor_4 g00525(new_n2872, new_n2871, new_n2874);
xnor_4 g00526(new_n2833, new_n2812, new_n2875);
xor_4  g00527(new_n2864, new_n2843, new_n2876);
nor_5  g00528(new_n2876, new_n2875, new_n2877);
xnor_4 g00529(new_n2876, new_n2875, new_n2878);
xnor_4 g00530(new_n2831, new_n2814, new_n2879);
xor_4  g00531(new_n2862, new_n2845, new_n2880);
nor_5  g00532(new_n2880, new_n2879, new_n2881);
xnor_4 g00533(new_n2880, new_n2879, new_n2882);
xnor_4 g00534(new_n2829, new_n2816_1, new_n2883);
xor_4  g00535(new_n2860_1, new_n2847, new_n2884);
nor_5  g00536(new_n2884, new_n2883, new_n2885);
xnor_4 g00537(new_n2884, new_n2883, new_n2886_1);
xnor_4 g00538(new_n2827, new_n2818, new_n2887_1);
xor_4  g00539(new_n2858_1, new_n2849, new_n2888);
nor_5  g00540(new_n2888, new_n2887_1, new_n2889);
xor_4  g00541(new_n2888, new_n2887_1, new_n2890);
xnor_4 g00542(new_n2825, new_n2820, new_n2891);
xor_4  g00543(new_n2856, new_n2851, new_n2892);
and_5  g00544(new_n2892, new_n2891, new_n2893);
xor_4  g00545(new_n2892, new_n2891, new_n2894);
xnor_4 g00546(new_n2823, new_n2822, new_n2895);
xor_4  g00547(new_n2854, new_n2853_1, new_n2896);
nor_5  g00548(new_n2896, new_n2895, new_n2897);
xor_4  g00549(n15780, n1451, new_n2898);
xnor_4 g00550(n26979, n2088, new_n2899);
nor_5  g00551(new_n2899, new_n2898, new_n2900);
xor_4  g00552(new_n2896, new_n2895, new_n2901);
and_5  g00553(new_n2901, new_n2900, new_n2902);
nor_5  g00554(new_n2902, new_n2897, new_n2903);
and_5  g00555(new_n2903, new_n2894, new_n2904);
nor_5  g00556(new_n2904, new_n2893, new_n2905);
and_5  g00557(new_n2905, new_n2890, new_n2906);
nor_5  g00558(new_n2906, new_n2889, new_n2907);
nor_5  g00559(new_n2907, new_n2886_1, new_n2908);
nor_5  g00560(new_n2908, new_n2885, new_n2909);
nor_5  g00561(new_n2909, new_n2882, new_n2910);
nor_5  g00562(new_n2910, new_n2881, new_n2911);
nor_5  g00563(new_n2911, new_n2878, new_n2912);
or_5   g00564(new_n2912, new_n2877, new_n2913);
nor_5  g00565(new_n2913, new_n2874, new_n2914);
nor_5  g00566(new_n2914, new_n2873, new_n2915);
xor_4  g00567(new_n2915, new_n2870, new_n2916);
xnor_4 g00568(new_n2916, new_n2807, new_n2917);
xor_4  g00569(new_n2804, new_n2770, new_n2918);
xor_4  g00570(new_n2913, new_n2874, new_n2919);
nor_5  g00571(new_n2919, new_n2918, new_n2920);
xnor_4 g00572(new_n2919, new_n2918, new_n2921);
xnor_4 g00573(new_n2802, new_n2773, new_n2922);
xor_4  g00574(new_n2911, new_n2878, new_n2923);
and_5  g00575(new_n2923, new_n2922, new_n2924);
xnor_4 g00576(new_n2923, new_n2922, new_n2925);
xnor_4 g00577(new_n2800, new_n2776, new_n2926);
xor_4  g00578(new_n2909, new_n2882, new_n2927);
and_5  g00579(new_n2927, new_n2926, new_n2928);
xnor_4 g00580(new_n2927, new_n2926, new_n2929_1);
xnor_4 g00581(new_n2798, new_n2779_1, new_n2930);
xor_4  g00582(new_n2907, new_n2886_1, new_n2931);
and_5  g00583(new_n2931, new_n2930, new_n2932);
xnor_4 g00584(new_n2931, new_n2930, new_n2933);
xor_4  g00585(new_n2905, new_n2890, new_n2934);
not_10 g00586(new_n2934, new_n2935);
xor_4  g00587(new_n2796, new_n2782, new_n2936);
nor_5  g00588(new_n2936, new_n2935, new_n2937);
xnor_4 g00589(new_n2936, new_n2935, new_n2938);
xnor_4 g00590(new_n2903, new_n2894, new_n2939);
xnor_4 g00591(n19005, n7149, new_n2940);
xnor_4 g00592(new_n2940, new_n2794, new_n2941);
and_5  g00593(new_n2941, new_n2939, new_n2942);
xnor_4 g00594(new_n2941, new_n2939, new_n2943);
xnor_4 g00595(n5438, n1152, new_n2944_1);
xor_4  g00596(new_n2899, new_n2898, new_n2945);
or_5   g00597(new_n2945, new_n2944_1, new_n2946);
xor_4  g00598(n14148, n4326, new_n2947);
xnor_4 g00599(new_n2947, new_n2792, new_n2948_1);
and_5  g00600(new_n2948_1, new_n2946, new_n2949);
xor_4  g00601(new_n2901, new_n2900, new_n2950);
xor_4  g00602(new_n2948_1, new_n2946, new_n2951);
and_5  g00603(new_n2951, new_n2950, new_n2952);
nor_5  g00604(new_n2952, new_n2949, new_n2953);
nor_5  g00605(new_n2953, new_n2943, new_n2954);
nor_5  g00606(new_n2954, new_n2942, new_n2955);
nor_5  g00607(new_n2955, new_n2938, new_n2956);
nor_5  g00608(new_n2956, new_n2937, new_n2957);
nor_5  g00609(new_n2957, new_n2933, new_n2958);
nor_5  g00610(new_n2958, new_n2932, new_n2959);
nor_5  g00611(new_n2959, new_n2929_1, new_n2960);
nor_5  g00612(new_n2960, new_n2928, new_n2961_1);
nor_5  g00613(new_n2961_1, new_n2925, new_n2962);
nor_5  g00614(new_n2962, new_n2924, new_n2963);
nor_5  g00615(new_n2963, new_n2921, new_n2964);
nor_5  g00616(new_n2964, new_n2920, new_n2965);
xnor_4 g00617(new_n2965, new_n2917, n142);
xnor_4 g00618(n7335, n4319, new_n2967);
nor_5  g00619(n23463, n5696, new_n2968);
xnor_4 g00620(n23463, n5696, new_n2969);
nor_5  g00621(n13367, n13074, new_n2970);
xnor_4 g00622(n13367, n13074, new_n2971_1);
nor_5  g00623(n10739, n932, new_n2972);
xnor_4 g00624(n10739, n932, new_n2973);
nor_5  g00625(n21753, n6691, new_n2974);
xnor_4 g00626(n21753, n6691, new_n2975);
nor_5  g00627(n21832, n3260, new_n2976);
xnor_4 g00628(n21832, n3260, new_n2977);
nor_5  g00629(n26913, n20489, new_n2978_1);
xnor_4 g00630(n26913, n20489, new_n2979_1);
nor_5  g00631(n16223, n2355, new_n2980);
xnor_4 g00632(n16223, n2355, new_n2981);
nor_5  g00633(n19494, n11121, new_n2982);
and_5  g00634(n16217, n2387, new_n2983);
xnor_4 g00635(n19494, n11121, new_n2984);
nor_5  g00636(new_n2984, new_n2983, new_n2985_1);
nor_5  g00637(new_n2985_1, new_n2982, new_n2986);
nor_5  g00638(new_n2986, new_n2981, new_n2987);
nor_5  g00639(new_n2987, new_n2980, new_n2988);
nor_5  g00640(new_n2988, new_n2979_1, new_n2989);
nor_5  g00641(new_n2989, new_n2978_1, new_n2990);
nor_5  g00642(new_n2990, new_n2977, new_n2991);
nor_5  g00643(new_n2991, new_n2976, new_n2992);
nor_5  g00644(new_n2992, new_n2975, new_n2993);
nor_5  g00645(new_n2993, new_n2974, new_n2994);
nor_5  g00646(new_n2994, new_n2973, new_n2995);
nor_5  g00647(new_n2995, new_n2972, new_n2996);
nor_5  g00648(new_n2996, new_n2971_1, new_n2997);
nor_5  g00649(new_n2997, new_n2970, new_n2998);
nor_5  g00650(new_n2998, new_n2969, new_n2999_1);
nor_5  g00651(new_n2999_1, new_n2968, new_n3000);
xor_4  g00652(new_n3000, new_n2967, new_n3001);
nor_5  g00653(new_n3001, n5025, new_n3002);
xnor_4 g00654(new_n3001, n5025, new_n3003);
xor_4  g00655(new_n2998, new_n2969, new_n3004);
nor_5  g00656(new_n3004, n6485, new_n3005);
xnor_4 g00657(new_n3004, n6485, new_n3006);
xor_4  g00658(new_n2996, new_n2971_1, new_n3007);
nor_5  g00659(new_n3007, n26036, new_n3008);
xnor_4 g00660(new_n3007, n26036, new_n3009);
xor_4  g00661(new_n2994, new_n2973, new_n3010_1);
nor_5  g00662(new_n3010_1, n19770, new_n3011);
xnor_4 g00663(new_n3010_1, n19770, new_n3012);
xor_4  g00664(new_n2992, new_n2975, new_n3013);
nor_5  g00665(new_n3013, n8782, new_n3014);
xnor_4 g00666(new_n3013, n8782, new_n3015);
xor_4  g00667(new_n2990, new_n2977, new_n3016);
nor_5  g00668(new_n3016, n8678, new_n3017_1);
xnor_4 g00669(new_n3016, n8678, new_n3018_1);
xor_4  g00670(new_n2988, new_n2979_1, new_n3019);
nor_5  g00671(new_n3019, n1432, new_n3020_1);
xnor_4 g00672(new_n3019, n1432, new_n3021);
xor_4  g00673(new_n2986, new_n2981, new_n3022);
nor_5  g00674(new_n3022, n21599, new_n3023);
xnor_4 g00675(new_n3022, n21599, new_n3024);
not_10 g00676(n25336, new_n3025);
xnor_4 g00677(n16217, n2387, new_n3026);
nor_5  g00678(new_n3026, n11424, new_n3027);
and_5  g00679(new_n3027, new_n3025, new_n3028);
xnor_4 g00680(new_n3027, n25336, new_n3029);
xnor_4 g00681(new_n2984, new_n2983, new_n3030_1);
and_5  g00682(new_n3030_1, new_n3029, new_n3031);
nor_5  g00683(new_n3031, new_n3028, new_n3032);
nor_5  g00684(new_n3032, new_n3024, new_n3033);
nor_5  g00685(new_n3033, new_n3023, new_n3034);
nor_5  g00686(new_n3034, new_n3021, new_n3035);
nor_5  g00687(new_n3035, new_n3020_1, new_n3036);
nor_5  g00688(new_n3036, new_n3018_1, new_n3037);
nor_5  g00689(new_n3037, new_n3017_1, new_n3038);
nor_5  g00690(new_n3038, new_n3015, new_n3039);
nor_5  g00691(new_n3039, new_n3014, new_n3040);
nor_5  g00692(new_n3040, new_n3012, new_n3041);
nor_5  g00693(new_n3041, new_n3011, new_n3042);
nor_5  g00694(new_n3042, new_n3009, new_n3043);
nor_5  g00695(new_n3043, new_n3008, new_n3044);
nor_5  g00696(new_n3044, new_n3006, new_n3045);
nor_5  g00697(new_n3045, new_n3005, new_n3046);
nor_5  g00698(new_n3046, new_n3003, new_n3047);
nor_5  g00699(new_n3047, new_n3002, new_n3048);
nor_5  g00700(n7335, n4319, new_n3049);
nor_5  g00701(new_n3000, new_n2967, new_n3050);
nor_5  g00702(new_n3050, new_n3049, new_n3051);
not_10 g00703(new_n3051, new_n3052);
nand_5 g00704(new_n3052, new_n3048, new_n3053);
not_10 g00705(n9967, new_n3054);
not_10 g00706(n20946, new_n3055);
not_10 g00707(n7751, new_n3056);
not_10 g00708(n26823, new_n3057);
not_10 g00709(n4812, new_n3058);
not_10 g00710(n24278, new_n3059);
nor_5  g00711(n12315, n3952, new_n3060);
not_10 g00712(new_n3060, new_n3061);
nor_5  g00713(new_n3061, n24618, new_n3062);
and_5  g00714(new_n3062, new_n3059, new_n3063);
and_5  g00715(new_n3063, new_n3058, new_n3064);
and_5  g00716(new_n3064, new_n3057, new_n3065);
and_5  g00717(new_n3065, new_n3056, new_n3066);
and_5  g00718(new_n3066, new_n3055, new_n3067_1);
and_5  g00719(new_n3067_1, new_n3054, new_n3068);
xnor_4 g00720(new_n3068, n3425, new_n3069);
not_10 g00721(new_n3069, new_n3070);
xor_4  g00722(new_n3046, new_n3003, new_n3071);
nor_5  g00723(new_n3071, new_n3070, new_n3072);
not_10 g00724(n3425, new_n3073);
and_5  g00725(new_n3068, new_n3073, new_n3074);
xnor_4 g00726(new_n3071, new_n3070, new_n3075);
xnor_4 g00727(new_n3067_1, n9967, new_n3076_1);
xor_4  g00728(new_n3044, new_n3006, new_n3077);
not_10 g00729(new_n3077, new_n3078);
and_5  g00730(new_n3078, new_n3076_1, new_n3079);
xor_4  g00731(new_n3077, new_n3076_1, new_n3080);
xnor_4 g00732(new_n3066, n20946, new_n3081);
not_10 g00733(new_n3081, new_n3082);
xor_4  g00734(new_n3042, new_n3009, new_n3083);
nor_5  g00735(new_n3083, new_n3082, new_n3084);
xnor_4 g00736(new_n3083, new_n3082, new_n3085);
xnor_4 g00737(new_n3065, n7751, new_n3086);
not_10 g00738(new_n3086, new_n3087);
xor_4  g00739(new_n3040, new_n3012, new_n3088);
nor_5  g00740(new_n3088, new_n3087, new_n3089_1);
xnor_4 g00741(new_n3088, new_n3087, new_n3090);
xnor_4 g00742(new_n3064, n26823, new_n3091);
not_10 g00743(new_n3091, new_n3092);
xor_4  g00744(new_n3038, new_n3015, new_n3093);
nor_5  g00745(new_n3093, new_n3092, new_n3094);
xnor_4 g00746(new_n3093, new_n3092, new_n3095);
xnor_4 g00747(new_n3063, n4812, new_n3096);
xor_4  g00748(new_n3036, new_n3018_1, new_n3097);
not_10 g00749(new_n3097, new_n3098);
and_5  g00750(new_n3098, new_n3096, new_n3099);
xor_4  g00751(new_n3097, new_n3096, new_n3100);
xnor_4 g00752(new_n3062, n24278, new_n3101);
xor_4  g00753(new_n3034, new_n3021, new_n3102);
not_10 g00754(new_n3102, new_n3103);
and_5  g00755(new_n3103, new_n3101, new_n3104);
xor_4  g00756(new_n3102, new_n3101, new_n3105);
xnor_4 g00757(new_n3060, n24618, new_n3106);
xor_4  g00758(new_n3032, new_n3024, new_n3107);
not_10 g00759(new_n3107, new_n3108);
and_5  g00760(new_n3108, new_n3106, new_n3109);
xor_4  g00761(new_n3107, new_n3106, new_n3110);
not_10 g00762(n3952, new_n3111);
xor_4  g00763(new_n3026, n11424, new_n3112);
not_10 g00764(new_n3112, new_n3113);
and_5  g00765(new_n3113, n12315, new_n3114);
and_5  g00766(new_n3114, new_n3111, new_n3115);
xor_4  g00767(new_n3030_1, new_n3029, new_n3116);
not_10 g00768(new_n3116, new_n3117);
xor_4  g00769(n12315, n3952, new_n3118);
nor_5  g00770(new_n3118, new_n3114, new_n3119);
nor_5  g00771(new_n3119, new_n3115, new_n3120);
and_5  g00772(new_n3120, new_n3117, new_n3121);
nor_5  g00773(new_n3121, new_n3115, new_n3122);
nor_5  g00774(new_n3122, new_n3110, new_n3123);
nor_5  g00775(new_n3123, new_n3109, new_n3124);
nor_5  g00776(new_n3124, new_n3105, new_n3125_1);
nor_5  g00777(new_n3125_1, new_n3104, new_n3126_1);
nor_5  g00778(new_n3126_1, new_n3100, new_n3127);
nor_5  g00779(new_n3127, new_n3099, new_n3128);
nor_5  g00780(new_n3128, new_n3095, new_n3129);
nor_5  g00781(new_n3129, new_n3094, new_n3130);
nor_5  g00782(new_n3130, new_n3090, new_n3131);
nor_5  g00783(new_n3131, new_n3089_1, new_n3132);
nor_5  g00784(new_n3132, new_n3085, new_n3133);
nor_5  g00785(new_n3133, new_n3084, new_n3134);
nor_5  g00786(new_n3134, new_n3080, new_n3135);
nor_5  g00787(new_n3135, new_n3079, new_n3136_1);
nor_5  g00788(new_n3136_1, new_n3075, new_n3137);
or_5   g00789(new_n3137, new_n3074, new_n3138);
or_5   g00790(new_n3138, new_n3072, new_n3139);
or_5   g00791(new_n3139, new_n3053, new_n3140);
nor_5  g00792(n7593, n5101, new_n3141);
xnor_4 g00793(n7593, n5101, new_n3142);
nor_5  g00794(n16507, n337, new_n3143);
xnor_4 g00795(n16507, n337, new_n3144);
nor_5  g00796(n22470, n3228, new_n3145);
xnor_4 g00797(n22470, n3228, new_n3146);
nor_5  g00798(n19116, n5302, new_n3147);
xnor_4 g00799(n19116, n5302, new_n3148);
nor_5  g00800(n25738, n6861, new_n3149);
xnor_4 g00801(n25738, n6861, new_n3150);
nor_5  g00802(n21471, n19357, new_n3151);
xnor_4 g00803(n21471, n19357, new_n3152);
nor_5  g00804(n18737, n2328, new_n3153);
xnor_4 g00805(n18737, n2328, new_n3154);
nor_5  g00806(n15053, n14603, new_n3155);
xnor_4 g00807(n15053, n14603, new_n3156);
nor_5  g00808(n25471, n20794, new_n3157);
and_5  g00809(n23333, n16502, new_n3158);
xnor_4 g00810(n25471, n20794, new_n3159);
nor_5  g00811(new_n3159, new_n3158, new_n3160);
nor_5  g00812(new_n3160, new_n3157, new_n3161_1);
nor_5  g00813(new_n3161_1, new_n3156, new_n3162);
nor_5  g00814(new_n3162, new_n3155, new_n3163);
nor_5  g00815(new_n3163, new_n3154, new_n3164_1);
nor_5  g00816(new_n3164_1, new_n3153, new_n3165);
nor_5  g00817(new_n3165, new_n3152, new_n3166);
nor_5  g00818(new_n3166, new_n3151, new_n3167);
nor_5  g00819(new_n3167, new_n3150, new_n3168);
nor_5  g00820(new_n3168, new_n3149, new_n3169);
nor_5  g00821(new_n3169, new_n3148, new_n3170);
nor_5  g00822(new_n3170, new_n3147, new_n3171);
nor_5  g00823(new_n3171, new_n3146, new_n3172);
nor_5  g00824(new_n3172, new_n3145, new_n3173);
nor_5  g00825(new_n3173, new_n3144, new_n3174);
nor_5  g00826(new_n3174, new_n3143, new_n3175);
nor_5  g00827(new_n3175, new_n3142, new_n3176);
nor_5  g00828(new_n3176, new_n3141, new_n3177);
nor_5  g00829(new_n3138, new_n3072, new_n3178);
xnor_4 g00830(new_n3051, new_n3048, new_n3179);
xor_4  g00831(new_n3179, new_n3178, new_n3180);
and_5  g00832(new_n3180, new_n3177, new_n3181);
nor_5  g00833(new_n3180, new_n3177, new_n3182);
xnor_4 g00834(new_n3136_1, new_n3075, new_n3183);
xor_4  g00835(new_n3175, new_n3142, new_n3184);
and_5  g00836(new_n3184, new_n3183, new_n3185);
xnor_4 g00837(new_n3184, new_n3183, new_n3186);
xnor_4 g00838(new_n3134, new_n3080, new_n3187);
xor_4  g00839(new_n3173, new_n3144, new_n3188);
and_5  g00840(new_n3188, new_n3187, new_n3189);
xnor_4 g00841(new_n3188, new_n3187, new_n3190);
xnor_4 g00842(new_n3132, new_n3085, new_n3191);
xor_4  g00843(new_n3171, new_n3146, new_n3192);
and_5  g00844(new_n3192, new_n3191, new_n3193);
xnor_4 g00845(new_n3192, new_n3191, new_n3194);
xnor_4 g00846(new_n3130, new_n3090, new_n3195);
xor_4  g00847(new_n3169, new_n3148, new_n3196);
and_5  g00848(new_n3196, new_n3195, new_n3197);
xnor_4 g00849(new_n3196, new_n3195, new_n3198);
xnor_4 g00850(new_n3128, new_n3095, new_n3199);
xor_4  g00851(new_n3167, new_n3150, new_n3200);
and_5  g00852(new_n3200, new_n3199, new_n3201);
xnor_4 g00853(new_n3200, new_n3199, new_n3202);
xnor_4 g00854(new_n3126_1, new_n3100, new_n3203);
xor_4  g00855(new_n3165, new_n3152, new_n3204);
and_5  g00856(new_n3204, new_n3203, new_n3205);
xnor_4 g00857(new_n3204, new_n3203, new_n3206);
xnor_4 g00858(new_n3124, new_n3105, new_n3207);
xor_4  g00859(new_n3163, new_n3154, new_n3208_1);
and_5  g00860(new_n3208_1, new_n3207, new_n3209);
xnor_4 g00861(new_n3208_1, new_n3207, new_n3210);
xnor_4 g00862(new_n3122, new_n3110, new_n3211);
xor_4  g00863(new_n3161_1, new_n3156, new_n3212);
and_5  g00864(new_n3212, new_n3211, new_n3213);
xnor_4 g00865(new_n3212, new_n3211, new_n3214);
xnor_4 g00866(n23333, n16502, new_n3215);
xor_4  g00867(new_n3112, n12315, new_n3216);
nor_5  g00868(new_n3216, new_n3215, new_n3217);
xnor_4 g00869(new_n3159, new_n3158, new_n3218);
nor_5  g00870(new_n3218, new_n3217, new_n3219_1);
xnor_4 g00871(new_n3120, new_n3117, new_n3220);
xor_4  g00872(n25471, n20794, new_n3221);
and_5  g00873(new_n3217, new_n3221, new_n3222);
nor_5  g00874(new_n3222, new_n3219_1, new_n3223);
and_5  g00875(new_n3223, new_n3220, new_n3224);
nor_5  g00876(new_n3224, new_n3219_1, new_n3225);
nor_5  g00877(new_n3225, new_n3214, new_n3226);
nor_5  g00878(new_n3226, new_n3213, new_n3227);
nor_5  g00879(new_n3227, new_n3210, new_n3228_1);
nor_5  g00880(new_n3228_1, new_n3209, new_n3229);
nor_5  g00881(new_n3229, new_n3206, new_n3230);
nor_5  g00882(new_n3230, new_n3205, new_n3231);
nor_5  g00883(new_n3231, new_n3202, new_n3232);
nor_5  g00884(new_n3232, new_n3201, new_n3233);
nor_5  g00885(new_n3233, new_n3198, new_n3234);
nor_5  g00886(new_n3234, new_n3197, new_n3235_1);
nor_5  g00887(new_n3235_1, new_n3194, new_n3236);
nor_5  g00888(new_n3236, new_n3193, new_n3237);
nor_5  g00889(new_n3237, new_n3190, new_n3238);
nor_5  g00890(new_n3238, new_n3189, new_n3239);
nor_5  g00891(new_n3239, new_n3186, new_n3240);
or_5   g00892(new_n3240, new_n3185, new_n3241);
nor_5  g00893(new_n3241, new_n3182, new_n3242);
nor_5  g00894(new_n3242, new_n3181, new_n3243);
nor_5  g00895(new_n3243, new_n3140, new_n3244_1);
nor_5  g00896(new_n3178, new_n3053, new_n3245);
or_5   g00897(new_n3052, new_n3048, new_n3246);
nor_5  g00898(new_n3246, new_n3139, new_n3247);
or_5   g00899(new_n3247, new_n3245, new_n3248);
or_5   g00900(new_n3248, new_n3243, new_n3249);
and_5  g00901(new_n3249, new_n3140, new_n3250);
nor_5  g00902(new_n3250, new_n3244_1, n175);
or_5   g00903(n20138, n9251, new_n3252);
or_5   g00904(new_n3252, n6385, new_n3253_1);
or_5   g00905(new_n3253_1, n3136, new_n3254);
or_5   g00906(new_n3254, n9557, new_n3255);
or_5   g00907(new_n3255, n25643, new_n3256);
or_5   g00908(new_n3256, n9942, new_n3257);
or_5   g00909(new_n3257, n16482, new_n3258);
nor_5  g00910(new_n3258, n14130, new_n3259);
xnor_4 g00911(new_n3259, n8856, new_n3260_1);
xor_4  g00912(new_n3260_1, n25494, new_n3261);
xor_4  g00913(new_n3258, n14130, new_n3262);
nor_5  g00914(new_n3262, n10117, new_n3263_1);
xnor_4 g00915(new_n3262, n10117, new_n3264);
xor_4  g00916(new_n3257, n16482, new_n3265);
nor_5  g00917(new_n3265, n13460, new_n3266);
xnor_4 g00918(new_n3265, n13460, new_n3267);
xor_4  g00919(new_n3256, n9942, new_n3268);
nor_5  g00920(new_n3268, n6104, new_n3269);
xnor_4 g00921(new_n3268, n6104, new_n3270);
xor_4  g00922(new_n3255, n25643, new_n3271);
nor_5  g00923(new_n3271, n4119, new_n3272);
xnor_4 g00924(new_n3271, n4119, new_n3273);
xor_4  g00925(new_n3254, n9557, new_n3274);
nor_5  g00926(new_n3274, n14510, new_n3275);
xnor_4 g00927(new_n3274, n14510, new_n3276);
xor_4  g00928(new_n3253_1, n3136, new_n3277);
nor_5  g00929(new_n3277, n13263, new_n3278);
xor_4  g00930(new_n3252, n6385, new_n3279_1);
nor_5  g00931(new_n3279_1, n20455, new_n3280);
xnor_4 g00932(new_n3279_1, n20455, new_n3281);
not_10 g00933(n1639, new_n3282);
xnor_4 g00934(n20138, n9251, new_n3283);
and_5  g00935(new_n3283, new_n3282, new_n3284);
nand_5 g00936(n16968, n9251, new_n3285);
xnor_4 g00937(new_n3283, n1639, new_n3286);
and_5  g00938(new_n3286, new_n3285, new_n3287);
nor_5  g00939(new_n3287, new_n3284, new_n3288);
nor_5  g00940(new_n3288, new_n3281, new_n3289_1);
nor_5  g00941(new_n3289_1, new_n3280, new_n3290);
xnor_4 g00942(new_n3277, n13263, new_n3291);
nor_5  g00943(new_n3291, new_n3290, new_n3292);
nor_5  g00944(new_n3292, new_n3278, new_n3293);
nor_5  g00945(new_n3293, new_n3276, new_n3294);
nor_5  g00946(new_n3294, new_n3275, new_n3295);
nor_5  g00947(new_n3295, new_n3273, new_n3296);
nor_5  g00948(new_n3296, new_n3272, new_n3297);
nor_5  g00949(new_n3297, new_n3270, new_n3298);
nor_5  g00950(new_n3298, new_n3269, new_n3299);
nor_5  g00951(new_n3299, new_n3267, new_n3300);
nor_5  g00952(new_n3300, new_n3266, new_n3301_1);
nor_5  g00953(new_n3301_1, new_n3264, new_n3302);
nor_5  g00954(new_n3302, new_n3263_1, new_n3303);
xnor_4 g00955(new_n3303, new_n3261, new_n3304);
xor_4  g00956(new_n3304, n26180, new_n3305);
xnor_4 g00957(new_n3301_1, new_n3264, new_n3306_1);
nor_5  g00958(new_n3306_1, n24004, new_n3307);
xnor_4 g00959(new_n3306_1, n24004, new_n3308);
xor_4  g00960(new_n3299, new_n3267, new_n3309);
not_10 g00961(new_n3309, new_n3310);
nor_5  g00962(new_n3310, n12871, new_n3311);
xor_4  g00963(new_n3309, n12871, new_n3312);
xnor_4 g00964(new_n3297, new_n3270, new_n3313);
nor_5  g00965(new_n3313, n23304, new_n3314);
xnor_4 g00966(new_n3313, n23304, new_n3315);
xnor_4 g00967(new_n3295, new_n3273, new_n3316_1);
nor_5  g00968(new_n3316_1, n19361, new_n3317);
xnor_4 g00969(new_n3316_1, n19361, new_n3318);
xnor_4 g00970(new_n3293, new_n3276, new_n3319);
nor_5  g00971(new_n3319, n1437, new_n3320_1);
xnor_4 g00972(new_n3319, n1437, new_n3321);
xnor_4 g00973(new_n3291, new_n3290, new_n3322);
nor_5  g00974(new_n3322, n4722, new_n3323);
xor_4  g00975(new_n3322, n4722, new_n3324_1);
xnor_4 g00976(new_n3288, new_n3281, new_n3325);
and_5  g00977(new_n3325, n14633, new_n3326);
xnor_4 g00978(new_n3325, n14633, new_n3327);
not_10 g00979(n8721, new_n3328);
and_5  g00980(n16968, n9251, new_n3329);
xnor_4 g00981(new_n3286, new_n3329, new_n3330);
nor_5  g00982(new_n3330, new_n3328, new_n3331);
xor_4  g00983(n16968, n9251, new_n3332_1);
nand_5 g00984(new_n3332_1, n18578, new_n3333);
xor_4  g00985(new_n3330, n8721, new_n3334);
nor_5  g00986(new_n3334, new_n3333, new_n3335);
nor_5  g00987(new_n3335, new_n3331, new_n3336);
nor_5  g00988(new_n3336, new_n3327, new_n3337);
nor_5  g00989(new_n3337, new_n3326, new_n3338);
and_5  g00990(new_n3338, new_n3324_1, new_n3339);
nor_5  g00991(new_n3339, new_n3323, new_n3340_1);
nor_5  g00992(new_n3340_1, new_n3321, new_n3341);
nor_5  g00993(new_n3341, new_n3320_1, new_n3342);
nor_5  g00994(new_n3342, new_n3318, new_n3343_1);
nor_5  g00995(new_n3343_1, new_n3317, new_n3344);
nor_5  g00996(new_n3344, new_n3315, new_n3345);
nor_5  g00997(new_n3345, new_n3314, new_n3346);
nor_5  g00998(new_n3346, new_n3312, new_n3347);
nor_5  g00999(new_n3347, new_n3311, new_n3348);
nor_5  g01000(new_n3348, new_n3308, new_n3349_1);
nor_5  g01001(new_n3349_1, new_n3307, new_n3350);
xnor_4 g01002(new_n3350, new_n3305, new_n3351);
xor_4  g01003(n3506, n2743, new_n3352);
not_10 g01004(n7026, new_n3353);
nor_5  g01005(n14899, new_n3353, new_n3354);
xor_4  g01006(n14899, n7026, new_n3355);
not_10 g01007(n13719, new_n3356);
nor_5  g01008(n18444, new_n3356, new_n3357);
xor_4  g01009(n18444, n13719, new_n3358);
not_10 g01010(n442, new_n3359);
nor_5  g01011(n24638, new_n3359, new_n3360);
xor_4  g01012(n24638, n442, new_n3361);
not_10 g01013(n9172, new_n3362);
nor_5  g01014(n21674, new_n3362, new_n3363);
xor_4  g01015(n21674, n9172, new_n3364);
not_10 g01016(n4913, new_n3365);
or_5   g01017(n17251, new_n3365, new_n3366_1);
xor_4  g01018(n17251, n4913, new_n3367);
not_10 g01019(n604, new_n3368);
or_5   g01020(n14790, new_n3368, new_n3369);
xor_4  g01021(n14790, n604, new_n3370);
not_10 g01022(n16824, new_n3371);
and_5  g01023(new_n3371, n10096, new_n3372);
nor_5  g01024(new_n3371, n10096, new_n3373);
not_10 g01025(n16521, new_n3374);
and_5  g01026(n16994, new_n3374, new_n3375);
or_5   g01027(n16994, new_n3374, new_n3376);
not_10 g01028(n9246, new_n3377);
nor_5  g01029(new_n3377, n7139, new_n3378);
and_5  g01030(new_n3378, new_n3376, new_n3379);
nor_5  g01031(new_n3379, new_n3375, new_n3380);
nor_5  g01032(new_n3380, new_n3373, new_n3381);
nor_5  g01033(new_n3381, new_n3372, new_n3382);
not_10 g01034(new_n3382, new_n3383);
or_5   g01035(new_n3383, new_n3370, new_n3384);
and_5  g01036(new_n3384, new_n3369, new_n3385);
or_5   g01037(new_n3385, new_n3367, new_n3386);
and_5  g01038(new_n3386, new_n3366_1, new_n3387);
nor_5  g01039(new_n3387, new_n3364, new_n3388);
nor_5  g01040(new_n3388, new_n3363, new_n3389);
nor_5  g01041(new_n3389, new_n3361, new_n3390_1);
nor_5  g01042(new_n3390_1, new_n3360, new_n3391);
nor_5  g01043(new_n3391, new_n3358, new_n3392);
nor_5  g01044(new_n3392, new_n3357, new_n3393);
nor_5  g01045(new_n3393, new_n3355, new_n3394);
nor_5  g01046(new_n3394, new_n3354, new_n3395);
xor_4  g01047(new_n3395, new_n3352, new_n3396);
or_5   g01048(n25565, n21993, new_n3397);
or_5   g01049(new_n3397, n11273, new_n3398);
or_5   g01050(new_n3398, n22290, new_n3399);
or_5   g01051(new_n3399, n9598, new_n3400);
or_5   g01052(new_n3400, n7670, new_n3401);
or_5   g01053(new_n3401, n13912, new_n3402);
nor_5  g01054(new_n3402, n20213, new_n3403);
not_10 g01055(new_n3403, new_n3404);
nor_5  g01056(new_n3404, n21489, new_n3405);
xnor_4 g01057(new_n3405, n9259, new_n3406);
xnor_4 g01058(new_n3406, new_n3396, new_n3407);
xor_4  g01059(new_n3393, new_n3355, new_n3408);
xnor_4 g01060(new_n3403, n21489, new_n3409);
and_5  g01061(new_n3409, new_n3408, new_n3410);
xnor_4 g01062(new_n3409, new_n3408, new_n3411);
xor_4  g01063(new_n3391, new_n3358, new_n3412);
xor_4  g01064(new_n3402, n20213, new_n3413);
nor_5  g01065(new_n3413, new_n3412, new_n3414);
xnor_4 g01066(new_n3413, new_n3412, new_n3415);
xor_4  g01067(new_n3389, new_n3361, new_n3416);
xor_4  g01068(new_n3401, n13912, new_n3417);
nor_5  g01069(new_n3417, new_n3416, new_n3418);
xnor_4 g01070(new_n3417, new_n3416, new_n3419);
xor_4  g01071(new_n3387, new_n3364, new_n3420);
xor_4  g01072(new_n3400, n7670, new_n3421);
nor_5  g01073(new_n3421, new_n3420, new_n3422);
xnor_4 g01074(new_n3421, new_n3420, new_n3423);
xor_4  g01075(new_n3399, n9598, new_n3424);
xor_4  g01076(new_n3385, new_n3367, new_n3425_1);
nor_5  g01077(new_n3425_1, new_n3424, new_n3426_1);
xnor_4 g01078(new_n3425_1, new_n3424, new_n3427);
xor_4  g01079(new_n3398, n22290, new_n3428);
xnor_4 g01080(new_n3382, new_n3370, new_n3429);
nor_5  g01081(new_n3429, new_n3428, new_n3430);
xnor_4 g01082(new_n3397, n11273, new_n3431);
xnor_4 g01083(n16824, n10096, new_n3432);
xnor_4 g01084(new_n3432, new_n3380, new_n3433);
and_5  g01085(new_n3433, new_n3431, new_n3434);
xnor_4 g01086(new_n3433, new_n3431, new_n3435);
xor_4  g01087(n25565, n21993, new_n3436);
not_10 g01088(new_n3436, new_n3437);
xor_4  g01089(n16994, n16521, new_n3438);
xnor_4 g01090(new_n3438, new_n3378, new_n3439);
and_5  g01091(new_n3439, new_n3437, new_n3440);
not_10 g01092(n21993, new_n3441);
xnor_4 g01093(n9246, n7139, new_n3442);
or_5   g01094(new_n3442, new_n3441, new_n3443);
xnor_4 g01095(new_n3439, new_n3436, new_n3444);
and_5  g01096(new_n3444, new_n3443, new_n3445);
nor_5  g01097(new_n3445, new_n3440, new_n3446);
nor_5  g01098(new_n3446, new_n3435, new_n3447);
nor_5  g01099(new_n3447, new_n3434, new_n3448);
xnor_4 g01100(new_n3429, new_n3428, new_n3449);
nor_5  g01101(new_n3449, new_n3448, new_n3450);
nor_5  g01102(new_n3450, new_n3430, new_n3451_1);
nor_5  g01103(new_n3451_1, new_n3427, new_n3452);
nor_5  g01104(new_n3452, new_n3426_1, new_n3453);
nor_5  g01105(new_n3453, new_n3423, new_n3454);
nor_5  g01106(new_n3454, new_n3422, new_n3455);
nor_5  g01107(new_n3455, new_n3419, new_n3456);
nor_5  g01108(new_n3456, new_n3418, new_n3457);
nor_5  g01109(new_n3457, new_n3415, new_n3458);
or_5   g01110(new_n3458, new_n3414, new_n3459_1);
nor_5  g01111(new_n3459_1, new_n3411, new_n3460_1);
nor_5  g01112(new_n3460_1, new_n3410, new_n3461);
xor_4  g01113(new_n3461, new_n3407, new_n3462);
xnor_4 g01114(new_n3462, new_n3351, new_n3463);
xnor_4 g01115(new_n3348, new_n3308, new_n3464);
xor_4  g01116(new_n3459_1, new_n3411, new_n3465);
nor_5  g01117(new_n3465, new_n3464, new_n3466);
xnor_4 g01118(new_n3465, new_n3464, new_n3467);
xor_4  g01119(new_n3346, new_n3312, new_n3468_1);
xor_4  g01120(new_n3457, new_n3415, new_n3469);
and_5  g01121(new_n3469, new_n3468_1, new_n3470);
xnor_4 g01122(new_n3469, new_n3468_1, new_n3471);
xor_4  g01123(new_n3344, new_n3315, new_n3472);
xor_4  g01124(new_n3455, new_n3419, new_n3473);
and_5  g01125(new_n3473, new_n3472, new_n3474);
xnor_4 g01126(new_n3473, new_n3472, new_n3475);
xor_4  g01127(new_n3342, new_n3318, new_n3476);
xor_4  g01128(new_n3453, new_n3423, new_n3477);
and_5  g01129(new_n3477, new_n3476, new_n3478);
xnor_4 g01130(new_n3477, new_n3476, new_n3479);
xor_4  g01131(new_n3340_1, new_n3321, new_n3480_1);
xor_4  g01132(new_n3451_1, new_n3427, new_n3481);
and_5  g01133(new_n3481, new_n3480_1, new_n3482);
xnor_4 g01134(new_n3481, new_n3480_1, new_n3483);
xnor_4 g01135(new_n3322, n4722, new_n3484);
xnor_4 g01136(new_n3338, new_n3484, new_n3485);
xor_4  g01137(new_n3449, new_n3448, new_n3486);
and_5  g01138(new_n3486, new_n3485, new_n3487);
xnor_4 g01139(new_n3486, new_n3485, new_n3488);
xor_4  g01140(new_n3336, new_n3327, new_n3489);
not_10 g01141(new_n3489, new_n3490);
xor_4  g01142(new_n3446, new_n3435, new_n3491);
and_5  g01143(new_n3491, new_n3490, new_n3492);
xor_4  g01144(new_n3491, new_n3489, new_n3493);
xnor_4 g01145(new_n3444, new_n3443, new_n3494);
xor_4  g01146(new_n3334, new_n3333, new_n3495);
nor_5  g01147(new_n3495, new_n3494, new_n3496);
xnor_4 g01148(new_n3332_1, n18578, new_n3497);
xor_4  g01149(new_n3442, n21993, new_n3498);
or_5   g01150(new_n3498, new_n3497, new_n3499);
xor_4  g01151(new_n3495, new_n3494, new_n3500);
and_5  g01152(new_n3500, new_n3499, new_n3501);
nor_5  g01153(new_n3501, new_n3496, new_n3502_1);
nor_5  g01154(new_n3502_1, new_n3493, new_n3503);
nor_5  g01155(new_n3503, new_n3492, new_n3504);
nor_5  g01156(new_n3504, new_n3488, new_n3505);
nor_5  g01157(new_n3505, new_n3487, new_n3506_1);
nor_5  g01158(new_n3506_1, new_n3483, new_n3507);
nor_5  g01159(new_n3507, new_n3482, new_n3508);
nor_5  g01160(new_n3508, new_n3479, new_n3509);
nor_5  g01161(new_n3509, new_n3478, new_n3510);
nor_5  g01162(new_n3510, new_n3475, new_n3511);
nor_5  g01163(new_n3511, new_n3474, new_n3512);
nor_5  g01164(new_n3512, new_n3471, new_n3513);
nor_5  g01165(new_n3513, new_n3470, new_n3514);
nor_5  g01166(new_n3514, new_n3467, new_n3515);
nor_5  g01167(new_n3515, new_n3466, new_n3516_1);
xnor_4 g01168(new_n3516_1, new_n3463, n235);
or_5   g01169(n25435, n13319, new_n3518);
or_5   g01170(new_n3518, n15967, new_n3519);
or_5   g01171(new_n3519, n25797, new_n3520);
or_5   g01172(new_n3520, n6369, new_n3521);
or_5   g01173(new_n3521, n21134, new_n3522);
xor_4  g01174(new_n3522, n2113, new_n3523);
xnor_4 g01175(new_n3523, n19327, new_n3524);
xor_4  g01176(new_n3521, n21134, new_n3525);
nor_5  g01177(new_n3525, n22597, new_n3526);
xnor_4 g01178(new_n3525, n22597, new_n3527);
xor_4  g01179(new_n3520, n6369, new_n3528_1);
nor_5  g01180(new_n3528_1, n26107, new_n3529);
xnor_4 g01181(new_n3528_1, n26107, new_n3530);
xor_4  g01182(new_n3519, n25797, new_n3531);
nor_5  g01183(new_n3531, n342, new_n3532);
xor_4  g01184(new_n3518, n15967, new_n3533);
nor_5  g01185(new_n3533, n26553, new_n3534);
xnor_4 g01186(new_n3533, n26553, new_n3535);
xor_4  g01187(n25435, n13319, new_n3536);
nor_5  g01188(new_n3536, n4964, new_n3537);
nand_5 g01189(n25435, n7876, new_n3538);
xor_4  g01190(new_n3536, n4964, new_n3539);
and_5  g01191(new_n3539, new_n3538, new_n3540);
nor_5  g01192(new_n3540, new_n3537, new_n3541_1);
nor_5  g01193(new_n3541_1, new_n3535, new_n3542);
nor_5  g01194(new_n3542, new_n3534, new_n3543);
xnor_4 g01195(new_n3531, n342, new_n3544);
nor_5  g01196(new_n3544, new_n3543, new_n3545);
nor_5  g01197(new_n3545, new_n3532, new_n3546);
nor_5  g01198(new_n3546, new_n3530, new_n3547);
nor_5  g01199(new_n3547, new_n3529, new_n3548);
nor_5  g01200(new_n3548, new_n3527, new_n3549);
nor_5  g01201(new_n3549, new_n3526, new_n3550);
xnor_4 g01202(new_n3550, new_n3524, new_n3551);
xnor_4 g01203(new_n3551, n25749, new_n3552);
not_10 g01204(n3161, new_n3553);
xor_4  g01205(new_n3548, new_n3527, new_n3554);
nor_5  g01206(new_n3554, new_n3553, new_n3555_1);
xor_4  g01207(new_n3554, n3161, new_n3556);
xnor_4 g01208(new_n3546, new_n3530, new_n3557);
and_5  g01209(new_n3557, n9003, new_n3558);
xnor_4 g01210(new_n3557, n9003, new_n3559);
not_10 g01211(n4957, new_n3560);
xor_4  g01212(new_n3544, new_n3543, new_n3561_1);
nor_5  g01213(new_n3561_1, new_n3560, new_n3562);
xor_4  g01214(new_n3561_1, n4957, new_n3563_1);
xnor_4 g01215(new_n3541_1, new_n3535, new_n3564);
and_5  g01216(new_n3564, n7524, new_n3565);
xnor_4 g01217(new_n3564, n7524, new_n3566);
not_10 g01218(n15743, new_n3567);
xor_4  g01219(new_n3539, new_n3538, new_n3568);
nor_5  g01220(new_n3568, new_n3567, new_n3569);
xor_4  g01221(n25435, n7876, new_n3570_1);
nand_5 g01222(new_n3570_1, n20658, new_n3571);
xor_4  g01223(new_n3568, n15743, new_n3572);
nor_5  g01224(new_n3572, new_n3571, new_n3573);
nor_5  g01225(new_n3573, new_n3569, new_n3574);
nor_5  g01226(new_n3574, new_n3566, new_n3575);
nor_5  g01227(new_n3575, new_n3565, new_n3576);
nor_5  g01228(new_n3576, new_n3563_1, new_n3577);
nor_5  g01229(new_n3577, new_n3562, new_n3578);
nor_5  g01230(new_n3578, new_n3559, new_n3579);
nor_5  g01231(new_n3579, new_n3558, new_n3580);
nor_5  g01232(new_n3580, new_n3556, new_n3581);
nor_5  g01233(new_n3581, new_n3555_1, new_n3582_1);
xnor_4 g01234(new_n3582_1, new_n3552, new_n3583);
xor_4  g01235(n26510, n22332, new_n3584);
not_10 g01236(n18907, new_n3585);
nor_5  g01237(n23068, new_n3585, new_n3586);
xor_4  g01238(n23068, n18907, new_n3587);
not_10 g01239(n2731, new_n3588);
nor_5  g01240(n19514, new_n3588, new_n3589);
xor_4  g01241(n19514, n2731, new_n3590);
not_10 g01242(n19911, new_n3591);
nor_5  g01243(new_n3591, n10053, new_n3592);
xor_4  g01244(n19911, n10053, new_n3593);
not_10 g01245(n8399, new_n3594);
nor_5  g01246(n13708, new_n3594, new_n3595);
not_10 g01247(n13708, new_n3596);
nor_5  g01248(new_n3596, n8399, new_n3597);
not_10 g01249(n9507, new_n3598);
nor_5  g01250(n18409, new_n3598, new_n3599);
not_10 g01251(n18409, new_n3600);
or_5   g01252(new_n3600, n9507, new_n3601);
not_10 g01253(n26979, new_n3602);
nor_5  g01254(new_n3602, n5704, new_n3603);
and_5  g01255(new_n3603, new_n3601, new_n3604);
nor_5  g01256(new_n3604, new_n3599, new_n3605);
nor_5  g01257(new_n3605, new_n3597, new_n3606);
or_5   g01258(new_n3606, new_n3595, new_n3607);
nor_5  g01259(new_n3607, new_n3593, new_n3608);
nor_5  g01260(new_n3608, new_n3592, new_n3609);
nor_5  g01261(new_n3609, new_n3590, new_n3610);
nor_5  g01262(new_n3610, new_n3589, new_n3611);
nor_5  g01263(new_n3611, new_n3587, new_n3612);
nor_5  g01264(new_n3612, new_n3586, new_n3613);
xor_4  g01265(new_n3613, new_n3584, new_n3614);
nor_5  g01266(n22043, n12121, new_n3615);
not_10 g01267(new_n3615, new_n3616);
or_5   g01268(new_n3616, n19618, new_n3617_1);
or_5   g01269(new_n3617_1, n1204, new_n3618_1);
or_5   g01270(new_n3618_1, n626, new_n3619);
or_5   g01271(new_n3619, n5337, new_n3620);
xor_4  g01272(new_n3620, n4325, new_n3621);
xnor_4 g01273(new_n3621, new_n3614, new_n3622);
xor_4  g01274(new_n3611, new_n3587, new_n3623);
xor_4  g01275(new_n3619, n5337, new_n3624);
nor_5  g01276(new_n3624, new_n3623, new_n3625);
xnor_4 g01277(new_n3624, new_n3623, new_n3626);
xor_4  g01278(new_n3609, new_n3590, new_n3627);
xor_4  g01279(new_n3618_1, n626, new_n3628);
nor_5  g01280(new_n3628, new_n3627, new_n3629);
xnor_4 g01281(new_n3628, new_n3627, new_n3630);
xor_4  g01282(new_n3617_1, n1204, new_n3631);
xor_4  g01283(new_n3607, new_n3593, new_n3632);
nor_5  g01284(new_n3632, new_n3631, new_n3633);
xnor_4 g01285(new_n3632, new_n3631, new_n3634);
xor_4  g01286(new_n3615, n19618, new_n3635);
xnor_4 g01287(n13708, n8399, new_n3636);
xnor_4 g01288(new_n3636, new_n3605, new_n3637);
and_5  g01289(new_n3637, new_n3635, new_n3638);
xnor_4 g01290(new_n3637, new_n3635, new_n3639);
xnor_4 g01291(n22043, n12121, new_n3640);
xor_4  g01292(n18409, n9507, new_n3641);
xnor_4 g01293(new_n3641, new_n3603, new_n3642_1);
nor_5  g01294(new_n3642_1, new_n3640, new_n3643);
xor_4  g01295(n26979, n5704, new_n3644);
and_5  g01296(new_n3644, n12121, new_n3645);
xor_4  g01297(new_n3642_1, new_n3640, new_n3646);
and_5  g01298(new_n3646, new_n3645, new_n3647);
or_5   g01299(new_n3647, new_n3643, new_n3648);
nor_5  g01300(new_n3648, new_n3639, new_n3649_1);
nor_5  g01301(new_n3649_1, new_n3638, new_n3650);
nor_5  g01302(new_n3650, new_n3634, new_n3651);
nor_5  g01303(new_n3651, new_n3633, new_n3652);
nor_5  g01304(new_n3652, new_n3630, new_n3653);
nor_5  g01305(new_n3653, new_n3629, new_n3654);
nor_5  g01306(new_n3654, new_n3626, new_n3655);
nor_5  g01307(new_n3655, new_n3625, new_n3656);
xor_4  g01308(new_n3656, new_n3622, new_n3657);
xnor_4 g01309(new_n3657, new_n3583, new_n3658);
xor_4  g01310(new_n3654, new_n3626, new_n3659);
not_10 g01311(new_n3659, new_n3660);
xor_4  g01312(new_n3580, new_n3556, new_n3661);
nor_5  g01313(new_n3661, new_n3660, new_n3662);
xor_4  g01314(new_n3661, new_n3659, new_n3663);
xor_4  g01315(new_n3652, new_n3630, new_n3664);
not_10 g01316(new_n3664, new_n3665_1);
xor_4  g01317(new_n3578, new_n3559, new_n3666);
nor_5  g01318(new_n3666, new_n3665_1, new_n3667);
xor_4  g01319(new_n3666, new_n3664, new_n3668);
xor_4  g01320(new_n3650, new_n3634, new_n3669);
not_10 g01321(new_n3669, new_n3670);
xor_4  g01322(new_n3576, new_n3563_1, new_n3671);
nor_5  g01323(new_n3671, new_n3670, new_n3672);
xor_4  g01324(new_n3671, new_n3669, new_n3673);
xnor_4 g01325(new_n3648, new_n3639, new_n3674);
xor_4  g01326(new_n3574, new_n3566, new_n3675);
nor_5  g01327(new_n3675, new_n3674, new_n3676);
xnor_4 g01328(new_n3675, new_n3674, new_n3677);
xor_4  g01329(new_n3646, new_n3645, new_n3678);
xor_4  g01330(new_n3572, new_n3571, new_n3679_1);
nor_5  g01331(new_n3679_1, new_n3678, new_n3680);
xnor_4 g01332(new_n3570_1, n20658, new_n3681);
xnor_4 g01333(n26979, n5704, new_n3682);
xor_4  g01334(new_n3682, n12121, new_n3683);
or_5   g01335(new_n3683, new_n3681, new_n3684);
xor_4  g01336(new_n3679_1, new_n3678, new_n3685);
and_5  g01337(new_n3685, new_n3684, new_n3686);
nor_5  g01338(new_n3686, new_n3680, new_n3687);
nor_5  g01339(new_n3687, new_n3677, new_n3688);
nor_5  g01340(new_n3688, new_n3676, new_n3689);
nor_5  g01341(new_n3689, new_n3673, new_n3690);
nor_5  g01342(new_n3690, new_n3672, new_n3691);
nor_5  g01343(new_n3691, new_n3668, new_n3692);
nor_5  g01344(new_n3692, new_n3667, new_n3693);
nor_5  g01345(new_n3693, new_n3663, new_n3694);
nor_5  g01346(new_n3694, new_n3662, new_n3695);
xnor_4 g01347(new_n3695, new_n3658, n242);
or_5   g01348(n21398, n11667, new_n3697);
or_5   g01349(new_n3697, n26572, new_n3698);
or_5   g01350(new_n3698, n5115, new_n3699);
or_5   g01351(new_n3699, n11223, new_n3700);
xor_4  g01352(new_n3700, n19477, new_n3701);
xnor_4 g01353(new_n3701, n11011, new_n3702);
xor_4  g01354(new_n3699, n11223, new_n3703);
nor_5  g01355(new_n3703, n16029, new_n3704);
xnor_4 g01356(new_n3703, n16029, new_n3705);
xor_4  g01357(new_n3698, n5115, new_n3706);
and_5  g01358(new_n3706, n16476, new_n3707);
xnor_4 g01359(new_n3706, n16476, new_n3708);
xor_4  g01360(new_n3697, n26572, new_n3709);
nor_5  g01361(new_n3709, n11615, new_n3710_1);
xnor_4 g01362(new_n3709, n11615, new_n3711);
not_10 g01363(n22433, new_n3712);
xnor_4 g01364(n21398, n11667, new_n3713);
and_5  g01365(new_n3713, new_n3712, new_n3714);
nand_5 g01366(n21398, n14090, new_n3715);
xnor_4 g01367(new_n3713, n22433, new_n3716);
and_5  g01368(new_n3716, new_n3715, new_n3717);
nor_5  g01369(new_n3717, new_n3714, new_n3718);
nor_5  g01370(new_n3718, new_n3711, new_n3719);
or_5   g01371(new_n3719, new_n3710_1, new_n3720);
nor_5  g01372(new_n3720, new_n3708, new_n3721);
or_5   g01373(new_n3721, new_n3707, new_n3722);
nor_5  g01374(new_n3722, new_n3705, new_n3723);
nor_5  g01375(new_n3723, new_n3704, new_n3724);
xnor_4 g01376(new_n3724, new_n3702, new_n3725_1);
xnor_4 g01377(new_n3725_1, n13677, new_n3726);
xnor_4 g01378(new_n3722, new_n3705, new_n3727);
nor_5  g01379(new_n3727, n18926, new_n3728);
xor_4  g01380(new_n3720, new_n3708, new_n3729);
and_5  g01381(new_n3729, n5451, new_n3730);
xnor_4 g01382(new_n3729, n5451, new_n3731);
not_10 g01383(n5330, new_n3732);
xor_4  g01384(new_n3718, new_n3711, new_n3733_1);
nor_5  g01385(new_n3733_1, new_n3732, new_n3734);
xnor_4 g01386(new_n3733_1, new_n3732, new_n3735);
and_5  g01387(n21398, n14090, new_n3736);
xnor_4 g01388(new_n3716, new_n3736, new_n3737);
not_10 g01389(new_n3737, new_n3738);
and_5  g01390(new_n3738, n7657, new_n3739);
nand_5 g01391(new_n2530, n25926, new_n3740_1);
xor_4  g01392(new_n3737, n7657, new_n3741);
nor_5  g01393(new_n3741, new_n3740_1, new_n3742);
nor_5  g01394(new_n3742, new_n3739, new_n3743);
nor_5  g01395(new_n3743, new_n3735, new_n3744);
nor_5  g01396(new_n3744, new_n3734, new_n3745);
nor_5  g01397(new_n3745, new_n3731, new_n3746);
or_5   g01398(new_n3746, new_n3730, new_n3747);
xnor_4 g01399(new_n3727, n18926, new_n3748);
nor_5  g01400(new_n3748, new_n3747, new_n3749);
nor_5  g01401(new_n3749, new_n3728, new_n3750);
xnor_4 g01402(new_n3750, new_n3726, new_n3751);
not_10 g01403(n19789, new_n3752);
not_10 g01404(n8285, new_n3753);
nor_5  g01405(n21687, n6729, new_n3754);
nand_5 g01406(new_n3754, new_n3753, new_n3755_1);
nor_5  g01407(new_n3755_1, n20169, new_n3756);
and_5  g01408(new_n3756, new_n3752, new_n3757);
xnor_4 g01409(new_n3757, n12398, new_n3758_1);
or_5   g01410(n19922, n10792, new_n3759);
or_5   g01411(new_n3759, n9323, new_n3760_1);
or_5   g01412(new_n3760_1, n1949, new_n3761);
or_5   g01413(new_n3761, n15424, new_n3762);
xor_4  g01414(new_n3762, n25694, new_n3763);
xnor_4 g01415(new_n3763, n20151, new_n3764);
xor_4  g01416(new_n3761, n15424, new_n3765);
and_5  g01417(new_n3765, n7693, new_n3766);
xor_4  g01418(new_n3760_1, n1949, new_n3767);
and_5  g01419(new_n3767, n10405, new_n3768);
xnor_4 g01420(new_n3767, n10405, new_n3769);
xor_4  g01421(new_n3759, n9323, new_n3770);
nor_5  g01422(new_n3770, n11302, new_n3771);
xnor_4 g01423(new_n3770, n11302, new_n3772);
xor_4  g01424(n19922, n10792, new_n3773);
nor_5  g01425(new_n3773, n17090, new_n3774);
and_5  g01426(n19922, n6773, new_n3775);
xnor_4 g01427(new_n3773, n17090, new_n3776);
nor_5  g01428(new_n3776, new_n3775, new_n3777);
nor_5  g01429(new_n3777, new_n3774, new_n3778);
nor_5  g01430(new_n3778, new_n3772, new_n3779);
or_5   g01431(new_n3779, new_n3771, new_n3780);
nor_5  g01432(new_n3780, new_n3769, new_n3781_1);
nor_5  g01433(new_n3781_1, new_n3768, new_n3782);
xnor_4 g01434(new_n3765, n7693, new_n3783);
nor_5  g01435(new_n3783, new_n3782, new_n3784);
nor_5  g01436(new_n3784, new_n3766, new_n3785_1);
xor_4  g01437(new_n3785_1, new_n3764, new_n3786);
xnor_4 g01438(new_n3786, new_n3758_1, new_n3787);
xnor_4 g01439(new_n3756, n19789, new_n3788);
xor_4  g01440(new_n3783, new_n3782, new_n3789);
nand_5 g01441(new_n3789, new_n3788, new_n3790);
xnor_4 g01442(new_n3789, new_n3788, new_n3791);
xor_4  g01443(new_n3780, new_n3769, new_n3792);
xor_4  g01444(new_n3755_1, n20169, new_n3793);
nor_5  g01445(new_n3793, new_n3792, new_n3794_1);
xor_4  g01446(new_n3793, new_n3792, new_n3795_1);
xor_4  g01447(new_n3778, new_n3772, new_n3796);
xor_4  g01448(new_n3754, n8285, new_n3797);
nor_5  g01449(new_n3797, new_n3796, new_n3798);
xnor_4 g01450(new_n3797, new_n3796, new_n3799);
xnor_4 g01451(n21687, n6729, new_n3800);
xor_4  g01452(new_n3776, new_n3775, new_n3801);
nor_5  g01453(new_n3801, new_n3800, new_n3802);
nand_5 g01454(new_n2528, n21687, new_n3803);
xnor_4 g01455(new_n3801, new_n3800, new_n3804);
nor_5  g01456(new_n3804, new_n3803, new_n3805);
nor_5  g01457(new_n3805, new_n3802, new_n3806);
nor_5  g01458(new_n3806, new_n3799, new_n3807);
nor_5  g01459(new_n3807, new_n3798, new_n3808);
and_5  g01460(new_n3808, new_n3795_1, new_n3809);
nor_5  g01461(new_n3809, new_n3794_1, new_n3810);
not_10 g01462(new_n3810, new_n3811);
or_5   g01463(new_n3811, new_n3791, new_n3812);
and_5  g01464(new_n3812, new_n3790, new_n3813);
xor_4  g01465(new_n3813, new_n3787, new_n3814);
xnor_4 g01466(new_n3814, new_n3751, new_n3815);
xor_4  g01467(new_n3810, new_n3791, new_n3816);
xor_4  g01468(new_n3748, new_n3747, new_n3817);
and_5  g01469(new_n3817, new_n3816, new_n3818);
xnor_4 g01470(new_n3817, new_n3816, new_n3819);
xnor_4 g01471(new_n3808, new_n3795_1, new_n3820);
xor_4  g01472(new_n3745, new_n3731, new_n3821);
nor_5  g01473(new_n3821, new_n3820, new_n3822);
xnor_4 g01474(new_n3821, new_n3820, new_n3823);
xor_4  g01475(new_n3743, new_n3735, new_n3824);
xor_4  g01476(new_n3806, new_n3799, new_n3825);
nor_5  g01477(new_n3825, new_n3824, new_n3826);
xnor_4 g01478(new_n3825, new_n3824, new_n3827);
xor_4  g01479(new_n3804, new_n3803, new_n3828_1);
xor_4  g01480(new_n3741, new_n3740_1, new_n3829);
nor_5  g01481(new_n3829, new_n3828_1, new_n3830);
or_5   g01482(new_n2531, new_n2529, new_n3831);
xor_4  g01483(new_n3829, new_n3828_1, new_n3832);
and_5  g01484(new_n3832, new_n3831, new_n3833);
nor_5  g01485(new_n3833, new_n3830, new_n3834);
nor_5  g01486(new_n3834, new_n3827, new_n3835);
nor_5  g01487(new_n3835, new_n3826, new_n3836);
nor_5  g01488(new_n3836, new_n3823, new_n3837);
nor_5  g01489(new_n3837, new_n3822, new_n3838);
nor_5  g01490(new_n3838, new_n3819, new_n3839);
nor_5  g01491(new_n3839, new_n3818, new_n3840);
xnor_4 g01492(new_n3840, new_n3815, n243);
xnor_4 g01493(n24786, n11302, new_n3842_1);
nor_5  g01494(n27120, n17090, new_n3843);
and_5  g01495(n23065, n6773, new_n3844);
xnor_4 g01496(n27120, n17090, new_n3845);
nor_5  g01497(new_n3845, new_n3844, new_n3846);
nor_5  g01498(new_n3846, new_n3843, new_n3847);
xor_4  g01499(new_n3847, new_n3842_1, new_n3848);
not_10 g01500(new_n3848, new_n3849);
xor_4  g01501(n20036, n1689, new_n3850_1);
not_10 g01502(n11192, new_n3851);
and_5  g01503(n22274, new_n3851, new_n3852);
or_5   g01504(n22274, new_n3851, new_n3853);
not_10 g01505(n9380, new_n3854);
and_5  g01506(n24129, new_n3854, new_n3855);
and_5  g01507(new_n3855, new_n3853, new_n3856);
nor_5  g01508(new_n3856, new_n3852, new_n3857);
xor_4  g01509(new_n3857, new_n3850_1, new_n3858);
xnor_4 g01510(new_n3858, new_n3849, new_n3859);
xor_4  g01511(new_n3845, new_n3844, new_n3860);
xor_4  g01512(n22274, n11192, new_n3861);
xnor_4 g01513(new_n3861, new_n3855, new_n3862);
nor_5  g01514(new_n3862, new_n3860, new_n3863);
xor_4  g01515(n23065, n6773, new_n3864);
not_10 g01516(new_n3864, new_n3865);
xnor_4 g01517(n24129, n9380, new_n3866);
or_5   g01518(new_n3866, new_n3865, new_n3867);
xnor_4 g01519(new_n3862, new_n3860, new_n3868);
nor_5  g01520(new_n3868, new_n3867, new_n3869_1);
nor_5  g01521(new_n3869_1, new_n3863, new_n3870);
xnor_4 g01522(new_n3870, new_n3859, new_n3871_1);
xnor_4 g01523(n5330, n919, new_n3872);
nor_5  g01524(n25316, n7657, new_n3873);
and_5  g01525(n25926, n20385, new_n3874);
xnor_4 g01526(n25316, n7657, new_n3875);
nor_5  g01527(new_n3875, new_n3874, new_n3876);
nor_5  g01528(new_n3876, new_n3873, new_n3877);
xor_4  g01529(new_n3877, new_n3872, new_n3878);
xnor_4 g01530(new_n3878, new_n3871_1, new_n3879);
xor_4  g01531(new_n3868, new_n3867, new_n3880);
xor_4  g01532(new_n3875, new_n3874, new_n3881);
nor_5  g01533(new_n3881, new_n3880, new_n3882);
xnor_4 g01534(n25926, n20385, new_n3883);
xnor_4 g01535(new_n3866, new_n3864, new_n3884);
nor_5  g01536(new_n3884, new_n3883, new_n3885);
xor_4  g01537(new_n3881, new_n3880, new_n3886);
and_5  g01538(new_n3886, new_n3885, new_n3887);
nor_5  g01539(new_n3887, new_n3882, new_n3888);
xnor_4 g01540(new_n3888, new_n3879, n248);
or_5   g01541(n24732, n6631, new_n3890);
or_5   g01542(new_n3890, n14684, new_n3891_1);
or_5   g01543(new_n3891_1, n17035, new_n3892);
xor_4  g01544(new_n3892, n19905, new_n3893);
xor_4  g01545(new_n3893, n6369, new_n3894);
xor_4  g01546(new_n3891_1, n17035, new_n3895);
and_5  g01547(new_n3895, n25797, new_n3896);
xor_4  g01548(new_n3895, n25797, new_n3897);
xor_4  g01549(new_n3890, n14684, new_n3898);
nor_5  g01550(new_n3898, n15967, new_n3899);
xnor_4 g01551(new_n3898, n15967, new_n3900);
not_10 g01552(n13319, new_n3901);
xnor_4 g01553(n24732, n6631, new_n3902);
and_5  g01554(new_n3902, new_n3901, new_n3903);
nand_5 g01555(n25435, n24732, new_n3904);
xnor_4 g01556(new_n3902, n13319, new_n3905);
and_5  g01557(new_n3905, new_n3904, new_n3906);
nor_5  g01558(new_n3906, new_n3903, new_n3907);
nor_5  g01559(new_n3907, new_n3900, new_n3908);
nor_5  g01560(new_n3908, new_n3899, new_n3909_1);
and_5  g01561(new_n3909_1, new_n3897, new_n3910);
nor_5  g01562(new_n3910, new_n3896, new_n3911);
xor_4  g01563(new_n3911, new_n3894, new_n3912);
or_5   g01564(n14148, n1152, new_n3913);
or_5   g01565(new_n3913, n7149, new_n3914);
or_5   g01566(new_n3914, n18558, new_n3915);
xor_4  g01567(new_n3915, n3468, new_n3916);
xnor_4 g01568(new_n3916, n19514, new_n3917);
xor_4  g01569(new_n3914, n18558, new_n3918_1);
and_5  g01570(new_n3918_1, n10053, new_n3919);
xnor_4 g01571(new_n3918_1, n10053, new_n3920);
xor_4  g01572(new_n3913, n7149, new_n3921);
and_5  g01573(new_n3921, n8399, new_n3922);
xnor_4 g01574(new_n3921, n8399, new_n3923);
xor_4  g01575(n14148, n1152, new_n3924);
and_5  g01576(new_n3924, n9507, new_n3925_1);
and_5  g01577(n26979, n1152, new_n3926);
xor_4  g01578(new_n3924, n9507, new_n3927);
and_5  g01579(new_n3927, new_n3926, new_n3928);
nor_5  g01580(new_n3928, new_n3925_1, new_n3929);
nor_5  g01581(new_n3929, new_n3923, new_n3930);
nor_5  g01582(new_n3930, new_n3922, new_n3931);
nor_5  g01583(new_n3931, new_n3920, new_n3932_1);
nor_5  g01584(new_n3932_1, new_n3919, new_n3933);
xor_4  g01585(new_n3933, new_n3917, new_n3934_1);
or_5   g01586(n10057, n8920, new_n3935);
or_5   g01587(new_n3935, n26748, new_n3936);
or_5   g01588(new_n3936, n21276, new_n3937);
xor_4  g01589(new_n3937, n13668, new_n3938);
xnor_4 g01590(new_n3938, n626, new_n3939);
xor_4  g01591(new_n3936, n21276, new_n3940);
and_5  g01592(new_n3940, n1204, new_n3941);
xnor_4 g01593(new_n3940, n1204, new_n3942);
xor_4  g01594(new_n3935, n26748, new_n3943);
and_5  g01595(new_n3943, n19618, new_n3944);
xnor_4 g01596(new_n3943, n19618, new_n3945_1);
xor_4  g01597(n10057, n8920, new_n3946);
nor_5  g01598(new_n3946, n22043, new_n3947);
nand_5 g01599(n12121, n8920, new_n3948);
xor_4  g01600(new_n3946, n22043, new_n3949);
and_5  g01601(new_n3949, new_n3948, new_n3950);
or_5   g01602(new_n3950, new_n3947, new_n3951);
nor_5  g01603(new_n3951, new_n3945_1, new_n3952_1);
nor_5  g01604(new_n3952_1, new_n3944, new_n3953);
nor_5  g01605(new_n3953, new_n3942, new_n3954);
nor_5  g01606(new_n3954, new_n3941, new_n3955);
xor_4  g01607(new_n3955, new_n3939, new_n3956);
xnor_4 g01608(new_n3956, new_n3934_1, new_n3957);
xor_4  g01609(new_n3931, new_n3920, new_n3958);
not_10 g01610(new_n3958, new_n3959_1);
xnor_4 g01611(new_n3953, new_n3942, new_n3960);
nor_5  g01612(new_n3960, new_n3959_1, new_n3961);
xor_4  g01613(new_n3960, new_n3958, new_n3962_1);
xnor_4 g01614(new_n3951, new_n3945_1, new_n3963);
xnor_4 g01615(new_n3927, new_n3926, new_n3964);
xor_4  g01616(new_n3949, new_n3948, new_n3965);
nor_5  g01617(new_n3965, new_n3964, new_n3966);
xnor_4 g01618(n12121, n8920, new_n3967);
xnor_4 g01619(n26979, n1152, new_n3968);
or_5   g01620(new_n3968, new_n3967, new_n3969);
xnor_4 g01621(new_n3965, new_n3964, new_n3970);
nor_5  g01622(new_n3970, new_n3969, new_n3971_1);
nor_5  g01623(new_n3971_1, new_n3966, new_n3972);
nor_5  g01624(new_n3972, new_n3963, new_n3973);
xor_4  g01625(new_n3929, new_n3923, new_n3974);
xor_4  g01626(new_n3972, new_n3963, new_n3975);
and_5  g01627(new_n3975, new_n3974, new_n3976);
nor_5  g01628(new_n3976, new_n3973, new_n3977);
nor_5  g01629(new_n3977, new_n3962_1, new_n3978);
nor_5  g01630(new_n3978, new_n3961, new_n3979);
xor_4  g01631(new_n3979, new_n3957, new_n3980);
xnor_4 g01632(new_n3980, new_n3912, new_n3981);
xor_4  g01633(new_n3909_1, new_n3897, new_n3982);
xor_4  g01634(new_n3977, new_n3962_1, new_n3983_1);
and_5  g01635(new_n3983_1, new_n3982, new_n3984_1);
xnor_4 g01636(new_n3983_1, new_n3982, new_n3985);
xnor_4 g01637(new_n3975, new_n3974, new_n3986);
xor_4  g01638(new_n3907, new_n3900, new_n3987);
nor_5  g01639(new_n3987, new_n3986, new_n3988);
xnor_4 g01640(new_n3987, new_n3986, new_n3989);
xor_4  g01641(new_n3970, new_n3969, new_n3990);
nor_5  g01642(new_n3990, new_n3905, new_n3991);
not_10 g01643(new_n3990, new_n3992);
and_5  g01644(n25435, n24732, new_n3993);
xnor_4 g01645(new_n3905, new_n3993, new_n3994);
or_5   g01646(new_n3994, new_n3992, new_n3995);
xnor_4 g01647(n25435, n24732, new_n3996);
xnor_4 g01648(new_n3968, new_n3967, new_n3997);
or_5   g01649(new_n3997, new_n3996, new_n3998);
and_5  g01650(new_n3998, new_n3995, new_n3999);
or_5   g01651(new_n3999, new_n3991, new_n4000_1);
nor_5  g01652(new_n4000_1, new_n3989, new_n4001);
nor_5  g01653(new_n4001, new_n3988, new_n4002);
nor_5  g01654(new_n4002, new_n3985, new_n4003);
nor_5  g01655(new_n4003, new_n3984_1, new_n4004);
xnor_4 g01656(new_n4004, new_n3981, n266);
not_10 g01657(n21839, new_n4006);
nor_5  g01658(n22270, new_n4006, new_n4007);
xor_4  g01659(n22270, n21839, new_n4008);
not_10 g01660(n27089, new_n4009);
nor_5  g01661(new_n4009, n8806, new_n4010_1);
xor_4  g01662(n27089, n8806, new_n4011);
not_10 g01663(n11841, new_n4012);
nor_5  g01664(new_n4012, n2479, new_n4013);
xor_4  g01665(n11841, n2479, new_n4014_1);
not_10 g01666(n10710, new_n4015);
nor_5  g01667(new_n4015, n9372, new_n4016);
xor_4  g01668(n10710, n9372, new_n4017);
not_10 g01669(n20929, new_n4018);
nor_5  g01670(new_n4018, n6596, new_n4019);
xor_4  g01671(n20929, n6596, new_n4020);
not_10 g01672(n8006, new_n4021);
nor_5  g01673(n15289, new_n4021, new_n4022);
xor_4  g01674(n15289, n8006, new_n4023);
not_10 g01675(n25074, new_n4024);
nor_5  g01676(new_n4024, n6556, new_n4025);
xor_4  g01677(n25074, n6556, new_n4026);
not_10 g01678(n16396, new_n4027);
and_5  g01679(n22871, new_n4027, new_n4028);
nor_5  g01680(n22871, new_n4027, new_n4029);
not_10 g01681(n9399, new_n4030);
and_5  g01682(n14275, new_n4030, new_n4031);
or_5   g01683(n14275, new_n4030, new_n4032);
not_10 g01684(n2088, new_n4033);
and_5  g01685(n25023, new_n4033, new_n4034);
and_5  g01686(new_n4034, new_n4032, new_n4035);
nor_5  g01687(new_n4035, new_n4031, new_n4036);
nor_5  g01688(new_n4036, new_n4029, new_n4037);
or_5   g01689(new_n4037, new_n4028, new_n4038);
nor_5  g01690(new_n4038, new_n4026, new_n4039);
nor_5  g01691(new_n4039, new_n4025, new_n4040);
nor_5  g01692(new_n4040, new_n4023, new_n4041);
nor_5  g01693(new_n4041, new_n4022, new_n4042);
nor_5  g01694(new_n4042, new_n4020, new_n4043);
nor_5  g01695(new_n4043, new_n4019, new_n4044);
nor_5  g01696(new_n4044, new_n4017, new_n4045);
nor_5  g01697(new_n4045, new_n4016, new_n4046);
nor_5  g01698(new_n4046, new_n4014_1, new_n4047);
nor_5  g01699(new_n4047, new_n4013, new_n4048);
nor_5  g01700(new_n4048, new_n4011, new_n4049);
nor_5  g01701(new_n4049, new_n4010_1, new_n4050);
nor_5  g01702(new_n4050, new_n4008, new_n4051);
nor_5  g01703(new_n4051, new_n4007, new_n4052);
xor_4  g01704(new_n4050, new_n4008, new_n4053);
nor_5  g01705(new_n4053, n23272, new_n4054);
xnor_4 g01706(new_n4053, n23272, new_n4055);
xor_4  g01707(new_n4048, new_n4011, new_n4056);
nor_5  g01708(new_n4056, n11481, new_n4057);
xnor_4 g01709(new_n4056, n11481, new_n4058);
xor_4  g01710(new_n4046, new_n4014_1, new_n4059);
nor_5  g01711(new_n4059, n16439, new_n4060);
xnor_4 g01712(new_n4059, n16439, new_n4061);
xor_4  g01713(new_n4044, new_n4017, new_n4062);
nor_5  g01714(new_n4062, n15241, new_n4063);
xnor_4 g01715(new_n4062, n15241, new_n4064);
xor_4  g01716(new_n4042, new_n4020, new_n4065);
nor_5  g01717(new_n4065, n7678, new_n4066);
xnor_4 g01718(new_n4065, n7678, new_n4067);
xor_4  g01719(new_n4040, new_n4023, new_n4068);
nor_5  g01720(new_n4068, n3785, new_n4069);
xnor_4 g01721(new_n4068, n3785, new_n4070);
xor_4  g01722(new_n4038, new_n4026, new_n4071_1);
nor_5  g01723(new_n4071_1, n20250, new_n4072);
not_10 g01724(n20250, new_n4073);
xnor_4 g01725(new_n4071_1, new_n4073, new_n4074);
not_10 g01726(n5822, new_n4075);
xnor_4 g01727(n22871, n16396, new_n4076);
xnor_4 g01728(new_n4076, new_n4036, new_n4077);
nor_5  g01729(new_n4077, new_n4075, new_n4078);
and_5  g01730(new_n4077, new_n4075, new_n4079);
not_10 g01731(n26443, new_n4080);
xor_4  g01732(n14275, n9399, new_n4081);
xnor_4 g01733(new_n4081, new_n4034, new_n4082);
and_5  g01734(new_n4082, new_n4080, new_n4083);
not_10 g01735(n1681, new_n4084);
xnor_4 g01736(n25023, n2088, new_n4085_1);
or_5   g01737(new_n4085_1, new_n4084, new_n4086);
xnor_4 g01738(new_n4082, n26443, new_n4087);
and_5  g01739(new_n4087, new_n4086, new_n4088_1);
or_5   g01740(new_n4088_1, new_n4083, new_n4089_1);
nor_5  g01741(new_n4089_1, new_n4079, new_n4090);
nor_5  g01742(new_n4090, new_n4078, new_n4091);
and_5  g01743(new_n4091, new_n4074, new_n4092);
nor_5  g01744(new_n4092, new_n4072, new_n4093);
nor_5  g01745(new_n4093, new_n4070, new_n4094);
nor_5  g01746(new_n4094, new_n4069, new_n4095);
nor_5  g01747(new_n4095, new_n4067, new_n4096);
nor_5  g01748(new_n4096, new_n4066, new_n4097);
nor_5  g01749(new_n4097, new_n4064, new_n4098);
nor_5  g01750(new_n4098, new_n4063, new_n4099);
nor_5  g01751(new_n4099, new_n4061, new_n4100_1);
nor_5  g01752(new_n4100_1, new_n4060, new_n4101);
nor_5  g01753(new_n4101, new_n4058, new_n4102);
nor_5  g01754(new_n4102, new_n4057, new_n4103_1);
nor_5  g01755(new_n4103_1, new_n4055, new_n4104);
nor_5  g01756(new_n4104, new_n4054, new_n4105);
and_5  g01757(new_n4105, new_n4052, new_n4106);
or_5   g01758(new_n3700, n19477, new_n4107);
or_5   g01759(new_n4107, n9318, new_n4108);
or_5   g01760(new_n4108, n25168, new_n4109);
or_5   g01761(new_n4109, n1999, new_n4110);
nor_5  g01762(new_n4110, n9396, new_n4111);
xor_4  g01763(new_n4110, n9396, new_n4112);
nor_5  g01764(new_n4112, n18880, new_n4113);
xor_4  g01765(new_n4109, n1999, new_n4114);
nor_5  g01766(new_n4114, n25475, new_n4115);
xnor_4 g01767(new_n4114, n25475, new_n4116);
xor_4  g01768(new_n4108, n25168, new_n4117);
nor_5  g01769(new_n4117, n23849, new_n4118);
xnor_4 g01770(new_n4117, n23849, new_n4119_1);
xor_4  g01771(new_n4107, n9318, new_n4120);
nor_5  g01772(new_n4120, n12446, new_n4121);
nor_5  g01773(new_n3701, n11011, new_n4122);
nor_5  g01774(new_n3724, new_n3702, new_n4123_1);
nor_5  g01775(new_n4123_1, new_n4122, new_n4124);
xnor_4 g01776(new_n4120, n12446, new_n4125);
nor_5  g01777(new_n4125, new_n4124, new_n4126);
nor_5  g01778(new_n4126, new_n4121, new_n4127);
nor_5  g01779(new_n4127, new_n4119_1, new_n4128);
nor_5  g01780(new_n4128, new_n4118, new_n4129);
nor_5  g01781(new_n4129, new_n4116, new_n4130);
nor_5  g01782(new_n4130, new_n4115, new_n4131);
and_5  g01783(new_n4112, n18880, new_n4132);
nor_5  g01784(new_n4132, new_n4131, new_n4133);
nor_5  g01785(new_n4133, new_n4113, new_n4134_1);
nor_5  g01786(new_n4134_1, new_n4111, new_n4135);
not_10 g01787(new_n4135, new_n4136);
not_10 g01788(n6785, new_n4137);
nor_5  g01789(n24032, n22843, new_n4138);
nand_5 g01790(new_n4138, new_n4137, new_n4139);
or_5   g01791(new_n4139, n24879, new_n4140);
or_5   g01792(new_n4140, n268, new_n4141);
or_5   g01793(new_n4141, n12587, new_n4142);
or_5   g01794(new_n4142, n25381, new_n4143);
or_5   g01795(new_n4143, n16376, new_n4144);
or_5   g01796(new_n4144, n24196, new_n4145);
xnor_4 g01797(new_n4145, n18105, new_n4146_1);
xor_4  g01798(new_n4112, n18880, new_n4147);
xnor_4 g01799(new_n4147, new_n4131, new_n4148);
nor_5  g01800(new_n4148, new_n4146_1, new_n4149);
nor_5  g01801(new_n4145, n18105, new_n4150_1);
xor_4  g01802(new_n4148, new_n4146_1, new_n4151_1);
xor_4  g01803(new_n4144, n24196, new_n4152_1);
xnor_4 g01804(new_n4129, new_n4116, new_n4153_1);
nor_5  g01805(new_n4153_1, new_n4152_1, new_n4154);
xnor_4 g01806(new_n4153_1, new_n4152_1, new_n4155);
xor_4  g01807(new_n4143, n16376, new_n4156);
xnor_4 g01808(new_n4127, new_n4119_1, new_n4157);
nor_5  g01809(new_n4157, new_n4156, new_n4158);
xnor_4 g01810(new_n4157, new_n4156, new_n4159);
xor_4  g01811(new_n4142, n25381, new_n4160);
xnor_4 g01812(new_n4125, new_n4124, new_n4161);
nor_5  g01813(new_n4161, new_n4160, new_n4162);
xnor_4 g01814(new_n4161, new_n4160, new_n4163);
xor_4  g01815(new_n4141, n12587, new_n4164);
nor_5  g01816(new_n4164, new_n3725_1, new_n4165_1);
xnor_4 g01817(new_n4164, new_n3725_1, new_n4166);
xor_4  g01818(new_n4140, n268, new_n4167);
nor_5  g01819(new_n4167, new_n3727, new_n4168);
xor_4  g01820(new_n4139, n24879, new_n4169);
nor_5  g01821(new_n4169, new_n3729, new_n4170);
xnor_4 g01822(new_n4169, new_n3729, new_n4171);
xor_4  g01823(new_n4138, n6785, new_n4172_1);
nor_5  g01824(new_n4172_1, new_n3733_1, new_n4173_1);
xnor_4 g01825(new_n4172_1, new_n3733_1, new_n4174);
xor_4  g01826(n24032, n22843, new_n4175);
nor_5  g01827(new_n4175, new_n3738, new_n4176_1);
nand_5 g01828(new_n2530, n22843, new_n4177);
xnor_4 g01829(new_n4175, new_n3737, new_n4178);
and_5  g01830(new_n4178, new_n4177, new_n4179);
or_5   g01831(new_n4179, new_n4176_1, new_n4180);
nor_5  g01832(new_n4180, new_n4174, new_n4181);
or_5   g01833(new_n4181, new_n4173_1, new_n4182);
nor_5  g01834(new_n4182, new_n4171, new_n4183);
nor_5  g01835(new_n4183, new_n4170, new_n4184);
xnor_4 g01836(new_n4167, new_n3727, new_n4185);
nor_5  g01837(new_n4185, new_n4184, new_n4186_1);
nor_5  g01838(new_n4186_1, new_n4168, new_n4187);
nor_5  g01839(new_n4187, new_n4166, new_n4188);
nor_5  g01840(new_n4188, new_n4165_1, new_n4189);
nor_5  g01841(new_n4189, new_n4163, new_n4190);
nor_5  g01842(new_n4190, new_n4162, new_n4191);
nor_5  g01843(new_n4191, new_n4159, new_n4192);
nor_5  g01844(new_n4192, new_n4158, new_n4193);
nor_5  g01845(new_n4193, new_n4155, new_n4194);
nor_5  g01846(new_n4194, new_n4154, new_n4195);
and_5  g01847(new_n4195, new_n4151_1, new_n4196);
or_5   g01848(new_n4196, new_n4150_1, new_n4197);
nor_5  g01849(new_n4197, new_n4149, new_n4198);
and_5  g01850(new_n4198, new_n4136, new_n4199);
xnor_4 g01851(new_n4199, new_n4106, new_n4200);
xor_4  g01852(new_n4105, new_n4052, new_n4201);
not_10 g01853(new_n4201, new_n4202);
xnor_4 g01854(new_n4198, new_n4135, new_n4203);
and_5  g01855(new_n4203, new_n4202, new_n4204_1);
xor_4  g01856(new_n4203, new_n4201, new_n4205_1);
xnor_4 g01857(new_n4195, new_n4151_1, new_n4206);
xor_4  g01858(new_n4103_1, new_n4055, new_n4207);
and_5  g01859(new_n4207, new_n4206, new_n4208);
xnor_4 g01860(new_n4207, new_n4206, new_n4209);
xor_4  g01861(new_n4193, new_n4155, new_n4210);
xor_4  g01862(new_n4101, new_n4058, new_n4211);
and_5  g01863(new_n4211, new_n4210, new_n4212);
xnor_4 g01864(new_n4211, new_n4210, new_n4213);
xor_4  g01865(new_n4191, new_n4159, new_n4214);
xor_4  g01866(new_n4099, new_n4061, new_n4215_1);
and_5  g01867(new_n4215_1, new_n4214, new_n4216);
xnor_4 g01868(new_n4215_1, new_n4214, new_n4217);
xor_4  g01869(new_n4189, new_n4163, new_n4218);
xor_4  g01870(new_n4097, new_n4064, new_n4219);
and_5  g01871(new_n4219, new_n4218, new_n4220);
xnor_4 g01872(new_n4219, new_n4218, new_n4221_1);
xor_4  g01873(new_n4187, new_n4166, new_n4222);
xor_4  g01874(new_n4095, new_n4067, new_n4223);
and_5  g01875(new_n4223, new_n4222, new_n4224_1);
xnor_4 g01876(new_n4223, new_n4222, new_n4225);
xor_4  g01877(new_n4093, new_n4070, new_n4226);
xor_4  g01878(new_n4185, new_n4184, new_n4227);
and_5  g01879(new_n4227, new_n4226, new_n4228);
xnor_4 g01880(new_n4227, new_n4226, new_n4229);
xor_4  g01881(new_n4182, new_n4171, new_n4230);
xor_4  g01882(new_n4091, new_n4074, new_n4231_1);
and_5  g01883(new_n4231_1, new_n4230, new_n4232);
xor_4  g01884(new_n4231_1, new_n4230, new_n4233);
xnor_4 g01885(new_n4180, new_n4174, new_n4234);
xnor_4 g01886(new_n4077, n5822, new_n4235);
xnor_4 g01887(new_n4235, new_n4089_1, new_n4236);
not_10 g01888(new_n4236, new_n4237);
nor_5  g01889(new_n4237, new_n4234, new_n4238);
xor_4  g01890(new_n4087, new_n4086, new_n4239);
xor_4  g01891(new_n4178, new_n4177, new_n4240);
and_5  g01892(new_n4240, new_n4239, new_n4241);
xor_4  g01893(new_n2530, n22843, new_n4242);
xnor_4 g01894(new_n4085_1, n1681, new_n4243);
nand_5 g01895(new_n4243, new_n4242, new_n4244);
xor_4  g01896(new_n4240, new_n4239, new_n4245);
and_5  g01897(new_n4245, new_n4244, new_n4246);
or_5   g01898(new_n4246, new_n4241, new_n4247);
xor_4  g01899(new_n4236, new_n4234, new_n4248);
nor_5  g01900(new_n4248, new_n4247, new_n4249);
nor_5  g01901(new_n4249, new_n4238, new_n4250);
and_5  g01902(new_n4250, new_n4233, new_n4251);
nor_5  g01903(new_n4251, new_n4232, new_n4252);
nor_5  g01904(new_n4252, new_n4229, new_n4253);
nor_5  g01905(new_n4253, new_n4228, new_n4254);
nor_5  g01906(new_n4254, new_n4225, new_n4255);
nor_5  g01907(new_n4255, new_n4224_1, new_n4256_1);
nor_5  g01908(new_n4256_1, new_n4221_1, new_n4257);
nor_5  g01909(new_n4257, new_n4220, new_n4258);
nor_5  g01910(new_n4258, new_n4217, new_n4259);
nor_5  g01911(new_n4259, new_n4216, new_n4260);
nor_5  g01912(new_n4260, new_n4213, new_n4261);
nor_5  g01913(new_n4261, new_n4212, new_n4262);
nor_5  g01914(new_n4262, new_n4209, new_n4263);
nor_5  g01915(new_n4263, new_n4208, new_n4264);
nor_5  g01916(new_n4264, new_n4205_1, new_n4265);
nor_5  g01917(new_n4265, new_n4204_1, new_n4266_1);
xnor_4 g01918(new_n4266_1, new_n4200, n298);
xor_4  g01919(n21735, n20604, new_n4268);
not_10 g01920(n24085, new_n4269);
nor_5  g01921(new_n4269, n16158, new_n4270);
xor_4  g01922(n24085, n16158, new_n4271);
not_10 g01923(n14071, new_n4272_1);
nor_5  g01924(new_n4272_1, n5752, new_n4273);
xor_4  g01925(n14071, n5752, new_n4274);
not_10 g01926(n1738, new_n4275);
and_5  g01927(n18171, new_n4275, new_n4276);
nor_5  g01928(n18171, new_n4275, new_n4277);
not_10 g01929(n12152, new_n4278);
and_5  g01930(n25073, new_n4278, new_n4279);
or_5   g01931(n25073, new_n4278, new_n4280);
not_10 g01932(n22309, new_n4281);
nor_5  g01933(new_n4281, n19107, new_n4282);
and_5  g01934(new_n4282, new_n4280, new_n4283);
nor_5  g01935(new_n4283, new_n4279, new_n4284);
nor_5  g01936(new_n4284, new_n4277, new_n4285);
or_5   g01937(new_n4285, new_n4276, new_n4286);
nor_5  g01938(new_n4286, new_n4274, new_n4287);
nor_5  g01939(new_n4287, new_n4273, new_n4288);
nor_5  g01940(new_n4288, new_n4271, new_n4289);
nor_5  g01941(new_n4289, new_n4270, new_n4290);
xor_4  g01942(new_n4290, new_n4268, new_n4291);
xor_4  g01943(n4119, n1525, new_n4292);
not_10 g01944(n16988, new_n4293);
nor_5  g01945(new_n4293, n14510, new_n4294);
xor_4  g01946(n16988, n14510, new_n4295);
not_10 g01947(n21779, new_n4296);
nor_5  g01948(new_n4296, n13263, new_n4297);
xor_4  g01949(n21779, n13263, new_n4298);
not_10 g01950(n20455, new_n4299);
nor_5  g01951(new_n4299, n5376, new_n4300);
and_5  g01952(new_n4299, n5376, new_n4301);
nor_5  g01953(n5128, new_n3282, new_n4302);
nand_5 g01954(n5128, new_n3282, new_n4303);
not_10 g01955(n16968, new_n4304);
nor_5  g01956(n23120, new_n4304, new_n4305);
and_5  g01957(new_n4305, new_n4303, new_n4306_1);
nor_5  g01958(new_n4306_1, new_n4302, new_n4307);
nor_5  g01959(new_n4307, new_n4301, new_n4308);
or_5   g01960(new_n4308, new_n4300, new_n4309);
nor_5  g01961(new_n4309, new_n4298, new_n4310);
nor_5  g01962(new_n4310, new_n4297, new_n4311);
nor_5  g01963(new_n4311, new_n4295, new_n4312);
nor_5  g01964(new_n4312, new_n4294, new_n4313);
xor_4  g01965(new_n4313, new_n4292, new_n4314);
xor_4  g01966(n12626, n4272, new_n4315);
not_10 g01967(n24319, new_n4316);
nor_5  g01968(new_n4316, n6971, new_n4317);
xor_4  g01969(n24319, n6971, new_n4318);
not_10 g01970(n7460, new_n4319_1);
nor_5  g01971(n22068, new_n4319_1, new_n4320);
xor_4  g01972(n22068, n7460, new_n4321);
not_10 g01973(n196, new_n4322);
and_5  g01974(n9460, new_n4322, new_n4323);
nor_5  g01975(n9460, new_n4322, new_n4324);
not_10 g01976(n11749, new_n4325_1);
and_5  g01977(n14954, new_n4325_1, new_n4326_1);
or_5   g01978(n14954, new_n4325_1, new_n4327);
not_10 g01979(n23831, new_n4328);
nor_5  g01980(new_n4328, n13424, new_n4329);
and_5  g01981(new_n4329, new_n4327, new_n4330);
nor_5  g01982(new_n4330, new_n4326_1, new_n4331);
nor_5  g01983(new_n4331, new_n4324, new_n4332);
or_5   g01984(new_n4332, new_n4323, new_n4333);
nor_5  g01985(new_n4333, new_n4321, new_n4334);
nor_5  g01986(new_n4334, new_n4320, new_n4335);
nor_5  g01987(new_n4335, new_n4318, new_n4336);
nor_5  g01988(new_n4336, new_n4317, new_n4337);
xor_4  g01989(new_n4337, new_n4315, new_n4338);
xnor_4 g01990(new_n4338, new_n4314, new_n4339);
xnor_4 g01991(new_n4311, new_n4295, new_n4340_1);
xnor_4 g01992(new_n4335, new_n4318, new_n4341);
nor_5  g01993(new_n4341, new_n4340_1, new_n4342);
xnor_4 g01994(new_n4341, new_n4340_1, new_n4343);
xor_4  g01995(new_n4309, new_n4298, new_n4344);
xor_4  g01996(new_n4333, new_n4321, new_n4345);
nor_5  g01997(new_n4345, new_n4344, new_n4346);
xnor_4 g01998(new_n4345, new_n4344, new_n4347);
xor_4  g01999(n20455, n5376, new_n4348);
xnor_4 g02000(new_n4348, new_n4307, new_n4349);
xnor_4 g02001(n9460, n196, new_n4350);
xnor_4 g02002(new_n4350, new_n4331, new_n4351);
not_10 g02003(new_n4351, new_n4352);
nor_5  g02004(new_n4352, new_n4349, new_n4353);
xnor_4 g02005(new_n4351, new_n4349, new_n4354);
xor_4  g02006(n5128, n1639, new_n4355);
xnor_4 g02007(new_n4355, new_n4305, new_n4356);
xor_4  g02008(n14954, n11749, new_n4357);
xnor_4 g02009(new_n4357, new_n4329, new_n4358);
nor_5  g02010(new_n4358, new_n4356, new_n4359);
xnor_4 g02011(n23120, n16968, new_n4360);
xnor_4 g02012(n23831, n13424, new_n4361);
nor_5  g02013(new_n4361, new_n4360, new_n4362);
xor_4  g02014(new_n4358, new_n4356, new_n4363);
and_5  g02015(new_n4363, new_n4362, new_n4364);
nor_5  g02016(new_n4364, new_n4359, new_n4365);
and_5  g02017(new_n4365, new_n4354, new_n4366);
nor_5  g02018(new_n4366, new_n4353, new_n4367);
nor_5  g02019(new_n4367, new_n4347, new_n4368);
or_5   g02020(new_n4368, new_n4346, new_n4369);
nor_5  g02021(new_n4369, new_n4343, new_n4370);
nor_5  g02022(new_n4370, new_n4342, new_n4371);
xor_4  g02023(new_n4371, new_n4339, new_n4372);
xnor_4 g02024(new_n4372, new_n4291, new_n4373);
xor_4  g02025(new_n4288, new_n4271, new_n4374_1);
xor_4  g02026(new_n4369, new_n4343, new_n4375);
nor_5  g02027(new_n4375, new_n4374_1, new_n4376_1);
xnor_4 g02028(new_n4375, new_n4374_1, new_n4377);
xnor_4 g02029(new_n4367, new_n4347, new_n4378);
xor_4  g02030(new_n4286, new_n4274, new_n4379);
nor_5  g02031(new_n4379, new_n4378, new_n4380);
xor_4  g02032(new_n4365, new_n4354, new_n4381);
xnor_4 g02033(n18171, n1738, new_n4382);
xnor_4 g02034(new_n4382, new_n4284, new_n4383);
and_5  g02035(new_n4383, new_n4381, new_n4384);
xnor_4 g02036(new_n4383, new_n4381, new_n4385);
xnor_4 g02037(n22309, n19107, new_n4386);
xnor_4 g02038(new_n4361, new_n4360, new_n4387);
or_5   g02039(new_n4387, new_n4386, new_n4388);
xor_4  g02040(n25073, n12152, new_n4389);
xnor_4 g02041(new_n4389, new_n4282, new_n4390);
and_5  g02042(new_n4390, new_n4388, new_n4391);
xnor_4 g02043(new_n4363, new_n4362, new_n4392);
xor_4  g02044(new_n4390, new_n4388, new_n4393);
and_5  g02045(new_n4393, new_n4392, new_n4394);
nor_5  g02046(new_n4394, new_n4391, new_n4395);
nor_5  g02047(new_n4395, new_n4385, new_n4396);
nor_5  g02048(new_n4396, new_n4384, new_n4397);
xnor_4 g02049(new_n4379, new_n4378, new_n4398);
nor_5  g02050(new_n4398, new_n4397, new_n4399);
nor_5  g02051(new_n4399, new_n4380, new_n4400);
nor_5  g02052(new_n4400, new_n4377, new_n4401_1);
or_5   g02053(new_n4401_1, new_n4376_1, new_n4402);
xor_4  g02054(new_n4402, new_n4373, n317);
nor_5  g02055(n9934, n3506, new_n4404);
xnor_4 g02056(n9934, n3506, new_n4405);
nor_5  g02057(n18496, n14899, new_n4406);
xnor_4 g02058(n18496, n14899, new_n4407);
nor_5  g02059(n26224, n18444, new_n4408);
xnor_4 g02060(n26224, n18444, new_n4409_1);
nor_5  g02061(n24638, n19327, new_n4410);
xnor_4 g02062(n24638, n19327, new_n4411);
nor_5  g02063(n22597, n21674, new_n4412);
xnor_4 g02064(n22597, n21674, new_n4413);
nor_5  g02065(n26107, n17251, new_n4414);
xnor_4 g02066(n26107, n17251, new_n4415);
nor_5  g02067(n14790, n342, new_n4416);
xnor_4 g02068(n14790, n342, new_n4417);
nor_5  g02069(n26553, n10096, new_n4418);
xnor_4 g02070(n26553, n10096, new_n4419);
nor_5  g02071(n16994, n4964, new_n4420);
and_5  g02072(n9246, n7876, new_n4421);
xnor_4 g02073(n16994, n4964, new_n4422);
nor_5  g02074(new_n4422, new_n4421, new_n4423);
nor_5  g02075(new_n4423, new_n4420, new_n4424_1);
nor_5  g02076(new_n4424_1, new_n4419, new_n4425);
nor_5  g02077(new_n4425, new_n4418, new_n4426_1);
nor_5  g02078(new_n4426_1, new_n4417, new_n4427);
nor_5  g02079(new_n4427, new_n4416, new_n4428);
nor_5  g02080(new_n4428, new_n4415, new_n4429);
nor_5  g02081(new_n4429, new_n4414, new_n4430);
nor_5  g02082(new_n4430, new_n4413, new_n4431);
nor_5  g02083(new_n4431, new_n4412, new_n4432_1);
nor_5  g02084(new_n4432_1, new_n4411, new_n4433);
nor_5  g02085(new_n4433, new_n4410, new_n4434);
nor_5  g02086(new_n4434, new_n4409_1, new_n4435);
nor_5  g02087(new_n4435, new_n4408, new_n4436);
nor_5  g02088(new_n4436, new_n4407, new_n4437);
nor_5  g02089(new_n4437, new_n4406, new_n4438);
nor_5  g02090(new_n4438, new_n4405, new_n4439);
nor_5  g02091(new_n4439, new_n4404, new_n4440);
not_10 g02092(n9259, new_n4441_1);
xnor_4 g02093(n9554, n2979, new_n4442);
nor_5  g02094(n26408, n647, new_n4443);
xnor_4 g02095(n26408, n647, new_n4444);
nor_5  g02096(n20409, n18227, new_n4445);
xnor_4 g02097(n20409, n18227, new_n4446);
nor_5  g02098(n25749, n7377, new_n4447);
xnor_4 g02099(n25749, n7377, new_n4448);
nor_5  g02100(n11630, n3161, new_n4449);
xnor_4 g02101(n11630, n3161, new_n4450);
nor_5  g02102(n13453, n9003, new_n4451_1);
xnor_4 g02103(n13453, n9003, new_n4452);
nor_5  g02104(n7421, n4957, new_n4453);
xnor_4 g02105(n7421, n4957, new_n4454);
nor_5  g02106(n19680, n7524, new_n4455);
xnor_4 g02107(n19680, n7524, new_n4456);
nor_5  g02108(n15743, n2809, new_n4457);
and_5  g02109(n20658, n15508, new_n4458);
xnor_4 g02110(n15743, n2809, new_n4459);
nor_5  g02111(new_n4459, new_n4458, new_n4460);
nor_5  g02112(new_n4460, new_n4457, new_n4461);
nor_5  g02113(new_n4461, new_n4456, new_n4462);
nor_5  g02114(new_n4462, new_n4455, new_n4463);
nor_5  g02115(new_n4463, new_n4454, new_n4464);
nor_5  g02116(new_n4464, new_n4453, new_n4465);
nor_5  g02117(new_n4465, new_n4452, new_n4466);
nor_5  g02118(new_n4466, new_n4451_1, new_n4467);
nor_5  g02119(new_n4467, new_n4450, new_n4468);
nor_5  g02120(new_n4468, new_n4449, new_n4469);
nor_5  g02121(new_n4469, new_n4448, new_n4470);
nor_5  g02122(new_n4470, new_n4447, new_n4471);
nor_5  g02123(new_n4471, new_n4446, new_n4472);
nor_5  g02124(new_n4472, new_n4445, new_n4473);
nor_5  g02125(new_n4473, new_n4444, new_n4474);
nor_5  g02126(new_n4474, new_n4443, new_n4475);
xor_4  g02127(new_n4475, new_n4442, new_n4476_1);
nor_5  g02128(new_n4476_1, new_n4441_1, new_n4477);
xor_4  g02129(new_n4476_1, n9259, new_n4478_1);
xor_4  g02130(new_n4473, new_n4444, new_n4479);
not_10 g02131(new_n4479, new_n4480);
and_5  g02132(new_n4480, n21489, new_n4481);
xor_4  g02133(new_n4479, n21489, new_n4482);
xor_4  g02134(new_n4471, new_n4446, new_n4483);
not_10 g02135(new_n4483, new_n4484);
and_5  g02136(new_n4484, n20213, new_n4485);
xor_4  g02137(new_n4483, n20213, new_n4486);
xor_4  g02138(new_n4469, new_n4448, new_n4487);
not_10 g02139(new_n4487, new_n4488);
and_5  g02140(new_n4488, n13912, new_n4489);
xor_4  g02141(new_n4487, n13912, new_n4490);
xor_4  g02142(new_n4467, new_n4450, new_n4491);
not_10 g02143(new_n4491, new_n4492);
and_5  g02144(new_n4492, n7670, new_n4493);
xor_4  g02145(new_n4491, n7670, new_n4494);
xor_4  g02146(new_n4465, new_n4452, new_n4495);
not_10 g02147(new_n4495, new_n4496);
and_5  g02148(new_n4496, n9598, new_n4497);
xor_4  g02149(new_n4495, n9598, new_n4498);
xor_4  g02150(new_n4463, new_n4454, new_n4499);
not_10 g02151(new_n4499, new_n4500);
and_5  g02152(new_n4500, n22290, new_n4501);
xor_4  g02153(new_n4499, n22290, new_n4502);
xor_4  g02154(new_n4461, new_n4456, new_n4503);
not_10 g02155(new_n4503, new_n4504);
nand_5 g02156(new_n4504, n11273, new_n4505);
xnor_4 g02157(new_n4459, new_n4458, new_n4506);
nor_5  g02158(new_n4506, n25565, new_n4507);
xnor_4 g02159(n20658, n15508, new_n4508);
nor_5  g02160(new_n4508, new_n3441, new_n4509);
xnor_4 g02161(new_n4506, n25565, new_n4510);
nor_5  g02162(new_n4510, new_n4509, new_n4511);
nor_5  g02163(new_n4511, new_n4507, new_n4512);
not_10 g02164(new_n4512, new_n4513);
xor_4  g02165(new_n4503, n11273, new_n4514_1);
or_5   g02166(new_n4514_1, new_n4513, new_n4515);
and_5  g02167(new_n4515, new_n4505, new_n4516);
nor_5  g02168(new_n4516, new_n4502, new_n4517);
nor_5  g02169(new_n4517, new_n4501, new_n4518);
nor_5  g02170(new_n4518, new_n4498, new_n4519);
nor_5  g02171(new_n4519, new_n4497, new_n4520);
nor_5  g02172(new_n4520, new_n4494, new_n4521);
nor_5  g02173(new_n4521, new_n4493, new_n4522);
nor_5  g02174(new_n4522, new_n4490, new_n4523);
nor_5  g02175(new_n4523, new_n4489, new_n4524);
nor_5  g02176(new_n4524, new_n4486, new_n4525);
nor_5  g02177(new_n4525, new_n4485, new_n4526);
nor_5  g02178(new_n4526, new_n4482, new_n4527);
nor_5  g02179(new_n4527, new_n4481, new_n4528);
nor_5  g02180(new_n4528, new_n4478_1, new_n4529_1);
nor_5  g02181(new_n4529_1, new_n4477, new_n4530);
nor_5  g02182(n9554, n2979, new_n4531);
nor_5  g02183(new_n4475, new_n4442, new_n4532);
or_5   g02184(new_n4532, new_n4531, new_n4533);
xnor_4 g02185(new_n4533, new_n4530, new_n4534);
xnor_4 g02186(new_n4528, new_n4478_1, new_n4535);
nor_5  g02187(new_n4535, n3740, new_n4536);
xor_4  g02188(new_n4528, new_n4478_1, new_n4537);
xnor_4 g02189(new_n4537, n3740, new_n4538);
xnor_4 g02190(new_n4526, new_n4482, new_n4539);
and_5  g02191(new_n4539, n2858, new_n4540);
xnor_4 g02192(new_n4539, n2858, new_n4541);
xnor_4 g02193(new_n4524, new_n4486, new_n4542);
and_5  g02194(new_n4542, n2659, new_n4543);
xnor_4 g02195(new_n4542, n2659, new_n4544);
xnor_4 g02196(new_n4522, new_n4490, new_n4545);
and_5  g02197(new_n4545, n24327, new_n4546);
xnor_4 g02198(new_n4545, n24327, new_n4547);
xnor_4 g02199(new_n4520, new_n4494, new_n4548);
and_5  g02200(new_n4548, n22198, new_n4549);
xnor_4 g02201(new_n4548, n22198, new_n4550);
xnor_4 g02202(new_n4518, new_n4498, new_n4551);
and_5  g02203(new_n4551, n20826, new_n4552_1);
xnor_4 g02204(new_n4551, n20826, new_n4553);
xnor_4 g02205(new_n4516, new_n4502, new_n4554);
and_5  g02206(new_n4554, n7305, new_n4555);
xor_4  g02207(new_n4514_1, new_n4512, new_n4556);
nor_5  g02208(new_n4556, n25872, new_n4557);
xor_4  g02209(new_n4556, n25872, new_n4558);
xor_4  g02210(new_n4510, new_n4509, new_n4559);
and_5  g02211(new_n4559, n20259, new_n4560);
xnor_4 g02212(new_n4508, n21993, new_n4561);
not_10 g02213(new_n4561, new_n4562);
or_5   g02214(new_n4562, n3925, new_n4563);
xor_4  g02215(new_n4559, n20259, new_n4564);
and_5  g02216(new_n4564, new_n4563, new_n4565);
nor_5  g02217(new_n4565, new_n4560, new_n4566);
and_5  g02218(new_n4566, new_n4558, new_n4567);
or_5   g02219(new_n4567, new_n4557, new_n4568);
xnor_4 g02220(new_n4554, n7305, new_n4569);
nor_5  g02221(new_n4569, new_n4568, new_n4570);
nor_5  g02222(new_n4570, new_n4555, new_n4571);
nor_5  g02223(new_n4571, new_n4553, new_n4572);
nor_5  g02224(new_n4572, new_n4552_1, new_n4573);
nor_5  g02225(new_n4573, new_n4550, new_n4574);
nor_5  g02226(new_n4574, new_n4549, new_n4575);
nor_5  g02227(new_n4575, new_n4547, new_n4576);
nor_5  g02228(new_n4576, new_n4546, new_n4577);
nor_5  g02229(new_n4577, new_n4544, new_n4578);
nor_5  g02230(new_n4578, new_n4543, new_n4579);
nor_5  g02231(new_n4579, new_n4541, new_n4580);
nor_5  g02232(new_n4580, new_n4540, new_n4581);
and_5  g02233(new_n4581, new_n4538, new_n4582);
nor_5  g02234(new_n4582, new_n4536, new_n4583);
xor_4  g02235(new_n4583, new_n4534, new_n4584);
xnor_4 g02236(new_n4584, new_n4440, new_n4585);
xor_4  g02237(new_n4438, new_n4405, new_n4586);
xor_4  g02238(new_n4581, new_n4538, new_n4587);
and_5  g02239(new_n4587, new_n4586, new_n4588_1);
xnor_4 g02240(new_n4587, new_n4586, new_n4589);
xor_4  g02241(new_n4436, new_n4407, new_n4590_1);
not_10 g02242(new_n4590_1, new_n4591);
xor_4  g02243(new_n4579, new_n4541, new_n4592);
nor_5  g02244(new_n4592, new_n4591, new_n4593);
xnor_4 g02245(new_n4592, new_n4591, new_n4594);
xor_4  g02246(new_n4434, new_n4409_1, new_n4595_1);
not_10 g02247(new_n4595_1, new_n4596);
xor_4  g02248(new_n4577, new_n4544, new_n4597);
nor_5  g02249(new_n4597, new_n4596, new_n4598);
xnor_4 g02250(new_n4597, new_n4596, new_n4599);
xor_4  g02251(new_n4432_1, new_n4411, new_n4600);
not_10 g02252(new_n4600, new_n4601);
xor_4  g02253(new_n4575, new_n4547, new_n4602);
nor_5  g02254(new_n4602, new_n4601, new_n4603);
xnor_4 g02255(new_n4602, new_n4601, new_n4604);
xor_4  g02256(new_n4430, new_n4413, new_n4605);
not_10 g02257(new_n4605, new_n4606);
xor_4  g02258(new_n4573, new_n4550, new_n4607);
nor_5  g02259(new_n4607, new_n4606, new_n4608);
xnor_4 g02260(new_n4607, new_n4606, new_n4609);
xor_4  g02261(new_n4428, new_n4415, new_n4610);
not_10 g02262(new_n4610, new_n4611);
xor_4  g02263(new_n4571, new_n4553, new_n4612);
nor_5  g02264(new_n4612, new_n4611, new_n4613);
xnor_4 g02265(new_n4612, new_n4611, new_n4614);
xnor_4 g02266(new_n4426_1, new_n4417, new_n4615);
xor_4  g02267(new_n4569, new_n4568, new_n4616);
nor_5  g02268(new_n4616, new_n4615, new_n4617);
xnor_4 g02269(new_n4616, new_n4615, new_n4618);
xnor_4 g02270(new_n4566, new_n4558, new_n4619);
xor_4  g02271(new_n4424_1, new_n4419, new_n4620);
not_10 g02272(new_n4620, new_n4621);
nor_5  g02273(new_n4621, new_n4619, new_n4622);
xnor_4 g02274(new_n4620, new_n4619, new_n4623);
xor_4  g02275(n16994, n4964, new_n4624_1);
xnor_4 g02276(new_n4561, n3925, new_n4625);
xnor_4 g02277(n9246, n7876, new_n4626);
nor_5  g02278(new_n4626, new_n4625, new_n4627);
and_5  g02279(new_n4627, new_n4624_1, new_n4628);
xnor_4 g02280(new_n4564, new_n4563, new_n4629);
xnor_4 g02281(new_n4422, new_n4421, new_n4630);
nor_5  g02282(new_n4630, new_n4627, new_n4631);
or_5   g02283(new_n4631, new_n4628, new_n4632);
nor_5  g02284(new_n4632, new_n4629, new_n4633);
nor_5  g02285(new_n4633, new_n4628, new_n4634);
and_5  g02286(new_n4634, new_n4623, new_n4635);
nor_5  g02287(new_n4635, new_n4622, new_n4636);
nor_5  g02288(new_n4636, new_n4618, new_n4637);
nor_5  g02289(new_n4637, new_n4617, new_n4638);
nor_5  g02290(new_n4638, new_n4614, new_n4639);
nor_5  g02291(new_n4639, new_n4613, new_n4640);
nor_5  g02292(new_n4640, new_n4609, new_n4641);
nor_5  g02293(new_n4641, new_n4608, new_n4642);
nor_5  g02294(new_n4642, new_n4604, new_n4643);
nor_5  g02295(new_n4643, new_n4603, new_n4644);
nor_5  g02296(new_n4644, new_n4599, new_n4645);
nor_5  g02297(new_n4645, new_n4598, new_n4646_1);
nor_5  g02298(new_n4646_1, new_n4594, new_n4647);
nor_5  g02299(new_n4647, new_n4593, new_n4648);
nor_5  g02300(new_n4648, new_n4589, new_n4649);
or_5   g02301(new_n4649, new_n4588_1, new_n4650);
xor_4  g02302(new_n4650, new_n4585, n332);
xnor_4 g02303(n18295, n16223, new_n4652);
nor_5  g02304(n19494, n6502, new_n4653);
and_5  g02305(n15780, n2387, new_n4654);
xnor_4 g02306(n19494, n6502, new_n4655);
nor_5  g02307(new_n4655, new_n4654, new_n4656);
nor_5  g02308(new_n4656, new_n4653, new_n4657);
xor_4  g02309(new_n4657, new_n4652, new_n4658);
xnor_4 g02310(new_n4658, n8381, new_n4659);
not_10 g02311(n20235, new_n4660);
xnor_4 g02312(n15780, n2387, new_n4661);
nor_5  g02313(new_n4661, n12495, new_n4662);
and_5  g02314(new_n4662, new_n4660, new_n4663);
xnor_4 g02315(new_n4662, n20235, new_n4664);
xor_4  g02316(new_n4655, new_n4654, new_n4665_1);
not_10 g02317(new_n4665_1, new_n4666);
and_5  g02318(new_n4666, new_n4664, new_n4667);
nor_5  g02319(new_n4667, new_n4663, new_n4668);
xnor_4 g02320(new_n4668, new_n4659, new_n4669);
not_10 g02321(n23146, new_n4670);
not_10 g02322(n16502, new_n4671);
nor_5  g02323(n21654, new_n4671, new_n4672);
xor_4  g02324(n25471, n23842, new_n4673);
xnor_4 g02325(new_n4673, new_n4672, new_n4674_1);
nor_5  g02326(new_n4674_1, new_n4670, new_n4675);
xor_4  g02327(n21654, n16502, new_n4676);
and_5  g02328(new_n4676, n17968, new_n4677);
xnor_4 g02329(new_n4674_1, n23146, new_n4678);
and_5  g02330(new_n4678, new_n4677, new_n4679);
nor_5  g02331(new_n4679, new_n4675, new_n4680);
xnor_4 g02332(n15053, n3828, new_n4681);
not_10 g02333(n25471, new_n4682);
nor_5  g02334(new_n4682, n23842, new_n4683);
or_5   g02335(n21654, new_n4671, new_n4684);
nor_5  g02336(new_n4673, new_n4684, new_n4685);
nor_5  g02337(new_n4685, new_n4683, new_n4686);
xnor_4 g02338(new_n4686, new_n4681, new_n4687);
xnor_4 g02339(new_n4687, n11184, new_n4688);
xnor_4 g02340(new_n4688, new_n4680, new_n4689);
xnor_4 g02341(new_n4689, new_n4669, new_n4690);
xor_4  g02342(new_n4678, new_n4677, new_n4691);
xnor_4 g02343(new_n4665_1, new_n4664, new_n4692);
not_10 g02344(new_n4692, new_n4693_1);
nor_5  g02345(new_n4693_1, new_n4691, new_n4694);
xor_4  g02346(new_n4661, n12495, new_n4695);
xnor_4 g02347(n21654, n16502, new_n4696);
xor_4  g02348(new_n4696, n17968, new_n4697);
or_5   g02349(new_n4697, new_n4695, new_n4698);
xnor_4 g02350(new_n4692, new_n4691, new_n4699);
and_5  g02351(new_n4699, new_n4698, new_n4700);
nor_5  g02352(new_n4700, new_n4694, new_n4701);
xnor_4 g02353(new_n4701, new_n4690, n357);
not_10 g02354(new_n3013, new_n4703);
xor_4  g02355(n22309, n9251, new_n4704);
and_5  g02356(n22309, n9251, new_n4705);
xnor_4 g02357(n25073, n20138, new_n4706);
xnor_4 g02358(new_n4706, new_n4705, new_n4707);
nor_5  g02359(new_n4707, new_n4704, new_n4708);
not_10 g02360(new_n4708, new_n4709);
xnor_4 g02361(n18171, n6385, new_n4710);
or_5   g02362(n25073, n20138, new_n4711);
or_5   g02363(new_n4706, new_n4705, new_n4712);
and_5  g02364(new_n4712, new_n4711, new_n4713);
xnor_4 g02365(new_n4713, new_n4710, new_n4714);
or_5   g02366(new_n4714, new_n4709, new_n4715);
xnor_4 g02367(n5752, n3136, new_n4716);
nor_5  g02368(n18171, n6385, new_n4717);
nor_5  g02369(new_n4713, new_n4710, new_n4718);
nor_5  g02370(new_n4718, new_n4717, new_n4719);
xor_4  g02371(new_n4719, new_n4716, new_n4720);
not_10 g02372(new_n4720, new_n4721);
or_5   g02373(new_n4721, new_n4715, new_n4722_1);
xnor_4 g02374(n16158, n9557, new_n4723);
nor_5  g02375(n5752, n3136, new_n4724);
nor_5  g02376(new_n4719, new_n4716, new_n4725);
nor_5  g02377(new_n4725, new_n4724, new_n4726);
xor_4  g02378(new_n4726, new_n4723, new_n4727);
not_10 g02379(new_n4727, new_n4728);
or_5   g02380(new_n4728, new_n4722_1, new_n4729);
xnor_4 g02381(n25643, n20604, new_n4730);
nor_5  g02382(n16158, n9557, new_n4731_1);
nor_5  g02383(new_n4726, new_n4723, new_n4732);
nor_5  g02384(new_n4732, new_n4731_1, new_n4733);
xor_4  g02385(new_n4733, new_n4730, new_n4734);
xnor_4 g02386(new_n4734, new_n4729, new_n4735);
xnor_4 g02387(new_n4735, new_n4703, new_n4736);
not_10 g02388(new_n3016, new_n4737);
xnor_4 g02389(new_n4727, new_n4722_1, new_n4738);
nor_5  g02390(new_n4738, new_n4737, new_n4739);
xnor_4 g02391(new_n4738, new_n4737, new_n4740);
not_10 g02392(new_n3019, new_n4741);
xnor_4 g02393(new_n4720, new_n4715, new_n4742);
nor_5  g02394(new_n4742, new_n4741, new_n4743);
xnor_4 g02395(new_n4742, new_n4741, new_n4744);
xor_4  g02396(new_n4714, new_n4708, new_n4745_1);
or_5   g02397(new_n4745_1, new_n3022, new_n4746);
not_10 g02398(new_n4704, new_n4747_1);
nor_5  g02399(new_n4747_1, new_n3026, new_n4748);
nor_5  g02400(new_n4748, new_n3030_1, new_n4749);
nor_5  g02401(n22309, n9251, new_n4750);
nor_5  g02402(new_n4712, new_n4750, new_n4751);
nor_5  g02403(new_n4751, new_n4708, new_n4752);
xor_4  g02404(n19494, n11121, new_n4753);
and_5  g02405(new_n4748, new_n4753, new_n4754);
or_5   g02406(new_n4754, new_n4749, new_n4755);
nor_5  g02407(new_n4755, new_n4752, new_n4756);
nor_5  g02408(new_n4756, new_n4749, new_n4757);
not_10 g02409(new_n4757, new_n4758);
xnor_4 g02410(new_n4745_1, new_n3022, new_n4759);
or_5   g02411(new_n4759, new_n4758, new_n4760);
nand_5 g02412(new_n4760, new_n4746, new_n4761);
nor_5  g02413(new_n4761, new_n4744, new_n4762);
nor_5  g02414(new_n4762, new_n4743, new_n4763);
nor_5  g02415(new_n4763, new_n4740, new_n4764);
nor_5  g02416(new_n4764, new_n4739, new_n4765);
xnor_4 g02417(new_n4765, new_n4736, new_n4766_1);
xor_4  g02418(n5255, n4119, new_n4767);
not_10 g02419(n21649, new_n4768);
nor_5  g02420(new_n4768, n14510, new_n4769);
xor_4  g02421(n21649, n14510, new_n4770_1);
not_10 g02422(n18274, new_n4771);
nor_5  g02423(new_n4771, n13263, new_n4772);
xor_4  g02424(n18274, n13263, new_n4773);
nor_5  g02425(new_n4299, n3828, new_n4774);
and_5  g02426(new_n4299, n3828, new_n4775);
nor_5  g02427(n23842, new_n3282, new_n4776);
nand_5 g02428(n23842, new_n3282, new_n4777_1);
nor_5  g02429(n21654, new_n4304, new_n4778);
and_5  g02430(new_n4778, new_n4777_1, new_n4779);
nor_5  g02431(new_n4779, new_n4776, new_n4780);
nor_5  g02432(new_n4780, new_n4775, new_n4781);
or_5   g02433(new_n4781, new_n4774, new_n4782);
nor_5  g02434(new_n4782, new_n4773, new_n4783);
nor_5  g02435(new_n4783, new_n4772, new_n4784);
nor_5  g02436(new_n4784, new_n4770_1, new_n4785_1);
nor_5  g02437(new_n4785_1, new_n4769, new_n4786);
xor_4  g02438(new_n4786, new_n4767, new_n4787);
xnor_4 g02439(new_n4787, new_n4766_1, new_n4788);
xnor_4 g02440(new_n4784, new_n4770_1, new_n4789);
xor_4  g02441(new_n4763, new_n4740, new_n4790);
and_5  g02442(new_n4790, new_n4789, new_n4791);
xnor_4 g02443(new_n4790, new_n4789, new_n4792);
xnor_4 g02444(new_n4761, new_n4744, new_n4793);
xor_4  g02445(new_n4782, new_n4773, new_n4794);
nor_5  g02446(new_n4794, new_n4793, new_n4795);
xnor_4 g02447(new_n4794, new_n4793, new_n4796);
xor_4  g02448(new_n4759, new_n4757, new_n4797);
xnor_4 g02449(n20455, n3828, new_n4798);
xnor_4 g02450(new_n4798, new_n4780, new_n4799);
and_5  g02451(new_n4799, new_n4797, new_n4800);
xnor_4 g02452(new_n4799, new_n4797, new_n4801);
xnor_4 g02453(n21654, n16968, new_n4802);
xor_4  g02454(new_n4704, new_n3026, new_n4803);
or_5   g02455(new_n4803, new_n4802, new_n4804_1);
xor_4  g02456(n23842, n1639, new_n4805);
xnor_4 g02457(new_n4805, new_n4778, new_n4806);
and_5  g02458(new_n4806, new_n4804_1, new_n4807);
xor_4  g02459(new_n4755, new_n4752, new_n4808);
xor_4  g02460(new_n4806, new_n4804_1, new_n4809);
and_5  g02461(new_n4809, new_n4808, new_n4810_1);
nor_5  g02462(new_n4810_1, new_n4807, new_n4811);
nor_5  g02463(new_n4811, new_n4801, new_n4812_1);
nor_5  g02464(new_n4812_1, new_n4800, new_n4813);
nor_5  g02465(new_n4813, new_n4796, new_n4814_1);
nor_5  g02466(new_n4814_1, new_n4795, new_n4815);
nor_5  g02467(new_n4815, new_n4792, new_n4816);
or_5   g02468(new_n4816, new_n4791, new_n4817);
xor_4  g02469(new_n4817, new_n4788, n422);
or_5   g02470(n23333, n20794, new_n4819);
or_5   g02471(new_n4819, n14603, new_n4820);
or_5   g02472(new_n4820, n18737, new_n4821);
or_5   g02473(new_n4821, n21471, new_n4822);
or_5   g02474(new_n4822, n25738, new_n4823);
or_5   g02475(new_n4823, n5302, new_n4824);
or_5   g02476(new_n4824, n3228, new_n4825);
xor_4  g02477(new_n4825, n337, new_n4826);
xnor_4 g02478(new_n4826, n6485, new_n4827);
xor_4  g02479(new_n4824, n3228, new_n4828);
nor_5  g02480(new_n4828, n26036, new_n4829);
xnor_4 g02481(new_n4828, n26036, new_n4830);
xor_4  g02482(new_n4823, n5302, new_n4831);
nor_5  g02483(new_n4831, n19770, new_n4832);
xnor_4 g02484(new_n4831, n19770, new_n4833);
xor_4  g02485(new_n4822, n25738, new_n4834);
nor_5  g02486(new_n4834, n8782, new_n4835);
xnor_4 g02487(new_n4834, n8782, new_n4836);
xor_4  g02488(new_n4821, n21471, new_n4837);
nor_5  g02489(new_n4837, n8678, new_n4838);
xnor_4 g02490(new_n4837, n8678, new_n4839);
xor_4  g02491(new_n4820, n18737, new_n4840);
nor_5  g02492(new_n4840, n1432, new_n4841);
xor_4  g02493(new_n4819, n14603, new_n4842);
nor_5  g02494(new_n4842, n21599, new_n4843);
xnor_4 g02495(new_n4842, n21599, new_n4844);
xor_4  g02496(n23333, n20794, new_n4845);
nor_5  g02497(new_n4845, n25336, new_n4846);
nand_5 g02498(n23333, n11424, new_n4847);
xor_4  g02499(new_n4845, n25336, new_n4848);
and_5  g02500(new_n4848, new_n4847, new_n4849);
nor_5  g02501(new_n4849, new_n4846, new_n4850_1);
nor_5  g02502(new_n4850_1, new_n4844, new_n4851);
nor_5  g02503(new_n4851, new_n4843, new_n4852);
xnor_4 g02504(new_n4840, n1432, new_n4853);
nor_5  g02505(new_n4853, new_n4852, new_n4854);
nor_5  g02506(new_n4854, new_n4841, new_n4855);
nor_5  g02507(new_n4855, new_n4839, new_n4856);
nor_5  g02508(new_n4856, new_n4838, new_n4857);
nor_5  g02509(new_n4857, new_n4836, new_n4858_1);
nor_5  g02510(new_n4858_1, new_n4835, new_n4859);
nor_5  g02511(new_n4859, new_n4833, new_n4860);
nor_5  g02512(new_n4860, new_n4832, new_n4861);
nor_5  g02513(new_n4861, new_n4830, new_n4862);
nor_5  g02514(new_n4862, new_n4829, new_n4863);
xnor_4 g02515(new_n4863, new_n4827, new_n4864);
xnor_4 g02516(n22379, n9967, new_n4865);
nor_5  g02517(n20946, n1662, new_n4866);
xnor_4 g02518(n20946, n1662, new_n4867);
nor_5  g02519(n12875, n7751, new_n4868);
xnor_4 g02520(n12875, n7751, new_n4869);
nor_5  g02521(n26823, n2035, new_n4870);
xnor_4 g02522(n26823, n2035, new_n4871);
nor_5  g02523(n5213, n4812, new_n4872);
xnor_4 g02524(n5213, n4812, new_n4873);
nor_5  g02525(n24278, n4665, new_n4874);
xnor_4 g02526(n24278, n4665, new_n4875);
nor_5  g02527(n24618, n19005, new_n4876);
xnor_4 g02528(n24618, n19005, new_n4877);
nor_5  g02529(n4326, n3952, new_n4878);
and_5  g02530(n12315, n5438, new_n4879);
xnor_4 g02531(n4326, n3952, new_n4880);
nor_5  g02532(new_n4880, new_n4879, new_n4881);
nor_5  g02533(new_n4881, new_n4878, new_n4882);
nor_5  g02534(new_n4882, new_n4877, new_n4883);
nor_5  g02535(new_n4883, new_n4876, new_n4884);
nor_5  g02536(new_n4884, new_n4875, new_n4885);
nor_5  g02537(new_n4885, new_n4874, new_n4886);
nor_5  g02538(new_n4886, new_n4873, new_n4887);
nor_5  g02539(new_n4887, new_n4872, new_n4888);
nor_5  g02540(new_n4888, new_n4871, new_n4889);
nor_5  g02541(new_n4889, new_n4870, new_n4890);
nor_5  g02542(new_n4890, new_n4869, new_n4891_1);
nor_5  g02543(new_n4891_1, new_n4868, new_n4892);
nor_5  g02544(new_n4892, new_n4867, new_n4893);
nor_5  g02545(new_n4893, new_n4866, new_n4894);
xnor_4 g02546(new_n4894, new_n4865, new_n4895);
xnor_4 g02547(n10763, n5696, new_n4896);
nor_5  g02548(n13367, n7437, new_n4897);
xnor_4 g02549(n13367, n7437, new_n4898);
nor_5  g02550(n20700, n932, new_n4899);
xnor_4 g02551(n20700, n932, new_n4900);
nor_5  g02552(n7099, n6691, new_n4901);
xnor_4 g02553(n7099, n6691, new_n4902);
nor_5  g02554(n12811, n3260, new_n4903);
xnor_4 g02555(n12811, n3260, new_n4904);
nor_5  g02556(n20489, n1118, new_n4905);
xnor_4 g02557(n20489, n1118, new_n4906);
nor_5  g02558(n25974, n2355, new_n4907);
xnor_4 g02559(n25974, n2355, new_n4908);
nor_5  g02560(n11121, n1630, new_n4909);
and_5  g02561(n16217, n1451, new_n4910);
xnor_4 g02562(n11121, n1630, new_n4911);
nor_5  g02563(new_n4911, new_n4910, new_n4912);
nor_5  g02564(new_n4912, new_n4909, new_n4913_1);
nor_5  g02565(new_n4913_1, new_n4908, new_n4914);
nor_5  g02566(new_n4914, new_n4907, new_n4915);
nor_5  g02567(new_n4915, new_n4906, new_n4916);
nor_5  g02568(new_n4916, new_n4905, new_n4917);
nor_5  g02569(new_n4917, new_n4904, new_n4918);
nor_5  g02570(new_n4918, new_n4903, new_n4919);
nor_5  g02571(new_n4919, new_n4902, new_n4920);
nor_5  g02572(new_n4920, new_n4901, new_n4921);
nor_5  g02573(new_n4921, new_n4900, new_n4922);
nor_5  g02574(new_n4922, new_n4899, new_n4923);
nor_5  g02575(new_n4923, new_n4898, new_n4924);
nor_5  g02576(new_n4924, new_n4897, new_n4925_1);
xor_4  g02577(new_n4925_1, new_n4896, new_n4926);
xnor_4 g02578(new_n4926, new_n4895, new_n4927);
xor_4  g02579(new_n4923, new_n4898, new_n4928);
xnor_4 g02580(new_n4892, new_n4867, new_n4929);
nor_5  g02581(new_n4929, new_n4928, new_n4930);
xnor_4 g02582(new_n4929, new_n4928, new_n4931);
xnor_4 g02583(new_n4921, new_n4900, new_n4932);
xor_4  g02584(new_n4890, new_n4869, new_n4933);
nor_5  g02585(new_n4933, new_n4932, new_n4934);
xnor_4 g02586(new_n4933, new_n4932, new_n4935);
xnor_4 g02587(new_n4919, new_n4902, new_n4936);
xor_4  g02588(new_n4888, new_n4871, new_n4937);
or_5   g02589(new_n4937, new_n4936, new_n4938);
xnor_4 g02590(new_n4915, new_n4906, new_n4939_1);
xor_4  g02591(new_n4884, new_n4875, new_n4940);
nor_5  g02592(new_n4940, new_n4939_1, new_n4941);
xnor_4 g02593(new_n4940, new_n4939_1, new_n4942);
xnor_4 g02594(new_n4913_1, new_n4908, new_n4943);
xor_4  g02595(new_n4882, new_n4877, new_n4944);
nor_5  g02596(new_n4944, new_n4943, new_n4945);
xor_4  g02597(new_n4880, new_n4879, new_n4946);
not_10 g02598(new_n4946, new_n4947_1);
xor_4  g02599(new_n4911, new_n4910, new_n4948);
and_5  g02600(new_n4948, new_n4947_1, new_n4949);
xnor_4 g02601(n12315, n5438, new_n4950);
xor_4  g02602(n16217, n1451, new_n4951);
nor_5  g02603(new_n4951, new_n4950, new_n4952_1);
xnor_4 g02604(new_n4948, new_n4946, new_n4953);
and_5  g02605(new_n4953, new_n4952_1, new_n4954);
nor_5  g02606(new_n4954, new_n4949, new_n4955);
xnor_4 g02607(new_n4944, new_n4943, new_n4956);
nor_5  g02608(new_n4956, new_n4955, new_n4957_1);
nor_5  g02609(new_n4957_1, new_n4945, new_n4958);
nor_5  g02610(new_n4958, new_n4942, new_n4959);
nor_5  g02611(new_n4959, new_n4941, new_n4960);
xnor_4 g02612(new_n4917, new_n4904, new_n4961);
and_5  g02613(new_n4961, new_n4960, new_n4962);
xnor_4 g02614(new_n4961, new_n4960, new_n4963);
xnor_4 g02615(new_n4886, new_n4873, new_n4964_1);
nor_5  g02616(new_n4964_1, new_n4963, new_n4965);
nor_5  g02617(new_n4965, new_n4962, new_n4966_1);
not_10 g02618(new_n4966_1, new_n4967_1);
xnor_4 g02619(new_n4937, new_n4936, new_n4968);
or_5   g02620(new_n4968, new_n4967_1, new_n4969);
and_5  g02621(new_n4969, new_n4938, new_n4970);
nor_5  g02622(new_n4970, new_n4935, new_n4971);
or_5   g02623(new_n4971, new_n4934, new_n4972_1);
nor_5  g02624(new_n4972_1, new_n4931, new_n4973);
nor_5  g02625(new_n4973, new_n4930, new_n4974);
xor_4  g02626(new_n4974, new_n4927, new_n4975);
xnor_4 g02627(new_n4975, new_n4864, new_n4976);
xnor_4 g02628(new_n4861, new_n4830, new_n4977);
xor_4  g02629(new_n4972_1, new_n4931, new_n4978);
nor_5  g02630(new_n4978, new_n4977, new_n4979);
xnor_4 g02631(new_n4978, new_n4977, new_n4980);
xor_4  g02632(new_n4859, new_n4833, new_n4981);
xor_4  g02633(new_n4970, new_n4935, new_n4982);
and_5  g02634(new_n4982, new_n4981, new_n4983);
xnor_4 g02635(new_n4982, new_n4981, new_n4984);
xor_4  g02636(new_n4857, new_n4836, new_n4985);
xnor_4 g02637(new_n4968, new_n4966_1, new_n4986);
and_5  g02638(new_n4986, new_n4985, new_n4987);
xnor_4 g02639(new_n4986, new_n4985, new_n4988);
xnor_4 g02640(new_n4855, new_n4839, new_n4989);
xor_4  g02641(new_n4964_1, new_n4963, new_n4990);
nor_5  g02642(new_n4990, new_n4989, new_n4991);
xnor_4 g02643(new_n4990, new_n4989, new_n4992);
xor_4  g02644(new_n4958, new_n4942, new_n4993);
xor_4  g02645(new_n4853, new_n4852, new_n4994);
and_5  g02646(new_n4994, new_n4993, new_n4995);
xor_4  g02647(new_n4994, new_n4993, new_n4996);
xor_4  g02648(new_n4850_1, new_n4844, new_n4997);
xor_4  g02649(new_n4956, new_n4955, new_n4998);
nor_5  g02650(new_n4998, new_n4997, new_n4999);
xnor_4 g02651(new_n4998, new_n4997, new_n5000);
xor_4  g02652(new_n4953, new_n4952_1, new_n5001);
not_10 g02653(new_n5001, new_n5002);
nor_5  g02654(new_n5002, new_n4848, new_n5003);
xor_4  g02655(new_n4848, new_n4847, new_n5004);
or_5   g02656(new_n5004, new_n5001, new_n5005);
xnor_4 g02657(n23333, n11424, new_n5006);
xor_4  g02658(new_n4951, new_n4950, new_n5007);
or_5   g02659(new_n5007, new_n5006, new_n5008);
and_5  g02660(new_n5008, new_n5005, new_n5009);
or_5   g02661(new_n5009, new_n5003, new_n5010);
nor_5  g02662(new_n5010, new_n5000, new_n5011_1);
nor_5  g02663(new_n5011_1, new_n4999, new_n5012);
and_5  g02664(new_n5012, new_n4996, new_n5013);
nor_5  g02665(new_n5013, new_n4995, new_n5014);
nor_5  g02666(new_n5014, new_n4992, new_n5015);
nor_5  g02667(new_n5015, new_n4991, new_n5016);
nor_5  g02668(new_n5016, new_n4988, new_n5017);
nor_5  g02669(new_n5017, new_n4987, new_n5018);
nor_5  g02670(new_n5018, new_n4984, new_n5019);
nor_5  g02671(new_n5019, new_n4983, new_n5020_1);
nor_5  g02672(new_n5020_1, new_n4980, new_n5021);
or_5   g02673(new_n5021, new_n4979, new_n5022);
xor_4  g02674(new_n5022, new_n4976, n431);
not_10 g02675(n23895, new_n5024_1);
nor_5  g02676(new_n5024_1, n8614, new_n5025_1);
xor_4  g02677(n23895, n8614, new_n5026_1);
not_10 g02678(n17351, new_n5027);
nor_5  g02679(new_n5027, n15182, new_n5028);
xor_4  g02680(n17351, n15182, new_n5029);
not_10 g02681(n11736, new_n5030);
nor_5  g02682(n27037, new_n5030, new_n5031_1);
xor_4  g02683(n27037, n11736, new_n5032);
not_10 g02684(n23200, new_n5033);
nor_5  g02685(new_n5033, n8964, new_n5034);
xor_4  g02686(n23200, n8964, new_n5035);
not_10 g02687(n17959, new_n5036);
nor_5  g02688(n20151, new_n5036, new_n5037);
xor_4  g02689(n20151, n17959, new_n5038);
not_10 g02690(n7566, new_n5039);
nor_5  g02691(n7693, new_n5039, new_n5040);
xor_4  g02692(n7693, n7566, new_n5041);
not_10 g02693(n7731, new_n5042);
nor_5  g02694(n10405, new_n5042, new_n5043);
xor_4  g02695(n10405, n7731, new_n5044);
not_10 g02696(n12341, new_n5045);
and_5  g02697(new_n5045, n11302, new_n5046_1);
nor_5  g02698(new_n5045, n11302, new_n5047);
not_10 g02699(n20986, new_n5048);
and_5  g02700(new_n5048, n17090, new_n5049);
or_5   g02701(new_n5048, n17090, new_n5050);
not_10 g02702(n6773, new_n5051);
nor_5  g02703(n12384, new_n5051, new_n5052);
and_5  g02704(new_n5052, new_n5050, new_n5053);
nor_5  g02705(new_n5053, new_n5049, new_n5054);
nor_5  g02706(new_n5054, new_n5047, new_n5055);
or_5   g02707(new_n5055, new_n5046_1, new_n5056);
nor_5  g02708(new_n5056, new_n5044, new_n5057);
nor_5  g02709(new_n5057, new_n5043, new_n5058);
nor_5  g02710(new_n5058, new_n5041, new_n5059);
nor_5  g02711(new_n5059, new_n5040, new_n5060_1);
nor_5  g02712(new_n5060_1, new_n5038, new_n5061);
nor_5  g02713(new_n5061, new_n5037, new_n5062_1);
nor_5  g02714(new_n5062_1, new_n5035, new_n5063);
nor_5  g02715(new_n5063, new_n5034, new_n5064_1);
nor_5  g02716(new_n5064_1, new_n5032, new_n5065);
nor_5  g02717(new_n5065, new_n5031_1, new_n5066);
nor_5  g02718(new_n5066, new_n5029, new_n5067);
nor_5  g02719(new_n5067, new_n5028, new_n5068);
nor_5  g02720(new_n5068, new_n5026_1, new_n5069);
nor_5  g02721(new_n5069, new_n5025_1, new_n5070);
not_10 g02722(n13494, new_n5071);
nor_5  g02723(n18880, new_n5071, new_n5072);
xor_4  g02724(n18880, n13494, new_n5073);
not_10 g02725(n25345, new_n5074);
nor_5  g02726(n25475, new_n5074, new_n5075);
xor_4  g02727(n25475, n25345, new_n5076);
not_10 g02728(n9655, new_n5077_1);
nor_5  g02729(n23849, new_n5077_1, new_n5078);
xor_4  g02730(n23849, n9655, new_n5079);
not_10 g02731(n13490, new_n5080);
nor_5  g02732(new_n5080, n12446, new_n5081);
xor_4  g02733(n13490, n12446, new_n5082_1);
not_10 g02734(n22660, new_n5083);
nor_5  g02735(new_n5083, n11011, new_n5084);
xor_4  g02736(n22660, n11011, new_n5085);
not_10 g02737(n1777, new_n5086);
nor_5  g02738(n16029, new_n5086, new_n5087);
xor_4  g02739(n16029, n1777, new_n5088);
not_10 g02740(n8745, new_n5089);
nor_5  g02741(n16476, new_n5089, new_n5090);
xor_4  g02742(n16476, n8745, new_n5091);
not_10 g02743(n15636, new_n5092);
and_5  g02744(new_n5092, n11615, new_n5093);
nor_5  g02745(new_n5092, n11615, new_n5094);
nor_5  g02746(new_n3712, n20077, new_n5095);
not_10 g02747(n20077, new_n5096);
or_5   g02748(n22433, new_n5096, new_n5097);
not_10 g02749(n6794, new_n5098_1);
and_5  g02750(n14090, new_n5098_1, new_n5099);
and_5  g02751(new_n5099, new_n5097, new_n5100);
nor_5  g02752(new_n5100, new_n5095, new_n5101_1);
nor_5  g02753(new_n5101_1, new_n5094, new_n5102);
or_5   g02754(new_n5102, new_n5093, new_n5103);
nor_5  g02755(new_n5103, new_n5091, new_n5104);
nor_5  g02756(new_n5104, new_n5090, new_n5105);
nor_5  g02757(new_n5105, new_n5088, new_n5106);
nor_5  g02758(new_n5106, new_n5087, new_n5107);
nor_5  g02759(new_n5107, new_n5085, new_n5108);
nor_5  g02760(new_n5108, new_n5084, new_n5109);
nor_5  g02761(new_n5109, new_n5082_1, new_n5110);
nor_5  g02762(new_n5110, new_n5081, new_n5111);
nor_5  g02763(new_n5111, new_n5079, new_n5112);
nor_5  g02764(new_n5112, new_n5078, new_n5113);
nor_5  g02765(new_n5113, new_n5076, new_n5114);
nor_5  g02766(new_n5114, new_n5075, new_n5115_1);
nor_5  g02767(new_n5115_1, new_n5073, new_n5116);
or_5   g02768(new_n5116, new_n5072, new_n5117);
xor_4  g02769(new_n5115_1, new_n5073, new_n5118);
or_5   g02770(n22173, n583, new_n5119);
or_5   g02771(new_n5119, n2146, new_n5120_1);
or_5   g02772(new_n5120_1, n23974, new_n5121);
or_5   g02773(new_n5121, n3909, new_n5122);
or_5   g02774(new_n5122, n20429, new_n5123);
or_5   g02775(new_n5123, n22554, new_n5124);
or_5   g02776(new_n5124, n23913, new_n5125);
xor_4  g02777(new_n5125, n26797, new_n5126);
nor_5  g02778(new_n5126, n10201, new_n5127);
xnor_4 g02779(new_n5126, n10201, new_n5128_1);
xor_4  g02780(new_n5124, n23913, new_n5129);
nor_5  g02781(new_n5129, n10593, new_n5130);
xnor_4 g02782(new_n5129, n10593, new_n5131_1);
xor_4  g02783(new_n5123, n22554, new_n5132);
nor_5  g02784(new_n5132, n18290, new_n5133);
xnor_4 g02785(new_n5132, n18290, new_n5134);
xor_4  g02786(new_n5122, n20429, new_n5135);
nor_5  g02787(new_n5135, n11580, new_n5136);
xnor_4 g02788(new_n5135, n11580, new_n5137);
xor_4  g02789(new_n5121, n3909, new_n5138);
nor_5  g02790(new_n5138, n15884, new_n5139);
xnor_4 g02791(new_n5138, n15884, new_n5140_1);
xor_4  g02792(new_n5120_1, n23974, new_n5141);
nor_5  g02793(new_n5141, n6356, new_n5142);
xor_4  g02794(new_n5119, n2146, new_n5143);
nor_5  g02795(new_n5143, n27104, new_n5144);
xnor_4 g02796(new_n5143, n27104, new_n5145);
not_10 g02797(n27188, new_n5146);
xnor_4 g02798(n22173, n583, new_n5147);
and_5  g02799(new_n5147, new_n5146, new_n5148);
nand_5 g02800(n6611, n583, new_n5149);
xnor_4 g02801(new_n5147, n27188, new_n5150);
and_5  g02802(new_n5150, new_n5149, new_n5151);
nor_5  g02803(new_n5151, new_n5148, new_n5152);
nor_5  g02804(new_n5152, new_n5145, new_n5153);
nor_5  g02805(new_n5153, new_n5144, new_n5154);
xnor_4 g02806(new_n5141, n6356, new_n5155);
nor_5  g02807(new_n5155, new_n5154, new_n5156);
nor_5  g02808(new_n5156, new_n5142, new_n5157);
nor_5  g02809(new_n5157, new_n5140_1, new_n5158_1);
nor_5  g02810(new_n5158_1, new_n5139, new_n5159);
nor_5  g02811(new_n5159, new_n5137, new_n5160);
nor_5  g02812(new_n5160, new_n5136, new_n5161);
nor_5  g02813(new_n5161, new_n5134, new_n5162);
nor_5  g02814(new_n5162, new_n5133, new_n5163);
nor_5  g02815(new_n5163, new_n5131_1, new_n5164);
nor_5  g02816(new_n5164, new_n5130, new_n5165);
nor_5  g02817(new_n5165, new_n5128_1, new_n5166);
or_5   g02818(new_n5166, new_n5127, new_n5167);
nor_5  g02819(new_n5125, n26797, new_n5168_1);
xnor_4 g02820(new_n5168_1, n12702, new_n5169);
xor_4  g02821(new_n5169, n12650, new_n5170);
xnor_4 g02822(new_n5170, new_n5167, new_n5171);
nor_5  g02823(new_n5171, new_n5118, new_n5172);
xnor_4 g02824(new_n5171, new_n5118, new_n5173);
xor_4  g02825(new_n5113, new_n5076, new_n5174);
xnor_4 g02826(new_n5165, new_n5128_1, new_n5175);
nor_5  g02827(new_n5175, new_n5174, new_n5176);
xnor_4 g02828(new_n5175, new_n5174, new_n5177);
xor_4  g02829(new_n5111, new_n5079, new_n5178);
xnor_4 g02830(new_n5163, new_n5131_1, new_n5179);
nor_5  g02831(new_n5179, new_n5178, new_n5180);
xnor_4 g02832(new_n5179, new_n5178, new_n5181);
xor_4  g02833(new_n5109, new_n5082_1, new_n5182);
not_10 g02834(new_n5182, new_n5183);
xor_4  g02835(new_n5161, new_n5134, new_n5184_1);
and_5  g02836(new_n5184_1, new_n5183, new_n5185);
xor_4  g02837(new_n5184_1, new_n5182, new_n5186);
xor_4  g02838(new_n5107, new_n5085, new_n5187);
xnor_4 g02839(new_n5159, new_n5137, new_n5188);
nor_5  g02840(new_n5188, new_n5187, new_n5189);
xnor_4 g02841(new_n5188, new_n5187, new_n5190);
xor_4  g02842(new_n5105, new_n5088, new_n5191);
not_10 g02843(new_n5191, new_n5192);
xor_4  g02844(new_n5157, new_n5140_1, new_n5193);
and_5  g02845(new_n5193, new_n5192, new_n5194);
xor_4  g02846(new_n5193, new_n5191, new_n5195);
xor_4  g02847(new_n5103, new_n5091, new_n5196);
xnor_4 g02848(new_n5155, new_n5154, new_n5197);
nor_5  g02849(new_n5197, new_n5196, new_n5198);
xor_4  g02850(new_n5197, new_n5196, new_n5199);
xor_4  g02851(new_n5152, new_n5145, new_n5200);
xnor_4 g02852(n15636, n11615, new_n5201);
xnor_4 g02853(new_n5201, new_n5101_1, new_n5202);
nor_5  g02854(new_n5202, new_n5200, new_n5203);
xnor_4 g02855(new_n5202, new_n5200, new_n5204);
xor_4  g02856(new_n5150, new_n5149, new_n5205);
xor_4  g02857(n22433, n20077, new_n5206);
xnor_4 g02858(new_n5206, new_n5099, new_n5207);
nor_5  g02859(new_n5207, new_n5205, new_n5208);
xnor_4 g02860(n14090, n6794, new_n5209);
xnor_4 g02861(n6611, n583, new_n5210);
nor_5  g02862(new_n5210, new_n5209, new_n5211_1);
xor_4  g02863(new_n5207, new_n5205, new_n5212);
and_5  g02864(new_n5212, new_n5211_1, new_n5213_1);
nor_5  g02865(new_n5213_1, new_n5208, new_n5214);
nor_5  g02866(new_n5214, new_n5204, new_n5215);
nor_5  g02867(new_n5215, new_n5203, new_n5216);
and_5  g02868(new_n5216, new_n5199, new_n5217);
nor_5  g02869(new_n5217, new_n5198, new_n5218);
nor_5  g02870(new_n5218, new_n5195, new_n5219);
nor_5  g02871(new_n5219, new_n5194, new_n5220);
nor_5  g02872(new_n5220, new_n5190, new_n5221);
nor_5  g02873(new_n5221, new_n5189, new_n5222);
nor_5  g02874(new_n5222, new_n5186, new_n5223);
nor_5  g02875(new_n5223, new_n5185, new_n5224);
nor_5  g02876(new_n5224, new_n5181, new_n5225);
nor_5  g02877(new_n5225, new_n5180, new_n5226_1);
nor_5  g02878(new_n5226_1, new_n5177, new_n5227);
nor_5  g02879(new_n5227, new_n5176, new_n5228_1);
nor_5  g02880(new_n5228_1, new_n5173, new_n5229);
or_5   g02881(new_n5229, new_n5172, new_n5230);
not_10 g02882(n12702, new_n5231);
and_5  g02883(new_n5168_1, new_n5231, new_n5232);
and_5  g02884(new_n5169, n12650, new_n5233);
nor_5  g02885(new_n5169, n12650, new_n5234);
nor_5  g02886(new_n5234, new_n5167, new_n5235);
or_5   g02887(new_n5235, new_n5233, new_n5236);
nor_5  g02888(new_n5236, new_n5232, new_n5237);
or_5   g02889(new_n5237, new_n5230, new_n5238);
nor_5  g02890(new_n5238, new_n5117, new_n5239);
and_5  g02891(new_n5237, new_n5230, new_n5240);
and_5  g02892(new_n5240, new_n5117, new_n5241);
nor_5  g02893(new_n5241, new_n5239, new_n5242);
xnor_4 g02894(new_n5242, new_n5070, new_n5243);
xnor_4 g02895(new_n5237, new_n5230, new_n5244);
xnor_4 g02896(new_n5244, new_n5117, new_n5245);
and_5  g02897(new_n5245, new_n5070, new_n5246);
nor_5  g02898(new_n5245, new_n5070, new_n5247);
xnor_4 g02899(new_n5068, new_n5026_1, new_n5248);
xor_4  g02900(new_n5228_1, new_n5173, new_n5249);
and_5  g02901(new_n5249, new_n5248, new_n5250);
xnor_4 g02902(new_n5249, new_n5248, new_n5251);
xnor_4 g02903(new_n5066, new_n5029, new_n5252);
xor_4  g02904(new_n5226_1, new_n5177, new_n5253);
and_5  g02905(new_n5253, new_n5252, new_n5254);
xnor_4 g02906(new_n5253, new_n5252, new_n5255_1);
xnor_4 g02907(new_n5064_1, new_n5032, new_n5256_1);
xor_4  g02908(new_n5224, new_n5181, new_n5257);
and_5  g02909(new_n5257, new_n5256_1, new_n5258);
xnor_4 g02910(new_n5257, new_n5256_1, new_n5259);
xnor_4 g02911(new_n5062_1, new_n5035, new_n5260);
xor_4  g02912(new_n5222, new_n5186, new_n5261);
and_5  g02913(new_n5261, new_n5260, new_n5262);
xnor_4 g02914(new_n5261, new_n5260, new_n5263);
xnor_4 g02915(new_n5060_1, new_n5038, new_n5264);
xor_4  g02916(new_n5220, new_n5190, new_n5265_1);
and_5  g02917(new_n5265_1, new_n5264, new_n5266);
xnor_4 g02918(new_n5265_1, new_n5264, new_n5267);
xnor_4 g02919(new_n5058, new_n5041, new_n5268);
xor_4  g02920(new_n5218, new_n5195, new_n5269);
and_5  g02921(new_n5269, new_n5268, new_n5270);
xnor_4 g02922(new_n5269, new_n5268, new_n5271);
xnor_4 g02923(new_n5216, new_n5199, new_n5272);
xor_4  g02924(new_n5056, new_n5044, new_n5273_1);
nor_5  g02925(new_n5273_1, new_n5272, new_n5274_1);
xnor_4 g02926(new_n5273_1, new_n5272, new_n5275);
xnor_4 g02927(new_n5214, new_n5204, new_n5276);
xnor_4 g02928(n12341, n11302, new_n5277);
xnor_4 g02929(new_n5277, new_n5054, new_n5278);
and_5  g02930(new_n5278, new_n5276, new_n5279);
xnor_4 g02931(new_n5278, new_n5276, new_n5280);
xnor_4 g02932(new_n5210, new_n5209, new_n5281);
xnor_4 g02933(n12384, n6773, new_n5282);
or_5   g02934(new_n5282, new_n5281, new_n5283);
xor_4  g02935(n20986, n17090, new_n5284);
xnor_4 g02936(new_n5284, new_n5052, new_n5285);
and_5  g02937(new_n5285, new_n5283, new_n5286);
xnor_4 g02938(new_n5212, new_n5211_1, new_n5287);
xor_4  g02939(new_n5285, new_n5283, new_n5288);
and_5  g02940(new_n5288, new_n5287, new_n5289);
nor_5  g02941(new_n5289, new_n5286, new_n5290);
nor_5  g02942(new_n5290, new_n5280, new_n5291);
nor_5  g02943(new_n5291, new_n5279, new_n5292);
nor_5  g02944(new_n5292, new_n5275, new_n5293);
nor_5  g02945(new_n5293, new_n5274_1, new_n5294);
nor_5  g02946(new_n5294, new_n5271, new_n5295);
nor_5  g02947(new_n5295, new_n5270, new_n5296);
nor_5  g02948(new_n5296, new_n5267, new_n5297);
nor_5  g02949(new_n5297, new_n5266, new_n5298);
nor_5  g02950(new_n5298, new_n5263, new_n5299);
nor_5  g02951(new_n5299, new_n5262, new_n5300_1);
nor_5  g02952(new_n5300_1, new_n5259, new_n5301);
nor_5  g02953(new_n5301, new_n5258, new_n5302_1);
nor_5  g02954(new_n5302_1, new_n5255_1, new_n5303);
nor_5  g02955(new_n5303, new_n5254, new_n5304);
nor_5  g02956(new_n5304, new_n5251, new_n5305);
or_5   g02957(new_n5305, new_n5250, new_n5306);
nor_5  g02958(new_n5306, new_n5247, new_n5307);
nor_5  g02959(new_n5307, new_n5246, new_n5308);
xnor_4 g02960(new_n5308, new_n5243, n457);
xnor_4 g02961(n24323, n1681, new_n5310);
xnor_4 g02962(n13781, n2088, new_n5311);
xnor_4 g02963(new_n5311, new_n5310, new_n5312);
nor_5  g02964(new_n5312, new_n5209, new_n5313);
xor_4  g02965(new_n5313, new_n5207, new_n5314);
or_5   g02966(new_n5311, new_n5310, new_n5315);
nor_5  g02967(n24323, new_n4084, new_n5316);
xnor_4 g02968(n26443, n25877, new_n5317);
xor_4  g02969(new_n5317, new_n5316, new_n5318);
xnor_4 g02970(new_n5318, new_n5315, new_n5319);
xor_4  g02971(n9399, n2088, new_n5320);
and_5  g02972(n13781, n2088, new_n5321);
nor_5  g02973(new_n5321, n11486, new_n5322);
and_5  g02974(n13781, n11486, new_n5323);
and_5  g02975(new_n5323, n2088, new_n5324);
or_5   g02976(new_n5324, new_n5322, new_n5325_1);
xor_4  g02977(new_n5325_1, new_n5320, new_n5326);
xor_4  g02978(new_n5326, new_n5319, new_n5327);
xnor_4 g02979(new_n5327, new_n5314, n463);
xor_4  g02980(n12121, n6775, new_n5329);
xor_4  g02981(new_n5329, n8920, new_n5330_1);
xnor_4 g02982(new_n2898, n5438, new_n5331);
xnor_4 g02983(new_n5331, new_n5330_1, n491);
xnor_4 g02984(new_n5292, new_n5275, n496);
xnor_4 g02985(n25926, n12384, new_n5334);
xor_4  g02986(new_n5334, n6773, new_n5335);
xor_4  g02987(new_n5209, n16167, new_n5336);
or_5   g02988(new_n5336, new_n5335, new_n5337_1);
not_10 g02989(n16167, new_n5338);
nor_5  g02990(new_n5209, new_n5338, new_n5339);
xnor_4 g02991(new_n5207, n18745, new_n5340);
xnor_4 g02992(new_n5340, new_n5339, new_n5341);
and_5  g02993(n25926, n12384, new_n5342);
xor_4  g02994(n25926, n7657, new_n5343);
xor_4  g02995(new_n5343, n20986, new_n5344);
xor_4  g02996(new_n5344, new_n5342, new_n5345);
or_5   g02997(new_n5334, new_n5051, new_n5346);
nor_5  g02998(new_n5346, n17090, new_n5347);
nor_5  g02999(n17090, n6773, new_n5348);
and_5  g03000(n17090, n6773, new_n5349);
and_5  g03001(new_n5349, new_n5334, new_n5350);
or_5   g03002(new_n5350, new_n5348, new_n5351_1);
or_5   g03003(new_n5351_1, new_n5347, new_n5352);
xor_4  g03004(new_n5352, new_n5345, new_n5353_1);
xor_4  g03005(new_n5353_1, new_n5341, new_n5354);
xnor_4 g03006(new_n5354, new_n5337_1, n498);
xnor_4 g03007(n25872, n19618, new_n5356);
nor_5  g03008(n22043, n20259, new_n5357);
and_5  g03009(n12121, n3925, new_n5358);
xnor_4 g03010(n22043, n20259, new_n5359);
nor_5  g03011(new_n5359, new_n5358, new_n5360);
nor_5  g03012(new_n5360, new_n5357, new_n5361);
xor_4  g03013(new_n5361, new_n5356, new_n5362);
xor_4  g03014(new_n5362, new_n4503, new_n5363);
xor_4  g03015(new_n5359, new_n5358, new_n5364);
nor_5  g03016(new_n5364, new_n4506, new_n5365);
xor_4  g03017(n12121, n3925, new_n5366);
or_5   g03018(new_n5366, new_n4508, new_n5367);
xor_4  g03019(new_n5364, new_n4506, new_n5368);
and_5  g03020(new_n5368, new_n5367, new_n5369);
nor_5  g03021(new_n5369, new_n5365, new_n5370);
xor_4  g03022(new_n5370, new_n5363, new_n5371);
xnor_4 g03023(new_n5371, new_n3564, new_n5372);
xor_4  g03024(new_n5368, new_n5367, new_n5373);
nor_5  g03025(new_n5373, new_n3539, new_n5374);
not_10 g03026(new_n5373, new_n5375);
or_5   g03027(new_n5375, new_n3568, new_n5376_1);
xnor_4 g03028(new_n5366, new_n4508, new_n5377);
nand_5 g03029(new_n5377, new_n3570_1, new_n5378);
and_5  g03030(new_n5378, new_n5376_1, new_n5379);
or_5   g03031(new_n5379, new_n5374, new_n5380);
xor_4  g03032(new_n5380, new_n5372, n521);
xor_4  g03033(new_n5282, new_n5281, n548);
xor_4  g03034(new_n4002, new_n3985, n554);
not_10 g03035(n2979, new_n5384);
not_10 g03036(n647, new_n5385);
not_10 g03037(n7524, new_n5386_1);
nor_5  g03038(n20658, n15743, new_n5387);
nand_5 g03039(new_n5387, new_n5386_1, new_n5388);
or_5   g03040(new_n5388, n4957, new_n5389);
or_5   g03041(new_n5389, n9003, new_n5390);
or_5   g03042(new_n5390, n3161, new_n5391);
or_5   g03043(new_n5391, n25749, new_n5392);
nor_5  g03044(new_n5392, n20409, new_n5393);
nand_5 g03045(new_n5393, new_n5385, new_n5394);
xnor_4 g03046(new_n5394, new_n5384, new_n5395);
xnor_4 g03047(n9259, n6456, new_n5396);
nor_5  g03048(n21489, n4085, new_n5397);
xnor_4 g03049(n21489, n4085, new_n5398);
nor_5  g03050(n26725, n20213, new_n5399_1);
xnor_4 g03051(n26725, n20213, new_n5400_1);
nor_5  g03052(n13912, n11980, new_n5401);
xnor_4 g03053(n13912, n11980, new_n5402);
nor_5  g03054(n7670, n3253, new_n5403_1);
xnor_4 g03055(n7670, n3253, new_n5404);
nor_5  g03056(n9598, n7759, new_n5405);
xnor_4 g03057(n9598, n7759, new_n5406);
nor_5  g03058(n22290, n12562, new_n5407);
xnor_4 g03059(n22290, n12562, new_n5408);
nor_5  g03060(n11273, n7949, new_n5409);
xnor_4 g03061(n11273, n7949, new_n5410);
nor_5  g03062(n25565, n24374, new_n5411);
and_5  g03063(n21993, n14575, new_n5412);
xnor_4 g03064(n25565, n24374, new_n5413);
nor_5  g03065(new_n5413, new_n5412, new_n5414);
nor_5  g03066(new_n5414, new_n5411, new_n5415);
nor_5  g03067(new_n5415, new_n5410, new_n5416);
nor_5  g03068(new_n5416, new_n5409, new_n5417);
nor_5  g03069(new_n5417, new_n5408, new_n5418);
nor_5  g03070(new_n5418, new_n5407, new_n5419);
nor_5  g03071(new_n5419, new_n5406, new_n5420);
nor_5  g03072(new_n5420, new_n5405, new_n5421);
nor_5  g03073(new_n5421, new_n5404, new_n5422);
nor_5  g03074(new_n5422, new_n5403_1, new_n5423);
nor_5  g03075(new_n5423, new_n5402, new_n5424);
nor_5  g03076(new_n5424, new_n5401, new_n5425);
nor_5  g03077(new_n5425, new_n5400_1, new_n5426);
nor_5  g03078(new_n5426, new_n5399_1, new_n5427);
nor_5  g03079(new_n5427, new_n5398, new_n5428);
nor_5  g03080(new_n5428, new_n5397, new_n5429);
xor_4  g03081(new_n5429, new_n5396, new_n5430_1);
xnor_4 g03082(new_n5430_1, new_n5395, new_n5431);
xnor_4 g03083(new_n5393, n647, new_n5432);
not_10 g03084(new_n5432, new_n5433);
xnor_4 g03085(new_n5427, new_n5398, new_n5434);
nor_5  g03086(new_n5434, new_n5433, new_n5435);
xor_4  g03087(new_n5434, new_n5432, new_n5436);
not_10 g03088(n20409, new_n5437);
xnor_4 g03089(new_n5392, new_n5437, new_n5438_1);
xor_4  g03090(new_n5425, new_n5400_1, new_n5439_1);
nor_5  g03091(new_n5439_1, new_n5438_1, new_n5440);
xnor_4 g03092(new_n5439_1, new_n5438_1, new_n5441);
not_10 g03093(n25749, new_n5442);
xnor_4 g03094(new_n5391, new_n5442, new_n5443_1);
xor_4  g03095(new_n5423, new_n5402, new_n5444);
nor_5  g03096(new_n5444, new_n5443_1, new_n5445);
xnor_4 g03097(new_n5444, new_n5443_1, new_n5446);
xnor_4 g03098(new_n5390, new_n3553, new_n5447);
xor_4  g03099(new_n5421, new_n5404, new_n5448);
nor_5  g03100(new_n5448, new_n5447, new_n5449);
xnor_4 g03101(new_n5448, new_n5447, new_n5450);
not_10 g03102(n9003, new_n5451_1);
xnor_4 g03103(new_n5389, new_n5451_1, new_n5452);
xor_4  g03104(new_n5419, new_n5406, new_n5453);
nor_5  g03105(new_n5453, new_n5452, new_n5454);
xnor_4 g03106(new_n5453, new_n5452, new_n5455);
xnor_4 g03107(new_n5388, new_n3560, new_n5456);
xor_4  g03108(new_n5417, new_n5408, new_n5457);
nor_5  g03109(new_n5457, new_n5456, new_n5458);
not_10 g03110(new_n5457, new_n5459);
xnor_4 g03111(new_n5459, new_n5456, new_n5460);
xnor_4 g03112(new_n5387, n7524, new_n5461);
xor_4  g03113(new_n5415, new_n5410, new_n5462);
and_5  g03114(new_n5462, new_n5461, new_n5463);
xnor_4 g03115(new_n5462, new_n5461, new_n5464);
xor_4  g03116(n21993, n14575, new_n5465);
not_10 g03117(new_n5465, new_n5466);
nor_5  g03118(new_n5466, n20658, new_n5467);
and_5  g03119(new_n5467, new_n3567, new_n5468);
xor_4  g03120(new_n5413, new_n5412, new_n5469);
not_10 g03121(new_n5469, new_n5470);
xor_4  g03122(n20658, n15743, new_n5471);
not_10 g03123(new_n5471, new_n5472_1);
nor_5  g03124(new_n5472_1, new_n5467, new_n5473);
nor_5  g03125(new_n5473, new_n5468, new_n5474);
and_5  g03126(new_n5474, new_n5470, new_n5475);
or_5   g03127(new_n5475, new_n5468, new_n5476);
nor_5  g03128(new_n5476, new_n5464, new_n5477);
nor_5  g03129(new_n5477, new_n5463, new_n5478);
and_5  g03130(new_n5478, new_n5460, new_n5479);
nor_5  g03131(new_n5479, new_n5458, new_n5480);
nor_5  g03132(new_n5480, new_n5455, new_n5481);
nor_5  g03133(new_n5481, new_n5454, new_n5482);
nor_5  g03134(new_n5482, new_n5450, new_n5483);
nor_5  g03135(new_n5483, new_n5449, new_n5484);
nor_5  g03136(new_n5484, new_n5446, new_n5485_1);
nor_5  g03137(new_n5485_1, new_n5445, new_n5486);
nor_5  g03138(new_n5486, new_n5441, new_n5487);
or_5   g03139(new_n5487, new_n5440, new_n5488);
nor_5  g03140(new_n5488, new_n5436, new_n5489);
nor_5  g03141(new_n5489, new_n5435, new_n5490);
xor_4  g03142(new_n5490, new_n5431, new_n5491);
xnor_4 g03143(n21784, n3582, new_n5492);
nor_5  g03144(n5521, n2145, new_n5493);
xnor_4 g03145(n5521, n2145, new_n5494);
nor_5  g03146(n11926, n5031, new_n5495);
xnor_4 g03147(n11926, n5031, new_n5496);
nor_5  g03148(n11044, n4325, new_n5497);
xnor_4 g03149(n11044, n4325, new_n5498);
nor_5  g03150(n5337, n2421, new_n5499);
xnor_4 g03151(n5337, n2421, new_n5500);
nor_5  g03152(n987, n626, new_n5501);
xnor_4 g03153(n987, n626, new_n5502);
nor_5  g03154(n20478, n1204, new_n5503);
xnor_4 g03155(n20478, n1204, new_n5504);
nor_5  g03156(n26882, n19618, new_n5505);
xnor_4 g03157(n26882, n19618, new_n5506);
nor_5  g03158(n22619, n22043, new_n5507);
and_5  g03159(n12121, n6775, new_n5508);
xnor_4 g03160(n22619, n22043, new_n5509);
nor_5  g03161(new_n5509, new_n5508, new_n5510);
nor_5  g03162(new_n5510, new_n5507, new_n5511);
nor_5  g03163(new_n5511, new_n5506, new_n5512);
nor_5  g03164(new_n5512, new_n5505, new_n5513);
nor_5  g03165(new_n5513, new_n5504, new_n5514);
nor_5  g03166(new_n5514, new_n5503, new_n5515);
nor_5  g03167(new_n5515, new_n5502, new_n5516);
nor_5  g03168(new_n5516, new_n5501, new_n5517_1);
nor_5  g03169(new_n5517_1, new_n5500, new_n5518);
nor_5  g03170(new_n5518, new_n5499, new_n5519);
nor_5  g03171(new_n5519, new_n5498, new_n5520);
nor_5  g03172(new_n5520, new_n5497, new_n5521_1);
nor_5  g03173(new_n5521_1, new_n5496, new_n5522);
nor_5  g03174(new_n5522, new_n5495, new_n5523);
nor_5  g03175(new_n5523, new_n5494, new_n5524_1);
nor_5  g03176(new_n5524_1, new_n5493, new_n5525);
xnor_4 g03177(new_n5525, new_n5492, new_n5526);
xnor_4 g03178(new_n5526, n8526, new_n5527);
xnor_4 g03179(new_n5523, new_n5494, new_n5528);
and_5  g03180(new_n5528, n2816, new_n5529);
xnor_4 g03181(new_n5528, n2816, new_n5530);
xnor_4 g03182(new_n5521_1, new_n5496, new_n5531);
and_5  g03183(new_n5531, n20359, new_n5532_1);
xnor_4 g03184(new_n5531, n20359, new_n5533);
xnor_4 g03185(new_n5519, new_n5498, new_n5534);
and_5  g03186(new_n5534, n4409, new_n5535);
xnor_4 g03187(new_n5534, n4409, new_n5536);
xnor_4 g03188(new_n5517_1, new_n5500, new_n5537);
and_5  g03189(new_n5537, n3570, new_n5538);
xnor_4 g03190(new_n5537, n3570, new_n5539);
xnor_4 g03191(new_n5515, new_n5502, new_n5540);
and_5  g03192(new_n5540, n13668, new_n5541);
xnor_4 g03193(new_n5540, n13668, new_n5542);
xnor_4 g03194(new_n5513, new_n5504, new_n5543);
and_5  g03195(new_n5543, n21276, new_n5544);
xnor_4 g03196(new_n5543, n21276, new_n5545);
xnor_4 g03197(new_n5511, new_n5506, new_n5546);
and_5  g03198(new_n5546, n26748, new_n5547);
xor_4  g03199(new_n5509, new_n5508, new_n5548);
not_10 g03200(new_n5548, new_n5549);
nor_5  g03201(new_n5549, n10057, new_n5550);
nand_5 g03202(new_n5329, n8920, new_n5551);
xnor_4 g03203(new_n5548, n10057, new_n5552);
and_5  g03204(new_n5552, new_n5551, new_n5553);
nor_5  g03205(new_n5553, new_n5550, new_n5554);
xor_4  g03206(new_n5546, n26748, new_n5555);
and_5  g03207(new_n5555, new_n5554, new_n5556);
nor_5  g03208(new_n5556, new_n5547, new_n5557);
nor_5  g03209(new_n5557, new_n5545, new_n5558);
nor_5  g03210(new_n5558, new_n5544, new_n5559);
nor_5  g03211(new_n5559, new_n5542, new_n5560);
nor_5  g03212(new_n5560, new_n5541, new_n5561);
nor_5  g03213(new_n5561, new_n5539, new_n5562);
nor_5  g03214(new_n5562, new_n5538, new_n5563);
nor_5  g03215(new_n5563, new_n5536, new_n5564_1);
nor_5  g03216(new_n5564_1, new_n5535, new_n5565);
nor_5  g03217(new_n5565, new_n5533, new_n5566);
nor_5  g03218(new_n5566, new_n5532_1, new_n5567);
nor_5  g03219(new_n5567, new_n5530, new_n5568);
nor_5  g03220(new_n5568, new_n5529, new_n5569);
xor_4  g03221(new_n5569, new_n5527, new_n5570);
xnor_4 g03222(new_n5570, new_n5491, new_n5571);
xor_4  g03223(new_n5567, new_n5530, new_n5572);
xor_4  g03224(new_n5488, new_n5436, new_n5573);
nor_5  g03225(new_n5573, new_n5572, new_n5574);
xnor_4 g03226(new_n5573, new_n5572, new_n5575);
xnor_4 g03227(new_n5486, new_n5441, new_n5576);
xor_4  g03228(new_n5565, new_n5533, new_n5577);
nor_5  g03229(new_n5577, new_n5576, new_n5578);
xnor_4 g03230(new_n5577, new_n5576, new_n5579_1);
xnor_4 g03231(new_n5484, new_n5446, new_n5580);
xor_4  g03232(new_n5563, new_n5536, new_n5581);
nor_5  g03233(new_n5581, new_n5580, new_n5582);
xnor_4 g03234(new_n5581, new_n5580, new_n5583);
xnor_4 g03235(new_n5482, new_n5450, new_n5584);
xor_4  g03236(new_n5561, new_n5539, new_n5585);
nor_5  g03237(new_n5585, new_n5584, new_n5586);
xnor_4 g03238(new_n5585, new_n5584, new_n5587);
xnor_4 g03239(new_n5480, new_n5455, new_n5588);
xor_4  g03240(new_n5559, new_n5542, new_n5589);
nor_5  g03241(new_n5589, new_n5588, new_n5590);
xnor_4 g03242(new_n5589, new_n5588, new_n5591);
xnor_4 g03243(new_n5478, new_n5460, new_n5592);
xor_4  g03244(new_n5557, new_n5545, new_n5593_1);
nor_5  g03245(new_n5593_1, new_n5592, new_n5594);
xnor_4 g03246(new_n5593_1, new_n5592, new_n5595);
xor_4  g03247(new_n5476, new_n5464, new_n5596);
xor_4  g03248(new_n5555, new_n5554, new_n5597);
nor_5  g03249(new_n5597, new_n5596, new_n5598);
not_10 g03250(new_n5597, new_n5599);
xnor_4 g03251(new_n5599, new_n5596, new_n5600);
xor_4  g03252(new_n5552, new_n5551, new_n5601);
xnor_4 g03253(new_n5474, new_n5469, new_n5602);
nor_5  g03254(new_n5602, new_n5601, new_n5603_1);
xor_4  g03255(new_n5465, n20658, new_n5604);
nand_5 g03256(new_n5604, new_n5330_1, new_n5605_1);
xnor_4 g03257(new_n5602, new_n5601, new_n5606);
nor_5  g03258(new_n5606, new_n5605_1, new_n5607);
nor_5  g03259(new_n5607, new_n5603_1, new_n5608);
and_5  g03260(new_n5608, new_n5600, new_n5609_1);
nor_5  g03261(new_n5609_1, new_n5598, new_n5610);
nor_5  g03262(new_n5610, new_n5595, new_n5611);
nor_5  g03263(new_n5611, new_n5594, new_n5612);
nor_5  g03264(new_n5612, new_n5591, new_n5613);
nor_5  g03265(new_n5613, new_n5590, new_n5614);
nor_5  g03266(new_n5614, new_n5587, new_n5615);
nor_5  g03267(new_n5615, new_n5586, new_n5616);
nor_5  g03268(new_n5616, new_n5583, new_n5617);
nor_5  g03269(new_n5617, new_n5582, new_n5618);
nor_5  g03270(new_n5618, new_n5579_1, new_n5619);
nor_5  g03271(new_n5619, new_n5578, new_n5620);
nor_5  g03272(new_n5620, new_n5575, new_n5621);
nor_5  g03273(new_n5621, new_n5574, new_n5622);
xnor_4 g03274(new_n5622, new_n5571, n567);
nor_5  g03275(n10250, n1831, new_n5624);
xnor_4 g03276(n10250, n1831, new_n5625);
nor_5  g03277(n13137, n7674, new_n5626);
xnor_4 g03278(n13137, n7674, new_n5627);
nor_5  g03279(n18452, n6397, new_n5628);
xnor_4 g03280(n18452, n6397, new_n5629);
nor_5  g03281(n21317, n19196, new_n5630);
xnor_4 g03282(n21317, n19196, new_n5631);
nor_5  g03283(n23586, n12398, new_n5632);
xnor_4 g03284(n23586, n12398, new_n5633);
nor_5  g03285(n21226, n19789, new_n5634_1);
xnor_4 g03286(n21226, n19789, new_n5635);
nor_5  g03287(n20169, n4426, new_n5636);
xnor_4 g03288(n20169, n4426, new_n5637);
nor_5  g03289(n20036, n8285, new_n5638);
xnor_4 g03290(n20036, n8285, new_n5639);
nor_5  g03291(n11192, n6729, new_n5640);
and_5  g03292(n21687, n9380, new_n5641);
xnor_4 g03293(n11192, n6729, new_n5642);
nor_5  g03294(new_n5642, new_n5641, new_n5643_1);
nor_5  g03295(new_n5643_1, new_n5640, new_n5644);
nor_5  g03296(new_n5644, new_n5639, new_n5645);
nor_5  g03297(new_n5645, new_n5638, new_n5646);
nor_5  g03298(new_n5646, new_n5637, new_n5647);
nor_5  g03299(new_n5647, new_n5636, new_n5648);
nor_5  g03300(new_n5648, new_n5635, new_n5649);
nor_5  g03301(new_n5649, new_n5634_1, new_n5650);
nor_5  g03302(new_n5650, new_n5633, new_n5651);
nor_5  g03303(new_n5651, new_n5632, new_n5652);
nor_5  g03304(new_n5652, new_n5631, new_n5653);
nor_5  g03305(new_n5653, new_n5630, new_n5654);
nor_5  g03306(new_n5654, new_n5629, new_n5655);
nor_5  g03307(new_n5655, new_n5628, new_n5656);
nor_5  g03308(new_n5656, new_n5627, new_n5657);
nor_5  g03309(new_n5657, new_n5626, new_n5658);
nor_5  g03310(new_n5658, new_n5625, new_n5659);
nor_5  g03311(new_n5659, new_n5624, new_n5660);
or_5   g03312(new_n3762, n25694, new_n5661);
or_5   g03313(new_n5661, n13110, new_n5662);
or_5   g03314(new_n5662, n1752, new_n5663);
or_5   g03315(new_n5663, n1288, new_n5664);
xor_4  g03316(new_n5664, n3320, new_n5665);
and_5  g03317(new_n5665, n8614, new_n5666);
nor_5  g03318(new_n5664, n3320, new_n5667);
or_5   g03319(new_n5665, n8614, new_n5668);
xor_4  g03320(new_n5663, n1288, new_n5669);
nor_5  g03321(new_n5669, n15182, new_n5670);
xnor_4 g03322(new_n5669, n15182, new_n5671);
xor_4  g03323(new_n5662, n1752, new_n5672);
nor_5  g03324(new_n5672, n27037, new_n5673);
xnor_4 g03325(new_n5672, n27037, new_n5674);
xor_4  g03326(new_n5661, n13110, new_n5675);
and_5  g03327(new_n5675, n8964, new_n5676);
xnor_4 g03328(new_n5675, n8964, new_n5677);
and_5  g03329(new_n3763, n20151, new_n5678);
nor_5  g03330(new_n3785_1, new_n3764, new_n5679);
nor_5  g03331(new_n5679, new_n5678, new_n5680_1);
nor_5  g03332(new_n5680_1, new_n5677, new_n5681);
or_5   g03333(new_n5681, new_n5676, new_n5682);
nor_5  g03334(new_n5682, new_n5674, new_n5683);
nor_5  g03335(new_n5683, new_n5673, new_n5684);
nor_5  g03336(new_n5684, new_n5671, new_n5685);
nor_5  g03337(new_n5685, new_n5670, new_n5686);
and_5  g03338(new_n5686, new_n5668, new_n5687_1);
or_5   g03339(new_n5687_1, new_n5667, new_n5688);
nor_5  g03340(new_n5688, new_n5666, new_n5689);
or_5   g03341(new_n5689, new_n5660, new_n5690);
xnor_4 g03342(new_n5689, new_n5660, new_n5691);
xnor_4 g03343(new_n5658, new_n5625, new_n5692);
xnor_4 g03344(new_n5665, n8614, new_n5693);
xnor_4 g03345(new_n5693, new_n5686, new_n5694);
and_5  g03346(new_n5694, new_n5692, new_n5695);
xnor_4 g03347(new_n5684, new_n5671, new_n5696_1);
xnor_4 g03348(new_n5656, new_n5627, new_n5697);
nor_5  g03349(new_n5697, new_n5696_1, new_n5698);
xnor_4 g03350(new_n5697, new_n5696_1, new_n5699);
xnor_4 g03351(new_n5682, new_n5674, new_n5700_1);
xnor_4 g03352(new_n5654, new_n5629, new_n5701);
nor_5  g03353(new_n5701, new_n5700_1, new_n5702);
xor_4  g03354(new_n5701, new_n5700_1, new_n5703);
xnor_4 g03355(new_n5652, new_n5631, new_n5704_1);
xor_4  g03356(new_n5680_1, new_n5677, new_n5705);
and_5  g03357(new_n5705, new_n5704_1, new_n5706);
xnor_4 g03358(new_n5650, new_n5633, new_n5707);
nor_5  g03359(new_n5707, new_n3786, new_n5708);
xnor_4 g03360(new_n5707, new_n3786, new_n5709);
xnor_4 g03361(new_n5648, new_n5635, new_n5710);
xnor_4 g03362(new_n5646, new_n5637, new_n5711);
nor_5  g03363(new_n5711, new_n3792, new_n5712);
xor_4  g03364(new_n5644, new_n5639, new_n5713);
nor_5  g03365(new_n5713, new_n3796, new_n5714);
xnor_4 g03366(new_n5713, new_n3796, new_n5715);
xor_4  g03367(new_n5642, new_n5641, new_n5716);
nor_5  g03368(new_n5716, new_n3801, new_n5717);
xor_4  g03369(n21687, n9380, new_n5718);
nand_5 g03370(new_n5718, new_n2528, new_n5719);
xnor_4 g03371(new_n5716, new_n3801, new_n5720);
nor_5  g03372(new_n5720, new_n5719, new_n5721);
nor_5  g03373(new_n5721, new_n5717, new_n5722);
nor_5  g03374(new_n5722, new_n5715, new_n5723);
or_5   g03375(new_n5723, new_n5714, new_n5724);
xnor_4 g03376(new_n5711, new_n3792, new_n5725);
nor_5  g03377(new_n5725, new_n5724, new_n5726);
nor_5  g03378(new_n5726, new_n5712, new_n5727);
nor_5  g03379(new_n5727, new_n5710, new_n5728);
not_10 g03380(new_n3789, new_n5729);
xor_4  g03381(new_n5727, new_n5710, new_n5730);
and_5  g03382(new_n5730, new_n5729, new_n5731);
nor_5  g03383(new_n5731, new_n5728, new_n5732_1);
nor_5  g03384(new_n5732_1, new_n5709, new_n5733);
or_5   g03385(new_n5733, new_n5708, new_n5734);
xnor_4 g03386(new_n5705, new_n5704_1, new_n5735);
nor_5  g03387(new_n5735, new_n5734, new_n5736);
nor_5  g03388(new_n5736, new_n5706, new_n5737);
and_5  g03389(new_n5737, new_n5703, new_n5738);
nor_5  g03390(new_n5738, new_n5702, new_n5739);
nor_5  g03391(new_n5739, new_n5699, new_n5740);
or_5   g03392(new_n5740, new_n5698, new_n5741);
xnor_4 g03393(new_n5694, new_n5692, new_n5742_1);
nor_5  g03394(new_n5742_1, new_n5741, new_n5743);
nor_5  g03395(new_n5743, new_n5695, new_n5744);
not_10 g03396(new_n5744, new_n5745);
or_5   g03397(new_n5745, new_n5691, new_n5746);
and_5  g03398(new_n5746, new_n5690, new_n5747);
xnor_4 g03399(new_n5744, new_n5691, new_n5748);
nor_5  g03400(n15766, n6105, new_n5749);
xnor_4 g03401(n15766, n6105, new_n5750);
nor_5  g03402(n25629, n3795, new_n5751);
xnor_4 g03403(n25629, n3795, new_n5752_1);
nor_5  g03404(n25464, n7692, new_n5753);
xnor_4 g03405(n25464, n7692, new_n5754);
nor_5  g03406(n23039, n4590, new_n5755);
xnor_4 g03407(n23039, n4590, new_n5756);
nor_5  g03408(n26752, n13677, new_n5757);
xnor_4 g03409(n26752, n13677, new_n5758);
nor_5  g03410(n18926, n6513, new_n5759);
xor_4  g03411(n18926, n6513, new_n5760);
and_5  g03412(n5451, n3918, new_n5761);
or_5   g03413(n5451, n3918, new_n5762);
nor_5  g03414(n5330, n919, new_n5763);
nor_5  g03415(new_n3877, new_n3872, new_n5764);
nor_5  g03416(new_n5764, new_n5763, new_n5765_1);
and_5  g03417(new_n5765_1, new_n5762, new_n5766);
nor_5  g03418(new_n5766, new_n5761, new_n5767);
and_5  g03419(new_n5767, new_n5760, new_n5768);
nor_5  g03420(new_n5768, new_n5759, new_n5769);
nor_5  g03421(new_n5769, new_n5758, new_n5770);
nor_5  g03422(new_n5770, new_n5757, new_n5771);
nor_5  g03423(new_n5771, new_n5756, new_n5772);
nor_5  g03424(new_n5772, new_n5755, new_n5773);
nor_5  g03425(new_n5773, new_n5754, new_n5774);
nor_5  g03426(new_n5774, new_n5753, new_n5775);
nor_5  g03427(new_n5775, new_n5752_1, new_n5776_1);
nor_5  g03428(new_n5776_1, new_n5751, new_n5777);
nor_5  g03429(new_n5777, new_n5750, new_n5778);
nor_5  g03430(new_n5778, new_n5749, new_n5779);
and_5  g03431(new_n5779, new_n5748, new_n5780);
xnor_4 g03432(new_n5779, new_n5748, new_n5781);
xor_4  g03433(new_n5777, new_n5750, new_n5782_1);
xor_4  g03434(new_n5742_1, new_n5741, new_n5783);
nor_5  g03435(new_n5783, new_n5782_1, new_n5784);
xnor_4 g03436(new_n5783, new_n5782_1, new_n5785);
xnor_4 g03437(new_n5739, new_n5699, new_n5786);
xor_4  g03438(new_n5775, new_n5752_1, new_n5787);
nor_5  g03439(new_n5787, new_n5786, new_n5788);
xnor_4 g03440(new_n5787, new_n5786, new_n5789);
xnor_4 g03441(new_n5737, new_n5703, new_n5790);
xor_4  g03442(new_n5773, new_n5754, new_n5791);
nor_5  g03443(new_n5791, new_n5790, new_n5792);
xnor_4 g03444(new_n5791, new_n5790, new_n5793);
xor_4  g03445(new_n5771, new_n5756, new_n5794);
xor_4  g03446(new_n5735, new_n5734, new_n5795);
nor_5  g03447(new_n5795, new_n5794, new_n5796);
xnor_4 g03448(new_n5795, new_n5794, new_n5797);
xnor_4 g03449(new_n5732_1, new_n5709, new_n5798);
xor_4  g03450(new_n5769, new_n5758, new_n5799);
nor_5  g03451(new_n5799, new_n5798, new_n5800);
xnor_4 g03452(new_n5799, new_n5798, new_n5801);
xor_4  g03453(new_n5730, new_n3789, new_n5802);
xor_4  g03454(new_n5767, new_n5760, new_n5803);
nor_5  g03455(new_n5803, new_n5802, new_n5804);
xnor_4 g03456(new_n5803, new_n5802, new_n5805);
xor_4  g03457(new_n5725, new_n5724, new_n5806);
xnor_4 g03458(n5451, n3918, new_n5807);
xnor_4 g03459(new_n5807, new_n5765_1, new_n5808);
and_5  g03460(new_n5808, new_n5806, new_n5809);
xnor_4 g03461(new_n5808, new_n5806, new_n5810);
xor_4  g03462(new_n5722, new_n5715, new_n5811);
nor_5  g03463(new_n5811, new_n3878, new_n5812);
xnor_4 g03464(new_n5811, new_n3878, new_n5813);
xor_4  g03465(new_n5720, new_n5719, new_n5814);
nor_5  g03466(new_n5814, new_n3881, new_n5815);
xor_4  g03467(new_n5718, new_n2528, new_n5816);
nor_5  g03468(new_n5816, new_n3883, new_n5817);
xor_4  g03469(new_n5814, new_n3881, new_n5818);
and_5  g03470(new_n5818, new_n5817, new_n5819);
nor_5  g03471(new_n5819, new_n5815, new_n5820);
nor_5  g03472(new_n5820, new_n5813, new_n5821);
nor_5  g03473(new_n5821, new_n5812, new_n5822_1);
nor_5  g03474(new_n5822_1, new_n5810, new_n5823);
nor_5  g03475(new_n5823, new_n5809, new_n5824);
nor_5  g03476(new_n5824, new_n5805, new_n5825);
nor_5  g03477(new_n5825, new_n5804, new_n5826);
nor_5  g03478(new_n5826, new_n5801, new_n5827);
nor_5  g03479(new_n5827, new_n5800, new_n5828);
nor_5  g03480(new_n5828, new_n5797, new_n5829);
nor_5  g03481(new_n5829, new_n5796, new_n5830);
nor_5  g03482(new_n5830, new_n5793, new_n5831);
nor_5  g03483(new_n5831, new_n5792, new_n5832);
nor_5  g03484(new_n5832, new_n5789, new_n5833_1);
nor_5  g03485(new_n5833_1, new_n5788, new_n5834_1);
nor_5  g03486(new_n5834_1, new_n5785, new_n5835);
nor_5  g03487(new_n5835, new_n5784, new_n5836);
nor_5  g03488(new_n5836, new_n5781, new_n5837);
nor_5  g03489(new_n5837, new_n5780, new_n5838);
nor_5  g03490(new_n5838, new_n5747, n588);
xor_4  g03491(n19803, n18584, new_n5840_1);
not_10 g03492(n12626, new_n5841_1);
nor_5  g03493(new_n5841_1, n4272, new_n5842_1);
nor_5  g03494(new_n4337, new_n4315, new_n5843);
nor_5  g03495(new_n5843, new_n5842_1, new_n5844);
xnor_4 g03496(new_n5844, new_n5840_1, new_n5845);
xor_4  g03497(n16911, n7773, new_n5846);
not_10 g03498(n376, new_n5847);
nor_5  g03499(n7721, new_n5847, new_n5848);
xor_4  g03500(n7721, n376, new_n5849);
not_10 g03501(n5517, new_n5850_1);
or_5   g03502(n21981, new_n5850_1, new_n5851);
xor_4  g03503(n21981, n5517, new_n5852);
not_10 g03504(n12113, new_n5853);
or_5   g03505(n12917, new_n5853, new_n5854);
xor_4  g03506(n12917, n12113, new_n5855);
not_10 g03507(n10614, new_n5856);
and_5  g03508(n21898, new_n5856, new_n5857);
nor_5  g03509(n21898, new_n5856, new_n5858);
not_10 g03510(n11266, new_n5859);
and_5  g03511(new_n5859, n9926, new_n5860);
or_5   g03512(new_n5859, n9926, new_n5861);
not_10 g03513(n22072, new_n5862);
nor_5  g03514(new_n5862, n2646, new_n5863);
and_5  g03515(new_n5863, new_n5861, new_n5864);
nor_5  g03516(new_n5864, new_n5860, new_n5865);
nor_5  g03517(new_n5865, new_n5858, new_n5866);
nor_5  g03518(new_n5866, new_n5857, new_n5867);
not_10 g03519(new_n5867, new_n5868);
or_5   g03520(new_n5868, new_n5855, new_n5869);
and_5  g03521(new_n5869, new_n5854, new_n5870);
or_5   g03522(new_n5870, new_n5852, new_n5871);
and_5  g03523(new_n5871, new_n5851, new_n5872);
nor_5  g03524(new_n5872, new_n5849, new_n5873);
nor_5  g03525(new_n5873, new_n5848, new_n5874);
xnor_4 g03526(new_n5874, new_n5846, new_n5875);
not_10 g03527(n1269, new_n5876);
not_10 g03528(n14576, new_n5877);
not_10 g03529(n5605, new_n5878);
nor_5  g03530(n15652, n4939, new_n5879);
nand_5 g03531(new_n5879, new_n5878, new_n5880);
nor_5  g03532(new_n5880, n2985, new_n5881);
and_5  g03533(new_n5881, new_n5877, new_n5882_1);
and_5  g03534(new_n5882_1, new_n5876, new_n5883);
xnor_4 g03535(new_n5883, n16818, new_n5884);
xnor_4 g03536(new_n5884, n1742, new_n5885);
xnor_4 g03537(new_n5882_1, n1269, new_n5886);
nor_5  g03538(new_n5886, n4858, new_n5887);
xnor_4 g03539(new_n5886, n4858, new_n5888);
xnor_4 g03540(new_n5881, n14576, new_n5889);
nor_5  g03541(new_n5889, n8244, new_n5890);
xnor_4 g03542(new_n5889, n8244, new_n5891);
not_10 g03543(n2985, new_n5892);
xnor_4 g03544(new_n5880, new_n5892, new_n5893);
nor_5  g03545(new_n5893, n9493, new_n5894);
xnor_4 g03546(new_n5879, n5605, new_n5895);
nor_5  g03547(new_n5895, n15167, new_n5896);
xnor_4 g03548(new_n5895, n15167, new_n5897);
xor_4  g03549(n15652, n4939, new_n5898);
nor_5  g03550(new_n5898, n21095, new_n5899);
nand_5 g03551(n8656, n4939, new_n5900);
xor_4  g03552(new_n5898, n21095, new_n5901);
and_5  g03553(new_n5901, new_n5900, new_n5902);
nor_5  g03554(new_n5902, new_n5899, new_n5903_1);
nor_5  g03555(new_n5903_1, new_n5897, new_n5904_1);
nor_5  g03556(new_n5904_1, new_n5896, new_n5905);
xnor_4 g03557(new_n5893, n9493, new_n5906);
nor_5  g03558(new_n5906, new_n5905, new_n5907);
nor_5  g03559(new_n5907, new_n5894, new_n5908);
nor_5  g03560(new_n5908, new_n5891, new_n5909);
nor_5  g03561(new_n5909, new_n5890, new_n5910);
nor_5  g03562(new_n5910, new_n5888, new_n5911_1);
or_5   g03563(new_n5911_1, new_n5887, new_n5912);
xnor_4 g03564(new_n5912, new_n5885, new_n5913);
xnor_4 g03565(new_n5913, new_n5875, new_n5914);
xnor_4 g03566(new_n5872, new_n5849, new_n5915);
xor_4  g03567(new_n5910, new_n5888, new_n5916);
nor_5  g03568(new_n5916, new_n5915, new_n5917);
xnor_4 g03569(new_n5916, new_n5915, new_n5918);
xor_4  g03570(new_n5870, new_n5852, new_n5919);
xnor_4 g03571(new_n5908, new_n5891, new_n5920);
nor_5  g03572(new_n5920, new_n5919, new_n5921);
xnor_4 g03573(new_n5920, new_n5919, new_n5922);
xnor_4 g03574(new_n5867, new_n5855, new_n5923);
xnor_4 g03575(new_n5906, new_n5905, new_n5924);
and_5  g03576(new_n5924, new_n5923, new_n5925);
xor_4  g03577(new_n5903_1, new_n5897, new_n5926);
xnor_4 g03578(n21898, n10614, new_n5927);
xnor_4 g03579(new_n5927, new_n5865, new_n5928);
and_5  g03580(new_n5928, new_n5926, new_n5929);
xnor_4 g03581(new_n5928, new_n5926, new_n5930);
xnor_4 g03582(n8656, n4939, new_n5931);
xnor_4 g03583(n22072, n2646, new_n5932);
nor_5  g03584(new_n5932, new_n5931, new_n5933);
xor_4  g03585(n11266, n9926, new_n5934);
xnor_4 g03586(new_n5934, new_n5863, new_n5935);
not_10 g03587(new_n5935, new_n5936_1);
nor_5  g03588(new_n5936_1, new_n5933, new_n5937);
xor_4  g03589(new_n5901, new_n5900, new_n5938);
xnor_4 g03590(new_n5935, new_n5933, new_n5939);
and_5  g03591(new_n5939, new_n5938, new_n5940);
nor_5  g03592(new_n5940, new_n5937, new_n5941);
nor_5  g03593(new_n5941, new_n5930, new_n5942);
or_5   g03594(new_n5942, new_n5929, new_n5943_1);
xnor_4 g03595(new_n5924, new_n5923, new_n5944);
nor_5  g03596(new_n5944, new_n5943_1, new_n5945);
or_5   g03597(new_n5945, new_n5925, new_n5946);
nor_5  g03598(new_n5946, new_n5922, new_n5947);
or_5   g03599(new_n5947, new_n5921, new_n5948);
nor_5  g03600(new_n5948, new_n5918, new_n5949);
nor_5  g03601(new_n5949, new_n5917, new_n5950);
xnor_4 g03602(new_n5950, new_n5914, new_n5951);
xnor_4 g03603(new_n5951, new_n5845, new_n5952);
xor_4  g03604(new_n5948, new_n5918, new_n5953);
nor_5  g03605(new_n5953, new_n4338, new_n5954);
xnor_4 g03606(new_n5953, new_n4338, new_n5955);
nor_5  g03607(new_n5945, new_n5925, new_n5956);
xnor_4 g03608(new_n5956, new_n5922, new_n5957);
and_5  g03609(new_n5957, new_n4341, new_n5958);
xnor_4 g03610(new_n5957, new_n4341, new_n5959);
nor_5  g03611(new_n5942, new_n5929, new_n5960);
xnor_4 g03612(new_n5944, new_n5960, new_n5961);
nor_5  g03613(new_n5961, new_n4345, new_n5962);
xnor_4 g03614(new_n5961, new_n4345, new_n5963);
xnor_4 g03615(new_n5941, new_n5930, new_n5964_1);
nor_5  g03616(new_n5964_1, new_n4352, new_n5965);
xnor_4 g03617(new_n5964_1, new_n4352, new_n5966);
xnor_4 g03618(new_n5932, new_n5931, new_n5967);
or_5   g03619(new_n5967, new_n4361, new_n5968);
and_5  g03620(new_n5968, new_n4358, new_n5969);
xor_4  g03621(new_n5939, new_n5938, new_n5970);
xor_4  g03622(new_n5968, new_n4358, new_n5971);
and_5  g03623(new_n5971, new_n5970, new_n5972);
nor_5  g03624(new_n5972, new_n5969, new_n5973);
nor_5  g03625(new_n5973, new_n5966, new_n5974);
nor_5  g03626(new_n5974, new_n5965, new_n5975);
nor_5  g03627(new_n5975, new_n5963, new_n5976);
nor_5  g03628(new_n5976, new_n5962, new_n5977);
nor_5  g03629(new_n5977, new_n5959, new_n5978);
nor_5  g03630(new_n5978, new_n5958, new_n5979);
nor_5  g03631(new_n5979, new_n5955, new_n5980_1);
or_5   g03632(new_n5980_1, new_n5954, new_n5981);
xor_4  g03633(new_n5981, new_n5952, n597);
xnor_4 g03634(n25926, n9646, new_n5983);
xor_4  g03635(new_n5983, n14230, new_n5984);
xor_4  g03636(new_n5984, new_n5336, n637);
xnor_4 g03637(n25797, n10611, new_n5986);
nor_5  g03638(n15967, n2783, new_n5987);
xnor_4 g03639(n15967, n2783, new_n5988);
nor_5  g03640(n15490, n13319, new_n5989);
and_5  g03641(n25435, n18, new_n5990);
xnor_4 g03642(n15490, n13319, new_n5991);
nor_5  g03643(new_n5991, new_n5990, new_n5992);
nor_5  g03644(new_n5992, new_n5989, new_n5993);
nor_5  g03645(new_n5993, new_n5988, new_n5994);
nor_5  g03646(new_n5994, new_n5987, new_n5995);
xnor_4 g03647(new_n5995, new_n5986, new_n5996);
xnor_4 g03648(new_n5996, n7421, new_n5997);
xnor_4 g03649(new_n5993, new_n5988, new_n5998);
and_5  g03650(new_n5998, n19680, new_n5999);
xor_4  g03651(new_n5998, n19680, new_n6000);
xor_4  g03652(new_n5991, new_n5990, new_n6001);
not_10 g03653(new_n6001, new_n6002);
nor_5  g03654(new_n6002, n2809, new_n6003);
xor_4  g03655(n25435, n18, new_n6004);
nand_5 g03656(new_n6004, n15508, new_n6005);
xnor_4 g03657(new_n6001, n2809, new_n6006);
and_5  g03658(new_n6006, new_n6005, new_n6007);
nor_5  g03659(new_n6007, new_n6003, new_n6008);
and_5  g03660(new_n6008, new_n6000, new_n6009);
nor_5  g03661(new_n6009, new_n5999, new_n6010);
xnor_4 g03662(new_n6010, new_n5997, new_n6011);
xnor_4 g03663(n18157, n11056, new_n6012_1);
nor_5  g03664(n15271, n12161, new_n6013);
xnor_4 g03665(n15271, n12161, new_n6014);
nor_5  g03666(n25877, n5026, new_n6015);
and_5  g03667(n24323, n8581, new_n6016);
xnor_4 g03668(n25877, n5026, new_n6017);
nor_5  g03669(new_n6017, new_n6016, new_n6018);
nor_5  g03670(new_n6018, new_n6015, new_n6019);
nor_5  g03671(new_n6019, new_n6014, new_n6020);
nor_5  g03672(new_n6020, new_n6013, new_n6021);
xnor_4 g03673(new_n6021, new_n6012_1, new_n6022_1);
xnor_4 g03674(new_n6022_1, n20250, new_n6023);
xnor_4 g03675(new_n6019, new_n6014, new_n6024);
nor_5  g03676(new_n6024, n5822, new_n6025);
xnor_4 g03677(new_n6017, new_n6016, new_n6026);
nor_5  g03678(new_n6026, n26443, new_n6027);
xor_4  g03679(n24323, n8581, new_n6028);
nand_5 g03680(new_n6028, n1681, new_n6029);
xor_4  g03681(new_n6026, n26443, new_n6030);
and_5  g03682(new_n6030, new_n6029, new_n6031_1);
nor_5  g03683(new_n6031_1, new_n6027, new_n6032);
xnor_4 g03684(new_n6024, n5822, new_n6033);
nor_5  g03685(new_n6033, new_n6032, new_n6034);
nor_5  g03686(new_n6034, new_n6025, new_n6035);
xor_4  g03687(new_n6035, new_n6023, new_n6036);
xnor_4 g03688(new_n6036, new_n6011, new_n6037);
xor_4  g03689(new_n6008, new_n6000, new_n6038);
xor_4  g03690(new_n6033, new_n6032, new_n6039);
nor_5  g03691(new_n6039, new_n6038, new_n6040);
xnor_4 g03692(new_n6039, new_n6038, new_n6041);
xor_4  g03693(new_n6006, new_n6005, new_n6042);
xnor_4 g03694(new_n6030, new_n6029, new_n6043);
nor_5  g03695(new_n6043, new_n6042, new_n6044_1);
xor_4  g03696(new_n6004, n15508, new_n6045);
not_10 g03697(new_n6045, new_n6046_1);
xor_4  g03698(new_n6028, n1681, new_n6047);
nor_5  g03699(new_n6047, new_n6046_1, new_n6048);
xor_4  g03700(new_n6043, new_n6042, new_n6049);
and_5  g03701(new_n6049, new_n6048, new_n6050);
or_5   g03702(new_n6050, new_n6044_1, new_n6051);
nor_5  g03703(new_n6051, new_n6041, new_n6052);
nor_5  g03704(new_n6052, new_n6040, new_n6053);
xnor_4 g03705(new_n6053, new_n6037, n646);
not_10 g03706(new_n3204, new_n6055);
nor_5  g03707(n19494, n2387, new_n6056);
not_10 g03708(new_n6056, new_n6057);
nor_5  g03709(new_n6057, n16223, new_n6058);
nand_5 g03710(new_n6058, new_n2356, new_n6059);
xnor_4 g03711(new_n6059, new_n2353, new_n6060);
xnor_4 g03712(new_n2447, n7566, new_n6061);
and_5  g03713(new_n2452, n7731, new_n6062);
xnor_4 g03714(new_n2452, n7731, new_n6063);
and_5  g03715(new_n2457, n12341, new_n6064);
xor_4  g03716(new_n2457, n12341, new_n6065);
nor_5  g03717(new_n2462, n12384, new_n6066);
and_5  g03718(new_n6066, new_n5048, new_n6067);
xnor_4 g03719(new_n6066, n20986, new_n6068);
and_5  g03720(new_n6068, new_n2465, new_n6069);
nor_5  g03721(new_n6069, new_n6067, new_n6070);
and_5  g03722(new_n6070, new_n6065, new_n6071);
nor_5  g03723(new_n6071, new_n6064, new_n6072);
nor_5  g03724(new_n6072, new_n6063, new_n6073);
nor_5  g03725(new_n6073, new_n6062, new_n6074);
xor_4  g03726(new_n6074, new_n6061, new_n6075);
xnor_4 g03727(new_n6075, new_n6060, new_n6076);
xnor_4 g03728(new_n6058, n26913, new_n6077);
not_10 g03729(new_n6077, new_n6078);
xnor_4 g03730(new_n6072, new_n6063, new_n6079);
nor_5  g03731(new_n6079, new_n6078, new_n6080);
xnor_4 g03732(new_n6079, new_n6078, new_n6081);
xor_4  g03733(new_n2462, n12384, new_n6082);
not_10 g03734(new_n6082, new_n6083);
and_5  g03735(new_n6083, n2387, new_n6084_1);
and_5  g03736(new_n6084_1, new_n2364, new_n6085);
xor_4  g03737(new_n6068, new_n2465, new_n6086);
not_10 g03738(new_n6086, new_n6087);
xor_4  g03739(n19494, n2387, new_n6088);
nor_5  g03740(new_n6088, new_n6084_1, new_n6089);
nor_5  g03741(new_n6089, new_n6085, new_n6090);
and_5  g03742(new_n6090, new_n6087, new_n6091);
nor_5  g03743(new_n6091, new_n6085, new_n6092);
xnor_4 g03744(new_n6056, n16223, new_n6093);
not_10 g03745(new_n6093, new_n6094);
nor_5  g03746(new_n6094, new_n6092, new_n6095);
xor_4  g03747(new_n6070, new_n6065, new_n6096);
xnor_4 g03748(new_n6093, new_n6092, new_n6097);
and_5  g03749(new_n6097, new_n6096, new_n6098);
nor_5  g03750(new_n6098, new_n6095, new_n6099);
nor_5  g03751(new_n6099, new_n6081, new_n6100);
nor_5  g03752(new_n6100, new_n6080, new_n6101);
xor_4  g03753(new_n6101, new_n6076, new_n6102);
xnor_4 g03754(new_n6102, new_n6055, new_n6103);
not_10 g03755(new_n3208_1, new_n6104_1);
xor_4  g03756(new_n6099, new_n6081, new_n6105_1);
nor_5  g03757(new_n6105_1, new_n6104_1, new_n6106);
not_10 g03758(new_n3212, new_n6107);
not_10 g03759(new_n6096, new_n6108);
xnor_4 g03760(new_n6097, new_n6108, new_n6109);
and_5  g03761(new_n6109, new_n6107, new_n6110);
xnor_4 g03762(new_n6109, new_n6107, new_n6111);
xor_4  g03763(new_n6082, n2387, new_n6112);
nor_5  g03764(new_n6112, new_n3215, new_n6113);
nor_5  g03765(new_n6113, new_n3218, new_n6114);
xnor_4 g03766(new_n6090, new_n6087, new_n6115);
and_5  g03767(new_n6113, new_n3221, new_n6116);
nor_5  g03768(new_n6116, new_n6114, new_n6117);
and_5  g03769(new_n6117, new_n6115, new_n6118);
or_5   g03770(new_n6118, new_n6114, new_n6119);
nor_5  g03771(new_n6119, new_n6111, new_n6120);
nor_5  g03772(new_n6120, new_n6110, new_n6121);
xnor_4 g03773(new_n6105_1, new_n3208_1, new_n6122);
and_5  g03774(new_n6122, new_n6121, new_n6123);
nor_5  g03775(new_n6123, new_n6106, new_n6124);
xnor_4 g03776(new_n6124, new_n6103, n696);
xnor_4 g03777(n25475, n23697, new_n6126);
nor_5  g03778(n23849, n2289, new_n6127);
xnor_4 g03779(n23849, n2289, new_n6128);
nor_5  g03780(n12446, n1112, new_n6129);
xnor_4 g03781(n12446, n1112, new_n6130);
nor_5  g03782(n20179, n11011, new_n6131);
xnor_4 g03783(n20179, n11011, new_n6132);
nor_5  g03784(n19228, n16029, new_n6133);
xnor_4 g03785(n19228, n16029, new_n6134);
nor_5  g03786(n16476, n15539, new_n6135);
xnor_4 g03787(n16476, n15539, new_n6136);
nor_5  g03788(n11615, n8052, new_n6137);
xnor_4 g03789(n11615, n8052, new_n6138);
nor_5  g03790(n22433, n10158, new_n6139);
and_5  g03791(n18962, n14090, new_n6140);
xnor_4 g03792(n22433, n10158, new_n6141);
nor_5  g03793(new_n6141, new_n6140, new_n6142);
nor_5  g03794(new_n6142, new_n6139, new_n6143);
nor_5  g03795(new_n6143, new_n6138, new_n6144);
nor_5  g03796(new_n6144, new_n6137, new_n6145);
nor_5  g03797(new_n6145, new_n6136, new_n6146);
nor_5  g03798(new_n6146, new_n6135, new_n6147);
nor_5  g03799(new_n6147, new_n6134, new_n6148);
nor_5  g03800(new_n6148, new_n6133, new_n6149);
nor_5  g03801(new_n6149, new_n6132, new_n6150);
nor_5  g03802(new_n6150, new_n6131, new_n6151);
nor_5  g03803(new_n6151, new_n6130, new_n6152);
nor_5  g03804(new_n6152, new_n6129, new_n6153);
nor_5  g03805(new_n6153, new_n6128, new_n6154);
nor_5  g03806(new_n6154, new_n6127, new_n6155);
xnor_4 g03807(new_n6155, new_n6126, new_n6156);
xnor_4 g03808(new_n6156, n25345, new_n6157);
xnor_4 g03809(new_n6153, new_n6128, new_n6158);
and_5  g03810(new_n6158, n9655, new_n6159);
xnor_4 g03811(new_n6158, n9655, new_n6160_1);
xnor_4 g03812(new_n6151, new_n6130, new_n6161);
nand_5 g03813(new_n6161, n13490, new_n6162);
xnor_4 g03814(new_n6161, n13490, new_n6163);
xnor_4 g03815(new_n6149, new_n6132, new_n6164);
nand_5 g03816(new_n6164, n22660, new_n6165);
xnor_4 g03817(new_n6147, new_n6134, new_n6166);
nor_5  g03818(new_n6166, n1777, new_n6167);
xnor_4 g03819(new_n6166, n1777, new_n6168);
xnor_4 g03820(new_n6145, new_n6136, new_n6169);
nor_5  g03821(new_n6169, n8745, new_n6170);
xor_4  g03822(new_n6169, n8745, new_n6171_1);
xnor_4 g03823(new_n6143, new_n6138, new_n6172);
and_5  g03824(new_n6172, n15636, new_n6173);
xor_4  g03825(new_n6172, n15636, new_n6174);
xor_4  g03826(n18962, n14090, new_n6175);
and_5  g03827(new_n6175, n6794, new_n6176);
nor_5  g03828(new_n6176, n20077, new_n6177);
xor_4  g03829(new_n6141, new_n6140, new_n6178);
not_10 g03830(new_n6178, new_n6179);
xnor_4 g03831(new_n6176, n20077, new_n6180);
nor_5  g03832(new_n6180, new_n6179, new_n6181);
nor_5  g03833(new_n6181, new_n6177, new_n6182);
and_5  g03834(new_n6182, new_n6174, new_n6183_1);
nor_5  g03835(new_n6183_1, new_n6173, new_n6184);
and_5  g03836(new_n6184, new_n6171_1, new_n6185);
nor_5  g03837(new_n6185, new_n6170, new_n6186);
nor_5  g03838(new_n6186, new_n6168, new_n6187);
nor_5  g03839(new_n6187, new_n6167, new_n6188);
not_10 g03840(new_n6188, new_n6189_1);
xnor_4 g03841(new_n6164, n22660, new_n6190);
or_5   g03842(new_n6190, new_n6189_1, new_n6191);
and_5  g03843(new_n6191, new_n6165, new_n6192);
or_5   g03844(new_n6192, new_n6163, new_n6193);
and_5  g03845(new_n6193, new_n6162, new_n6194);
nor_5  g03846(new_n6194, new_n6160_1, new_n6195);
nor_5  g03847(new_n6195, new_n6159, new_n6196);
xnor_4 g03848(new_n6196, new_n6157, new_n6197);
xnor_4 g03849(n21915, n15182, new_n6198);
nor_5  g03850(n27037, n13775, new_n6199);
xnor_4 g03851(n27037, n13775, new_n6200);
nor_5  g03852(n8964, n1293, new_n6201);
xnor_4 g03853(n8964, n1293, new_n6202);
nor_5  g03854(n20151, n19042, new_n6203);
xnor_4 g03855(n20151, n19042, new_n6204_1);
nor_5  g03856(n19472, n7693, new_n6205);
xor_4  g03857(n19472, n7693, new_n6206);
and_5  g03858(n25370, n10405, new_n6207);
or_5   g03859(n25370, n10405, new_n6208);
nor_5  g03860(n24786, n11302, new_n6209);
nor_5  g03861(new_n3847, new_n3842_1, new_n6210);
nor_5  g03862(new_n6210, new_n6209, new_n6211);
and_5  g03863(new_n6211, new_n6208, new_n6212);
nor_5  g03864(new_n6212, new_n6207, new_n6213);
and_5  g03865(new_n6213, new_n6206, new_n6214);
nor_5  g03866(new_n6214, new_n6205, new_n6215);
nor_5  g03867(new_n6215, new_n6204_1, new_n6216);
nor_5  g03868(new_n6216, new_n6203, new_n6217);
nor_5  g03869(new_n6217, new_n6202, new_n6218_1);
nor_5  g03870(new_n6218_1, new_n6201, new_n6219);
nor_5  g03871(new_n6219, new_n6200, new_n6220);
nor_5  g03872(new_n6220, new_n6199, new_n6221);
xnor_4 g03873(new_n6221, new_n6198, new_n6222);
xnor_4 g03874(new_n6222, n17351, new_n6223_1);
xnor_4 g03875(new_n6219, new_n6200, new_n6224);
and_5  g03876(new_n6224, n11736, new_n6225);
xnor_4 g03877(new_n6224, n11736, new_n6226);
xnor_4 g03878(new_n6217, new_n6202, new_n6227);
and_5  g03879(new_n6227, n23200, new_n6228);
xnor_4 g03880(new_n6227, n23200, new_n6229);
xnor_4 g03881(new_n6215, new_n6204_1, new_n6230);
and_5  g03882(new_n6230, n17959, new_n6231);
xnor_4 g03883(new_n6230, n17959, new_n6232);
xnor_4 g03884(new_n6213, new_n6206, new_n6233_1);
and_5  g03885(new_n6233_1, n7566, new_n6234);
xnor_4 g03886(new_n6233_1, n7566, new_n6235);
xnor_4 g03887(n25370, n10405, new_n6236);
xnor_4 g03888(new_n6236, new_n6211, new_n6237);
and_5  g03889(new_n6237, n7731, new_n6238);
xnor_4 g03890(new_n6237, n7731, new_n6239);
nor_5  g03891(new_n3848, new_n5045, new_n6240);
and_5  g03892(new_n3860, new_n5048, new_n6241);
nand_5 g03893(new_n3864, n12384, new_n6242);
xnor_4 g03894(new_n3860, n20986, new_n6243);
and_5  g03895(new_n6243, new_n6242, new_n6244);
nor_5  g03896(new_n6244, new_n6241, new_n6245_1);
xnor_4 g03897(new_n3848, n12341, new_n6246);
and_5  g03898(new_n6246, new_n6245_1, new_n6247);
nor_5  g03899(new_n6247, new_n6240, new_n6248_1);
nor_5  g03900(new_n6248_1, new_n6239, new_n6249);
nor_5  g03901(new_n6249, new_n6238, new_n6250);
nor_5  g03902(new_n6250, new_n6235, new_n6251);
nor_5  g03903(new_n6251, new_n6234, new_n6252);
nor_5  g03904(new_n6252, new_n6232, new_n6253);
nor_5  g03905(new_n6253, new_n6231, new_n6254);
nor_5  g03906(new_n6254, new_n6229, new_n6255);
nor_5  g03907(new_n6255, new_n6228, new_n6256_1);
nor_5  g03908(new_n6256_1, new_n6226, new_n6257);
nor_5  g03909(new_n6257, new_n6225, new_n6258);
xor_4  g03910(new_n6258, new_n6223_1, new_n6259);
xnor_4 g03911(new_n6259, new_n6197, new_n6260);
xnor_4 g03912(new_n6256_1, new_n6226, new_n6261);
xor_4  g03913(new_n6194, new_n6160_1, new_n6262);
and_5  g03914(new_n6262, new_n6261, new_n6263);
xnor_4 g03915(new_n6262, new_n6261, new_n6264);
xnor_4 g03916(new_n6254, new_n6229, new_n6265);
xor_4  g03917(new_n6192, new_n6163, new_n6266);
and_5  g03918(new_n6266, new_n6265, new_n6267);
xnor_4 g03919(new_n6266, new_n6265, new_n6268);
xnor_4 g03920(new_n6252, new_n6232, new_n6269);
xnor_4 g03921(new_n6190, new_n6188, new_n6270);
and_5  g03922(new_n6270, new_n6269, new_n6271_1);
xnor_4 g03923(new_n6270, new_n6269, new_n6272);
xor_4  g03924(new_n6186, new_n6168, new_n6273);
xor_4  g03925(new_n6250, new_n6235, new_n6274);
nor_5  g03926(new_n6274, new_n6273, new_n6275);
xnor_4 g03927(new_n6274, new_n6273, new_n6276_1);
xor_4  g03928(new_n6184, new_n6171_1, new_n6277);
xor_4  g03929(new_n6248_1, new_n6239, new_n6278);
nor_5  g03930(new_n6278, new_n6277, new_n6279);
xnor_4 g03931(new_n6278, new_n6277, new_n6280);
xnor_4 g03932(new_n6246, new_n6245_1, new_n6281);
xor_4  g03933(new_n6182, new_n6174, new_n6282);
and_5  g03934(new_n6282, new_n6281, new_n6283);
xnor_4 g03935(new_n6282, new_n6281, new_n6284);
xnor_4 g03936(new_n6243, new_n6242, new_n6285);
xnor_4 g03937(new_n6180, new_n6178, new_n6286);
nor_5  g03938(new_n6286, new_n6285, new_n6287);
xor_4  g03939(new_n6175, n6794, new_n6288);
not_10 g03940(new_n6288, new_n6289);
xor_4  g03941(new_n3864, n12384, new_n6290);
nor_5  g03942(new_n6290, new_n6289, new_n6291);
xor_4  g03943(new_n6286, new_n6285, new_n6292);
and_5  g03944(new_n6292, new_n6291, new_n6293);
nor_5  g03945(new_n6293, new_n6287, new_n6294);
nor_5  g03946(new_n6294, new_n6284, new_n6295);
nor_5  g03947(new_n6295, new_n6283, new_n6296);
nor_5  g03948(new_n6296, new_n6280, new_n6297);
nor_5  g03949(new_n6297, new_n6279, new_n6298);
nor_5  g03950(new_n6298, new_n6276_1, new_n6299);
nor_5  g03951(new_n6299, new_n6275, new_n6300);
nor_5  g03952(new_n6300, new_n6272, new_n6301);
nor_5  g03953(new_n6301, new_n6271_1, new_n6302);
nor_5  g03954(new_n6302, new_n6268, new_n6303);
nor_5  g03955(new_n6303, new_n6267, new_n6304);
nor_5  g03956(new_n6304, new_n6264, new_n6305);
nor_5  g03957(new_n6305, new_n6263, new_n6306);
xnor_4 g03958(new_n6306, new_n6260, n723);
xor_4  g03959(n26986, n2272, new_n6308_1);
not_10 g03960(n21287, new_n6309);
and_5  g03961(n25331, new_n6309, new_n6310);
xor_4  g03962(n25331, n21287, new_n6311_1);
not_10 g03963(n4256, new_n6312);
and_5  g03964(n18483, new_n6312, new_n6313);
xor_4  g03965(n18483, n4256, new_n6314);
not_10 g03966(n22332, new_n6315);
and_5  g03967(new_n6315, n21934, new_n6316);
xor_4  g03968(n22332, n21934, new_n6317);
and_5  g03969(new_n3585, n18901, new_n6318);
xor_4  g03970(n18907, n18901, new_n6319);
and_5  g03971(n4376, new_n3588, new_n6320);
xor_4  g03972(n4376, n2731, new_n6321);
and_5  g03973(new_n3591, n14570, new_n6322);
xor_4  g03974(n19911, n14570, new_n6323_1);
nor_5  g03975(n23775, new_n3596, new_n6324);
and_5  g03976(n23775, new_n3596, new_n6325);
nor_5  g03977(new_n3600, n8259, new_n6326);
and_5  g03978(new_n3600, n8259, new_n6327);
not_10 g03979(n5704, new_n6328);
or_5   g03980(n11479, new_n6328, new_n6329);
nor_5  g03981(new_n6329, new_n6327, new_n6330_1);
nor_5  g03982(new_n6330_1, new_n6326, new_n6331);
nor_5  g03983(new_n6331, new_n6325, new_n6332);
or_5   g03984(new_n6332, new_n6324, new_n6333);
nor_5  g03985(new_n6333, new_n6323_1, new_n6334);
nor_5  g03986(new_n6334, new_n6322, new_n6335);
nor_5  g03987(new_n6335, new_n6321, new_n6336);
nor_5  g03988(new_n6336, new_n6320, new_n6337);
nor_5  g03989(new_n6337, new_n6319, new_n6338);
nor_5  g03990(new_n6338, new_n6318, new_n6339_1);
nor_5  g03991(new_n6339_1, new_n6317, new_n6340);
nor_5  g03992(new_n6340, new_n6316, new_n6341);
nor_5  g03993(new_n6341, new_n6314, new_n6342);
nor_5  g03994(new_n6342, new_n6313, new_n6343);
nor_5  g03995(new_n6343, new_n6311_1, new_n6344);
nor_5  g03996(new_n6344, new_n6310, new_n6345);
xnor_4 g03997(new_n6345, new_n6308_1, new_n6346);
xnor_4 g03998(n1255, n468, new_n6347);
nor_5  g03999(n9512, n5400, new_n6348);
xnor_4 g04000(n9512, n5400, new_n6349);
nor_5  g04001(n23923, n16608, new_n6350);
xnor_4 g04002(n23923, n16608, new_n6351);
nor_5  g04003(n21735, n329, new_n6352);
xnor_4 g04004(n21735, n329, new_n6353);
nor_5  g04005(n24170, n24085, new_n6354_1);
xnor_4 g04006(n24170, n24085, new_n6355);
nor_5  g04007(n14071, n2409, new_n6356_1);
xnor_4 g04008(n14071, n2409, new_n6357);
nor_5  g04009(n8869, n1738, new_n6358);
xnor_4 g04010(n8869, n1738, new_n6359);
nor_5  g04011(n12152, n10372, new_n6360);
and_5  g04012(n19107, n7428, new_n6361);
xnor_4 g04013(n12152, n10372, new_n6362);
nor_5  g04014(new_n6362, new_n6361, new_n6363);
nor_5  g04015(new_n6363, new_n6360, new_n6364);
nor_5  g04016(new_n6364, new_n6359, new_n6365);
nor_5  g04017(new_n6365, new_n6358, new_n6366);
nor_5  g04018(new_n6366, new_n6357, new_n6367);
nor_5  g04019(new_n6367, new_n6356_1, new_n6368);
nor_5  g04020(new_n6368, new_n6355, new_n6369_1);
nor_5  g04021(new_n6369_1, new_n6354_1, new_n6370);
nor_5  g04022(new_n6370, new_n6353, new_n6371);
nor_5  g04023(new_n6371, new_n6352, new_n6372);
nor_5  g04024(new_n6372, new_n6351, new_n6373);
nor_5  g04025(new_n6373, new_n6350, new_n6374);
nor_5  g04026(new_n6374, new_n6349, new_n6375_1);
nor_5  g04027(new_n6375_1, new_n6348, new_n6376);
xnor_4 g04028(new_n6376, new_n6347, new_n6377);
xnor_4 g04029(n14130, n12861, new_n6378);
nor_5  g04030(n16482, n13333, new_n6379_1);
xnor_4 g04031(n16482, n13333, new_n6380);
nor_5  g04032(n9942, n2210, new_n6381_1);
xnor_4 g04033(n9942, n2210, new_n6382);
nor_5  g04034(n25643, n20604, new_n6383_1);
nor_5  g04035(new_n4733, new_n4730, new_n6384);
nor_5  g04036(new_n6384, new_n6383_1, new_n6385_1);
nor_5  g04037(new_n6385_1, new_n6382, new_n6386);
nor_5  g04038(new_n6386, new_n6381_1, new_n6387);
nor_5  g04039(new_n6387, new_n6380, new_n6388);
nor_5  g04040(new_n6388, new_n6379_1, new_n6389);
xor_4  g04041(new_n6389, new_n6378, new_n6390);
nor_5  g04042(new_n6390, new_n6377, new_n6391);
xnor_4 g04043(new_n6390, new_n6377, new_n6392);
xnor_4 g04044(new_n6374, new_n6349, new_n6393);
xor_4  g04045(new_n6387, new_n6380, new_n6394);
nor_5  g04046(new_n6394, new_n6393, new_n6395);
xnor_4 g04047(new_n6394, new_n6393, new_n6396);
xnor_4 g04048(new_n6385_1, new_n6382, new_n6397_1);
xor_4  g04049(new_n6372, new_n6351, new_n6398);
and_5  g04050(new_n6398, new_n6397_1, new_n6399);
xnor_4 g04051(new_n6398, new_n6397_1, new_n6400);
not_10 g04052(new_n4734, new_n6401);
xor_4  g04053(new_n6370, new_n6353, new_n6402);
and_5  g04054(new_n6402, new_n6401, new_n6403);
xor_4  g04055(new_n6402, new_n4734, new_n6404);
xor_4  g04056(new_n6368, new_n6355, new_n6405);
and_5  g04057(new_n6405, new_n4728, new_n6406);
xor_4  g04058(new_n6405, new_n4727, new_n6407_1);
xor_4  g04059(new_n6366, new_n6357, new_n6408);
and_5  g04060(new_n6408, new_n4721, new_n6409);
xor_4  g04061(new_n6408, new_n4720, new_n6410);
xor_4  g04062(new_n6364, new_n6359, new_n6411);
and_5  g04063(new_n6411, new_n4714, new_n6412);
xnor_4 g04064(new_n6411, new_n4714, new_n6413);
xor_4  g04065(new_n6362, new_n6361, new_n6414);
and_5  g04066(new_n6414, new_n4707, new_n6415);
xnor_4 g04067(n19107, n7428, new_n6416);
nand_5 g04068(new_n6416, new_n4704, new_n6417);
xnor_4 g04069(new_n6414, new_n4707, new_n6418);
nor_5  g04070(new_n6418, new_n6417, new_n6419);
nor_5  g04071(new_n6419, new_n6415, new_n6420);
nor_5  g04072(new_n6420, new_n6413, new_n6421);
nor_5  g04073(new_n6421, new_n6412, new_n6422);
nor_5  g04074(new_n6422, new_n6410, new_n6423);
nor_5  g04075(new_n6423, new_n6409, new_n6424);
nor_5  g04076(new_n6424, new_n6407_1, new_n6425);
nor_5  g04077(new_n6425, new_n6406, new_n6426);
nor_5  g04078(new_n6426, new_n6404, new_n6427_1);
nor_5  g04079(new_n6427_1, new_n6403, new_n6428);
nor_5  g04080(new_n6428, new_n6400, new_n6429);
nor_5  g04081(new_n6429, new_n6399, new_n6430);
nor_5  g04082(new_n6430, new_n6396, new_n6431_1);
nor_5  g04083(new_n6431_1, new_n6395, new_n6432);
nor_5  g04084(new_n6432, new_n6392, new_n6433);
nor_5  g04085(new_n6433, new_n6391, new_n6434);
xnor_4 g04086(n22442, n22253, new_n6435);
nor_5  g04087(n1255, n468, new_n6436);
nor_5  g04088(new_n6376, new_n6347, new_n6437_1);
nor_5  g04089(new_n6437_1, new_n6436, new_n6438);
xnor_4 g04090(new_n6438, new_n6435, new_n6439);
xnor_4 g04091(n8856, n8305, new_n6440);
nor_5  g04092(n14130, n12861, new_n6441);
nor_5  g04093(new_n6389, new_n6378, new_n6442);
nor_5  g04094(new_n6442, new_n6441, new_n6443);
xor_4  g04095(new_n6443, new_n6440, new_n6444);
xnor_4 g04096(new_n6444, new_n6439, new_n6445);
xor_4  g04097(new_n6445, new_n6434, new_n6446);
and_5  g04098(new_n6446, new_n6346, new_n6447);
xnor_4 g04099(new_n6446, new_n6346, new_n6448);
xnor_4 g04100(new_n6343, new_n6311_1, new_n6449);
xor_4  g04101(new_n6432, new_n6392, new_n6450);
and_5  g04102(new_n6450, new_n6449, new_n6451);
xnor_4 g04103(new_n6450, new_n6449, new_n6452);
xnor_4 g04104(new_n6341, new_n6314, new_n6453);
xor_4  g04105(new_n6430, new_n6396, new_n6454);
and_5  g04106(new_n6454, new_n6453, new_n6455);
xnor_4 g04107(new_n6454, new_n6453, new_n6456_1);
xnor_4 g04108(new_n6339_1, new_n6317, new_n6457_1);
xor_4  g04109(new_n6428, new_n6400, new_n6458);
and_5  g04110(new_n6458, new_n6457_1, new_n6459);
xnor_4 g04111(new_n6458, new_n6457_1, new_n6460);
xnor_4 g04112(new_n6337, new_n6319, new_n6461);
xor_4  g04113(new_n6426, new_n6404, new_n6462);
and_5  g04114(new_n6462, new_n6461, new_n6463);
xnor_4 g04115(new_n6462, new_n6461, new_n6464);
xnor_4 g04116(new_n6335, new_n6321, new_n6465_1);
xor_4  g04117(new_n6424, new_n6407_1, new_n6466);
and_5  g04118(new_n6466, new_n6465_1, new_n6467);
xnor_4 g04119(new_n6466, new_n6465_1, new_n6468);
xnor_4 g04120(new_n6422, new_n6410, new_n6469);
xor_4  g04121(new_n6333, new_n6323_1, new_n6470_1);
nor_5  g04122(new_n6470_1, new_n6469, new_n6471);
xor_4  g04123(new_n6420, new_n6413, new_n6472);
xnor_4 g04124(n23775, n13708, new_n6473);
xnor_4 g04125(new_n6473, new_n6331, new_n6474);
and_5  g04126(new_n6474, new_n6472, new_n6475);
not_10 g04127(new_n6472, new_n6476_1);
xnor_4 g04128(new_n6474, new_n6476_1, new_n6477);
xor_4  g04129(new_n6416, new_n4704, new_n6478);
xnor_4 g04130(n11479, n5704, new_n6479);
or_5   g04131(new_n6479, new_n6478, new_n6480);
xnor_4 g04132(n18409, n8259, new_n6481);
xnor_4 g04133(new_n6481, new_n6329, new_n6482);
nor_5  g04134(new_n6482, new_n6480, new_n6483);
xor_4  g04135(new_n6418, new_n6417, new_n6484);
xnor_4 g04136(new_n6482, new_n6480, new_n6485_1);
nor_5  g04137(new_n6485_1, new_n6484, new_n6486);
nor_5  g04138(new_n6486, new_n6483, new_n6487);
and_5  g04139(new_n6487, new_n6477, new_n6488);
nor_5  g04140(new_n6488, new_n6475, new_n6489);
xnor_4 g04141(new_n6470_1, new_n6469, new_n6490);
nor_5  g04142(new_n6490, new_n6489, new_n6491);
nor_5  g04143(new_n6491, new_n6471, new_n6492);
nor_5  g04144(new_n6492, new_n6468, new_n6493);
nor_5  g04145(new_n6493, new_n6467, new_n6494);
nor_5  g04146(new_n6494, new_n6464, new_n6495);
nor_5  g04147(new_n6495, new_n6463, new_n6496);
nor_5  g04148(new_n6496, new_n6460, new_n6497);
nor_5  g04149(new_n6497, new_n6459, new_n6498);
nor_5  g04150(new_n6498, new_n6456_1, new_n6499);
nor_5  g04151(new_n6499, new_n6455, new_n6500);
nor_5  g04152(new_n6500, new_n6452, new_n6501);
nor_5  g04153(new_n6501, new_n6451, new_n6502_1);
nor_5  g04154(new_n6502_1, new_n6448, new_n6503);
nor_5  g04155(new_n6503, new_n6447, new_n6504);
not_10 g04156(n26986, new_n6505);
and_5  g04157(new_n6505, n2272, new_n6506_1);
nor_5  g04158(new_n6345, new_n6308_1, new_n6507);
nor_5  g04159(new_n6507, new_n6506_1, new_n6508);
nor_5  g04160(n22442, n22253, new_n6509);
nor_5  g04161(new_n6438, new_n6435, new_n6510);
nor_5  g04162(new_n6510, new_n6509, new_n6511);
nor_5  g04163(n8856, n8305, new_n6512);
nor_5  g04164(new_n6443, new_n6440, new_n6513_1);
or_5   g04165(new_n6513_1, new_n6512, new_n6514_1);
xor_4  g04166(new_n6514_1, new_n6511, new_n6515);
nor_5  g04167(new_n6444, new_n6439, new_n6516);
nor_5  g04168(new_n6445, new_n6434, new_n6517);
nor_5  g04169(new_n6517, new_n6516, new_n6518);
xor_4  g04170(new_n6518, new_n6515, new_n6519);
xnor_4 g04171(new_n6519, new_n6508, new_n6520);
xnor_4 g04172(new_n6520, new_n6504, n735);
xnor_4 g04173(n21138, n14230, new_n6522);
xor_4  g04174(new_n6175, n19234, new_n6523);
xor_4  g04175(new_n6523, n26167, new_n6524);
xnor_4 g04176(new_n6524, new_n6522, n779);
not_10 g04177(n17458, new_n6526);
and_5  g04178(new_n6526, n8526, new_n6527);
xor_4  g04179(n17458, n8526, new_n6528);
not_10 g04180(n1222, new_n6529);
and_5  g04181(n2816, new_n6529, new_n6530);
xor_4  g04182(n2816, n1222, new_n6531);
not_10 g04183(n25240, new_n6532);
and_5  g04184(new_n6532, n20359, new_n6533);
xor_4  g04185(n25240, n20359, new_n6534);
not_10 g04186(n10125, new_n6535);
and_5  g04187(new_n6535, n4409, new_n6536);
xor_4  g04188(n10125, n4409, new_n6537);
not_10 g04189(n8067, new_n6538);
and_5  g04190(new_n6538, n3570, new_n6539);
xor_4  g04191(n8067, n3570, new_n6540);
not_10 g04192(n20923, new_n6541);
nand_5 g04193(new_n6541, n13668, new_n6542_1);
xor_4  g04194(n20923, n13668, new_n6543);
not_10 g04195(n18157, new_n6544);
nand_5 g04196(n21276, new_n6544, new_n6545);
xor_4  g04197(n21276, n18157, new_n6546);
not_10 g04198(n12161, new_n6547);
nor_5  g04199(n26748, new_n6547, new_n6548);
and_5  g04200(n26748, new_n6547, new_n6549);
not_10 g04201(n5026, new_n6550);
nor_5  g04202(n10057, new_n6550, new_n6551);
nand_5 g04203(n10057, new_n6550, new_n6552);
not_10 g04204(n8581, new_n6553);
nor_5  g04205(n8920, new_n6553, new_n6554);
and_5  g04206(new_n6554, new_n6552, new_n6555);
nor_5  g04207(new_n6555, new_n6551, new_n6556_1);
nor_5  g04208(new_n6556_1, new_n6549, new_n6557);
nor_5  g04209(new_n6557, new_n6548, new_n6558_1);
not_10 g04210(new_n6558_1, new_n6559);
or_5   g04211(new_n6559, new_n6546, new_n6560_1);
and_5  g04212(new_n6560_1, new_n6545, new_n6561);
or_5   g04213(new_n6561, new_n6543, new_n6562);
and_5  g04214(new_n6562, new_n6542_1, new_n6563);
nor_5  g04215(new_n6563, new_n6540, new_n6564);
nor_5  g04216(new_n6564, new_n6539, new_n6565);
nor_5  g04217(new_n6565, new_n6537, new_n6566);
nor_5  g04218(new_n6566, new_n6536, new_n6567_1);
nor_5  g04219(new_n6567_1, new_n6534, new_n6568);
nor_5  g04220(new_n6568, new_n6533, new_n6569);
nor_5  g04221(new_n6569, new_n6531, new_n6570);
nor_5  g04222(new_n6570, new_n6530, new_n6571);
nor_5  g04223(new_n6571, new_n6528, new_n6572);
nor_5  g04224(new_n6572, new_n6527, new_n6573);
nor_5  g04225(new_n6505, n19282, new_n6574);
xor_4  g04226(n26986, n19282, new_n6575);
nor_5  g04227(new_n6309, n12657, new_n6576_1);
xor_4  g04228(n21287, n12657, new_n6577);
nor_5  g04229(n17077, new_n6312, new_n6578);
xor_4  g04230(n17077, n4256, new_n6579);
nor_5  g04231(n26510, new_n6315, new_n6580);
nor_5  g04232(new_n3613, new_n3584, new_n6581);
nor_5  g04233(new_n6581, new_n6580, new_n6582);
nor_5  g04234(new_n6582, new_n6579, new_n6583);
nor_5  g04235(new_n6583, new_n6578, new_n6584);
nor_5  g04236(new_n6584, new_n6577, new_n6585);
nor_5  g04237(new_n6585, new_n6576_1, new_n6586);
nor_5  g04238(new_n6586, new_n6575, new_n6587_1);
nor_5  g04239(new_n6587_1, new_n6574, new_n6588);
xnor_4 g04240(new_n6588, new_n6573, new_n6589);
xor_4  g04241(new_n6571, new_n6528, new_n6590_1);
xor_4  g04242(new_n6586, new_n6575, new_n6591);
and_5  g04243(new_n6591, new_n6590_1, new_n6592);
xnor_4 g04244(new_n6591, new_n6590_1, new_n6593);
xor_4  g04245(new_n6569, new_n6531, new_n6594);
xor_4  g04246(new_n6584, new_n6577, new_n6595);
nor_5  g04247(new_n6595, new_n6594, new_n6596_1);
xnor_4 g04248(new_n6595, new_n6594, new_n6597);
xor_4  g04249(new_n6567_1, new_n6534, new_n6598);
xor_4  g04250(new_n6582, new_n6579, new_n6599);
nor_5  g04251(new_n6599, new_n6598, new_n6600);
xnor_4 g04252(new_n6599, new_n6598, new_n6601);
xor_4  g04253(new_n6565, new_n6537, new_n6602);
nor_5  g04254(new_n6602, new_n3614, new_n6603);
xnor_4 g04255(new_n6602, new_n3614, new_n6604);
xor_4  g04256(new_n6563, new_n6540, new_n6605);
nor_5  g04257(new_n6605, new_n3623, new_n6606);
xnor_4 g04258(new_n6605, new_n3623, new_n6607);
xor_4  g04259(new_n6561, new_n6543, new_n6608);
nor_5  g04260(new_n6608, new_n3627, new_n6609);
xnor_4 g04261(new_n6608, new_n3627, new_n6610);
xnor_4 g04262(new_n6558_1, new_n6546, new_n6611_1);
nor_5  g04263(new_n6611_1, new_n3632, new_n6612_1);
xnor_4 g04264(new_n6611_1, new_n3632, new_n6613);
xnor_4 g04265(n26748, n12161, new_n6614);
xnor_4 g04266(new_n6614, new_n6556_1, new_n6615);
and_5  g04267(new_n6615, new_n3637, new_n6616);
xnor_4 g04268(new_n6615, new_n3637, new_n6617);
xor_4  g04269(n10057, n5026, new_n6618);
xnor_4 g04270(new_n6618, new_n6554, new_n6619);
nor_5  g04271(new_n6619, new_n3642_1, new_n6620);
xnor_4 g04272(n8920, n8581, new_n6621);
nor_5  g04273(new_n6621, new_n3682, new_n6622);
xor_4  g04274(new_n6619, new_n3642_1, new_n6623);
and_5  g04275(new_n6623, new_n6622, new_n6624);
nor_5  g04276(new_n6624, new_n6620, new_n6625);
not_10 g04277(new_n6625, new_n6626);
nor_5  g04278(new_n6626, new_n6617, new_n6627);
nor_5  g04279(new_n6627, new_n6616, new_n6628_1);
nor_5  g04280(new_n6628_1, new_n6613, new_n6629);
nor_5  g04281(new_n6629, new_n6612_1, new_n6630_1);
nor_5  g04282(new_n6630_1, new_n6610, new_n6631_1);
nor_5  g04283(new_n6631_1, new_n6609, new_n6632);
nor_5  g04284(new_n6632, new_n6607, new_n6633);
nor_5  g04285(new_n6633, new_n6606, new_n6634_1);
nor_5  g04286(new_n6634_1, new_n6604, new_n6635);
nor_5  g04287(new_n6635, new_n6603, new_n6636);
nor_5  g04288(new_n6636, new_n6601, new_n6637);
nor_5  g04289(new_n6637, new_n6600, new_n6638);
nor_5  g04290(new_n6638, new_n6597, new_n6639);
or_5   g04291(new_n6639, new_n6596_1, new_n6640);
nor_5  g04292(new_n6640, new_n6593, new_n6641);
nor_5  g04293(new_n6641, new_n6592, new_n6642);
xnor_4 g04294(new_n6642, new_n6589, new_n6643);
nor_5  g04295(n11898, new_n5384, new_n6644);
xor_4  g04296(n11898, n2979, new_n6645);
nor_5  g04297(n19941, new_n5385, new_n6646);
xor_4  g04298(n19941, n647, new_n6647);
nor_5  g04299(new_n5437, n1099, new_n6648);
xor_4  g04300(n20409, n1099, new_n6649);
nor_5  g04301(new_n5442, n2113, new_n6650);
xor_4  g04302(n25749, n2113, new_n6651);
nor_5  g04303(n21134, new_n3553, new_n6652_1);
xor_4  g04304(n21134, n3161, new_n6653);
nor_5  g04305(new_n5451_1, n6369, new_n6654);
xor_4  g04306(n9003, n6369, new_n6655_1);
nor_5  g04307(n25797, new_n3560, new_n6656);
xor_4  g04308(n25797, n4957, new_n6657);
and_5  g04309(n15967, new_n5386_1, new_n6658);
nor_5  g04310(n15967, new_n5386_1, new_n6659_1);
nor_5  g04311(n15743, new_n3901, new_n6660);
or_5   g04312(new_n3567, n13319, new_n6661);
not_10 g04313(n25435, new_n6662);
nor_5  g04314(new_n6662, n20658, new_n6663);
and_5  g04315(new_n6663, new_n6661, new_n6664);
nor_5  g04316(new_n6664, new_n6660, new_n6665);
nor_5  g04317(new_n6665, new_n6659_1, new_n6666);
or_5   g04318(new_n6666, new_n6658, new_n6667);
nor_5  g04319(new_n6667, new_n6657, new_n6668);
nor_5  g04320(new_n6668, new_n6656, new_n6669_1);
nor_5  g04321(new_n6669_1, new_n6655_1, new_n6670);
nor_5  g04322(new_n6670, new_n6654, new_n6671_1);
nor_5  g04323(new_n6671_1, new_n6653, new_n6672);
nor_5  g04324(new_n6672, new_n6652_1, new_n6673_1);
nor_5  g04325(new_n6673_1, new_n6651, new_n6674_1);
nor_5  g04326(new_n6674_1, new_n6650, new_n6675);
nor_5  g04327(new_n6675, new_n6649, new_n6676);
nor_5  g04328(new_n6676, new_n6648, new_n6677);
nor_5  g04329(new_n6677, new_n6647, new_n6678);
nor_5  g04330(new_n6678, new_n6646, new_n6679);
nor_5  g04331(new_n6679, new_n6645, new_n6680);
nor_5  g04332(new_n6680, new_n6644, new_n6681);
not_10 g04333(new_n6681, new_n6682);
xnor_4 g04334(new_n6682, new_n6643, new_n6683);
xor_4  g04335(new_n6679, new_n6645, new_n6684_1);
xor_4  g04336(new_n6640, new_n6593, new_n6685);
nor_5  g04337(new_n6685, new_n6684_1, new_n6686);
xnor_4 g04338(new_n6685, new_n6684_1, new_n6687);
xnor_4 g04339(new_n6677, new_n6647, new_n6688);
xor_4  g04340(new_n6638, new_n6597, new_n6689);
and_5  g04341(new_n6689, new_n6688, new_n6690);
xnor_4 g04342(new_n6689, new_n6688, new_n6691_1);
xnor_4 g04343(new_n6675, new_n6649, new_n6692);
xor_4  g04344(new_n6636, new_n6601, new_n6693);
and_5  g04345(new_n6693, new_n6692, new_n6694);
xnor_4 g04346(new_n6693, new_n6692, new_n6695);
xnor_4 g04347(new_n6673_1, new_n6651, new_n6696);
xor_4  g04348(new_n6634_1, new_n6604, new_n6697);
and_5  g04349(new_n6697, new_n6696, new_n6698);
xnor_4 g04350(new_n6697, new_n6696, new_n6699);
xnor_4 g04351(new_n6671_1, new_n6653, new_n6700);
xor_4  g04352(new_n6632, new_n6607, new_n6701);
and_5  g04353(new_n6701, new_n6700, new_n6702);
xnor_4 g04354(new_n6701, new_n6700, new_n6703);
xnor_4 g04355(new_n6669_1, new_n6655_1, new_n6704);
xor_4  g04356(new_n6630_1, new_n6610, new_n6705);
and_5  g04357(new_n6705, new_n6704, new_n6706_1);
xnor_4 g04358(new_n6705, new_n6704, new_n6707_1);
xnor_4 g04359(new_n6628_1, new_n6613, new_n6708);
xor_4  g04360(new_n6667, new_n6657, new_n6709);
nor_5  g04361(new_n6709, new_n6708, new_n6710);
xnor_4 g04362(new_n6625, new_n6617, new_n6711);
xnor_4 g04363(n15967, n7524, new_n6712);
xnor_4 g04364(new_n6712, new_n6665, new_n6713);
and_5  g04365(new_n6713, new_n6711, new_n6714);
xnor_4 g04366(new_n6713, new_n6711, new_n6715);
xnor_4 g04367(n25435, n20658, new_n6716);
xnor_4 g04368(new_n6621, new_n3682, new_n6717);
or_5   g04369(new_n6717, new_n6716, new_n6718);
xor_4  g04370(n15743, n13319, new_n6719);
xnor_4 g04371(new_n6719, new_n6663, new_n6720);
and_5  g04372(new_n6720, new_n6718, new_n6721);
xnor_4 g04373(new_n6623, new_n6622, new_n6722);
xor_4  g04374(new_n6720, new_n6718, new_n6723);
and_5  g04375(new_n6723, new_n6722, new_n6724);
nor_5  g04376(new_n6724, new_n6721, new_n6725);
nor_5  g04377(new_n6725, new_n6715, new_n6726);
nor_5  g04378(new_n6726, new_n6714, new_n6727);
xnor_4 g04379(new_n6709, new_n6708, new_n6728);
nor_5  g04380(new_n6728, new_n6727, new_n6729_1);
nor_5  g04381(new_n6729_1, new_n6710, new_n6730);
nor_5  g04382(new_n6730, new_n6707_1, new_n6731);
nor_5  g04383(new_n6731, new_n6706_1, new_n6732);
nor_5  g04384(new_n6732, new_n6703, new_n6733);
nor_5  g04385(new_n6733, new_n6702, new_n6734);
nor_5  g04386(new_n6734, new_n6699, new_n6735);
nor_5  g04387(new_n6735, new_n6698, new_n6736_1);
nor_5  g04388(new_n6736_1, new_n6695, new_n6737);
nor_5  g04389(new_n6737, new_n6694, new_n6738);
nor_5  g04390(new_n6738, new_n6691_1, new_n6739);
nor_5  g04391(new_n6739, new_n6690, new_n6740);
nor_5  g04392(new_n6740, new_n6687, new_n6741);
nor_5  g04393(new_n6741, new_n6686, new_n6742);
xnor_4 g04394(new_n6742, new_n6683, n809);
not_10 g04395(n2978, new_n6744);
nor_5  g04396(n19282, new_n6744, new_n6745);
xor_4  g04397(n19282, n2978, new_n6746);
not_10 g04398(n23697, new_n6747);
nor_5  g04399(new_n6747, n12657, new_n6748);
xor_4  g04400(n23697, n12657, new_n6749);
not_10 g04401(n2289, new_n6750);
nor_5  g04402(n17077, new_n6750, new_n6751);
xor_4  g04403(n17077, n2289, new_n6752);
not_10 g04404(n1112, new_n6753);
nor_5  g04405(n26510, new_n6753, new_n6754);
xor_4  g04406(n26510, n1112, new_n6755);
not_10 g04407(n20179, new_n6756);
nor_5  g04408(n23068, new_n6756, new_n6757);
xor_4  g04409(n23068, n20179, new_n6758);
not_10 g04410(n19228, new_n6759);
nor_5  g04411(n19514, new_n6759, new_n6760);
xor_4  g04412(n19514, n19228, new_n6761);
not_10 g04413(n15539, new_n6762);
nor_5  g04414(new_n6762, n10053, new_n6763);
xor_4  g04415(n15539, n10053, new_n6764);
nor_5  g04416(new_n3594, n8052, new_n6765);
not_10 g04417(n8052, new_n6766);
nor_5  g04418(n8399, new_n6766, new_n6767);
nor_5  g04419(n10158, new_n3598, new_n6768);
not_10 g04420(n10158, new_n6769);
or_5   g04421(new_n6769, n9507, new_n6770);
nor_5  g04422(new_n3602, n18962, new_n6771);
and_5  g04423(new_n6771, new_n6770, new_n6772);
nor_5  g04424(new_n6772, new_n6768, new_n6773_1);
nor_5  g04425(new_n6773_1, new_n6767, new_n6774);
or_5   g04426(new_n6774, new_n6765, new_n6775_1);
nor_5  g04427(new_n6775_1, new_n6764, new_n6776);
nor_5  g04428(new_n6776, new_n6763, new_n6777);
nor_5  g04429(new_n6777, new_n6761, new_n6778);
nor_5  g04430(new_n6778, new_n6760, new_n6779);
nor_5  g04431(new_n6779, new_n6758, new_n6780);
nor_5  g04432(new_n6780, new_n6757, new_n6781);
nor_5  g04433(new_n6781, new_n6755, new_n6782);
nor_5  g04434(new_n6782, new_n6754, new_n6783);
nor_5  g04435(new_n6783, new_n6752, new_n6784);
nor_5  g04436(new_n6784, new_n6751, new_n6785_1);
nor_5  g04437(new_n6785_1, new_n6749, new_n6786);
nor_5  g04438(new_n6786, new_n6748, new_n6787);
nor_5  g04439(new_n6787, new_n6746, new_n6788);
nor_5  g04440(new_n6788, new_n6745, new_n6789);
nor_5  g04441(n26986, n22626, new_n6790_1);
not_10 g04442(new_n2415, new_n6791_1);
or_5   g04443(new_n6791_1, new_n2410, new_n6792);
xnor_4 g04444(n4256, n1654, new_n6793);
nor_5  g04445(n22332, n13783, new_n6794_1);
nor_5  g04446(new_n2414, new_n2411, new_n6795);
nor_5  g04447(new_n6795, new_n6794_1, new_n6796);
xnor_4 g04448(new_n6796, new_n6793, new_n6797);
or_5   g04449(new_n6797, new_n6792, new_n6798);
xnor_4 g04450(n21287, n14440, new_n6799);
nor_5  g04451(n4256, n1654, new_n6800);
nor_5  g04452(new_n6796, new_n6793, new_n6801);
nor_5  g04453(new_n6801, new_n6800, new_n6802_1);
xnor_4 g04454(new_n6802_1, new_n6799, new_n6803);
or_5   g04455(new_n6803, new_n6798, new_n6804);
xnor_4 g04456(n26986, n22626, new_n6805);
nor_5  g04457(n21287, n14440, new_n6806);
nor_5  g04458(new_n6802_1, new_n6799, new_n6807);
nor_5  g04459(new_n6807, new_n6806, new_n6808);
xnor_4 g04460(new_n6808, new_n6805, new_n6809);
nor_5  g04461(new_n6809, new_n6804, new_n6810);
and_5  g04462(new_n6810, new_n6790_1, new_n6811);
nor_5  g04463(new_n6808, new_n6805, new_n6812);
or_5   g04464(new_n6812, new_n6790_1, new_n6813);
nor_5  g04465(new_n6813, new_n6810, new_n6814_1);
nor_5  g04466(new_n6814_1, new_n6811, new_n6815);
nor_5  g04467(n13494, n3425, new_n6816);
xnor_4 g04468(n13494, n3425, new_n6817);
nor_5  g04469(n25345, n9967, new_n6818);
xor_4  g04470(n25345, n9967, new_n6819);
and_5  g04471(n20946, n9655, new_n6820);
or_5   g04472(n20946, n9655, new_n6821);
nor_5  g04473(n13490, n7751, new_n6822);
nor_5  g04474(new_n2438, new_n2417, new_n6823);
nor_5  g04475(new_n6823, new_n6822, new_n6824);
and_5  g04476(new_n6824, new_n6821, new_n6825);
nor_5  g04477(new_n6825, new_n6820, new_n6826_1);
and_5  g04478(new_n6826_1, new_n6819, new_n6827);
nor_5  g04479(new_n6827, new_n6818, new_n6828);
nor_5  g04480(new_n6828, new_n6817, new_n6829);
nor_5  g04481(new_n6829, new_n6816, new_n6830);
and_5  g04482(new_n6830, new_n6815, new_n6831);
or_5   g04483(new_n6830, new_n6815, new_n6832);
xor_4  g04484(new_n6809, new_n6804, new_n6833);
xor_4  g04485(new_n6828, new_n6817, new_n6834);
not_10 g04486(new_n6834, new_n6835_1);
nor_5  g04487(new_n6835_1, new_n6833, new_n6836);
xnor_4 g04488(new_n6835_1, new_n6833, new_n6837);
xor_4  g04489(new_n6803, new_n6798, new_n6838);
xor_4  g04490(new_n6826_1, new_n6819, new_n6839);
not_10 g04491(new_n6839, new_n6840);
nor_5  g04492(new_n6840, new_n6838, new_n6841);
xnor_4 g04493(new_n6840, new_n6838, new_n6842);
xor_4  g04494(new_n6797, new_n6792, new_n6843);
xnor_4 g04495(n20946, n9655, new_n6844);
xnor_4 g04496(new_n6844, new_n6824, new_n6845);
nor_5  g04497(new_n6845, new_n6843, new_n6846);
xnor_4 g04498(new_n6845, new_n6843, new_n6847);
nor_5  g04499(new_n2440_1, new_n2416_1, new_n6848);
nor_5  g04500(new_n2484, new_n2441, new_n6849);
nor_5  g04501(new_n6849, new_n6848, new_n6850);
nor_5  g04502(new_n6850, new_n6847, new_n6851);
nor_5  g04503(new_n6851, new_n6846, new_n6852);
nor_5  g04504(new_n6852, new_n6842, new_n6853_1);
nor_5  g04505(new_n6853_1, new_n6841, new_n6854);
nor_5  g04506(new_n6854, new_n6837, new_n6855);
nor_5  g04507(new_n6855, new_n6836, new_n6856);
and_5  g04508(new_n6856, new_n6832, new_n6857);
or_5   g04509(new_n6857, new_n6811, new_n6858);
nor_5  g04510(new_n6858, new_n6831, new_n6859);
xnor_4 g04511(new_n6859, new_n6789, new_n6860);
xnor_4 g04512(new_n6830, new_n6815, new_n6861_1);
xnor_4 g04513(new_n6861_1, new_n6856, new_n6862_1);
nor_5  g04514(new_n6862_1, new_n6789, new_n6863_1);
xnor_4 g04515(new_n6862_1, new_n6789, new_n6864);
xnor_4 g04516(new_n6787, new_n6746, new_n6865);
xor_4  g04517(new_n6854, new_n6837, new_n6866);
and_5  g04518(new_n6866, new_n6865, new_n6867_1);
xnor_4 g04519(new_n6866, new_n6865, new_n6868);
xnor_4 g04520(new_n6785_1, new_n6749, new_n6869);
xor_4  g04521(new_n6852, new_n6842, new_n6870);
and_5  g04522(new_n6870, new_n6869, new_n6871);
xnor_4 g04523(new_n6870, new_n6869, new_n6872);
xnor_4 g04524(new_n6783, new_n6752, new_n6873);
xor_4  g04525(new_n6850, new_n6847, new_n6874);
and_5  g04526(new_n6874, new_n6873, new_n6875);
xnor_4 g04527(new_n6874, new_n6873, new_n6876);
not_10 g04528(new_n2485, new_n6877);
xor_4  g04529(new_n6781, new_n6755, new_n6878);
nor_5  g04530(new_n6878, new_n6877, new_n6879);
xor_4  g04531(new_n6878, new_n2485, new_n6880);
not_10 g04532(new_n2488, new_n6881);
xor_4  g04533(new_n6779, new_n6758, new_n6882);
nor_5  g04534(new_n6882, new_n6881, new_n6883);
xor_4  g04535(new_n6882, new_n2488, new_n6884);
not_10 g04536(new_n2492, new_n6885);
xor_4  g04537(new_n6777, new_n6761, new_n6886);
nor_5  g04538(new_n6886, new_n6885, new_n6887);
xor_4  g04539(new_n6886, new_n2492, new_n6888);
not_10 g04540(new_n2496, new_n6889);
xor_4  g04541(new_n6775_1, new_n6764, new_n6890);
nor_5  g04542(new_n6890, new_n6889, new_n6891);
xor_4  g04543(new_n6890, new_n2496, new_n6892);
xnor_4 g04544(n8399, n8052, new_n6893);
xnor_4 g04545(new_n6893, new_n6773_1, new_n6894);
and_5  g04546(new_n6894, new_n2499, new_n6895);
xnor_4 g04547(new_n6894, new_n2499, new_n6896);
xnor_4 g04548(n26979, n18962, new_n6897);
or_5   g04549(new_n6897, new_n2505, new_n6898);
xor_4  g04550(n10158, n9507, new_n6899);
xnor_4 g04551(new_n6899, new_n6771, new_n6900);
and_5  g04552(new_n6900, new_n6898, new_n6901);
xor_4  g04553(new_n6900, new_n6898, new_n6902);
and_5  g04554(new_n6902, new_n2510, new_n6903);
nor_5  g04555(new_n6903, new_n6901, new_n6904);
nor_5  g04556(new_n6904, new_n6896, new_n6905);
nor_5  g04557(new_n6905, new_n6895, new_n6906);
nor_5  g04558(new_n6906, new_n6892, new_n6907);
nor_5  g04559(new_n6907, new_n6891, new_n6908);
nor_5  g04560(new_n6908, new_n6888, new_n6909);
nor_5  g04561(new_n6909, new_n6887, new_n6910);
nor_5  g04562(new_n6910, new_n6884, new_n6911);
nor_5  g04563(new_n6911, new_n6883, new_n6912);
nor_5  g04564(new_n6912, new_n6880, new_n6913);
nor_5  g04565(new_n6913, new_n6879, new_n6914);
nor_5  g04566(new_n6914, new_n6876, new_n6915);
nor_5  g04567(new_n6915, new_n6875, new_n6916);
nor_5  g04568(new_n6916, new_n6872, new_n6917);
nor_5  g04569(new_n6917, new_n6871, new_n6918);
nor_5  g04570(new_n6918, new_n6868, new_n6919);
nor_5  g04571(new_n6919, new_n6867_1, new_n6920);
nor_5  g04572(new_n6920, new_n6864, new_n6921);
nor_5  g04573(new_n6921, new_n6863_1, new_n6922);
xnor_4 g04574(new_n6922, new_n6860, n819);
not_10 g04575(n8856, new_n6924);
nor_5  g04576(n22626, new_n6924, new_n6925);
xor_4  g04577(n22626, n8856, new_n6926);
not_10 g04578(n14130, new_n6927);
nor_5  g04579(n14440, new_n6927, new_n6928);
xor_4  g04580(n14440, n14130, new_n6929);
not_10 g04581(n16482, new_n6930);
nor_5  g04582(new_n6930, n1654, new_n6931);
xor_4  g04583(n16482, n1654, new_n6932);
not_10 g04584(n9942, new_n6933);
nor_5  g04585(n13783, new_n6933, new_n6934);
xor_4  g04586(n13783, n9942, new_n6935);
not_10 g04587(n25643, new_n6936);
nor_5  g04588(n26660, new_n6936, new_n6937);
xor_4  g04589(n26660, n25643, new_n6938);
not_10 g04590(n3018, new_n6939);
and_5  g04591(n9557, new_n6939, new_n6940);
xor_4  g04592(n9557, n3018, new_n6941);
not_10 g04593(n3136, new_n6942);
nor_5  g04594(n3480, new_n6942, new_n6943);
xor_4  g04595(n3480, n3136, new_n6944);
not_10 g04596(n16722, new_n6945);
nor_5  g04597(new_n6945, n6385, new_n6946);
nor_5  g04598(n16722, new_n2359, new_n6947);
not_10 g04599(n11486, new_n6948);
nor_5  g04600(n20138, new_n6948, new_n6949);
or_5   g04601(new_n2362, n11486, new_n6950);
not_10 g04602(n13781, new_n6951);
nor_5  g04603(new_n6951, n9251, new_n6952);
and_5  g04604(new_n6952, new_n6950, new_n6953);
nor_5  g04605(new_n6953, new_n6949, new_n6954);
nor_5  g04606(new_n6954, new_n6947, new_n6955);
or_5   g04607(new_n6955, new_n6946, new_n6956);
nor_5  g04608(new_n6956, new_n6944, new_n6957);
nor_5  g04609(new_n6957, new_n6943, new_n6958);
nor_5  g04610(new_n6958, new_n6941, new_n6959);
nor_5  g04611(new_n6959, new_n6940, new_n6960);
nor_5  g04612(new_n6960, new_n6938, new_n6961);
nor_5  g04613(new_n6961, new_n6937, new_n6962);
nor_5  g04614(new_n6962, new_n6935, new_n6963);
nor_5  g04615(new_n6963, new_n6934, new_n6964);
nor_5  g04616(new_n6964, new_n6932, new_n6965_1);
nor_5  g04617(new_n6965_1, new_n6931, new_n6966);
nor_5  g04618(new_n6966, new_n6929, new_n6967_1);
nor_5  g04619(new_n6967_1, new_n6928, new_n6968);
nor_5  g04620(new_n6968, new_n6926, new_n6969);
nor_5  g04621(new_n6969, new_n6925, new_n6970);
not_10 g04622(n25120, new_n6971_1);
and_5  g04623(new_n6971_1, n3582, new_n6972);
xor_4  g04624(n25120, n3582, new_n6973);
not_10 g04625(n8363, new_n6974);
and_5  g04626(new_n6974, n2145, new_n6975_1);
xor_4  g04627(n8363, n2145, new_n6976);
not_10 g04628(n14680, new_n6977);
and_5  g04629(new_n6977, n5031, new_n6978);
xor_4  g04630(n14680, n5031, new_n6979);
not_10 g04631(n17250, new_n6980);
and_5  g04632(new_n6980, n11044, new_n6981);
xor_4  g04633(n17250, n11044, new_n6982);
not_10 g04634(n23160, new_n6983_1);
and_5  g04635(new_n6983_1, n2421, new_n6984);
xor_4  g04636(n23160, n2421, new_n6985_1);
not_10 g04637(n16524, new_n6986);
nand_5 g04638(new_n6986, n987, new_n6987);
xor_4  g04639(n16524, n987, new_n6988);
not_10 g04640(n20478, new_n6989);
or_5   g04641(new_n6989, n11056, new_n6990);
xor_4  g04642(n20478, n11056, new_n6991);
not_10 g04643(n26882, new_n6992);
and_5  g04644(new_n6992, n15271, new_n6993);
nor_5  g04645(new_n6992, n15271, new_n6994);
not_10 g04646(n22619, new_n6995);
and_5  g04647(n25877, new_n6995, new_n6996);
or_5   g04648(n25877, new_n6995, new_n6997);
not_10 g04649(n24323, new_n6998_1);
nor_5  g04650(new_n6998_1, n6775, new_n6999);
and_5  g04651(new_n6999, new_n6997, new_n7000);
nor_5  g04652(new_n7000, new_n6996, new_n7001);
nor_5  g04653(new_n7001, new_n6994, new_n7002);
nor_5  g04654(new_n7002, new_n6993, new_n7003);
not_10 g04655(new_n7003, new_n7004);
or_5   g04656(new_n7004, new_n6991, new_n7005);
and_5  g04657(new_n7005, new_n6990, new_n7006);
or_5   g04658(new_n7006, new_n6988, new_n7007);
and_5  g04659(new_n7007, new_n6987, new_n7008);
nor_5  g04660(new_n7008, new_n6985_1, new_n7009);
nor_5  g04661(new_n7009, new_n6984, new_n7010);
nor_5  g04662(new_n7010, new_n6982, new_n7011);
nor_5  g04663(new_n7011, new_n6981, new_n7012);
nor_5  g04664(new_n7012, new_n6979, new_n7013);
nor_5  g04665(new_n7013, new_n6978, new_n7014);
nor_5  g04666(new_n7014, new_n6976, new_n7015);
nor_5  g04667(new_n7015, new_n6975_1, new_n7016);
nor_5  g04668(new_n7016, new_n6973, new_n7017);
nor_5  g04669(new_n7017, new_n6972, new_n7018);
xnor_4 g04670(new_n7018, new_n6970, new_n7019);
xor_4  g04671(new_n7016, new_n6973, new_n7020);
xor_4  g04672(new_n6968, new_n6926, new_n7021);
nor_5  g04673(new_n7021, new_n7020, new_n7022);
xnor_4 g04674(new_n7021, new_n7020, new_n7023);
xor_4  g04675(new_n7014, new_n6976, new_n7024);
xor_4  g04676(new_n6966, new_n6929, new_n7025);
nor_5  g04677(new_n7025, new_n7024, new_n7026_1);
xnor_4 g04678(new_n7025, new_n7024, new_n7027);
xor_4  g04679(new_n7012, new_n6979, new_n7028);
xor_4  g04680(new_n6964, new_n6932, new_n7029);
nor_5  g04681(new_n7029, new_n7028, new_n7030);
xnor_4 g04682(new_n7029, new_n7028, new_n7031);
xor_4  g04683(new_n7010, new_n6982, new_n7032_1);
xor_4  g04684(new_n6962, new_n6935, new_n7033);
nor_5  g04685(new_n7033, new_n7032_1, new_n7034);
xnor_4 g04686(new_n7033, new_n7032_1, new_n7035);
xor_4  g04687(new_n7008, new_n6985_1, new_n7036);
xor_4  g04688(new_n6960, new_n6938, new_n7037);
nor_5  g04689(new_n7037, new_n7036, new_n7038_1);
xnor_4 g04690(new_n7037, new_n7036, new_n7039);
xor_4  g04691(new_n7006, new_n6988, new_n7040);
xor_4  g04692(new_n6958, new_n6941, new_n7041);
nor_5  g04693(new_n7041, new_n7040, new_n7042);
xnor_4 g04694(new_n7041, new_n7040, new_n7043);
xnor_4 g04695(new_n7003, new_n6991, new_n7044);
xor_4  g04696(new_n6956, new_n6944, new_n7045);
nor_5  g04697(new_n7045, new_n7044, new_n7046);
xnor_4 g04698(new_n7045, new_n7044, new_n7047);
xnor_4 g04699(n26882, n15271, new_n7048);
xnor_4 g04700(new_n7048, new_n7001, new_n7049);
xnor_4 g04701(n16722, n6385, new_n7050);
xnor_4 g04702(new_n7050, new_n6954, new_n7051);
and_5  g04703(new_n7051, new_n7049, new_n7052);
xnor_4 g04704(new_n7051, new_n7049, new_n7053);
xor_4  g04705(n25877, n22619, new_n7054);
xnor_4 g04706(new_n7054, new_n6999, new_n7055);
xor_4  g04707(n20138, n11486, new_n7056);
xnor_4 g04708(new_n7056, new_n6952, new_n7057_1);
and_5  g04709(new_n7057_1, new_n7055, new_n7058);
xnor_4 g04710(n24323, n6775, new_n7059);
xnor_4 g04711(n13781, n9251, new_n7060);
or_5   g04712(new_n7060, new_n7059, new_n7061);
xor_4  g04713(new_n7057_1, new_n7055, new_n7062);
and_5  g04714(new_n7062, new_n7061, new_n7063);
nor_5  g04715(new_n7063, new_n7058, new_n7064);
nor_5  g04716(new_n7064, new_n7053, new_n7065);
nor_5  g04717(new_n7065, new_n7052, new_n7066);
nor_5  g04718(new_n7066, new_n7047, new_n7067);
nor_5  g04719(new_n7067, new_n7046, new_n7068);
nor_5  g04720(new_n7068, new_n7043, new_n7069);
nor_5  g04721(new_n7069, new_n7042, new_n7070);
nor_5  g04722(new_n7070, new_n7039, new_n7071);
nor_5  g04723(new_n7071, new_n7038_1, new_n7072);
nor_5  g04724(new_n7072, new_n7035, new_n7073);
nor_5  g04725(new_n7073, new_n7034, new_n7074);
nor_5  g04726(new_n7074, new_n7031, new_n7075);
nor_5  g04727(new_n7075, new_n7030, new_n7076);
nor_5  g04728(new_n7076, new_n7027, new_n7077);
nor_5  g04729(new_n7077, new_n7026_1, new_n7078);
nor_5  g04730(new_n7078, new_n7023, new_n7079_1);
nor_5  g04731(new_n7079_1, new_n7022, new_n7080);
xnor_4 g04732(new_n7080, new_n7019, new_n7081);
or_5   g04733(n15508, n2809, new_n7082);
or_5   g04734(new_n7082, n19680, new_n7083);
or_5   g04735(new_n7083, n7421, new_n7084);
or_5   g04736(new_n7084, n13453, new_n7085);
or_5   g04737(new_n7085, n11630, new_n7086);
or_5   g04738(new_n7086, n7377, new_n7087);
or_5   g04739(new_n7087, n18227, new_n7088);
or_5   g04740(new_n7088, n26408, new_n7089);
nor_5  g04741(new_n7089, n9554, new_n7090);
xor_4  g04742(new_n7089, n9554, new_n7091);
nor_5  g04743(new_n7091, n9259, new_n7092);
xor_4  g04744(new_n7088, n26408, new_n7093);
nor_5  g04745(new_n7093, n21489, new_n7094);
xnor_4 g04746(new_n7093, n21489, new_n7095);
xor_4  g04747(new_n7087, n18227, new_n7096);
nor_5  g04748(new_n7096, n20213, new_n7097);
xnor_4 g04749(new_n7096, n20213, new_n7098);
xor_4  g04750(new_n7086, n7377, new_n7099_1);
nor_5  g04751(new_n7099_1, n13912, new_n7100);
xnor_4 g04752(new_n7099_1, n13912, new_n7101);
xor_4  g04753(new_n7085, n11630, new_n7102);
nor_5  g04754(new_n7102, n7670, new_n7103);
xnor_4 g04755(new_n7102, n7670, new_n7104);
xor_4  g04756(new_n7084, n13453, new_n7105);
nor_5  g04757(new_n7105, n9598, new_n7106);
xnor_4 g04758(new_n7105, n9598, new_n7107);
xor_4  g04759(new_n7083, n7421, new_n7108);
nor_5  g04760(new_n7108, n22290, new_n7109);
xor_4  g04761(new_n7082, n19680, new_n7110);
nor_5  g04762(new_n7110, n11273, new_n7111);
xnor_4 g04763(new_n7110, n11273, new_n7112);
xor_4  g04764(n15508, n2809, new_n7113);
nor_5  g04765(new_n7113, n25565, new_n7114);
nand_5 g04766(n21993, n15508, new_n7115);
xor_4  g04767(new_n7113, n25565, new_n7116);
and_5  g04768(new_n7116, new_n7115, new_n7117);
nor_5  g04769(new_n7117, new_n7114, new_n7118);
nor_5  g04770(new_n7118, new_n7112, new_n7119);
nor_5  g04771(new_n7119, new_n7111, new_n7120);
xnor_4 g04772(new_n7108, n22290, new_n7121);
nor_5  g04773(new_n7121, new_n7120, new_n7122);
nor_5  g04774(new_n7122, new_n7109, new_n7123);
nor_5  g04775(new_n7123, new_n7107, new_n7124);
nor_5  g04776(new_n7124, new_n7106, new_n7125);
nor_5  g04777(new_n7125, new_n7104, new_n7126);
nor_5  g04778(new_n7126, new_n7103, new_n7127);
nor_5  g04779(new_n7127, new_n7101, new_n7128);
nor_5  g04780(new_n7128, new_n7100, new_n7129);
nor_5  g04781(new_n7129, new_n7098, new_n7130);
nor_5  g04782(new_n7130, new_n7097, new_n7131);
nor_5  g04783(new_n7131, new_n7095, new_n7132);
nor_5  g04784(new_n7132, new_n7094, new_n7133);
and_5  g04785(new_n7091, n9259, new_n7134);
nor_5  g04786(new_n7134, new_n7133, new_n7135);
nor_5  g04787(new_n7135, new_n7092, new_n7136);
nor_5  g04788(new_n7136, new_n7090, new_n7137);
xnor_4 g04789(new_n7137, new_n7081, new_n7138);
xnor_4 g04790(new_n7078, new_n7023, new_n7139_1);
xnor_4 g04791(new_n7091, n9259, new_n7140);
xnor_4 g04792(new_n7140, new_n7133, new_n7141);
nor_5  g04793(new_n7141, new_n7139_1, new_n7142);
xor_4  g04794(new_n7141, new_n7139_1, new_n7143);
xnor_4 g04795(new_n7076, new_n7027, new_n7144);
xor_4  g04796(new_n7131, new_n7095, new_n7145);
not_10 g04797(new_n7145, new_n7146);
and_5  g04798(new_n7146, new_n7144, new_n7147);
xnor_4 g04799(new_n7146, new_n7144, new_n7148);
xnor_4 g04800(new_n7074, new_n7031, new_n7149_1);
xor_4  g04801(new_n7129, new_n7098, new_n7150);
not_10 g04802(new_n7150, new_n7151);
and_5  g04803(new_n7151, new_n7149_1, new_n7152);
xnor_4 g04804(new_n7151, new_n7149_1, new_n7153);
xnor_4 g04805(new_n7072, new_n7035, new_n7154);
xnor_4 g04806(new_n7127, new_n7101, new_n7155);
nor_5  g04807(new_n7155, new_n7154, new_n7156);
and_5  g04808(new_n7155, new_n7154, new_n7157);
xnor_4 g04809(new_n7070, new_n7039, new_n7158);
xor_4  g04810(new_n7125, new_n7104, new_n7159);
not_10 g04811(new_n7159, new_n7160);
nor_5  g04812(new_n7160, new_n7158, new_n7161);
xnor_4 g04813(new_n7160, new_n7158, new_n7162);
xor_4  g04814(new_n7123, new_n7107, new_n7163);
not_10 g04815(new_n7163, new_n7164);
xnor_4 g04816(new_n7068, new_n7043, new_n7165);
nor_5  g04817(new_n7165, new_n7164, new_n7166);
xnor_4 g04818(new_n7165, new_n7164, new_n7167);
xnor_4 g04819(new_n7066, new_n7047, new_n7168);
xor_4  g04820(new_n7121, new_n7120, new_n7169);
not_10 g04821(new_n7169, new_n7170);
nor_5  g04822(new_n7170, new_n7168, new_n7171);
nand_5 g04823(new_n7170, new_n7168, new_n7172);
xor_4  g04824(new_n7064, new_n7053, new_n7173);
xor_4  g04825(new_n7062, new_n7061, new_n7174);
and_5  g04826(n21993, n15508, new_n7175);
xnor_4 g04827(new_n7116, new_n7175, new_n7176);
and_5  g04828(new_n7176, new_n7174, new_n7177);
xnor_4 g04829(n21993, n15508, new_n7178);
xnor_4 g04830(new_n7060, new_n7059, new_n7179);
or_5   g04831(new_n7179, new_n7178, new_n7180);
xor_4  g04832(new_n7176, new_n7174, new_n7181);
and_5  g04833(new_n7181, new_n7180, new_n7182);
or_5   g04834(new_n7182, new_n7177, new_n7183);
nor_5  g04835(new_n7183, new_n7173, new_n7184);
xnor_4 g04836(new_n7118, new_n7112, new_n7185);
xor_4  g04837(new_n7183, new_n7173, new_n7186);
and_5  g04838(new_n7186, new_n7185, new_n7187);
nor_5  g04839(new_n7187, new_n7184, new_n7188);
and_5  g04840(new_n7188, new_n7172, new_n7189);
nor_5  g04841(new_n7189, new_n7171, new_n7190_1);
nor_5  g04842(new_n7190_1, new_n7167, new_n7191);
nor_5  g04843(new_n7191, new_n7166, new_n7192);
nor_5  g04844(new_n7192, new_n7162, new_n7193);
nor_5  g04845(new_n7193, new_n7161, new_n7194);
nor_5  g04846(new_n7194, new_n7157, new_n7195);
or_5   g04847(new_n7195, new_n7156, new_n7196);
nor_5  g04848(new_n7196, new_n7153, new_n7197);
nor_5  g04849(new_n7197, new_n7152, new_n7198);
nor_5  g04850(new_n7198, new_n7148, new_n7199);
nor_5  g04851(new_n7199, new_n7147, new_n7200);
and_5  g04852(new_n7200, new_n7143, new_n7201);
or_5   g04853(new_n7201, new_n7142, new_n7202);
xor_4  g04854(new_n7202, new_n7138, n829);
not_10 g04855(n22764, new_n7204);
xnor_4 g04856(n23272, n14826, new_n7205);
nor_5  g04857(n23493, n11481, new_n7206);
xnor_4 g04858(n23493, n11481, new_n7207);
nor_5  g04859(n16439, n10275, new_n7208);
xnor_4 g04860(n16439, n10275, new_n7209);
nor_5  g04861(n15241, n15146, new_n7210);
xnor_4 g04862(n15241, n15146, new_n7211);
nor_5  g04863(n11579, n7678, new_n7212);
xnor_4 g04864(n11579, n7678, new_n7213);
nor_5  g04865(n3785, n21, new_n7214);
xnor_4 g04866(n3785, n21, new_n7215);
nor_5  g04867(n20250, n1682, new_n7216);
xnor_4 g04868(n20250, n1682, new_n7217);
nor_5  g04869(n7963, n5822, new_n7218);
xnor_4 g04870(n7963, n5822, new_n7219);
nor_5  g04871(n26443, n10017, new_n7220);
and_5  g04872(n3618, n1681, new_n7221);
xnor_4 g04873(n26443, n10017, new_n7222);
nor_5  g04874(new_n7222, new_n7221, new_n7223);
nor_5  g04875(new_n7223, new_n7220, new_n7224);
nor_5  g04876(new_n7224, new_n7219, new_n7225);
nor_5  g04877(new_n7225, new_n7218, new_n7226);
nor_5  g04878(new_n7226, new_n7217, new_n7227);
nor_5  g04879(new_n7227, new_n7216, new_n7228);
nor_5  g04880(new_n7228, new_n7215, new_n7229_1);
nor_5  g04881(new_n7229_1, new_n7214, new_n7230_1);
nor_5  g04882(new_n7230_1, new_n7213, new_n7231);
nor_5  g04883(new_n7231, new_n7212, new_n7232);
nor_5  g04884(new_n7232, new_n7211, new_n7233_1);
nor_5  g04885(new_n7233_1, new_n7210, new_n7234);
nor_5  g04886(new_n7234, new_n7209, new_n7235);
nor_5  g04887(new_n7235, new_n7208, new_n7236_1);
nor_5  g04888(new_n7236_1, new_n7207, new_n7237);
nor_5  g04889(new_n7237, new_n7206, new_n7238);
xnor_4 g04890(new_n7238, new_n7205, new_n7239);
and_5  g04891(new_n7239, new_n7204, new_n7240);
xor_4  g04892(new_n7239, n22764, new_n7241);
not_10 g04893(n26264, new_n7242);
xnor_4 g04894(new_n7236_1, new_n7207, new_n7243);
and_5  g04895(new_n7243, new_n7242, new_n7244);
xor_4  g04896(new_n7243, n26264, new_n7245);
not_10 g04897(n7841, new_n7246);
xnor_4 g04898(new_n7234, new_n7209, new_n7247);
and_5  g04899(new_n7247, new_n7246, new_n7248);
xor_4  g04900(new_n7247, n7841, new_n7249);
not_10 g04901(n16812, new_n7250);
xnor_4 g04902(new_n7232, new_n7211, new_n7251);
and_5  g04903(new_n7251, new_n7250, new_n7252);
xor_4  g04904(new_n7251, n16812, new_n7253_1);
not_10 g04905(n25068, new_n7254);
xnor_4 g04906(new_n7230_1, new_n7213, new_n7255);
and_5  g04907(new_n7255, new_n7254, new_n7256_1);
xor_4  g04908(new_n7255, n25068, new_n7257);
not_10 g04909(n2331, new_n7258);
xnor_4 g04910(new_n7228, new_n7215, new_n7259);
and_5  g04911(new_n7259, new_n7258, new_n7260);
xor_4  g04912(new_n7259, n2331, new_n7261);
not_10 g04913(n22631, new_n7262);
xnor_4 g04914(new_n7226, new_n7217, new_n7263);
nand_5 g04915(new_n7263, new_n7262, new_n7264);
xor_4  g04916(new_n7263, n22631, new_n7265);
not_10 g04917(n16743, new_n7266);
xnor_4 g04918(new_n7224, new_n7219, new_n7267);
nor_5  g04919(new_n7267, new_n7266, new_n7268_1);
xor_4  g04920(new_n7267, n16743, new_n7269);
not_10 g04921(n15258, new_n7270);
nor_5  g04922(new_n2523, n4588, new_n7271);
and_5  g04923(new_n7271, new_n7270, new_n7272);
xor_4  g04924(new_n7222, new_n7221, new_n7273);
not_10 g04925(new_n7273, new_n7274);
xnor_4 g04926(new_n7271, n15258, new_n7275);
and_5  g04927(new_n7275, new_n7274, new_n7276);
or_5   g04928(new_n7276, new_n7272, new_n7277_1);
nor_5  g04929(new_n7277_1, new_n7269, new_n7278);
nor_5  g04930(new_n7278, new_n7268_1, new_n7279);
not_10 g04931(new_n7279, new_n7280_1);
or_5   g04932(new_n7280_1, new_n7265, new_n7281);
and_5  g04933(new_n7281, new_n7264, new_n7282);
nor_5  g04934(new_n7282, new_n7261, new_n7283);
nor_5  g04935(new_n7283, new_n7260, new_n7284);
nor_5  g04936(new_n7284, new_n7257, new_n7285);
nor_5  g04937(new_n7285, new_n7256_1, new_n7286);
nor_5  g04938(new_n7286, new_n7253_1, new_n7287);
nor_5  g04939(new_n7287, new_n7252, new_n7288);
nor_5  g04940(new_n7288, new_n7249, new_n7289);
nor_5  g04941(new_n7289, new_n7248, new_n7290);
nor_5  g04942(new_n7290, new_n7245, new_n7291);
nor_5  g04943(new_n7291, new_n7244, new_n7292);
nor_5  g04944(new_n7292, new_n7241, new_n7293);
nor_5  g04945(new_n7293, new_n7240, new_n7294);
nor_5  g04946(n23272, n14826, new_n7295);
nor_5  g04947(new_n7238, new_n7205, new_n7296);
nor_5  g04948(new_n7296, new_n7295, new_n7297);
not_10 g04949(new_n7297, new_n7298_1);
and_5  g04950(new_n7298_1, new_n7294, new_n7299);
nor_5  g04951(n18105, new_n5231, new_n7300);
xor_4  g04952(n18105, n12702, new_n7301);
not_10 g04953(n26797, new_n7302);
nor_5  g04954(new_n7302, n24196, new_n7303);
xor_4  g04955(n26797, n24196, new_n7304);
not_10 g04956(n23913, new_n7305_1);
nor_5  g04957(new_n7305_1, n16376, new_n7306);
xor_4  g04958(n23913, n16376, new_n7307);
not_10 g04959(n22554, new_n7308_1);
nor_5  g04960(n25381, new_n7308_1, new_n7309);
xor_4  g04961(n25381, n22554, new_n7310);
not_10 g04962(n20429, new_n7311);
nor_5  g04963(new_n7311, n12587, new_n7312);
xor_4  g04964(n20429, n12587, new_n7313_1);
not_10 g04965(n3909, new_n7314);
nor_5  g04966(new_n7314, n268, new_n7315);
xor_4  g04967(n3909, n268, new_n7316);
not_10 g04968(n23974, new_n7317);
nor_5  g04969(n24879, new_n7317, new_n7318);
xor_4  g04970(n24879, n23974, new_n7319);
nor_5  g04971(new_n4137, n2146, new_n7320);
and_5  g04972(new_n4137, n2146, new_n7321);
not_10 g04973(n24032, new_n7322);
nor_5  g04974(new_n7322, n22173, new_n7323);
not_10 g04975(n22843, new_n7324);
nor_5  g04976(new_n7324, n583, new_n7325);
nand_5 g04977(new_n7322, n22173, new_n7326);
and_5  g04978(new_n7326, new_n7325, new_n7327);
nor_5  g04979(new_n7327, new_n7323, new_n7328);
nor_5  g04980(new_n7328, new_n7321, new_n7329);
or_5   g04981(new_n7329, new_n7320, new_n7330_1);
nor_5  g04982(new_n7330_1, new_n7319, new_n7331);
nor_5  g04983(new_n7331, new_n7318, new_n7332);
nor_5  g04984(new_n7332, new_n7316, new_n7333);
nor_5  g04985(new_n7333, new_n7315, new_n7334);
nor_5  g04986(new_n7334, new_n7313_1, new_n7335_1);
nor_5  g04987(new_n7335_1, new_n7312, new_n7336);
nor_5  g04988(new_n7336, new_n7310, new_n7337);
nor_5  g04989(new_n7337, new_n7309, new_n7338);
nor_5  g04990(new_n7338, new_n7307, new_n7339_1);
nor_5  g04991(new_n7339_1, new_n7306, new_n7340);
nor_5  g04992(new_n7340, new_n7304, new_n7341);
nor_5  g04993(new_n7341, new_n7303, new_n7342);
nor_5  g04994(new_n7342, new_n7301, new_n7343);
or_5   g04995(new_n7343, new_n7300, new_n7344);
xor_4  g04996(new_n7342, new_n7301, new_n7345);
nor_5  g04997(new_n7345, n1536, new_n7346_1);
xnor_4 g04998(new_n7345, n1536, new_n7347);
xor_4  g04999(new_n7340, new_n7304, new_n7348);
nor_5  g05000(new_n7348, n19454, new_n7349_1);
xnor_4 g05001(new_n7348, n19454, new_n7350);
xor_4  g05002(new_n7338, new_n7307, new_n7351);
nor_5  g05003(new_n7351, n9445, new_n7352);
xnor_4 g05004(new_n7351, n9445, new_n7353);
xor_4  g05005(new_n7336, new_n7310, new_n7354);
nor_5  g05006(new_n7354, n1279, new_n7355);
xnor_4 g05007(new_n7354, n1279, new_n7356);
xor_4  g05008(new_n7334, new_n7313_1, new_n7357);
nor_5  g05009(new_n7357, n8324, new_n7358);
xnor_4 g05010(new_n7357, n8324, new_n7359);
xor_4  g05011(new_n7332, new_n7316, new_n7360);
nor_5  g05012(new_n7360, n12546, new_n7361);
xnor_4 g05013(new_n7360, n12546, new_n7362);
xor_4  g05014(new_n7330_1, new_n7319, new_n7363_1);
nor_5  g05015(new_n7363_1, n21078, new_n7364);
xnor_4 g05016(new_n7363_1, n21078, new_n7365);
xnor_4 g05017(n6785, n2146, new_n7366);
xnor_4 g05018(new_n7366, new_n7328, new_n7367);
not_10 g05019(new_n7367, new_n7368);
and_5  g05020(new_n7368, n24485, new_n7369);
nor_5  g05021(new_n7368, n24485, new_n7370);
xor_4  g05022(n24032, n22173, new_n7371);
xnor_4 g05023(new_n7371, new_n7325, new_n7372);
not_10 g05024(new_n7372, new_n7373);
nor_5  g05025(new_n7373, n2420, new_n7374);
not_10 g05026(new_n2525, new_n7375);
nand_5 g05027(new_n7375, n22201, new_n7376);
xnor_4 g05028(new_n7372, n2420, new_n7377_1);
and_5  g05029(new_n7377_1, new_n7376, new_n7378);
or_5   g05030(new_n7378, new_n7374, new_n7379);
nor_5  g05031(new_n7379, new_n7370, new_n7380);
or_5   g05032(new_n7380, new_n7369, new_n7381);
nor_5  g05033(new_n7381, new_n7365, new_n7382);
nor_5  g05034(new_n7382, new_n7364, new_n7383);
nor_5  g05035(new_n7383, new_n7362, new_n7384);
nor_5  g05036(new_n7384, new_n7361, new_n7385);
nor_5  g05037(new_n7385, new_n7359, new_n7386);
nor_5  g05038(new_n7386, new_n7358, new_n7387);
nor_5  g05039(new_n7387, new_n7356, new_n7388);
nor_5  g05040(new_n7388, new_n7355, new_n7389);
nor_5  g05041(new_n7389, new_n7353, new_n7390_1);
nor_5  g05042(new_n7390_1, new_n7352, new_n7391);
nor_5  g05043(new_n7391, new_n7350, new_n7392);
nor_5  g05044(new_n7392, new_n7349_1, new_n7393);
nor_5  g05045(new_n7393, new_n7347, new_n7394);
or_5   g05046(new_n7394, new_n7346_1, new_n7395);
nor_5  g05047(new_n7395, new_n7344, new_n7396);
xnor_4 g05048(new_n7297, new_n7294, new_n7397);
xor_4  g05049(new_n7395, new_n7344, new_n7398);
nor_5  g05050(new_n7398, new_n7397, new_n7399);
xnor_4 g05051(new_n7398, new_n7397, new_n7400);
xor_4  g05052(new_n7292, new_n7241, new_n7401);
xor_4  g05053(new_n7393, new_n7347, new_n7402);
and_5  g05054(new_n7402, new_n7401, new_n7403_1);
xnor_4 g05055(new_n7402, new_n7401, new_n7404);
xor_4  g05056(new_n7290, new_n7245, new_n7405);
xor_4  g05057(new_n7391, new_n7350, new_n7406);
and_5  g05058(new_n7406, new_n7405, new_n7407);
xnor_4 g05059(new_n7406, new_n7405, new_n7408_1);
xor_4  g05060(new_n7288, new_n7249, new_n7409);
xor_4  g05061(new_n7389, new_n7353, new_n7410);
and_5  g05062(new_n7410, new_n7409, new_n7411);
xnor_4 g05063(new_n7410, new_n7409, new_n7412);
xor_4  g05064(new_n7286, new_n7253_1, new_n7413);
xor_4  g05065(new_n7387, new_n7356, new_n7414);
and_5  g05066(new_n7414, new_n7413, new_n7415);
xnor_4 g05067(new_n7414, new_n7413, new_n7416);
xor_4  g05068(new_n7284, new_n7257, new_n7417);
xor_4  g05069(new_n7385, new_n7359, new_n7418);
and_5  g05070(new_n7418, new_n7417, new_n7419);
xnor_4 g05071(new_n7418, new_n7417, new_n7420);
xor_4  g05072(new_n7282, new_n7261, new_n7421_1);
xor_4  g05073(new_n7383, new_n7362, new_n7422);
and_5  g05074(new_n7422, new_n7421_1, new_n7423);
xnor_4 g05075(new_n7422, new_n7421_1, new_n7424);
xnor_4 g05076(new_n7279, new_n7265, new_n7425);
xor_4  g05077(new_n7381, new_n7365, new_n7426);
and_5  g05078(new_n7426, new_n7425, new_n7427);
xnor_4 g05079(new_n7426, new_n7425, new_n7428_1);
xor_4  g05080(new_n7277_1, new_n7269, new_n7429);
xnor_4 g05081(new_n7367, n24485, new_n7430);
xnor_4 g05082(new_n7430, new_n7379, new_n7431);
nor_5  g05083(new_n7431, new_n7429, new_n7432_1);
xor_4  g05084(new_n7431, new_n7429, new_n7433);
xor_4  g05085(new_n7377_1, new_n7376, new_n7434);
xnor_4 g05086(new_n7275, new_n7273, new_n7435);
nor_5  g05087(new_n7435, new_n7434, new_n7436);
not_10 g05088(new_n2524, new_n7437_1);
nand_5 g05089(new_n2526, new_n7437_1, new_n7438);
xnor_4 g05090(new_n7435, new_n7434, new_n7439);
nor_5  g05091(new_n7439, new_n7438, new_n7440);
nor_5  g05092(new_n7440, new_n7436, new_n7441);
and_5  g05093(new_n7441, new_n7433, new_n7442);
nor_5  g05094(new_n7442, new_n7432_1, new_n7443);
nor_5  g05095(new_n7443, new_n7428_1, new_n7444);
nor_5  g05096(new_n7444, new_n7427, new_n7445);
nor_5  g05097(new_n7445, new_n7424, new_n7446);
nor_5  g05098(new_n7446, new_n7423, new_n7447);
nor_5  g05099(new_n7447, new_n7420, new_n7448);
nor_5  g05100(new_n7448, new_n7419, new_n7449);
nor_5  g05101(new_n7449, new_n7416, new_n7450);
nor_5  g05102(new_n7450, new_n7415, new_n7451);
nor_5  g05103(new_n7451, new_n7412, new_n7452);
nor_5  g05104(new_n7452, new_n7411, new_n7453);
nor_5  g05105(new_n7453, new_n7408_1, new_n7454);
nor_5  g05106(new_n7454, new_n7407, new_n7455);
nor_5  g05107(new_n7455, new_n7404, new_n7456);
nor_5  g05108(new_n7456, new_n7403_1, new_n7457);
nor_5  g05109(new_n7457, new_n7400, new_n7458);
nor_5  g05110(new_n7458, new_n7399, new_n7459);
xor_4  g05111(new_n7459, new_n7396, new_n7460_1);
xnor_4 g05112(new_n7460_1, new_n7299, n849);
xnor_4 g05113(new_n2511, new_n2510, n858);
or_5   g05114(n16994, n9246, new_n7463);
or_5   g05115(new_n7463, n10096, new_n7464);
or_5   g05116(new_n7464, n14790, new_n7465);
or_5   g05117(new_n7465, n17251, new_n7466);
or_5   g05118(new_n7466, n21674, new_n7467);
or_5   g05119(new_n7467, n24638, new_n7468);
or_5   g05120(new_n7468, n18444, new_n7469);
or_5   g05121(new_n7469, n14899, new_n7470);
xor_4  g05122(new_n7470, n3506, new_n7471);
xnor_4 g05123(new_n7471, n1314, new_n7472);
xor_4  g05124(new_n7469, n14899, new_n7473);
and_5  g05125(new_n7473, n3306, new_n7474);
or_5   g05126(new_n7473, n3306, new_n7475_1);
xor_4  g05127(new_n7468, n18444, new_n7476);
nor_5  g05128(new_n7476, n22335, new_n7477_1);
xnor_4 g05129(new_n7476, n22335, new_n7478);
xor_4  g05130(new_n7467, n24638, new_n7479);
nor_5  g05131(new_n7479, n24048, new_n7480);
xnor_4 g05132(new_n7479, n24048, new_n7481);
xor_4  g05133(new_n7466, n21674, new_n7482);
nor_5  g05134(new_n7482, n1525, new_n7483);
xnor_4 g05135(new_n7482, n1525, new_n7484);
xor_4  g05136(new_n7465, n17251, new_n7485);
nor_5  g05137(new_n7485, n16988, new_n7486);
xnor_4 g05138(new_n7485, n16988, new_n7487);
xor_4  g05139(new_n7464, n14790, new_n7488);
nor_5  g05140(new_n7488, n21779, new_n7489);
xor_4  g05141(new_n7463, n10096, new_n7490);
nor_5  g05142(new_n7490, n5376, new_n7491);
xnor_4 g05143(new_n7490, n5376, new_n7492);
xor_4  g05144(n16994, n9246, new_n7493);
nor_5  g05145(new_n7493, n5128, new_n7494);
and_5  g05146(n23120, n9246, new_n7495);
xnor_4 g05147(new_n7493, n5128, new_n7496);
nor_5  g05148(new_n7496, new_n7495, new_n7497);
nor_5  g05149(new_n7497, new_n7494, new_n7498);
nor_5  g05150(new_n7498, new_n7492, new_n7499);
nor_5  g05151(new_n7499, new_n7491, new_n7500);
xnor_4 g05152(new_n7488, n21779, new_n7501);
nor_5  g05153(new_n7501, new_n7500, new_n7502);
nor_5  g05154(new_n7502, new_n7489, new_n7503);
nor_5  g05155(new_n7503, new_n7487, new_n7504);
nor_5  g05156(new_n7504, new_n7486, new_n7505);
nor_5  g05157(new_n7505, new_n7484, new_n7506);
nor_5  g05158(new_n7506, new_n7483, new_n7507_1);
nor_5  g05159(new_n7507_1, new_n7481, new_n7508);
nor_5  g05160(new_n7508, new_n7480, new_n7509);
nor_5  g05161(new_n7509, new_n7478, new_n7510);
nor_5  g05162(new_n7510, new_n7477_1, new_n7511);
and_5  g05163(new_n7511, new_n7475_1, new_n7512);
nor_5  g05164(new_n7512, new_n7474, new_n7513);
xnor_4 g05165(new_n7513, new_n7472, new_n7514_1);
nor_5  g05166(new_n7514_1, n22442, new_n7515);
xnor_4 g05167(new_n7514_1, n22442, new_n7516);
xor_4  g05168(new_n7473, n3306, new_n7517);
xnor_4 g05169(new_n7517, new_n7511, new_n7518);
and_5  g05170(new_n7518, n468, new_n7519);
xor_4  g05171(new_n7518, n468, new_n7520);
xor_4  g05172(new_n7509, new_n7478, new_n7521);
nor_5  g05173(new_n7521, n5400, new_n7522);
xnor_4 g05174(new_n7521, n5400, new_n7523);
xor_4  g05175(new_n7507_1, new_n7481, new_n7524_1);
nor_5  g05176(new_n7524_1, n23923, new_n7525);
xnor_4 g05177(new_n7524_1, n23923, new_n7526);
xor_4  g05178(new_n7505, new_n7484, new_n7527);
and_5  g05179(new_n7527, n329, new_n7528);
or_5   g05180(new_n7527, n329, new_n7529);
xor_4  g05181(new_n7501, new_n7500, new_n7530);
nor_5  g05182(new_n7530, n2409, new_n7531);
xnor_4 g05183(new_n7530, n2409, new_n7532);
xor_4  g05184(new_n7498, new_n7492, new_n7533);
nor_5  g05185(new_n7533, n8869, new_n7534);
xor_4  g05186(new_n7496, new_n7495, new_n7535);
nor_5  g05187(new_n7535, n10372, new_n7536);
xnor_4 g05188(n23120, n9246, new_n7537);
and_5  g05189(new_n7537, n7428, new_n7538);
xnor_4 g05190(new_n7535, n10372, new_n7539);
nor_5  g05191(new_n7539, new_n7538, new_n7540);
nor_5  g05192(new_n7540, new_n7536, new_n7541);
xnor_4 g05193(new_n7533, n8869, new_n7542);
nor_5  g05194(new_n7542, new_n7541, new_n7543);
nor_5  g05195(new_n7543, new_n7534, new_n7544);
nor_5  g05196(new_n7544, new_n7532, new_n7545);
nor_5  g05197(new_n7545, new_n7531, new_n7546);
nor_5  g05198(new_n7546, n24170, new_n7547);
xor_4  g05199(new_n7503, new_n7487, new_n7548);
xnor_4 g05200(new_n7546, n24170, new_n7549);
nor_5  g05201(new_n7549, new_n7548, new_n7550);
nor_5  g05202(new_n7550, new_n7547, new_n7551);
and_5  g05203(new_n7551, new_n7529, new_n7552);
or_5   g05204(new_n7552, new_n7528, new_n7553);
nor_5  g05205(new_n7553, new_n7526, new_n7554);
nor_5  g05206(new_n7554, new_n7525, new_n7555);
nor_5  g05207(new_n7555, new_n7523, new_n7556);
nor_5  g05208(new_n7556, new_n7522, new_n7557);
and_5  g05209(new_n7557, new_n7520, new_n7558_1);
or_5   g05210(new_n7558_1, new_n7519, new_n7559);
nor_5  g05211(new_n7559, new_n7516, new_n7560);
nor_5  g05212(new_n7560, new_n7515, new_n7561);
nor_5  g05213(new_n7471, n1314, new_n7562);
nor_5  g05214(new_n7513, new_n7562, new_n7563);
nor_5  g05215(new_n7470, n3506, new_n7564);
and_5  g05216(new_n7471, n1314, new_n7565);
or_5   g05217(new_n7565, new_n7564, new_n7566_1);
nor_5  g05218(new_n7566_1, new_n7563, new_n7567);
xor_4  g05219(new_n7567, new_n7561, new_n7568);
not_10 g05220(new_n3304, new_n7569_1);
nor_5  g05221(new_n7569_1, n26180, new_n7570);
nor_5  g05222(new_n3350, new_n3305, new_n7571);
nor_5  g05223(new_n7571, new_n7570, new_n7572_1);
and_5  g05224(new_n3259, new_n6924, new_n7573);
nor_5  g05225(new_n3260_1, n25494, new_n7574);
and_5  g05226(new_n3260_1, n25494, new_n7575_1);
nor_5  g05227(new_n3303, new_n7575_1, new_n7576);
nor_5  g05228(new_n7576, new_n7574, new_n7577);
or_5   g05229(new_n7577, new_n7573, new_n7578);
xnor_4 g05230(new_n7578, new_n7572_1, new_n7579);
xor_4  g05231(new_n7579, new_n7568, new_n7580);
xor_4  g05232(new_n7559, new_n7516, new_n7581);
nor_5  g05233(new_n7581, new_n3351, new_n7582);
xnor_4 g05234(new_n7581, new_n3351, new_n7583);
xor_4  g05235(new_n3348, new_n3308, new_n7584);
xor_4  g05236(new_n7557, new_n7520, new_n7585_1);
and_5  g05237(new_n7585_1, new_n7584, new_n7586);
xnor_4 g05238(new_n7585_1, new_n7584, new_n7587);
not_10 g05239(new_n3468_1, new_n7588_1);
xor_4  g05240(new_n7555, new_n7523, new_n7589);
nor_5  g05241(new_n7589, new_n7588_1, new_n7590);
xor_4  g05242(new_n7589, new_n3468_1, new_n7591);
not_10 g05243(new_n3472, new_n7592);
xor_4  g05244(new_n7553, new_n7526, new_n7593_1);
nor_5  g05245(new_n7593_1, new_n7592, new_n7594);
not_10 g05246(new_n3476, new_n7595);
xor_4  g05247(new_n7527, n329, new_n7596);
xnor_4 g05248(new_n7596, new_n7551, new_n7597);
nor_5  g05249(new_n7597, new_n7595, new_n7598_1);
xor_4  g05250(new_n7597, new_n3476, new_n7599);
not_10 g05251(new_n3480_1, new_n7600);
xor_4  g05252(new_n7549, new_n7548, new_n7601);
nor_5  g05253(new_n7601, new_n7600, new_n7602);
not_10 g05254(new_n3485, new_n7603);
xor_4  g05255(new_n7544, new_n7532, new_n7604);
nor_5  g05256(new_n7604, new_n7603, new_n7605);
xor_4  g05257(new_n7604, new_n3485, new_n7606);
xor_4  g05258(new_n7542, new_n7541, new_n7607_1);
nor_5  g05259(new_n7607_1, new_n3489, new_n7608);
xor_4  g05260(new_n7539, new_n7538, new_n7609);
nor_5  g05261(new_n7609, new_n3495, new_n7610_1);
xor_4  g05262(new_n7537, n7428, new_n7611);
or_5   g05263(new_n7611, new_n3497, new_n7612);
xor_4  g05264(new_n7609, new_n3495, new_n7613);
and_5  g05265(new_n7613, new_n7612, new_n7614);
nor_5  g05266(new_n7614, new_n7610_1, new_n7615);
xnor_4 g05267(new_n7607_1, new_n3489, new_n7616_1);
nor_5  g05268(new_n7616_1, new_n7615, new_n7617);
nor_5  g05269(new_n7617, new_n7608, new_n7618);
nor_5  g05270(new_n7618, new_n7606, new_n7619);
or_5   g05271(new_n7619, new_n7605, new_n7620);
xnor_4 g05272(new_n7601, new_n3480_1, new_n7621);
and_5  g05273(new_n7621, new_n7620, new_n7622);
nor_5  g05274(new_n7622, new_n7602, new_n7623);
nor_5  g05275(new_n7623, new_n7599, new_n7624);
or_5   g05276(new_n7624, new_n7598_1, new_n7625);
xnor_4 g05277(new_n7593_1, new_n3472, new_n7626);
and_5  g05278(new_n7626, new_n7625, new_n7627);
nor_5  g05279(new_n7627, new_n7594, new_n7628);
nor_5  g05280(new_n7628, new_n7591, new_n7629);
nor_5  g05281(new_n7629, new_n7590, new_n7630_1);
nor_5  g05282(new_n7630_1, new_n7587, new_n7631);
nor_5  g05283(new_n7631, new_n7586, new_n7632);
nor_5  g05284(new_n7632, new_n7583, new_n7633);
or_5   g05285(new_n7633, new_n7582, new_n7634);
xnor_4 g05286(new_n7634, new_n7580, n873);
xnor_4 g05287(new_n4763, new_n4740, new_n7636);
xor_4  g05288(n4812, n2731, new_n7637);
nor_5  g05289(new_n3059, n19911, new_n7638);
xor_4  g05290(n24278, n19911, new_n7639);
nor_5  g05291(n24618, new_n3596, new_n7640);
not_10 g05292(n24618, new_n7641);
nor_5  g05293(new_n7641, n13708, new_n7642);
nor_5  g05294(new_n3600, n3952, new_n7643_1);
or_5   g05295(n18409, new_n3111, new_n7644);
nor_5  g05296(n12315, new_n6328, new_n7645);
and_5  g05297(new_n7645, new_n7644, new_n7646);
nor_5  g05298(new_n7646, new_n7643_1, new_n7647_1);
nor_5  g05299(new_n7647_1, new_n7642, new_n7648);
or_5   g05300(new_n7648, new_n7640, new_n7649);
nor_5  g05301(new_n7649, new_n7639, new_n7650);
nor_5  g05302(new_n7650, new_n7638, new_n7651);
xor_4  g05303(new_n7651, new_n7637, new_n7652);
xnor_4 g05304(new_n7652, new_n7636, new_n7653);
xor_4  g05305(new_n7649, new_n7639, new_n7654);
nor_5  g05306(new_n7654, new_n4793, new_n7655);
xnor_4 g05307(n24618, n13708, new_n7656);
xnor_4 g05308(new_n7656, new_n7647_1, new_n7657_1);
nor_5  g05309(new_n7657_1, new_n4797, new_n7658);
xnor_4 g05310(new_n7657_1, new_n4797, new_n7659);
xnor_4 g05311(n12315, n5704, new_n7660);
or_5   g05312(new_n7660, new_n4803, new_n7661);
nor_5  g05313(new_n7661, new_n4808, new_n7662);
xnor_4 g05314(new_n7661, new_n4808, new_n7663);
xor_4  g05315(n18409, n3952, new_n7664);
xnor_4 g05316(new_n7664, new_n7645, new_n7665);
nor_5  g05317(new_n7665, new_n7663, new_n7666);
nor_5  g05318(new_n7666, new_n7662, new_n7667);
nor_5  g05319(new_n7667, new_n7659, new_n7668);
nor_5  g05320(new_n7668, new_n7658, new_n7669);
xor_4  g05321(new_n7654, new_n4793, new_n7670_1);
and_5  g05322(new_n7670_1, new_n7669, new_n7671);
or_5   g05323(new_n7671, new_n7655, new_n7672);
xor_4  g05324(new_n7672, new_n7653, n879);
xnor_4 g05325(new_n7263, n18157, new_n7674_1);
nor_5  g05326(new_n7267, n12161, new_n7675);
nor_5  g05327(new_n7273, new_n6550, new_n7676);
or_5   g05328(new_n2523, new_n6553, new_n7677);
xor_4  g05329(new_n7273, n5026, new_n7678_1);
nor_5  g05330(new_n7678_1, new_n7677, new_n7679_1);
nor_5  g05331(new_n7679_1, new_n7676, new_n7680);
xor_4  g05332(new_n7267, n12161, new_n7681);
and_5  g05333(new_n7681, new_n7680, new_n7682);
nor_5  g05334(new_n7682, new_n7675, new_n7683);
xnor_4 g05335(new_n7683, new_n7674_1, new_n7684);
xnor_4 g05336(new_n7681, new_n7680, new_n7685);
xnor_4 g05337(new_n5998, n14684, new_n7686_1);
not_10 g05338(n6631, new_n7687);
and_5  g05339(new_n6001, new_n7687, new_n7688);
and_5  g05340(new_n6004, n24732, new_n7689);
xor_4  g05341(new_n6001, n6631, new_n7690);
nor_5  g05342(new_n7690, new_n7689, new_n7691);
nor_5  g05343(new_n7691, new_n7688, new_n7692_1);
xor_4  g05344(new_n7692_1, new_n7686_1, new_n7693_1);
nor_5  g05345(new_n7693_1, new_n7685, new_n7694);
xnor_4 g05346(new_n7693_1, new_n7685, new_n7695);
xor_4  g05347(new_n7690, new_n7689, new_n7696);
xor_4  g05348(new_n7678_1, new_n7677, new_n7697);
nor_5  g05349(new_n7697, new_n7696, new_n7698_1);
xnor_4 g05350(new_n6004, n24732, new_n7699);
xnor_4 g05351(new_n2523, n8581, new_n7700);
nor_5  g05352(new_n7700, new_n7699, new_n7701);
xor_4  g05353(new_n7697, new_n7696, new_n7702);
and_5  g05354(new_n7702, new_n7701, new_n7703);
nor_5  g05355(new_n7703, new_n7698_1, new_n7704);
nor_5  g05356(new_n7704, new_n7695, new_n7705);
nor_5  g05357(new_n7705, new_n7694, new_n7706);
xor_4  g05358(new_n7706, new_n7684, new_n7707);
xor_4  g05359(new_n5996, n17035, new_n7708_1);
nor_5  g05360(new_n5998, n14684, new_n7709);
nor_5  g05361(new_n7692_1, new_n7686_1, new_n7710);
nor_5  g05362(new_n7710, new_n7709, new_n7711);
xor_4  g05363(new_n7711, new_n7708_1, new_n7712);
xnor_4 g05364(new_n7712, new_n7707, n887);
xnor_4 g05365(new_n5534, n24327, new_n7714);
and_5  g05366(new_n5537, n22198, new_n7715);
xnor_4 g05367(new_n5537, n22198, new_n7716);
and_5  g05368(new_n5540, n20826, new_n7717);
xnor_4 g05369(new_n5540, n20826, new_n7718);
and_5  g05370(new_n5543, n7305, new_n7719);
xnor_4 g05371(new_n5543, n7305, new_n7720);
and_5  g05372(new_n5546, n25872, new_n7721_1);
nor_5  g05373(new_n5549, n20259, new_n7722);
nand_5 g05374(new_n5329, n3925, new_n7723);
xnor_4 g05375(new_n5548, n20259, new_n7724);
and_5  g05376(new_n7724, new_n7723, new_n7725);
nor_5  g05377(new_n7725, new_n7722, new_n7726);
xor_4  g05378(new_n5546, n25872, new_n7727);
and_5  g05379(new_n7727, new_n7726, new_n7728);
nor_5  g05380(new_n7728, new_n7721_1, new_n7729);
nor_5  g05381(new_n7729, new_n7720, new_n7730);
nor_5  g05382(new_n7730, new_n7719, new_n7731_1);
nor_5  g05383(new_n7731_1, new_n7718, new_n7732);
nor_5  g05384(new_n7732, new_n7717, new_n7733);
nor_5  g05385(new_n7733, new_n7716, new_n7734);
nor_5  g05386(new_n7734, new_n7715, new_n7735);
xor_4  g05387(new_n7735, new_n7714, new_n7736);
xor_4  g05388(new_n2875, n25119, new_n7737);
and_5  g05389(new_n2879, n1163, new_n7738);
nor_5  g05390(new_n2883, n18537, new_n7739);
xnor_4 g05391(new_n2883, n18537, new_n7740);
nor_5  g05392(new_n2887_1, n7057, new_n7741);
xor_4  g05393(new_n2887_1, n7057, new_n7742);
and_5  g05394(new_n2891, n8381, new_n7743);
xor_4  g05395(new_n2891, n8381, new_n7744);
and_5  g05396(new_n2898, n12495, new_n7745);
nor_5  g05397(new_n7745, n20235, new_n7746);
xnor_4 g05398(new_n7745, n20235, new_n7747);
nor_5  g05399(new_n7747, new_n2895, new_n7748);
nor_5  g05400(new_n7748, new_n7746, new_n7749);
and_5  g05401(new_n7749, new_n7744, new_n7750);
nor_5  g05402(new_n7750, new_n7743, new_n7751_1);
and_5  g05403(new_n7751_1, new_n7742, new_n7752);
nor_5  g05404(new_n7752, new_n7741, new_n7753);
nor_5  g05405(new_n7753, new_n7740, new_n7754);
or_5   g05406(new_n7754, new_n7739, new_n7755);
xnor_4 g05407(new_n2879, n1163, new_n7756);
nor_5  g05408(new_n7756, new_n7755, new_n7757);
nor_5  g05409(new_n7757, new_n7738, new_n7758);
xor_4  g05410(new_n7758, new_n7737, new_n7759_1);
xnor_4 g05411(new_n7759_1, new_n7736, new_n7760);
xnor_4 g05412(new_n7733, new_n7716, new_n7761);
xor_4  g05413(new_n7756, new_n7755, new_n7762);
nor_5  g05414(new_n7762, new_n7761, new_n7763);
xnor_4 g05415(new_n7762, new_n7761, new_n7764);
xor_4  g05416(new_n7753, new_n7740, new_n7765);
xor_4  g05417(new_n7731_1, new_n7718, new_n7766);
and_5  g05418(new_n7766, new_n7765, new_n7767);
xnor_4 g05419(new_n7766, new_n7765, new_n7768);
xor_4  g05420(new_n7751_1, new_n7742, new_n7769_1);
xor_4  g05421(new_n7729, new_n7720, new_n7770);
and_5  g05422(new_n7770, new_n7769_1, new_n7771);
xnor_4 g05423(new_n7770, new_n7769_1, new_n7772);
xnor_4 g05424(new_n7749, new_n7744, new_n7773_1);
xor_4  g05425(new_n7727, new_n7726, new_n7774);
and_5  g05426(new_n7774, new_n7773_1, new_n7775);
xnor_4 g05427(new_n7774, new_n7773_1, new_n7776);
xor_4  g05428(new_n7724, new_n7723, new_n7777);
not_10 g05429(new_n7777, new_n7778);
xor_4  g05430(new_n7747, new_n2895, new_n7779);
and_5  g05431(new_n7779, new_n7778, new_n7780_1);
xor_4  g05432(new_n5329, n3925, new_n7781);
not_10 g05433(new_n7781, new_n7782);
xor_4  g05434(new_n2898, n12495, new_n7783);
nor_5  g05435(new_n7783, new_n7782, new_n7784);
xnor_4 g05436(new_n7779, new_n7777, new_n7785);
and_5  g05437(new_n7785, new_n7784, new_n7786);
nor_5  g05438(new_n7786, new_n7780_1, new_n7787);
nor_5  g05439(new_n7787, new_n7776, new_n7788_1);
nor_5  g05440(new_n7788_1, new_n7775, new_n7789);
nor_5  g05441(new_n7789, new_n7772, new_n7790);
nor_5  g05442(new_n7790, new_n7771, new_n7791);
nor_5  g05443(new_n7791, new_n7768, new_n7792);
nor_5  g05444(new_n7792, new_n7767, new_n7793);
nor_5  g05445(new_n7793, new_n7764, new_n7794_1);
nor_5  g05446(new_n7794_1, new_n7763, new_n7795);
xnor_4 g05447(new_n7795, new_n7760, n904);
nor_5  g05448(n18962, n10158, new_n7797);
nand_5 g05449(new_n7797, new_n6766, new_n7798);
or_5   g05450(new_n7798, n15539, new_n7799);
xnor_4 g05451(new_n7799, new_n6759, new_n7800);
xor_4  g05452(new_n7800, n21471, new_n7801);
xnor_4 g05453(new_n7798, new_n6762, new_n7802);
and_5  g05454(new_n7802, n18737, new_n7803);
xnor_4 g05455(new_n7802, n18737, new_n7804);
xnor_4 g05456(new_n7797, n8052, new_n7805);
and_5  g05457(new_n7805, n14603, new_n7806);
xnor_4 g05458(new_n7805, n14603, new_n7807);
xor_4  g05459(n18962, n10158, new_n7808);
nor_5  g05460(new_n7808, n20794, new_n7809);
nand_5 g05461(n23333, n18962, new_n7810);
xor_4  g05462(new_n7808, n20794, new_n7811_1);
and_5  g05463(new_n7811_1, new_n7810, new_n7812);
or_5   g05464(new_n7812, new_n7809, new_n7813);
nor_5  g05465(new_n7813, new_n7807, new_n7814);
nor_5  g05466(new_n7814, new_n7806, new_n7815);
nor_5  g05467(new_n7815, new_n7804, new_n7816);
nor_5  g05468(new_n7816, new_n7803, new_n7817);
xnor_4 g05469(new_n7817, new_n7801, new_n7818);
xnor_4 g05470(new_n7818, n19472, new_n7819);
xor_4  g05471(new_n7815, new_n7804, new_n7820);
nor_5  g05472(new_n7820, n25370, new_n7821);
xor_4  g05473(new_n7813, new_n7807, new_n7822);
and_5  g05474(new_n7822, n24786, new_n7823);
xnor_4 g05475(new_n7822, n24786, new_n7824);
xor_4  g05476(n23333, n18962, new_n7825);
and_5  g05477(new_n7825, n23065, new_n7826);
and_5  g05478(new_n7826, new_n7811_1, new_n7827);
xnor_4 g05479(new_n7811_1, new_n7810, new_n7828);
nor_5  g05480(new_n7828, new_n7826, new_n7829);
nor_5  g05481(new_n7829, new_n7827, new_n7830_1);
and_5  g05482(new_n7830_1, n27120, new_n7831);
nor_5  g05483(new_n7831, new_n7827, new_n7832);
nor_5  g05484(new_n7832, new_n7824, new_n7833);
nor_5  g05485(new_n7833, new_n7823, new_n7834_1);
not_10 g05486(new_n7834_1, new_n7835);
xnor_4 g05487(new_n7820, n25370, new_n7836);
nor_5  g05488(new_n7836, new_n7835, new_n7837);
or_5   g05489(new_n7837, new_n7821, new_n7838);
xor_4  g05490(new_n7838, new_n7819, new_n7839);
xnor_4 g05491(new_n7839, new_n6075, new_n7840);
xnor_4 g05492(new_n7836, new_n7834_1, new_n7841_1);
and_5  g05493(new_n7841_1, new_n6079, new_n7842);
xnor_4 g05494(new_n7841_1, new_n6079, new_n7843);
xnor_4 g05495(new_n7830_1, n27120, new_n7844);
and_5  g05496(new_n7844, new_n6086, new_n7845);
xnor_4 g05497(new_n7825, n23065, new_n7846);
or_5   g05498(new_n7846, new_n6082, new_n7847);
xor_4  g05499(new_n7844, new_n6086, new_n7848);
and_5  g05500(new_n7848, new_n7847, new_n7849);
nor_5  g05501(new_n7849, new_n7845, new_n7850);
nor_5  g05502(new_n7850, new_n6096, new_n7851);
xnor_4 g05503(new_n7832, new_n7824, new_n7852);
xor_4  g05504(new_n7850, new_n6096, new_n7853);
and_5  g05505(new_n7853, new_n7852, new_n7854);
nor_5  g05506(new_n7854, new_n7851, new_n7855);
nor_5  g05507(new_n7855, new_n7843, new_n7856);
nor_5  g05508(new_n7856, new_n7842, new_n7857);
xnor_4 g05509(new_n7857, new_n7840, n948);
xor_4  g05510(n25972, n10250, new_n7859);
not_10 g05511(n21915, new_n7860);
nor_5  g05512(new_n7860, n7674, new_n7861);
xor_4  g05513(n21915, n7674, new_n7862);
not_10 g05514(n13775, new_n7863);
nor_5  g05515(new_n7863, n6397, new_n7864);
xor_4  g05516(n13775, n6397, new_n7865);
not_10 g05517(n1293, new_n7866);
nor_5  g05518(n19196, new_n7866, new_n7867);
xor_4  g05519(n19196, n1293, new_n7868);
not_10 g05520(n19042, new_n7869);
nor_5  g05521(n23586, new_n7869, new_n7870);
xor_4  g05522(n23586, n19042, new_n7871);
not_10 g05523(n19472, new_n7872);
nor_5  g05524(n21226, new_n7872, new_n7873);
xor_4  g05525(n21226, n19472, new_n7874);
not_10 g05526(n25370, new_n7875);
nor_5  g05527(new_n7875, n4426, new_n7876_1);
xor_4  g05528(n25370, n4426, new_n7877);
not_10 g05529(n20036, new_n7878);
nor_5  g05530(n24786, new_n7878, new_n7879);
and_5  g05531(n24786, new_n7878, new_n7880);
nor_5  g05532(n27120, new_n3851, new_n7881);
nand_5 g05533(n27120, new_n3851, new_n7882);
nor_5  g05534(n23065, new_n3854, new_n7883);
and_5  g05535(new_n7883, new_n7882, new_n7884_1);
nor_5  g05536(new_n7884_1, new_n7881, new_n7885);
nor_5  g05537(new_n7885, new_n7880, new_n7886);
or_5   g05538(new_n7886, new_n7879, new_n7887);
nor_5  g05539(new_n7887, new_n7877, new_n7888);
nor_5  g05540(new_n7888, new_n7876_1, new_n7889);
nor_5  g05541(new_n7889, new_n7874, new_n7890);
nor_5  g05542(new_n7890, new_n7873, new_n7891);
nor_5  g05543(new_n7891, new_n7871, new_n7892);
nor_5  g05544(new_n7892, new_n7870, new_n7893);
nor_5  g05545(new_n7893, new_n7868, new_n7894);
nor_5  g05546(new_n7894, new_n7867, new_n7895);
nor_5  g05547(new_n7895, new_n7865, new_n7896);
nor_5  g05548(new_n7896, new_n7864, new_n7897);
nor_5  g05549(new_n7897, new_n7862, new_n7898);
nor_5  g05550(new_n7898, new_n7861, new_n7899);
xor_4  g05551(new_n7899, new_n7859, new_n7900);
xor_4  g05552(n20040, n2978, new_n7901);
nor_5  g05553(new_n6747, n19531, new_n7902);
xor_4  g05554(n23697, n19531, new_n7903);
nor_5  g05555(n18345, new_n6750, new_n7904);
xor_4  g05556(n18345, n2289, new_n7905);
nor_5  g05557(n13190, new_n6753, new_n7906);
xor_4  g05558(n13190, n1112, new_n7907);
nor_5  g05559(new_n6756, n3460, new_n7908);
xor_4  g05560(n20179, n3460, new_n7909);
or_5   g05561(new_n6759, n5226, new_n7910);
xor_4  g05562(n19228, n5226, new_n7911);
or_5   g05563(n17664, new_n6762, new_n7912);
xor_4  g05564(n17664, n15539, new_n7913);
and_5  g05565(n23369, new_n6766, new_n7914);
nor_5  g05566(n23369, new_n6766, new_n7915);
and_5  g05567(new_n6769, n1136, new_n7916);
or_5   g05568(new_n6769, n1136, new_n7917_1);
not_10 g05569(n18962, new_n7918);
and_5  g05570(n19234, new_n7918, new_n7919);
and_5  g05571(new_n7919, new_n7917_1, new_n7920);
nor_5  g05572(new_n7920, new_n7916, new_n7921);
nor_5  g05573(new_n7921, new_n7915, new_n7922);
nor_5  g05574(new_n7922, new_n7914, new_n7923);
not_10 g05575(new_n7923, new_n7924);
or_5   g05576(new_n7924, new_n7913, new_n7925);
and_5  g05577(new_n7925, new_n7912, new_n7926);
or_5   g05578(new_n7926, new_n7911, new_n7927);
and_5  g05579(new_n7927, new_n7910, new_n7928);
nor_5  g05580(new_n7928, new_n7909, new_n7929);
nor_5  g05581(new_n7929, new_n7908, new_n7930);
nor_5  g05582(new_n7930, new_n7907, new_n7931);
nor_5  g05583(new_n7931, new_n7906, new_n7932);
nor_5  g05584(new_n7932, new_n7905, new_n7933);
nor_5  g05585(new_n7933, new_n7904, new_n7934);
nor_5  g05586(new_n7934, new_n7903, new_n7935);
nor_5  g05587(new_n7935, new_n7902, new_n7936);
xor_4  g05588(new_n7936, new_n7901, new_n7937_1);
or_5   g05589(n15258, n4588, new_n7938);
or_5   g05590(new_n7938, n16743, new_n7939);
or_5   g05591(new_n7939, n22631, new_n7940);
or_5   g05592(new_n7940, n2331, new_n7941);
or_5   g05593(new_n7941, n25068, new_n7942);
or_5   g05594(new_n7942, n16812, new_n7943_1);
or_5   g05595(new_n7943_1, n7841, new_n7944);
nor_5  g05596(new_n7944, n26264, new_n7945);
xnor_4 g05597(new_n7945, n22764, new_n7946);
xor_4  g05598(new_n7946, n12507, new_n7947);
xor_4  g05599(new_n7944, n26264, new_n7948);
and_5  g05600(new_n7948, n15077, new_n7949_1);
nor_5  g05601(new_n7948, n15077, new_n7950_1);
xor_4  g05602(new_n7943_1, n7841, new_n7951);
and_5  g05603(new_n7951, n3710, new_n7952);
or_5   g05604(new_n7951, n3710, new_n7953);
xor_4  g05605(new_n7942, n16812, new_n7954);
nor_5  g05606(new_n7954, n26318, new_n7955);
xnor_4 g05607(new_n7954, n26318, new_n7956);
xor_4  g05608(new_n7941, n25068, new_n7957);
nor_5  g05609(new_n7957, n26054, new_n7958);
xnor_4 g05610(new_n7957, n26054, new_n7959_1);
xor_4  g05611(new_n7940, n2331, new_n7960);
nor_5  g05612(new_n7960, n19081, new_n7961);
xnor_4 g05613(new_n7960, n19081, new_n7962);
xor_4  g05614(new_n7939, n22631, new_n7963_1);
nor_5  g05615(new_n7963_1, n8309, new_n7964);
xor_4  g05616(new_n7938, n16743, new_n7965);
nor_5  g05617(new_n7965, n19144, new_n7966);
xnor_4 g05618(new_n7965, n19144, new_n7967);
not_10 g05619(n12593, new_n7968_1);
xnor_4 g05620(n15258, n4588, new_n7969);
and_5  g05621(new_n7969, new_n7968_1, new_n7970);
and_5  g05622(n13714, n4588, new_n7971);
xor_4  g05623(new_n7969, n12593, new_n7972);
nor_5  g05624(new_n7972, new_n7971, new_n7973);
nor_5  g05625(new_n7973, new_n7970, new_n7974);
nor_5  g05626(new_n7974, new_n7967, new_n7975);
nor_5  g05627(new_n7975, new_n7966, new_n7976);
xnor_4 g05628(new_n7963_1, n8309, new_n7977);
nor_5  g05629(new_n7977, new_n7976, new_n7978);
nor_5  g05630(new_n7978, new_n7964, new_n7979);
nor_5  g05631(new_n7979, new_n7962, new_n7980);
nor_5  g05632(new_n7980, new_n7961, new_n7981);
nor_5  g05633(new_n7981, new_n7959_1, new_n7982);
nor_5  g05634(new_n7982, new_n7958, new_n7983);
nor_5  g05635(new_n7983, new_n7956, new_n7984);
nor_5  g05636(new_n7984, new_n7955, new_n7985);
and_5  g05637(new_n7985, new_n7953, new_n7986);
nor_5  g05638(new_n7986, new_n7952, new_n7987);
nor_5  g05639(new_n7987, new_n7950_1, new_n7988);
nor_5  g05640(new_n7988, new_n7949_1, new_n7989);
xnor_4 g05641(new_n7989, new_n7947, new_n7990);
xnor_4 g05642(new_n7990, new_n7937_1, new_n7991);
xor_4  g05643(new_n7934, new_n7903, new_n7992_1);
xor_4  g05644(new_n7948, n15077, new_n7993);
xnor_4 g05645(new_n7993, new_n7987, new_n7994);
and_5  g05646(new_n7994, new_n7992_1, new_n7995);
xnor_4 g05647(new_n7994, new_n7992_1, new_n7996);
xor_4  g05648(new_n7932, new_n7905, new_n7997);
xnor_4 g05649(new_n7951, n3710, new_n7998);
xnor_4 g05650(new_n7998, new_n7985, new_n7999_1);
nor_5  g05651(new_n7999_1, new_n7997, new_n8000);
xnor_4 g05652(new_n7999_1, new_n7997, new_n8001);
xor_4  g05653(new_n7930, new_n7907, new_n8002);
xnor_4 g05654(new_n7983, new_n7956, new_n8003);
nor_5  g05655(new_n8003, new_n8002, new_n8004);
xnor_4 g05656(new_n8003, new_n8002, new_n8005);
xnor_4 g05657(new_n7928, new_n7909, new_n8006_1);
xor_4  g05658(new_n7981, new_n7959_1, new_n8007);
and_5  g05659(new_n8007, new_n8006_1, new_n8008);
xnor_4 g05660(new_n8007, new_n8006_1, new_n8009);
xnor_4 g05661(new_n7926, new_n7911, new_n8010);
xor_4  g05662(new_n7979, new_n7962, new_n8011);
and_5  g05663(new_n8011, new_n8010, new_n8012);
xor_4  g05664(new_n7926, new_n7911, new_n8013);
xor_4  g05665(new_n8011, new_n8013, new_n8014);
xnor_4 g05666(new_n7923, new_n7913, new_n8015);
xnor_4 g05667(new_n7977, new_n7976, new_n8016);
nor_5  g05668(new_n8016, new_n8015, new_n8017);
xor_4  g05669(new_n8016, new_n8015, new_n8018);
xor_4  g05670(new_n7974, new_n7967, new_n8019);
xnor_4 g05671(n23369, n8052, new_n8020);
xnor_4 g05672(new_n8020, new_n7921, new_n8021);
nor_5  g05673(new_n8021, new_n8019, new_n8022);
xnor_4 g05674(new_n8021, new_n8019, new_n8023);
xor_4  g05675(new_n7972, new_n7971, new_n8024);
xor_4  g05676(n10158, n1136, new_n8025);
xnor_4 g05677(new_n8025, new_n7919, new_n8026);
nor_5  g05678(new_n8026, new_n8024, new_n8027_1);
xnor_4 g05679(n19234, n18962, new_n8028);
xnor_4 g05680(n13714, n4588, new_n8029);
nor_5  g05681(new_n8029, new_n8028, new_n8030);
xor_4  g05682(new_n8026, new_n8024, new_n8031_1);
and_5  g05683(new_n8031_1, new_n8030, new_n8032);
nor_5  g05684(new_n8032, new_n8027_1, new_n8033);
nor_5  g05685(new_n8033, new_n8023, new_n8034);
nor_5  g05686(new_n8034, new_n8022, new_n8035);
and_5  g05687(new_n8035, new_n8018, new_n8036);
nor_5  g05688(new_n8036, new_n8017, new_n8037);
nor_5  g05689(new_n8037, new_n8014, new_n8038);
nor_5  g05690(new_n8038, new_n8012, new_n8039);
nor_5  g05691(new_n8039, new_n8009, new_n8040);
nor_5  g05692(new_n8040, new_n8008, new_n8041);
nor_5  g05693(new_n8041, new_n8005, new_n8042_1);
nor_5  g05694(new_n8042_1, new_n8004, new_n8043);
nor_5  g05695(new_n8043, new_n8001, new_n8044);
or_5   g05696(new_n8044, new_n8000, new_n8045);
nor_5  g05697(new_n8045, new_n7996, new_n8046);
nor_5  g05698(new_n8046, new_n7995, new_n8047);
xor_4  g05699(new_n8047, new_n7991, new_n8048);
xnor_4 g05700(new_n8048, new_n7900, new_n8049);
xor_4  g05701(new_n7897, new_n7862, new_n8050);
xor_4  g05702(new_n8045, new_n7996, new_n8051);
nor_5  g05703(new_n8051, new_n8050, new_n8052_1);
xnor_4 g05704(new_n8051, new_n8050, new_n8053);
xnor_4 g05705(new_n7895, new_n7865, new_n8054);
xor_4  g05706(new_n8043, new_n8001, new_n8055);
and_5  g05707(new_n8055, new_n8054, new_n8056);
xnor_4 g05708(new_n8055, new_n8054, new_n8057);
xnor_4 g05709(new_n7893, new_n7868, new_n8058);
xor_4  g05710(new_n8041, new_n8005, new_n8059);
and_5  g05711(new_n8059, new_n8058, new_n8060);
xnor_4 g05712(new_n8059, new_n8058, new_n8061);
xnor_4 g05713(new_n7891, new_n7871, new_n8062);
xor_4  g05714(new_n8039, new_n8009, new_n8063);
and_5  g05715(new_n8063, new_n8062, new_n8064);
xnor_4 g05716(new_n8063, new_n8062, new_n8065);
xnor_4 g05717(new_n7889, new_n7874, new_n8066);
xor_4  g05718(new_n8037, new_n8014, new_n8067_1);
and_5  g05719(new_n8067_1, new_n8066, new_n8068);
xnor_4 g05720(new_n8067_1, new_n8066, new_n8069);
xnor_4 g05721(new_n8035, new_n8018, new_n8070);
xor_4  g05722(new_n7887, new_n7877, new_n8071);
nor_5  g05723(new_n8071, new_n8070, new_n8072);
xnor_4 g05724(new_n8071, new_n8070, new_n8073);
xnor_4 g05725(new_n8033, new_n8023, new_n8074);
xnor_4 g05726(n24786, n20036, new_n8075);
xnor_4 g05727(new_n8075, new_n7885, new_n8076);
and_5  g05728(new_n8076, new_n8074, new_n8077);
xnor_4 g05729(new_n8076, new_n8074, new_n8078);
xnor_4 g05730(n23065, n9380, new_n8079);
xnor_4 g05731(new_n8029, new_n8028, new_n8080);
or_5   g05732(new_n8080, new_n8079, new_n8081);
xor_4  g05733(n27120, n11192, new_n8082);
xnor_4 g05734(new_n8082, new_n7883, new_n8083);
and_5  g05735(new_n8083, new_n8081, new_n8084);
xnor_4 g05736(new_n8031_1, new_n8030, new_n8085);
xor_4  g05737(new_n8083, new_n8081, new_n8086);
and_5  g05738(new_n8086, new_n8085, new_n8087);
nor_5  g05739(new_n8087, new_n8084, new_n8088);
nor_5  g05740(new_n8088, new_n8078, new_n8089);
nor_5  g05741(new_n8089, new_n8077, new_n8090);
nor_5  g05742(new_n8090, new_n8073, new_n8091);
nor_5  g05743(new_n8091, new_n8072, new_n8092);
nor_5  g05744(new_n8092, new_n8069, new_n8093);
nor_5  g05745(new_n8093, new_n8068, new_n8094);
nor_5  g05746(new_n8094, new_n8065, new_n8095_1);
nor_5  g05747(new_n8095_1, new_n8064, new_n8096);
nor_5  g05748(new_n8096, new_n8061, new_n8097);
nor_5  g05749(new_n8097, new_n8060, new_n8098);
nor_5  g05750(new_n8098, new_n8057, new_n8099);
nor_5  g05751(new_n8099, new_n8056, new_n8100);
nor_5  g05752(new_n8100, new_n8053, new_n8101);
or_5   g05753(new_n8101, new_n8052_1, new_n8102);
xor_4  g05754(new_n8102, new_n8049, n957);
xnor_4 g05755(new_n8028, n20385, new_n8104);
xnor_4 g05756(n26167, n24129, new_n8105);
xnor_4 g05757(new_n8105, n21138, new_n8106);
xor_4  g05758(new_n8106, new_n8104, n980);
and_5  g05759(new_n7020, new_n4053, new_n8108);
xnor_4 g05760(new_n7020, new_n4053, new_n8109_1);
nor_5  g05761(new_n7024, new_n4056, new_n8110);
xnor_4 g05762(new_n7024, new_n4056, new_n8111);
nor_5  g05763(new_n7028, new_n4059, new_n8112);
xnor_4 g05764(new_n7028, new_n4059, new_n8113);
nor_5  g05765(new_n7032_1, new_n4062, new_n8114);
xnor_4 g05766(new_n7032_1, new_n4062, new_n8115);
nor_5  g05767(new_n7036, new_n4065, new_n8116);
xnor_4 g05768(new_n7036, new_n4065, new_n8117);
nor_5  g05769(new_n7040, new_n4068, new_n8118);
xnor_4 g05770(new_n7040, new_n4068, new_n8119);
nor_5  g05771(new_n7044, new_n4071_1, new_n8120);
xnor_4 g05772(new_n7044, new_n4071_1, new_n8121);
and_5  g05773(new_n7049, new_n4077, new_n8122);
xor_4  g05774(new_n7049, new_n4077, new_n8123);
nor_5  g05775(new_n7055, new_n4082, new_n8124);
nor_5  g05776(new_n7059, new_n4085_1, new_n8125);
xor_4  g05777(new_n7055, new_n4082, new_n8126);
and_5  g05778(new_n8126, new_n8125, new_n8127_1);
nor_5  g05779(new_n8127_1, new_n8124, new_n8128);
and_5  g05780(new_n8128, new_n8123, new_n8129);
nor_5  g05781(new_n8129, new_n8122, new_n8130_1);
nor_5  g05782(new_n8130_1, new_n8121, new_n8131);
nor_5  g05783(new_n8131, new_n8120, new_n8132);
nor_5  g05784(new_n8132, new_n8119, new_n8133);
nor_5  g05785(new_n8133, new_n8118, new_n8134);
nor_5  g05786(new_n8134, new_n8117, new_n8135_1);
nor_5  g05787(new_n8135_1, new_n8116, new_n8136);
nor_5  g05788(new_n8136, new_n8115, new_n8137);
nor_5  g05789(new_n8137, new_n8114, new_n8138);
nor_5  g05790(new_n8138, new_n8113, new_n8139_1);
nor_5  g05791(new_n8139_1, new_n8112, new_n8140);
nor_5  g05792(new_n8140, new_n8111, new_n8141);
or_5   g05793(new_n8141, new_n8110, new_n8142);
nor_5  g05794(new_n8142, new_n8109_1, new_n8143);
nor_5  g05795(new_n8143, new_n8108, new_n8144);
xnor_4 g05796(new_n7018, new_n4052, new_n8145);
xor_4  g05797(new_n8145, new_n8144, new_n8146);
not_10 g05798(n16544, new_n8147);
nor_5  g05799(new_n8147, n12650, new_n8148_1);
xor_4  g05800(n16544, n12650, new_n8149_1);
not_10 g05801(n6814, new_n8150);
nor_5  g05802(n10201, new_n8150, new_n8151);
xor_4  g05803(n10201, n6814, new_n8152);
not_10 g05804(n19701, new_n8153);
nor_5  g05805(new_n8153, n10593, new_n8154);
xor_4  g05806(n19701, n10593, new_n8155);
not_10 g05807(n23529, new_n8156);
nor_5  g05808(new_n8156, n18290, new_n8157);
xor_4  g05809(n23529, n18290, new_n8158);
not_10 g05810(n24620, new_n8159_1);
nor_5  g05811(new_n8159_1, n11580, new_n8160);
xor_4  g05812(n24620, n11580, new_n8161);
not_10 g05813(n5211, new_n8162);
nor_5  g05814(n15884, new_n8162, new_n8163);
xor_4  g05815(n15884, n5211, new_n8164);
not_10 g05816(n12956, new_n8165);
nor_5  g05817(new_n8165, n6356, new_n8166);
xor_4  g05818(n12956, n6356, new_n8167);
not_10 g05819(n18295, new_n8168);
and_5  g05820(n27104, new_n8168, new_n8169);
nor_5  g05821(n27104, new_n8168, new_n8170);
nor_5  g05822(new_n5146, n6502, new_n8171);
not_10 g05823(n6502, new_n8172);
or_5   g05824(n27188, new_n8172, new_n8173);
not_10 g05825(n6611, new_n8174);
nor_5  g05826(n15780, new_n8174, new_n8175);
and_5  g05827(new_n8175, new_n8173, new_n8176);
nor_5  g05828(new_n8176, new_n8171, new_n8177);
nor_5  g05829(new_n8177, new_n8170, new_n8178);
or_5   g05830(new_n8178, new_n8169, new_n8179_1);
nor_5  g05831(new_n8179_1, new_n8167, new_n8180);
nor_5  g05832(new_n8180, new_n8166, new_n8181);
nor_5  g05833(new_n8181, new_n8164, new_n8182);
nor_5  g05834(new_n8182, new_n8163, new_n8183);
nor_5  g05835(new_n8183, new_n8161, new_n8184);
nor_5  g05836(new_n8184, new_n8160, new_n8185);
nor_5  g05837(new_n8185, new_n8158, new_n8186);
nor_5  g05838(new_n8186, new_n8157, new_n8187);
nor_5  g05839(new_n8187, new_n8155, new_n8188);
nor_5  g05840(new_n8188, new_n8154, new_n8189);
nor_5  g05841(new_n8189, new_n8152, new_n8190);
nor_5  g05842(new_n8190, new_n8151, new_n8191);
nor_5  g05843(new_n8191, new_n8149_1, new_n8192);
nor_5  g05844(new_n8192, new_n8148_1, new_n8193);
xnor_4 g05845(new_n8193, new_n8146, new_n8194_1);
xor_4  g05846(new_n8191, new_n8149_1, new_n8195);
xor_4  g05847(new_n8142, new_n8109_1, new_n8196);
nor_5  g05848(new_n8196, new_n8195, new_n8197);
xnor_4 g05849(new_n8196, new_n8195, new_n8198);
xnor_4 g05850(new_n8189, new_n8152, new_n8199);
xor_4  g05851(new_n8140, new_n8111, new_n8200);
and_5  g05852(new_n8200, new_n8199, new_n8201);
xnor_4 g05853(new_n8200, new_n8199, new_n8202);
xnor_4 g05854(new_n8187, new_n8155, new_n8203);
xor_4  g05855(new_n8138, new_n8113, new_n8204);
and_5  g05856(new_n8204, new_n8203, new_n8205);
xnor_4 g05857(new_n8204, new_n8203, new_n8206);
xnor_4 g05858(new_n8185, new_n8158, new_n8207);
xor_4  g05859(new_n8136, new_n8115, new_n8208);
and_5  g05860(new_n8208, new_n8207, new_n8209);
xnor_4 g05861(new_n8208, new_n8207, new_n8210);
xnor_4 g05862(new_n8183, new_n8161, new_n8211);
xor_4  g05863(new_n8134, new_n8117, new_n8212);
and_5  g05864(new_n8212, new_n8211, new_n8213);
xnor_4 g05865(new_n8212, new_n8211, new_n8214);
xnor_4 g05866(new_n8181, new_n8164, new_n8215_1);
xor_4  g05867(new_n8132, new_n8119, new_n8216);
and_5  g05868(new_n8216, new_n8215_1, new_n8217);
xnor_4 g05869(new_n8216, new_n8215_1, new_n8218);
xor_4  g05870(new_n8130_1, new_n8121, new_n8219);
not_10 g05871(new_n8219, new_n8220);
xor_4  g05872(new_n8179_1, new_n8167, new_n8221);
nor_5  g05873(new_n8221, new_n8220, new_n8222);
xor_4  g05874(new_n8128, new_n8123, new_n8223);
xnor_4 g05875(n27104, n18295, new_n8224);
xnor_4 g05876(new_n8224, new_n8177, new_n8225);
and_5  g05877(new_n8225, new_n8223, new_n8226);
xnor_4 g05878(new_n8225, new_n8223, new_n8227);
xnor_4 g05879(n15780, n6611, new_n8228);
xnor_4 g05880(new_n7059, new_n4085_1, new_n8229);
or_5   g05881(new_n8229, new_n8228, new_n8230);
xor_4  g05882(n27188, n6502, new_n8231);
xnor_4 g05883(new_n8231, new_n8175, new_n8232);
and_5  g05884(new_n8232, new_n8230, new_n8233);
xnor_4 g05885(new_n8126, new_n8125, new_n8234);
xor_4  g05886(new_n8232, new_n8230, new_n8235);
and_5  g05887(new_n8235, new_n8234, new_n8236);
nor_5  g05888(new_n8236, new_n8233, new_n8237);
nor_5  g05889(new_n8237, new_n8227, new_n8238);
nor_5  g05890(new_n8238, new_n8226, new_n8239);
xor_4  g05891(new_n8221, new_n8219, new_n8240);
nor_5  g05892(new_n8240, new_n8239, new_n8241);
nor_5  g05893(new_n8241, new_n8222, new_n8242);
nor_5  g05894(new_n8242, new_n8218, new_n8243);
nor_5  g05895(new_n8243, new_n8217, new_n8244_1);
nor_5  g05896(new_n8244_1, new_n8214, new_n8245);
nor_5  g05897(new_n8245, new_n8213, new_n8246);
nor_5  g05898(new_n8246, new_n8210, new_n8247);
nor_5  g05899(new_n8247, new_n8209, new_n8248);
nor_5  g05900(new_n8248, new_n8206, new_n8249);
nor_5  g05901(new_n8249, new_n8205, new_n8250);
nor_5  g05902(new_n8250, new_n8202, new_n8251);
nor_5  g05903(new_n8251, new_n8201, new_n8252);
nor_5  g05904(new_n8252, new_n8198, new_n8253);
nor_5  g05905(new_n8253, new_n8197, new_n8254);
xnor_4 g05906(new_n8254, new_n8194_1, n982);
nor_5  g05907(n26808, n7339, new_n8256_1);
not_10 g05908(new_n8256_1, new_n8257);
or_5   g05909(new_n8257, n1667, new_n8258);
or_5   g05910(new_n8258, n2680, new_n8259_1);
or_5   g05911(new_n8259_1, n2547, new_n8260);
or_5   g05912(new_n8260, n2999, new_n8261);
or_5   g05913(new_n8261, n14702, new_n8262);
nor_5  g05914(new_n8262, n13914, new_n8263);
not_10 g05915(new_n8263, new_n8264);
or_5   g05916(new_n8264, n3279, new_n8265);
xnor_4 g05917(new_n8265, n4306, new_n8266);
xor_4  g05918(n23166, n18105, new_n8267_1);
not_10 g05919(n10577, new_n8268);
nor_5  g05920(n24196, new_n8268, new_n8269);
xor_4  g05921(n24196, n10577, new_n8270);
not_10 g05922(n6381, new_n8271);
nor_5  g05923(n16376, new_n8271, new_n8272);
xor_4  g05924(n16376, n6381, new_n8273);
not_10 g05925(n14345, new_n8274);
nor_5  g05926(n25381, new_n8274, new_n8275);
xor_4  g05927(n25381, n14345, new_n8276_1);
not_10 g05928(n11356, new_n8277);
nor_5  g05929(n12587, new_n8277, new_n8278);
xor_4  g05930(n12587, n11356, new_n8279);
not_10 g05931(n3164, new_n8280);
or_5   g05932(new_n8280, n268, new_n8281);
xor_4  g05933(n3164, n268, new_n8282);
not_10 g05934(n10611, new_n8283);
or_5   g05935(n24879, new_n8283, new_n8284);
xor_4  g05936(n24879, n10611, new_n8285_1);
nor_5  g05937(new_n4137, n2783, new_n8286);
not_10 g05938(n2783, new_n8287);
nor_5  g05939(n6785, new_n8287, new_n8288_1);
nor_5  g05940(new_n7322, n15490, new_n8289);
not_10 g05941(n15490, new_n8290);
or_5   g05942(n24032, new_n8290, new_n8291);
nor_5  g05943(new_n7324, n18, new_n8292);
and_5  g05944(new_n8292, new_n8291, new_n8293);
nor_5  g05945(new_n8293, new_n8289, new_n8294);
nor_5  g05946(new_n8294, new_n8288_1, new_n8295);
nor_5  g05947(new_n8295, new_n8286, new_n8296);
not_10 g05948(new_n8296, new_n8297);
or_5   g05949(new_n8297, new_n8285_1, new_n8298);
and_5  g05950(new_n8298, new_n8284, new_n8299);
or_5   g05951(new_n8299, new_n8282, new_n8300);
and_5  g05952(new_n8300, new_n8281, new_n8301);
nor_5  g05953(new_n8301, new_n8279, new_n8302);
nor_5  g05954(new_n8302, new_n8278, new_n8303);
nor_5  g05955(new_n8303, new_n8276_1, new_n8304);
nor_5  g05956(new_n8304, new_n8275, new_n8305_1);
nor_5  g05957(new_n8305_1, new_n8273, new_n8306_1);
nor_5  g05958(new_n8306_1, new_n8272, new_n8307);
nor_5  g05959(new_n8307, new_n8270, new_n8308);
nor_5  g05960(new_n8308, new_n8269, new_n8309_1);
xnor_4 g05961(new_n8309_1, new_n8267_1, new_n8310);
xnor_4 g05962(new_n8310, new_n8266, new_n8311);
xnor_4 g05963(new_n8263, n3279, new_n8312);
xor_4  g05964(new_n8307, new_n8270, new_n8313);
and_5  g05965(new_n8313, new_n8312, new_n8314);
xnor_4 g05966(new_n8313, new_n8312, new_n8315);
xor_4  g05967(new_n8262, n13914, new_n8316);
xor_4  g05968(new_n8305_1, new_n8273, new_n8317);
nor_5  g05969(new_n8317, new_n8316, new_n8318);
xnor_4 g05970(new_n8317, new_n8316, new_n8319);
xor_4  g05971(new_n8261, n14702, new_n8320_1);
xor_4  g05972(new_n8303, new_n8276_1, new_n8321_1);
nor_5  g05973(new_n8321_1, new_n8320_1, new_n8322);
xnor_4 g05974(new_n8321_1, new_n8320_1, new_n8323);
xor_4  g05975(new_n8260, n2999, new_n8324_1);
xor_4  g05976(new_n8301, new_n8279, new_n8325);
nor_5  g05977(new_n8325, new_n8324_1, new_n8326);
xor_4  g05978(new_n8259_1, n2547, new_n8327);
xor_4  g05979(new_n8299, new_n8282, new_n8328);
nor_5  g05980(new_n8328, new_n8327, new_n8329);
xnor_4 g05981(new_n8328, new_n8327, new_n8330);
xor_4  g05982(new_n8258, n2680, new_n8331);
xnor_4 g05983(new_n8296, new_n8285_1, new_n8332);
nor_5  g05984(new_n8332, new_n8331, new_n8333);
xor_4  g05985(new_n8256_1, n1667, new_n8334);
xnor_4 g05986(n6785, n2783, new_n8335);
xnor_4 g05987(new_n8335, new_n8294, new_n8336);
and_5  g05988(new_n8336, new_n8334, new_n8337);
xnor_4 g05989(new_n8336, new_n8334, new_n8338);
xnor_4 g05990(n26808, n7339, new_n8339_1);
xor_4  g05991(n24032, n15490, new_n8340);
xnor_4 g05992(new_n8340, new_n8292, new_n8341);
nor_5  g05993(new_n8341, new_n8339_1, new_n8342);
not_10 g05994(n26808, new_n8343);
xnor_4 g05995(n22843, n18, new_n8344);
nor_5  g05996(new_n8344, new_n8343, new_n8345);
xor_4  g05997(new_n8341, new_n8339_1, new_n8346);
and_5  g05998(new_n8346, new_n8345, new_n8347);
or_5   g05999(new_n8347, new_n8342, new_n8348);
nor_5  g06000(new_n8348, new_n8338, new_n8349);
nor_5  g06001(new_n8349, new_n8337, new_n8350);
xnor_4 g06002(new_n8332, new_n8331, new_n8351);
nor_5  g06003(new_n8351, new_n8350, new_n8352);
nor_5  g06004(new_n8352, new_n8333, new_n8353);
nor_5  g06005(new_n8353, new_n8330, new_n8354);
nor_5  g06006(new_n8354, new_n8329, new_n8355);
xnor_4 g06007(new_n8325, new_n8324_1, new_n8356);
nor_5  g06008(new_n8356, new_n8355, new_n8357);
nor_5  g06009(new_n8357, new_n8326, new_n8358);
nor_5  g06010(new_n8358, new_n8323, new_n8359);
nor_5  g06011(new_n8359, new_n8322, new_n8360);
nor_5  g06012(new_n8360, new_n8319, new_n8361);
or_5   g06013(new_n8361, new_n8318, new_n8362);
nor_5  g06014(new_n8362, new_n8315, new_n8363_1);
nor_5  g06015(new_n8363_1, new_n8314, new_n8364);
xor_4  g06016(new_n8364, new_n8311, new_n8365);
xor_4  g06017(new_n8365, new_n4207, new_n8366);
not_10 g06018(new_n4211, new_n8367);
xor_4  g06019(new_n8362, new_n8315, new_n8368);
nor_5  g06020(new_n8368, new_n8367, new_n8369);
xor_4  g06021(new_n8368, new_n4211, new_n8370);
xor_4  g06022(new_n8360, new_n8319, new_n8371);
and_5  g06023(new_n8371, new_n4215_1, new_n8372);
xnor_4 g06024(new_n8371, new_n4215_1, new_n8373);
xor_4  g06025(new_n8358, new_n8323, new_n8374);
and_5  g06026(new_n8374, new_n4219, new_n8375);
xnor_4 g06027(new_n8374, new_n4219, new_n8376_1);
xor_4  g06028(new_n8356, new_n8355, new_n8377);
and_5  g06029(new_n8377, new_n4223, new_n8378);
xnor_4 g06030(new_n8377, new_n4223, new_n8379);
xor_4  g06031(new_n8353, new_n8330, new_n8380);
and_5  g06032(new_n8380, new_n4226, new_n8381_1);
xnor_4 g06033(new_n8380, new_n4226, new_n8382);
xor_4  g06034(new_n8351, new_n8350, new_n8383);
and_5  g06035(new_n8383, new_n4231_1, new_n8384);
xor_4  g06036(new_n8383, new_n4231_1, new_n8385);
xor_4  g06037(new_n8348, new_n8338, new_n8386);
nor_5  g06038(new_n8386, new_n4237, new_n8387);
xor_4  g06039(new_n8386, new_n4236, new_n8388);
not_10 g06040(new_n4239, new_n8389);
xor_4  g06041(new_n8346, new_n8345, new_n8390);
and_5  g06042(new_n8390, new_n8389, new_n8391);
xnor_4 g06043(new_n8344, n26808, new_n8392);
nand_5 g06044(new_n8392, new_n4243, new_n8393);
xor_4  g06045(new_n8390, new_n4239, new_n8394);
nor_5  g06046(new_n8394, new_n8393, new_n8395);
nor_5  g06047(new_n8395, new_n8391, new_n8396);
nor_5  g06048(new_n8396, new_n8388, new_n8397);
nor_5  g06049(new_n8397, new_n8387, new_n8398);
and_5  g06050(new_n8398, new_n8385, new_n8399_1);
nor_5  g06051(new_n8399_1, new_n8384, new_n8400);
nor_5  g06052(new_n8400, new_n8382, new_n8401);
nor_5  g06053(new_n8401, new_n8381_1, new_n8402);
nor_5  g06054(new_n8402, new_n8379, new_n8403);
nor_5  g06055(new_n8403, new_n8378, new_n8404);
nor_5  g06056(new_n8404, new_n8376_1, new_n8405_1);
nor_5  g06057(new_n8405_1, new_n8375, new_n8406);
nor_5  g06058(new_n8406, new_n8373, new_n8407);
nor_5  g06059(new_n8407, new_n8372, new_n8408_1);
nor_5  g06060(new_n8408_1, new_n8370, new_n8409);
nor_5  g06061(new_n8409, new_n8369, new_n8410);
xnor_4 g06062(new_n8410, new_n8366, n984);
xnor_4 g06063(new_n8404, new_n8376_1, n1005);
xnor_4 g06064(new_n3235_1, new_n3194, n1016);
xnor_4 g06065(new_n3836, new_n3823, n1020);
xnor_4 g06066(n18290, n12875, new_n8415);
nor_5  g06067(n11580, n2035, new_n8416);
xnor_4 g06068(n11580, n2035, new_n8417_1);
nor_5  g06069(n15884, n5213, new_n8418);
xnor_4 g06070(n15884, n5213, new_n8419);
nor_5  g06071(n6356, n4665, new_n8420);
xnor_4 g06072(n6356, n4665, new_n8421);
nor_5  g06073(n27104, n19005, new_n8422);
xnor_4 g06074(n27104, n19005, new_n8423);
nor_5  g06075(n27188, n4326, new_n8424);
and_5  g06076(n6611, n5438, new_n8425);
xnor_4 g06077(n27188, n4326, new_n8426);
nor_5  g06078(new_n8426, new_n8425, new_n8427);
nor_5  g06079(new_n8427, new_n8424, new_n8428);
nor_5  g06080(new_n8428, new_n8423, new_n8429);
nor_5  g06081(new_n8429, new_n8422, new_n8430);
nor_5  g06082(new_n8430, new_n8421, new_n8431);
nor_5  g06083(new_n8431, new_n8420, new_n8432_1);
nor_5  g06084(new_n8432_1, new_n8419, new_n8433);
nor_5  g06085(new_n8433, new_n8418, new_n8434);
nor_5  g06086(new_n8434, new_n8417_1, new_n8435);
nor_5  g06087(new_n8435, new_n8416, new_n8436);
xnor_4 g06088(new_n8436, new_n8415, new_n8437);
xnor_4 g06089(new_n8437, n23529, new_n8438);
xnor_4 g06090(new_n8434, new_n8417_1, new_n8439_1);
nor_5  g06091(new_n8439_1, n24620, new_n8440);
xnor_4 g06092(new_n8439_1, n24620, new_n8441);
xor_4  g06093(new_n8432_1, new_n8419, new_n8442);
and_5  g06094(new_n8442, new_n8162, new_n8443);
xor_4  g06095(new_n8442, n5211, new_n8444);
xnor_4 g06096(new_n8430, new_n8421, new_n8445);
nor_5  g06097(new_n8445, n12956, new_n8446);
xnor_4 g06098(new_n8445, n12956, new_n8447);
xnor_4 g06099(new_n8428, new_n8423, new_n8448);
nor_5  g06100(new_n8448, n18295, new_n8449);
xnor_4 g06101(new_n8426, new_n8425, new_n8450);
and_5  g06102(new_n8450, n6502, new_n8451);
xor_4  g06103(n6611, n5438, new_n8452);
nand_5 g06104(new_n8452, n15780, new_n8453_1);
xnor_4 g06105(new_n8450, n6502, new_n8454);
nor_5  g06106(new_n8454, new_n8453_1, new_n8455);
nor_5  g06107(new_n8455, new_n8451, new_n8456);
xor_4  g06108(new_n8448, n18295, new_n8457);
and_5  g06109(new_n8457, new_n8456, new_n8458);
nor_5  g06110(new_n8458, new_n8449, new_n8459);
nor_5  g06111(new_n8459, new_n8447, new_n8460);
nor_5  g06112(new_n8460, new_n8446, new_n8461);
nor_5  g06113(new_n8461, new_n8444, new_n8462);
nor_5  g06114(new_n8462, new_n8443, new_n8463);
nor_5  g06115(new_n8463, new_n8441, new_n8464);
nor_5  g06116(new_n8464, new_n8440, new_n8465);
xor_4  g06117(new_n8465, new_n8438, new_n8466);
xnor_4 g06118(n17250, n4409, new_n8467);
nor_5  g06119(n23160, n3570, new_n8468);
xnor_4 g06120(n23160, n3570, new_n8469);
nor_5  g06121(n16524, n13668, new_n8470);
xnor_4 g06122(n16524, n13668, new_n8471);
nor_5  g06123(n21276, n11056, new_n8472);
xnor_4 g06124(n21276, n11056, new_n8473);
nor_5  g06125(n26748, n15271, new_n8474);
xnor_4 g06126(n26748, n15271, new_n8475);
nor_5  g06127(n25877, n10057, new_n8476);
and_5  g06128(n24323, n8920, new_n8477);
xnor_4 g06129(n25877, n10057, new_n8478);
nor_5  g06130(new_n8478, new_n8477, new_n8479);
nor_5  g06131(new_n8479, new_n8476, new_n8480_1);
nor_5  g06132(new_n8480_1, new_n8475, new_n8481);
nor_5  g06133(new_n8481, new_n8474, new_n8482);
nor_5  g06134(new_n8482, new_n8473, new_n8483);
nor_5  g06135(new_n8483, new_n8472, new_n8484);
nor_5  g06136(new_n8484, new_n8471, new_n8485);
nor_5  g06137(new_n8485, new_n8470, new_n8486);
nor_5  g06138(new_n8486, new_n8469, new_n8487);
nor_5  g06139(new_n8487, new_n8468, new_n8488);
xnor_4 g06140(new_n8488, new_n8467, new_n8489_1);
xnor_4 g06141(new_n8489_1, n11044, new_n8490);
xnor_4 g06142(new_n8486, new_n8469, new_n8491);
and_5  g06143(new_n8491, n2421, new_n8492);
xnor_4 g06144(new_n8491, n2421, new_n8493);
xnor_4 g06145(new_n8484, new_n8471, new_n8494);
and_5  g06146(new_n8494, n987, new_n8495);
xnor_4 g06147(new_n8494, n987, new_n8496);
xnor_4 g06148(new_n8482, new_n8473, new_n8497);
and_5  g06149(new_n8497, n20478, new_n8498);
xnor_4 g06150(new_n8497, n20478, new_n8499);
xnor_4 g06151(new_n8480_1, new_n8475, new_n8500);
and_5  g06152(new_n8500, n26882, new_n8501);
xnor_4 g06153(new_n8478, new_n8477, new_n8502);
nor_5  g06154(new_n8502, n22619, new_n8503);
xor_4  g06155(n24323, n8920, new_n8504);
nand_5 g06156(new_n8504, n6775, new_n8505_1);
xor_4  g06157(new_n8502, n22619, new_n8506);
and_5  g06158(new_n8506, new_n8505_1, new_n8507);
nor_5  g06159(new_n8507, new_n8503, new_n8508);
xor_4  g06160(new_n8500, n26882, new_n8509);
and_5  g06161(new_n8509, new_n8508, new_n8510_1);
nor_5  g06162(new_n8510_1, new_n8501, new_n8511);
nor_5  g06163(new_n8511, new_n8499, new_n8512);
nor_5  g06164(new_n8512, new_n8498, new_n8513);
nor_5  g06165(new_n8513, new_n8496, new_n8514);
nor_5  g06166(new_n8514, new_n8495, new_n8515);
nor_5  g06167(new_n8515, new_n8493, new_n8516);
nor_5  g06168(new_n8516, new_n8492, new_n8517);
xor_4  g06169(new_n8517, new_n8490, new_n8518);
xnor_4 g06170(new_n8518, new_n8466, new_n8519_1);
xor_4  g06171(new_n8463, new_n8441, new_n8520);
xor_4  g06172(new_n8515, new_n8493, new_n8521);
and_5  g06173(new_n8521, new_n8520, new_n8522);
xnor_4 g06174(new_n8521, new_n8520, new_n8523);
xor_4  g06175(new_n8461, new_n8444, new_n8524);
xor_4  g06176(new_n8513, new_n8496, new_n8525);
and_5  g06177(new_n8525, new_n8524, new_n8526_1);
xnor_4 g06178(new_n8525, new_n8524, new_n8527);
xor_4  g06179(new_n8459, new_n8447, new_n8528);
xor_4  g06180(new_n8511, new_n8499, new_n8529);
and_5  g06181(new_n8529, new_n8528, new_n8530);
xnor_4 g06182(new_n8529, new_n8528, new_n8531);
xor_4  g06183(new_n8457, new_n8456, new_n8532);
xor_4  g06184(new_n8509, new_n8508, new_n8533);
and_5  g06185(new_n8533, new_n8532, new_n8534);
xnor_4 g06186(new_n8533, new_n8532, new_n8535_1);
xor_4  g06187(new_n8506, new_n8505_1, new_n8536);
xor_4  g06188(new_n8454, new_n8453_1, new_n8537);
nor_5  g06189(new_n8537, new_n8536, new_n8538);
xor_4  g06190(new_n8504, n6775, new_n8539);
not_10 g06191(new_n8539, new_n8540);
xor_4  g06192(new_n8452, n15780, new_n8541);
nor_5  g06193(new_n8541, new_n8540, new_n8542);
xor_4  g06194(new_n8537, new_n8536, new_n8543);
and_5  g06195(new_n8543, new_n8542, new_n8544);
nor_5  g06196(new_n8544, new_n8538, new_n8545);
nor_5  g06197(new_n8545, new_n8535_1, new_n8546);
nor_5  g06198(new_n8546, new_n8534, new_n8547);
nor_5  g06199(new_n8547, new_n8531, new_n8548);
nor_5  g06200(new_n8548, new_n8530, new_n8549);
nor_5  g06201(new_n8549, new_n8527, new_n8550_1);
nor_5  g06202(new_n8550_1, new_n8526_1, new_n8551);
nor_5  g06203(new_n8551, new_n8523, new_n8552);
nor_5  g06204(new_n8552, new_n8522, new_n8553);
xnor_4 g06205(new_n8553, new_n8519_1, n1044);
or_5   g06206(n22619, n6775, new_n8555);
or_5   g06207(new_n8555, n26882, new_n8556);
xor_4  g06208(new_n8556, n20478, new_n8557);
xnor_4 g06209(new_n8557, n7305, new_n8558);
xor_4  g06210(new_n8555, n26882, new_n8559);
and_5  g06211(new_n8559, n25872, new_n8560);
xnor_4 g06212(new_n8559, n25872, new_n8561);
xor_4  g06213(n22619, n6775, new_n8562);
and_5  g06214(new_n8562, n20259, new_n8563_1);
and_5  g06215(n6775, n3925, new_n8564);
xor_4  g06216(new_n8562, n20259, new_n8565);
and_5  g06217(new_n8565, new_n8564, new_n8566);
nor_5  g06218(new_n8566, new_n8563_1, new_n8567);
nor_5  g06219(new_n8567, new_n8561, new_n8568);
nor_5  g06220(new_n8568, new_n8560, new_n8569);
xor_4  g06221(new_n8569, new_n8558, new_n8570);
or_5   g06222(n9399, n2088, new_n8571);
or_5   g06223(new_n8571, n16396, new_n8572);
xor_4  g06224(new_n8572, n25074, new_n8573);
xnor_4 g06225(new_n8573, n3480, new_n8574);
xor_4  g06226(new_n8571, n16396, new_n8575);
and_5  g06227(new_n8575, n16722, new_n8576);
xnor_4 g06228(new_n8575, n16722, new_n8577);
nor_5  g06229(new_n5325_1, new_n5320, new_n8578);
or_5   g06230(new_n8578, new_n5322, new_n8579);
nor_5  g06231(new_n8579, new_n8577, new_n8580);
nor_5  g06232(new_n8580, new_n8576, new_n8581_1);
xor_4  g06233(new_n8581_1, new_n8574, new_n8582);
xnor_4 g06234(new_n8582, new_n8570, new_n8583);
xnor_4 g06235(new_n8579, new_n8577, new_n8584);
xor_4  g06236(new_n8567, new_n8561, new_n8585);
not_10 g06237(new_n8585, new_n8586);
nor_5  g06238(new_n8586, new_n8584, new_n8587);
xor_4  g06239(new_n8585, new_n8584, new_n8588);
xor_4  g06240(new_n8565, new_n8564, new_n8589);
not_10 g06241(new_n8589, new_n8590);
nor_5  g06242(new_n8590, new_n5326, new_n8591);
xnor_4 g06243(n6775, n3925, new_n8592);
or_5   g06244(new_n8592, new_n5311, new_n8593);
xor_4  g06245(new_n8589, new_n5326, new_n8594_1);
nor_5  g06246(new_n8594_1, new_n8593, new_n8595);
nor_5  g06247(new_n8595, new_n8591, new_n8596);
nor_5  g06248(new_n8596, new_n8588, new_n8597);
nor_5  g06249(new_n8597, new_n8587, new_n8598);
xor_4  g06250(new_n8598, new_n8583, new_n8599);
xor_4  g06251(n12956, n7057, new_n8600);
nor_5  g06252(new_n8168, n8381, new_n8601);
not_10 g06253(n8381, new_n8602);
nor_5  g06254(n18295, new_n8602, new_n8603);
nor_5  g06255(n20235, new_n8172, new_n8604);
or_5   g06256(new_n4660, n6502, new_n8605);
not_10 g06257(n12495, new_n8606);
and_5  g06258(n15780, new_n8606, new_n8607);
and_5  g06259(new_n8607, new_n8605, new_n8608_1);
nor_5  g06260(new_n8608_1, new_n8604, new_n8609);
nor_5  g06261(new_n8609, new_n8603, new_n8610);
nor_5  g06262(new_n8610, new_n8601, new_n8611);
xor_4  g06263(new_n8611, new_n8600, new_n8612);
xor_4  g06264(new_n8612, new_n8599, new_n8613);
xnor_4 g06265(new_n8596, new_n8588, new_n8614_1);
xnor_4 g06266(n18295, n8381, new_n8615);
xnor_4 g06267(new_n8615, new_n8609, new_n8616);
and_5  g06268(new_n8616, new_n8614_1, new_n8617);
xnor_4 g06269(new_n8616, new_n8614_1, new_n8618);
xnor_4 g06270(n15780, n12495, new_n8619);
xnor_4 g06271(new_n8592, new_n5311, new_n8620_1);
or_5   g06272(new_n8620_1, new_n8619, new_n8621);
xor_4  g06273(n20235, n6502, new_n8622);
xnor_4 g06274(new_n8622, new_n8607, new_n8623);
and_5  g06275(new_n8623, new_n8621, new_n8624);
xnor_4 g06276(new_n8594_1, new_n8593, new_n8625);
xor_4  g06277(new_n8623, new_n8621, new_n8626);
and_5  g06278(new_n8626, new_n8625, new_n8627);
nor_5  g06279(new_n8627, new_n8624, new_n8628);
nor_5  g06280(new_n8628, new_n8618, new_n8629);
or_5   g06281(new_n8629, new_n8617, new_n8630);
xor_4  g06282(new_n8630, new_n8613, n1060);
xnor_4 g06283(new_n3233, new_n3198, n1069);
xnor_4 g06284(n9832, n3959, new_n8633);
nor_5  g06285(n11566, n1558, new_n8634);
xnor_4 g06286(n11566, n1558, new_n8635);
nor_5  g06287(n26744, n21749, new_n8636);
xnor_4 g06288(n26744, n21749, new_n8637_1);
nor_5  g06289(n26625, n7769, new_n8638_1);
and_5  g06290(n21138, n14230, new_n8639);
xnor_4 g06291(n26625, n7769, new_n8640);
nor_5  g06292(new_n8640, new_n8639, new_n8641);
nor_5  g06293(new_n8641, new_n8638_1, new_n8642);
nor_5  g06294(new_n8642, new_n8637_1, new_n8643);
nor_5  g06295(new_n8643, new_n8636, new_n8644);
nor_5  g06296(new_n8644, new_n8635, new_n8645);
nor_5  g06297(new_n8645, new_n8634, new_n8646);
xnor_4 g06298(new_n8646, new_n8633, new_n8647);
or_5   g06299(n26167, n22591, new_n8648);
or_5   g06300(new_n8648, n17095, new_n8649);
or_5   g06301(new_n8649, n15378, new_n8650);
xor_4  g06302(new_n8650, n19575, new_n8651);
xnor_4 g06303(new_n6166, n5226, new_n8652);
and_5  g06304(new_n6169, n17664, new_n8653);
xnor_4 g06305(new_n6169, n17664, new_n8654);
and_5  g06306(new_n6172, n23369, new_n8655);
xor_4  g06307(new_n6172, n23369, new_n8656_1);
nor_5  g06308(new_n6179, n1136, new_n8657);
nand_5 g06309(new_n6175, n19234, new_n8658);
xnor_4 g06310(new_n6178, n1136, new_n8659);
and_5  g06311(new_n8659, new_n8658, new_n8660);
nor_5  g06312(new_n8660, new_n8657, new_n8661);
and_5  g06313(new_n8661, new_n8656_1, new_n8662_1);
nor_5  g06314(new_n8662_1, new_n8655, new_n8663);
nor_5  g06315(new_n8663, new_n8654, new_n8664);
nor_5  g06316(new_n8664, new_n8653, new_n8665);
xor_4  g06317(new_n8665, new_n8652, new_n8666);
xnor_4 g06318(new_n8666, new_n8651, new_n8667);
xor_4  g06319(new_n8663, new_n8654, new_n8668);
xor_4  g06320(new_n8649, n15378, new_n8669);
nor_5  g06321(new_n8669, new_n8668, new_n8670);
xnor_4 g06322(new_n8669, new_n8668, new_n8671);
xor_4  g06323(new_n8661, new_n8656_1, new_n8672);
xor_4  g06324(new_n8648, n17095, new_n8673);
nor_5  g06325(new_n8673, new_n8672, new_n8674);
xnor_4 g06326(new_n8673, new_n8672, new_n8675);
xor_4  g06327(new_n8659, new_n8658, new_n8676);
not_10 g06328(n26167, new_n8677);
nor_5  g06329(new_n6523, new_n8677, new_n8678_1);
xnor_4 g06330(new_n8678_1, n22591, new_n8679);
nor_5  g06331(new_n8679, new_n8676, new_n8680);
nand_5 g06332(new_n6523, n26167, new_n8681);
nor_5  g06333(new_n8681, n22591, new_n8682);
or_5   g06334(new_n8682, new_n8680, new_n8683);
nor_5  g06335(new_n8683, new_n8675, new_n8684);
nor_5  g06336(new_n8684, new_n8674, new_n8685);
nor_5  g06337(new_n8685, new_n8671, new_n8686);
nor_5  g06338(new_n8686, new_n8670, new_n8687_1);
xor_4  g06339(new_n8687_1, new_n8667, new_n8688);
xnor_4 g06340(new_n8688, new_n8647, new_n8689);
xnor_4 g06341(new_n8685, new_n8671, new_n8690);
xor_4  g06342(new_n8644, new_n8635, new_n8691);
nor_5  g06343(new_n8691, new_n8690, new_n8692);
xor_4  g06344(new_n8691, new_n8690, new_n8693);
xnor_4 g06345(new_n8683, new_n8675, new_n8694_1);
xor_4  g06346(new_n8642, new_n8637_1, new_n8695);
and_5  g06347(new_n8695, new_n8694_1, new_n8696);
xnor_4 g06348(new_n8695, new_n8694_1, new_n8697);
not_10 g06349(new_n8676, new_n8698);
xnor_4 g06350(new_n8679, new_n8698, new_n8699);
xor_4  g06351(new_n8640, new_n8639, new_n8700);
nor_5  g06352(new_n8700, new_n8699, new_n8701);
nor_5  g06353(new_n6524, new_n6522, new_n8702);
xor_4  g06354(new_n8700, new_n8699, new_n8703);
and_5  g06355(new_n8703, new_n8702, new_n8704);
or_5   g06356(new_n8704, new_n8701, new_n8705);
nor_5  g06357(new_n8705, new_n8697, new_n8706);
nor_5  g06358(new_n8706, new_n8696, new_n8707);
and_5  g06359(new_n8707, new_n8693, new_n8708);
or_5   g06360(new_n8708, new_n8692, new_n8709);
xor_4  g06361(new_n8709, new_n8689, n1111);
xnor_4 g06362(new_n2569, n25475, new_n8711);
and_5  g06363(new_n2572, n23849, new_n8712);
xnor_4 g06364(new_n2572, n23849, new_n8713);
and_5  g06365(new_n2575, n12446, new_n8714);
nor_5  g06366(new_n2577, n11011, new_n8715);
xnor_4 g06367(new_n2577, n11011, new_n8716_1);
or_5   g06368(new_n2580, n16029, new_n8717);
xnor_4 g06369(new_n2580, n16029, new_n8718);
and_5  g06370(new_n2583, n16476, new_n8719);
xnor_4 g06371(new_n2583, n16476, new_n8720);
and_5  g06372(new_n2586, n11615, new_n8721_1);
and_5  g06373(new_n2588, new_n3712, new_n8722);
nand_5 g06374(new_n2591, n14090, new_n8723);
xnor_4 g06375(new_n2588, n22433, new_n8724);
and_5  g06376(new_n8724, new_n8723, new_n8725);
nor_5  g06377(new_n8725, new_n8722, new_n8726);
xor_4  g06378(new_n2586, n11615, new_n8727);
and_5  g06379(new_n8727, new_n8726, new_n8728);
nor_5  g06380(new_n8728, new_n8721_1, new_n8729);
nor_5  g06381(new_n8729, new_n8720, new_n8730);
nor_5  g06382(new_n8730, new_n8719, new_n8731);
not_10 g06383(new_n8731, new_n8732);
or_5   g06384(new_n8732, new_n8718, new_n8733);
and_5  g06385(new_n8733, new_n8717, new_n8734);
nor_5  g06386(new_n8734, new_n8716_1, new_n8735);
or_5   g06387(new_n8735, new_n8715, new_n8736);
xnor_4 g06388(new_n2575, n12446, new_n8737);
nor_5  g06389(new_n8737, new_n8736, new_n8738);
nor_5  g06390(new_n8738, new_n8714, new_n8739);
nor_5  g06391(new_n8739, new_n8713, new_n8740);
nor_5  g06392(new_n8740, new_n8712, new_n8741);
xnor_4 g06393(new_n8741, new_n8711, new_n8742);
or_5   g06394(new_n8572, n25074, new_n8743);
or_5   g06395(new_n8743, n8006, new_n8744_1);
or_5   g06396(new_n8744_1, n20929, new_n8745_1);
or_5   g06397(new_n8745_1, n10710, new_n8746);
or_5   g06398(new_n8746, n11841, new_n8747);
xor_4  g06399(new_n8747, n27089, new_n8748);
xnor_4 g06400(new_n8748, new_n2660, new_n8749);
xor_4  g06401(new_n8746, n11841, new_n8750);
and_5  g06402(new_n8750, new_n2665, new_n8751);
xor_4  g06403(new_n8750, new_n2665, new_n8752);
xor_4  g06404(new_n8745_1, n10710, new_n8753);
nor_5  g06405(new_n8753, new_n2669, new_n8754);
xnor_4 g06406(new_n8753, new_n2669, new_n8755);
xor_4  g06407(new_n8744_1, n20929, new_n8756);
nor_5  g06408(new_n8756, new_n2673, new_n8757);
xnor_4 g06409(new_n8756, new_n2673, new_n8758);
xor_4  g06410(new_n8743, n8006, new_n8759);
nor_5  g06411(new_n8759, new_n2677, new_n8760);
nor_5  g06412(new_n8573, new_n2680_1, new_n8761);
xnor_4 g06413(new_n8573, new_n2680_1, new_n8762);
nor_5  g06414(new_n8575, new_n2684, new_n8763);
xnor_4 g06415(new_n8575, new_n2684, new_n8764);
nor_5  g06416(new_n5320, new_n2688, new_n8765);
nor_5  g06417(new_n2690, n2088, new_n8766);
xor_4  g06418(new_n5320, new_n2688, new_n8767);
and_5  g06419(new_n8767, new_n8766, new_n8768);
nor_5  g06420(new_n8768, new_n8765, new_n8769);
nor_5  g06421(new_n8769, new_n8764, new_n8770);
nor_5  g06422(new_n8770, new_n8763, new_n8771);
nor_5  g06423(new_n8771, new_n8762, new_n8772);
nor_5  g06424(new_n8772, new_n8761, new_n8773);
xnor_4 g06425(new_n8759, new_n2677, new_n8774);
nor_5  g06426(new_n8774, new_n8773, new_n8775);
nor_5  g06427(new_n8775, new_n8760, new_n8776);
nor_5  g06428(new_n8776, new_n8758, new_n8777);
nor_5  g06429(new_n8777, new_n8757, new_n8778);
nor_5  g06430(new_n8778, new_n8755, new_n8779);
nor_5  g06431(new_n8779, new_n8754, new_n8780);
and_5  g06432(new_n8780, new_n8752, new_n8781);
nor_5  g06433(new_n8781, new_n8751, new_n8782_1);
xor_4  g06434(new_n8782_1, new_n8749, new_n8783);
xnor_4 g06435(new_n8783, new_n8742, new_n8784);
xor_4  g06436(new_n8739, new_n8713, new_n8785);
xor_4  g06437(new_n8780, new_n8752, new_n8786);
and_5  g06438(new_n8786, new_n8785, new_n8787);
xnor_4 g06439(new_n8786, new_n8785, new_n8788);
xnor_4 g06440(new_n8737, new_n8736, new_n8789);
xor_4  g06441(new_n8778, new_n8755, new_n8790);
and_5  g06442(new_n8790, new_n8789, new_n8791);
xor_4  g06443(new_n8737, new_n8736, new_n8792);
xnor_4 g06444(new_n8790, new_n8792, new_n8793);
xor_4  g06445(new_n8734, new_n8716_1, new_n8794);
xor_4  g06446(new_n8776, new_n8758, new_n8795);
nor_5  g06447(new_n8795, new_n8794, new_n8796);
xnor_4 g06448(new_n8795, new_n8794, new_n8797);
xnor_4 g06449(new_n8731, new_n8718, new_n8798);
xor_4  g06450(new_n8774, new_n8773, new_n8799);
nor_5  g06451(new_n8799, new_n8798, new_n8800);
xnor_4 g06452(new_n8799, new_n8798, new_n8801);
xor_4  g06453(new_n8771, new_n8762, new_n8802);
xnor_4 g06454(new_n8729, new_n8720, new_n8803_1);
nor_5  g06455(new_n8803_1, new_n8802, new_n8804);
xnor_4 g06456(new_n8803_1, new_n8802, new_n8805);
xnor_4 g06457(new_n8769, new_n8764, new_n8806_1);
xor_4  g06458(new_n8727, new_n8726, new_n8807);
and_5  g06459(new_n8807, new_n8806_1, new_n8808);
xnor_4 g06460(new_n8807, new_n8806_1, new_n8809_1);
xnor_4 g06461(new_n8767, new_n8766, new_n8810);
xor_4  g06462(new_n8724, new_n8723, new_n8811);
not_10 g06463(new_n8811, new_n8812);
nor_5  g06464(new_n8812, new_n8810, new_n8813);
xor_4  g06465(new_n2591, n14090, new_n8814);
not_10 g06466(new_n8814, new_n8815);
xor_4  g06467(new_n2690, n2088, new_n8816);
or_5   g06468(new_n8816, new_n8815, new_n8817);
xnor_4 g06469(new_n8811, new_n8810, new_n8818);
and_5  g06470(new_n8818, new_n8817, new_n8819);
or_5   g06471(new_n8819, new_n8813, new_n8820);
nor_5  g06472(new_n8820, new_n8809_1, new_n8821_1);
nor_5  g06473(new_n8821_1, new_n8808, new_n8822);
nor_5  g06474(new_n8822, new_n8805, new_n8823);
nor_5  g06475(new_n8823, new_n8804, new_n8824_1);
nor_5  g06476(new_n8824_1, new_n8801, new_n8825);
nor_5  g06477(new_n8825, new_n8800, new_n8826);
nor_5  g06478(new_n8826, new_n8797, new_n8827_1);
nor_5  g06479(new_n8827_1, new_n8796, new_n8828);
and_5  g06480(new_n8828, new_n8793, new_n8829);
or_5   g06481(new_n8829, new_n8791, new_n8830);
nor_5  g06482(new_n8830, new_n8788, new_n8831);
nor_5  g06483(new_n8831, new_n8787, new_n8832);
xnor_4 g06484(new_n8832, new_n8784, n1119);
xnor_4 g06485(new_n7169, new_n7168, new_n8834);
xnor_4 g06486(new_n8834, new_n7188, n1120);
xnor_4 g06487(n9246, n3925, new_n8836);
xnor_4 g06488(new_n8836, new_n7060, new_n8837);
xnor_4 g06489(n12495, n7428, new_n8838);
xor_4  g06490(new_n8838, new_n8837, n1196);
xor_4  g06491(n16223, n15636, new_n8840);
nor_5  g06492(new_n5096, n19494, new_n8841);
or_5   g06493(n20077, new_n2364, new_n8842);
nor_5  g06494(new_n5098_1, n2387, new_n8843);
and_5  g06495(new_n8843, new_n8842, new_n8844);
nor_5  g06496(new_n8844, new_n8841, new_n8845);
xor_4  g06497(new_n8845, new_n8840, new_n8846);
xnor_4 g06498(new_n8846, new_n7173, new_n8847);
xnor_4 g06499(n6794, n2387, new_n8848);
or_5   g06500(new_n8848, new_n7179, new_n8849_1);
xor_4  g06501(n20077, n19494, new_n8850);
xnor_4 g06502(new_n8850, new_n8843, new_n8851);
and_5  g06503(new_n8851, new_n8849_1, new_n8852);
xor_4  g06504(new_n8851, new_n8849_1, new_n8853);
and_5  g06505(new_n8853, new_n7174, new_n8854);
nor_5  g06506(new_n8854, new_n8852, new_n8855);
xnor_4 g06507(new_n8855, new_n8847, n1237);
xor_4  g06508(new_n5245, new_n5070, new_n8857);
xnor_4 g06509(new_n8857, new_n5306, n1239);
xnor_4 g06510(n22764, n1536, new_n8859);
nor_5  g06511(n26264, n19454, new_n8860);
xnor_4 g06512(n26264, n19454, new_n8861_1);
nor_5  g06513(n9445, n7841, new_n8862_1);
xnor_4 g06514(n9445, n7841, new_n8863);
nor_5  g06515(n16812, n1279, new_n8864);
xnor_4 g06516(n16812, n1279, new_n8865);
nor_5  g06517(n25068, n8324, new_n8866);
xnor_4 g06518(n25068, n8324, new_n8867);
nor_5  g06519(n12546, n2331, new_n8868);
xnor_4 g06520(n12546, n2331, new_n8869_1);
nor_5  g06521(n22631, n21078, new_n8870);
xnor_4 g06522(n22631, n21078, new_n8871);
nor_5  g06523(n24485, n16743, new_n8872);
xnor_4 g06524(n24485, n16743, new_n8873);
nor_5  g06525(n15258, n2420, new_n8874);
and_5  g06526(n22201, n4588, new_n8875);
xnor_4 g06527(n15258, n2420, new_n8876);
nor_5  g06528(new_n8876, new_n8875, new_n8877);
nor_5  g06529(new_n8877, new_n8874, new_n8878);
nor_5  g06530(new_n8878, new_n8873, new_n8879);
nor_5  g06531(new_n8879, new_n8872, new_n8880);
nor_5  g06532(new_n8880, new_n8871, new_n8881);
nor_5  g06533(new_n8881, new_n8870, new_n8882);
nor_5  g06534(new_n8882, new_n8869_1, new_n8883);
nor_5  g06535(new_n8883, new_n8868, new_n8884_1);
nor_5  g06536(new_n8884_1, new_n8867, new_n8885);
nor_5  g06537(new_n8885, new_n8866, new_n8886);
nor_5  g06538(new_n8886, new_n8865, new_n8887);
nor_5  g06539(new_n8887, new_n8864, new_n8888);
nor_5  g06540(new_n8888, new_n8863, new_n8889);
nor_5  g06541(new_n8889, new_n8862_1, new_n8890);
nor_5  g06542(new_n8890, new_n8861_1, new_n8891);
nor_5  g06543(new_n8891, new_n8860, new_n8892);
xnor_4 g06544(new_n8892, new_n8859, new_n8893);
nor_5  g06545(new_n8893, n2416, new_n8894);
xnor_4 g06546(new_n8893, n2416, new_n8895);
xnor_4 g06547(new_n8890, new_n8861_1, new_n8896);
nor_5  g06548(new_n8896, n21905, new_n8897);
xnor_4 g06549(new_n8896, n21905, new_n8898);
xnor_4 g06550(new_n8888, new_n8863, new_n8899);
nor_5  g06551(new_n8899, n22918, new_n8900);
xnor_4 g06552(new_n8899, n22918, new_n8901);
xnor_4 g06553(new_n8886, new_n8865, new_n8902);
nor_5  g06554(new_n8902, n25923, new_n8903);
xnor_4 g06555(new_n8902, n25923, new_n8904);
xnor_4 g06556(new_n8884_1, new_n8867, new_n8905);
nor_5  g06557(new_n8905, n6790, new_n8906);
xnor_4 g06558(new_n8905, n6790, new_n8907);
xnor_4 g06559(new_n8882, new_n8869_1, new_n8908);
nor_5  g06560(new_n8908, n22879, new_n8909_1);
xnor_4 g06561(new_n8908, n22879, new_n8910);
xnor_4 g06562(new_n8880, new_n8871, new_n8911_1);
nor_5  g06563(new_n8911_1, n2117, new_n8912);
xnor_4 g06564(new_n8911_1, n2117, new_n8913);
xnor_4 g06565(new_n8878, new_n8873, new_n8914);
nor_5  g06566(new_n8914, n5882, new_n8915);
xnor_4 g06567(new_n8876, new_n8875, new_n8916);
nor_5  g06568(new_n8916, n11775, new_n8917);
xor_4  g06569(n22201, n4588, new_n8918);
nand_5 g06570(new_n8918, n27134, new_n8919);
xor_4  g06571(new_n8916, n11775, new_n8920_1);
and_5  g06572(new_n8920_1, new_n8919, new_n8921);
nor_5  g06573(new_n8921, new_n8917, new_n8922);
xnor_4 g06574(new_n8914, n5882, new_n8923);
nor_5  g06575(new_n8923, new_n8922, new_n8924);
nor_5  g06576(new_n8924, new_n8915, new_n8925);
nor_5  g06577(new_n8925, new_n8913, new_n8926);
nor_5  g06578(new_n8926, new_n8912, new_n8927);
nor_5  g06579(new_n8927, new_n8910, new_n8928);
nor_5  g06580(new_n8928, new_n8909_1, new_n8929);
nor_5  g06581(new_n8929, new_n8907, new_n8930);
nor_5  g06582(new_n8930, new_n8906, new_n8931);
nor_5  g06583(new_n8931, new_n8904, new_n8932);
nor_5  g06584(new_n8932, new_n8903, new_n8933);
nor_5  g06585(new_n8933, new_n8901, new_n8934);
nor_5  g06586(new_n8934, new_n8900, new_n8935);
nor_5  g06587(new_n8935, new_n8898, new_n8936);
nor_5  g06588(new_n8936, new_n8897, new_n8937);
nor_5  g06589(new_n8937, new_n8895, new_n8938);
nor_5  g06590(new_n8938, new_n8894, new_n8939);
nor_5  g06591(n22764, n1536, new_n8940);
nor_5  g06592(new_n8892, new_n8859, new_n8941);
nor_5  g06593(new_n8941, new_n8940, new_n8942);
and_5  g06594(new_n8942, new_n8939, new_n8943_1);
nor_5  g06595(n23493, n8405, new_n8944);
nor_5  g06596(n22359, n10275, new_n8945);
nor_5  g06597(n15146, n5532, new_n8946);
nor_5  g06598(n11579, n3962, new_n8947);
nor_5  g06599(n23513, n21, new_n8948);
xnor_4 g06600(n23513, n21, new_n8949);
nor_5  g06601(n6427, n1682, new_n8950);
and_5  g06602(n6427, n1682, new_n8951);
nor_5  g06603(n7963, n6590, new_n8952);
nor_5  g06604(n20349, n10017, new_n8953);
and_5  g06605(n15936, n3618, new_n8954);
and_5  g06606(n20349, n10017, new_n8955);
nor_5  g06607(new_n8955, new_n8954, new_n8956);
nor_5  g06608(new_n8956, new_n8953, new_n8957);
and_5  g06609(n7963, n6590, new_n8958);
nor_5  g06610(new_n8958, new_n8957, new_n8959);
nor_5  g06611(new_n8959, new_n8952, new_n8960);
nor_5  g06612(new_n8960, new_n8951, new_n8961);
nor_5  g06613(new_n8961, new_n8950, new_n8962);
nor_5  g06614(new_n8962, new_n8949, new_n8963);
nor_5  g06615(new_n8963, new_n8948, new_n8964_1);
xnor_4 g06616(n11579, n3962, new_n8965);
nor_5  g06617(new_n8965, new_n8964_1, new_n8966);
nor_5  g06618(new_n8966, new_n8947, new_n8967);
xnor_4 g06619(n15146, n5532, new_n8968);
nor_5  g06620(new_n8968, new_n8967, new_n8969);
nor_5  g06621(new_n8969, new_n8946, new_n8970);
xnor_4 g06622(n22359, n10275, new_n8971_1);
nor_5  g06623(new_n8971_1, new_n8970, new_n8972);
nor_5  g06624(new_n8972, new_n8945, new_n8973);
xnor_4 g06625(n23493, n8405, new_n8974);
nor_5  g06626(new_n8974, new_n8973, new_n8975);
nor_5  g06627(new_n8975, new_n8944, new_n8976);
xnor_4 g06628(n14826, n13549, new_n8977);
xnor_4 g06629(new_n8977, new_n8976, new_n8978);
nor_5  g06630(new_n8978, n18105, new_n8979);
xnor_4 g06631(new_n8978, n18105, new_n8980);
xnor_4 g06632(new_n8974, new_n8973, new_n8981);
nor_5  g06633(new_n8981, n24196, new_n8982_1);
xnor_4 g06634(new_n8981, n24196, new_n8983);
xnor_4 g06635(new_n8971_1, new_n8970, new_n8984);
nor_5  g06636(new_n8984, n16376, new_n8985);
xnor_4 g06637(new_n8984, n16376, new_n8986);
xnor_4 g06638(new_n8968, new_n8967, new_n8987);
nor_5  g06639(new_n8987, n25381, new_n8988);
xnor_4 g06640(new_n8987, n25381, new_n8989);
xnor_4 g06641(new_n8965, new_n8964_1, new_n8990);
nor_5  g06642(new_n8990, n12587, new_n8991);
xnor_4 g06643(new_n8990, n12587, new_n8992);
xnor_4 g06644(new_n8962, new_n8949, new_n8993_1);
nor_5  g06645(new_n8993_1, n268, new_n8994);
xnor_4 g06646(new_n8993_1, n268, new_n8995);
xnor_4 g06647(n6427, n1682, new_n8996);
xnor_4 g06648(new_n8996, new_n8960, new_n8997);
nor_5  g06649(new_n8997, n24879, new_n8998);
xnor_4 g06650(new_n8997, n24879, new_n8999);
xnor_4 g06651(n7963, n6590, new_n9000);
xnor_4 g06652(new_n9000, new_n8957, new_n9001);
nor_5  g06653(new_n9001, n6785, new_n9002);
xnor_4 g06654(n20349, n10017, new_n9003_1);
xnor_4 g06655(new_n9003_1, new_n8954, new_n9004);
nor_5  g06656(new_n9004, n24032, new_n9005);
xnor_4 g06657(n15936, n3618, new_n9006);
or_5   g06658(new_n9006, new_n7324, new_n9007);
xor_4  g06659(new_n9004, n24032, new_n9008);
and_5  g06660(new_n9008, new_n9007, new_n9009);
nor_5  g06661(new_n9009, new_n9005, new_n9010);
xnor_4 g06662(new_n9001, n6785, new_n9011);
nor_5  g06663(new_n9011, new_n9010, new_n9012_1);
nor_5  g06664(new_n9012_1, new_n9002, new_n9013);
nor_5  g06665(new_n9013, new_n8999, new_n9014);
nor_5  g06666(new_n9014, new_n8998, new_n9015);
nor_5  g06667(new_n9015, new_n8995, new_n9016);
nor_5  g06668(new_n9016, new_n8994, new_n9017);
nor_5  g06669(new_n9017, new_n8992, new_n9018);
nor_5  g06670(new_n9018, new_n8991, new_n9019);
nor_5  g06671(new_n9019, new_n8989, new_n9020);
nor_5  g06672(new_n9020, new_n8988, new_n9021);
nor_5  g06673(new_n9021, new_n8986, new_n9022);
nor_5  g06674(new_n9022, new_n8985, new_n9023);
nor_5  g06675(new_n9023, new_n8983, new_n9024);
nor_5  g06676(new_n9024, new_n8982_1, new_n9025);
nor_5  g06677(new_n9025, new_n8980, new_n9026);
nor_5  g06678(new_n9026, new_n8979, new_n9027);
nor_5  g06679(new_n8977, new_n8976, new_n9028);
nor_5  g06680(n14826, n13549, new_n9029);
nor_5  g06681(new_n9029, new_n9028, new_n9030);
nand_5 g06682(new_n9030, new_n9027, new_n9031);
xnor_4 g06683(new_n9031, new_n8943_1, new_n9032_1);
xnor_4 g06684(new_n8942, new_n8939, new_n9033);
xor_4  g06685(new_n9030, new_n9027, new_n9034);
and_5  g06686(new_n9034, new_n9033, new_n9035);
xnor_4 g06687(new_n9034, new_n9033, new_n9036);
xnor_4 g06688(new_n8937, new_n8895, new_n9037);
xor_4  g06689(new_n9025, new_n8980, new_n9038);
nor_5  g06690(new_n9038, new_n9037, new_n9039);
xnor_4 g06691(new_n9038, new_n9037, new_n9040);
xnor_4 g06692(new_n8935, new_n8898, new_n9041);
xor_4  g06693(new_n9023, new_n8983, new_n9042_1);
nor_5  g06694(new_n9042_1, new_n9041, new_n9043);
xnor_4 g06695(new_n9042_1, new_n9041, new_n9044);
xnor_4 g06696(new_n8933, new_n8901, new_n9045);
xor_4  g06697(new_n9021, new_n8986, new_n9046_1);
nor_5  g06698(new_n9046_1, new_n9045, new_n9047_1);
xnor_4 g06699(new_n9046_1, new_n9045, new_n9048);
xnor_4 g06700(new_n8931, new_n8904, new_n9049);
xor_4  g06701(new_n9019, new_n8989, new_n9050);
nor_5  g06702(new_n9050, new_n9049, new_n9051);
xnor_4 g06703(new_n9050, new_n9049, new_n9052);
xnor_4 g06704(new_n8929, new_n8907, new_n9053);
xor_4  g06705(new_n9017, new_n8992, new_n9054);
nor_5  g06706(new_n9054, new_n9053, new_n9055);
xnor_4 g06707(new_n9054, new_n9053, new_n9056);
xnor_4 g06708(new_n8927, new_n8910, new_n9057);
xor_4  g06709(new_n9015, new_n8995, new_n9058);
nor_5  g06710(new_n9058, new_n9057, new_n9059);
xnor_4 g06711(new_n9058, new_n9057, new_n9060);
xnor_4 g06712(new_n8925, new_n8913, new_n9061);
xor_4  g06713(new_n9013, new_n8999, new_n9062);
nor_5  g06714(new_n9062, new_n9061, new_n9063);
xnor_4 g06715(new_n9062, new_n9061, new_n9064);
xnor_4 g06716(new_n8923, new_n8922, new_n9065);
xor_4  g06717(new_n9011, new_n9010, new_n9066);
nor_5  g06718(new_n9066, new_n9065, new_n9067);
xnor_4 g06719(new_n9066, new_n9065, new_n9068);
xnor_4 g06720(new_n8920_1, new_n8919, new_n9069);
xor_4  g06721(new_n9008, new_n9007, new_n9070);
nor_5  g06722(new_n9070, new_n9069, new_n9071);
xor_4  g06723(new_n8918, n27134, new_n9072);
xnor_4 g06724(new_n9006, n22843, new_n9073);
not_10 g06725(new_n9073, new_n9074);
nor_5  g06726(new_n9074, new_n9072, new_n9075);
xor_4  g06727(new_n9070, new_n9069, new_n9076);
and_5  g06728(new_n9076, new_n9075, new_n9077);
nor_5  g06729(new_n9077, new_n9071, new_n9078);
nor_5  g06730(new_n9078, new_n9068, new_n9079);
nor_5  g06731(new_n9079, new_n9067, new_n9080);
nor_5  g06732(new_n9080, new_n9064, new_n9081);
nor_5  g06733(new_n9081, new_n9063, new_n9082);
nor_5  g06734(new_n9082, new_n9060, new_n9083);
nor_5  g06735(new_n9083, new_n9059, new_n9084);
nor_5  g06736(new_n9084, new_n9056, new_n9085);
nor_5  g06737(new_n9085, new_n9055, new_n9086);
nor_5  g06738(new_n9086, new_n9052, new_n9087);
nor_5  g06739(new_n9087, new_n9051, new_n9088);
nor_5  g06740(new_n9088, new_n9048, new_n9089);
nor_5  g06741(new_n9089, new_n9047_1, new_n9090_1);
nor_5  g06742(new_n9090_1, new_n9044, new_n9091);
nor_5  g06743(new_n9091, new_n9043, new_n9092);
nor_5  g06744(new_n9092, new_n9040, new_n9093);
nor_5  g06745(new_n9093, new_n9039, new_n9094);
nor_5  g06746(new_n9094, new_n9036, new_n9095);
nor_5  g06747(new_n9095, new_n9035, new_n9096);
xnor_4 g06748(new_n9096, new_n9032_1, n1302);
not_10 g06749(n12507, new_n9098);
nor_5  g06750(n13951, new_n9098, new_n9099);
xor_4  g06751(n13951, n12507, new_n9100);
not_10 g06752(n15077, new_n9101);
nor_5  g06753(n22793, new_n9101, new_n9102);
xor_4  g06754(n22793, n15077, new_n9103);
not_10 g06755(n3710, new_n9104_1);
nor_5  g06756(n8439, new_n9104_1, new_n9105);
xor_4  g06757(n8439, n3710, new_n9106);
not_10 g06758(n26318, new_n9107);
nor_5  g06759(new_n9107, n25523, new_n9108);
xor_4  g06760(n26318, n25523, new_n9109);
not_10 g06761(n26054, new_n9110);
nor_5  g06762(new_n9110, n5579, new_n9111);
xor_4  g06763(n26054, n5579, new_n9112);
not_10 g06764(n19081, new_n9113);
nor_5  g06765(n23430, new_n9113, new_n9114);
xor_4  g06766(n23430, n19081, new_n9115);
not_10 g06767(n8309, new_n9116);
nor_5  g06768(n10411, new_n9116, new_n9117);
xor_4  g06769(n10411, n8309, new_n9118);
not_10 g06770(n16971, new_n9119);
nor_5  g06771(n19144, new_n9119, new_n9120);
not_10 g06772(n19144, new_n9121);
nor_5  g06773(new_n9121, n16971, new_n9122);
not_10 g06774(n11503, new_n9123);
nor_5  g06775(n12593, new_n9123, new_n9124);
or_5   g06776(new_n7968_1, n11503, new_n9125);
not_10 g06777(n18151, new_n9126);
nor_5  g06778(new_n9126, n13714, new_n9127);
and_5  g06779(new_n9127, new_n9125, new_n9128);
nor_5  g06780(new_n9128, new_n9124, new_n9129_1);
nor_5  g06781(new_n9129_1, new_n9122, new_n9130);
or_5   g06782(new_n9130, new_n9120, new_n9131);
nor_5  g06783(new_n9131, new_n9118, new_n9132);
nor_5  g06784(new_n9132, new_n9117, new_n9133);
nor_5  g06785(new_n9133, new_n9115, new_n9134);
nor_5  g06786(new_n9134, new_n9114, new_n9135);
nor_5  g06787(new_n9135, new_n9112, new_n9136);
nor_5  g06788(new_n9136, new_n9111, new_n9137);
nor_5  g06789(new_n9137, new_n9109, new_n9138);
nor_5  g06790(new_n9138, new_n9108, new_n9139);
nor_5  g06791(new_n9139, new_n9106, new_n9140);
nor_5  g06792(new_n9140, new_n9105, new_n9141);
nor_5  g06793(new_n9141, new_n9103, new_n9142);
nor_5  g06794(new_n9142, new_n9102, new_n9143);
nor_5  g06795(new_n9143, new_n9100, new_n9144);
nor_5  g06796(new_n9144, new_n9099, new_n9145);
nor_5  g06797(n12650, n11220, new_n9146_1);
xnor_4 g06798(n12650, n11220, new_n9147);
nor_5  g06799(n22379, n10201, new_n9148);
xnor_4 g06800(n22379, n10201, new_n9149);
nor_5  g06801(n10593, n1662, new_n9150);
xnor_4 g06802(n10593, n1662, new_n9151);
nor_5  g06803(n18290, n12875, new_n9152);
nor_5  g06804(new_n8436, new_n8415, new_n9153);
nor_5  g06805(new_n9153, new_n9152, new_n9154);
nor_5  g06806(new_n9154, new_n9151, new_n9155);
nor_5  g06807(new_n9155, new_n9150, new_n9156);
nor_5  g06808(new_n9156, new_n9149, new_n9157);
nor_5  g06809(new_n9157, new_n9148, new_n9158);
nor_5  g06810(new_n9158, new_n9147, new_n9159);
nor_5  g06811(new_n9159, new_n9146_1, new_n9160);
nor_5  g06812(n22270, n2944, new_n9161);
nor_5  g06813(new_n2656, new_n2623, new_n9162);
nor_5  g06814(new_n9162, new_n9161, new_n9163);
xor_4  g06815(new_n9163, new_n9160, new_n9164_1);
not_10 g06816(new_n2657, new_n9165);
xor_4  g06817(new_n9158, new_n9147, new_n9166_1);
nor_5  g06818(new_n9166_1, new_n9165, new_n9167);
xnor_4 g06819(new_n9156, new_n9149, new_n9168);
nor_5  g06820(new_n9168, new_n2660, new_n9169);
xnor_4 g06821(new_n9168, new_n2660, new_n9170);
xnor_4 g06822(new_n9154, new_n9151, new_n9171);
nor_5  g06823(new_n9171, new_n2665, new_n9172_1);
xnor_4 g06824(new_n9171, new_n2665, new_n9173);
nor_5  g06825(new_n8437, new_n2669, new_n9174);
nor_5  g06826(new_n8439_1, new_n2673, new_n9175);
xor_4  g06827(new_n8439_1, new_n2673, new_n9176);
not_10 g06828(new_n2677, new_n9177);
nor_5  g06829(new_n8442, new_n9177, new_n9178);
nor_5  g06830(new_n8445, new_n2680_1, new_n9179);
xnor_4 g06831(new_n8445, new_n2680_1, new_n9180);
nor_5  g06832(new_n8448, new_n2684, new_n9181);
xnor_4 g06833(new_n8448, new_n2684, new_n9182_1);
nor_5  g06834(new_n8450, new_n2688, new_n9183);
nor_5  g06835(new_n8452, new_n2690, new_n9184);
xor_4  g06836(new_n8450, new_n2688, new_n9185);
and_5  g06837(new_n9185, new_n9184, new_n9186);
nor_5  g06838(new_n9186, new_n9183, new_n9187);
nor_5  g06839(new_n9187, new_n9182_1, new_n9188);
nor_5  g06840(new_n9188, new_n9181, new_n9189);
nor_5  g06841(new_n9189, new_n9180, new_n9190);
or_5   g06842(new_n9190, new_n9179, new_n9191_1);
xor_4  g06843(new_n8442, new_n2677, new_n9192);
nor_5  g06844(new_n9192, new_n9191_1, new_n9193);
nor_5  g06845(new_n9193, new_n9178, new_n9194);
and_5  g06846(new_n9194, new_n9176, new_n9195);
nor_5  g06847(new_n9195, new_n9175, new_n9196);
xnor_4 g06848(new_n8437, new_n2669, new_n9197);
nor_5  g06849(new_n9197, new_n9196, new_n9198);
nor_5  g06850(new_n9198, new_n9174, new_n9199);
nor_5  g06851(new_n9199, new_n9173, new_n9200);
nor_5  g06852(new_n9200, new_n9172_1, new_n9201);
nor_5  g06853(new_n9201, new_n9170, new_n9202);
or_5   g06854(new_n9202, new_n9169, new_n9203);
xor_4  g06855(new_n9166_1, new_n2657, new_n9204);
nor_5  g06856(new_n9204, new_n9203, new_n9205);
nor_5  g06857(new_n9205, new_n9167, new_n9206);
xor_4  g06858(new_n9206, new_n9164_1, new_n9207);
xnor_4 g06859(new_n9207, new_n9145, new_n9208);
xor_4  g06860(new_n9143, new_n9100, new_n9209);
xor_4  g06861(new_n9204, new_n9203, new_n9210);
nor_5  g06862(new_n9210, new_n9209, new_n9211);
xnor_4 g06863(new_n9210, new_n9209, new_n9212);
xnor_4 g06864(new_n9141, new_n9103, new_n9213);
xor_4  g06865(new_n9201, new_n9170, new_n9214);
and_5  g06866(new_n9214, new_n9213, new_n9215);
xnor_4 g06867(new_n9214, new_n9213, new_n9216);
xnor_4 g06868(new_n9139, new_n9106, new_n9217_1);
xor_4  g06869(new_n9199, new_n9173, new_n9218);
and_5  g06870(new_n9218, new_n9217_1, new_n9219);
xnor_4 g06871(new_n9218, new_n9217_1, new_n9220_1);
xnor_4 g06872(new_n9137, new_n9109, new_n9221);
xor_4  g06873(new_n9197, new_n9196, new_n9222);
and_5  g06874(new_n9222, new_n9221, new_n9223);
xnor_4 g06875(new_n9222, new_n9221, new_n9224);
xnor_4 g06876(new_n9135, new_n9112, new_n9225);
xor_4  g06877(new_n9194, new_n9176, new_n9226);
and_5  g06878(new_n9226, new_n9225, new_n9227);
xor_4  g06879(new_n9133, new_n9115, new_n9228);
xor_4  g06880(new_n9192, new_n9191_1, new_n9229);
nor_5  g06881(new_n9229, new_n9228, new_n9230);
xnor_4 g06882(new_n9229, new_n9228, new_n9231);
xnor_4 g06883(new_n9189, new_n9180, new_n9232);
xor_4  g06884(new_n9131, new_n9118, new_n9233);
nor_5  g06885(new_n9233, new_n9232, new_n9234);
xor_4  g06886(new_n9187, new_n9182_1, new_n9235);
xnor_4 g06887(n19144, n16971, new_n9236);
xnor_4 g06888(new_n9236, new_n9129_1, new_n9237);
and_5  g06889(new_n9237, new_n9235, new_n9238);
xnor_4 g06890(new_n9187, new_n9182_1, new_n9239);
xnor_4 g06891(new_n9237, new_n9239, new_n9240);
xor_4  g06892(new_n8452, new_n2690, new_n9241);
xnor_4 g06893(n18151, n13714, new_n9242);
or_5   g06894(new_n9242, new_n9241, new_n9243);
xor_4  g06895(n12593, n11503, new_n9244);
xnor_4 g06896(new_n9244, new_n9127, new_n9245);
nor_5  g06897(new_n9245, new_n9243, new_n9246_1);
xor_4  g06898(new_n9185, new_n9184, new_n9247);
xnor_4 g06899(new_n9245, new_n9243, new_n9248);
nor_5  g06900(new_n9248, new_n9247, new_n9249);
nor_5  g06901(new_n9249, new_n9246_1, new_n9250);
and_5  g06902(new_n9250, new_n9240, new_n9251_1);
nor_5  g06903(new_n9251_1, new_n9238, new_n9252);
xnor_4 g06904(new_n9233, new_n9232, new_n9253);
nor_5  g06905(new_n9253, new_n9252, new_n9254);
nor_5  g06906(new_n9254, new_n9234, new_n9255);
nor_5  g06907(new_n9255, new_n9231, new_n9256);
nor_5  g06908(new_n9256, new_n9230, new_n9257);
xnor_4 g06909(new_n9226, new_n9225, new_n9258);
nor_5  g06910(new_n9258, new_n9257, new_n9259_1);
nor_5  g06911(new_n9259_1, new_n9227, new_n9260);
nor_5  g06912(new_n9260, new_n9224, new_n9261_1);
nor_5  g06913(new_n9261_1, new_n9223, new_n9262);
nor_5  g06914(new_n9262, new_n9220_1, new_n9263);
nor_5  g06915(new_n9263, new_n9219, new_n9264);
nor_5  g06916(new_n9264, new_n9216, new_n9265);
nor_5  g06917(new_n9265, new_n9215, new_n9266);
nor_5  g06918(new_n9266, new_n9212, new_n9267);
nor_5  g06919(new_n9267, new_n9211, new_n9268);
xnor_4 g06920(new_n9268, new_n9208, n1332);
nor_5  g06921(new_n5118, n14692, new_n9270);
xnor_4 g06922(new_n5118, n14692, new_n9271);
nor_5  g06923(new_n5174, n4100, new_n9272);
xnor_4 g06924(new_n5174, n4100, new_n9273);
nor_5  g06925(new_n5178, n21957, new_n9274);
xnor_4 g06926(new_n5178, n21957, new_n9275);
nor_5  g06927(new_n5182, n15761, new_n9276);
xnor_4 g06928(new_n5182, n15761, new_n9277);
nor_5  g06929(new_n5187, n11201, new_n9278);
xnor_4 g06930(new_n5187, n11201, new_n9279);
nor_5  g06931(new_n5191, n18690, new_n9280);
xnor_4 g06932(new_n5191, n18690, new_n9281);
nor_5  g06933(new_n5196, n12153, new_n9282);
xnor_4 g06934(new_n5196, n12153, new_n9283);
not_10 g06935(n13044, new_n9284);
nor_5  g06936(new_n5202, new_n9284, new_n9285);
and_5  g06937(new_n5202, new_n9284, new_n9286);
not_10 g06938(new_n5207, new_n9287_1);
nor_5  g06939(new_n9287_1, n18745, new_n9288);
xor_4  g06940(new_n5207, n18745, new_n9289);
nor_5  g06941(new_n9289, new_n5339, new_n9290);
or_5   g06942(new_n9290, new_n9288, new_n9291);
nor_5  g06943(new_n9291, new_n9286, new_n9292);
or_5   g06944(new_n9292, new_n9285, new_n9293);
nor_5  g06945(new_n9293, new_n9283, new_n9294);
nor_5  g06946(new_n9294, new_n9282, new_n9295);
nor_5  g06947(new_n9295, new_n9281, new_n9296);
nor_5  g06948(new_n9296, new_n9280, new_n9297);
nor_5  g06949(new_n9297, new_n9279, new_n9298);
nor_5  g06950(new_n9298, new_n9278, new_n9299);
nor_5  g06951(new_n9299, new_n9277, new_n9300);
nor_5  g06952(new_n9300, new_n9276, new_n9301);
nor_5  g06953(new_n9301, new_n9275, new_n9302);
nor_5  g06954(new_n9302, new_n9274, new_n9303);
nor_5  g06955(new_n9303, new_n9273, new_n9304);
nor_5  g06956(new_n9304, new_n9272, new_n9305);
nor_5  g06957(new_n9305, new_n9271, new_n9306);
or_5   g06958(new_n9306, new_n9270, new_n9307);
nor_5  g06959(new_n9307, new_n5117, new_n9308_1);
not_10 g06960(n20151, new_n9309);
not_10 g06961(new_n5348, new_n9310);
or_5   g06962(new_n9310, n11302, new_n9311);
or_5   g06963(new_n9311, n10405, new_n9312);
nor_5  g06964(new_n9312, n7693, new_n9313);
nand_5 g06965(new_n9313, new_n9309, new_n9314);
or_5   g06966(new_n9314, n8964, new_n9315);
nor_5  g06967(new_n9315, n27037, new_n9316);
not_10 g06968(new_n9316, new_n9317);
or_5   g06969(new_n9317, n15182, new_n9318_1);
nor_5  g06970(new_n9318_1, n8614, new_n9319);
or_5   g06971(n25926, n7657, new_n9320);
or_5   g06972(new_n9320, n5330, new_n9321);
or_5   g06973(new_n9321, n5451, new_n9322);
or_5   g06974(new_n9322, n18926, new_n9323_1);
or_5   g06975(new_n9323_1, n13677, new_n9324);
or_5   g06976(new_n9324, n23039, new_n9325);
or_5   g06977(new_n9325, n7692, new_n9326);
or_5   g06978(new_n9326, n25629, new_n9327);
nor_5  g06979(new_n9327, n15766, new_n9328);
xor_4  g06980(new_n9327, n15766, new_n9329);
nor_5  g06981(new_n9329, n23895, new_n9330);
xor_4  g06982(new_n9326, n25629, new_n9331);
nor_5  g06983(new_n9331, n17351, new_n9332);
xnor_4 g06984(new_n9331, n17351, new_n9333);
xor_4  g06985(new_n9325, n7692, new_n9334);
nor_5  g06986(new_n9334, n11736, new_n9335);
xnor_4 g06987(new_n9334, n11736, new_n9336);
xor_4  g06988(new_n9324, n23039, new_n9337);
nor_5  g06989(new_n9337, n23200, new_n9338);
xnor_4 g06990(new_n9337, n23200, new_n9339);
xor_4  g06991(new_n9323_1, n13677, new_n9340);
nor_5  g06992(new_n9340, n17959, new_n9341);
xor_4  g06993(new_n9322, n18926, new_n9342);
nor_5  g06994(new_n9342, n7566, new_n9343);
xor_4  g06995(new_n9342, n7566, new_n9344_1);
xor_4  g06996(new_n9321, n5451, new_n9345);
and_5  g06997(new_n9345, n7731, new_n9346);
nor_5  g06998(new_n9345, n7731, new_n9347);
xor_4  g06999(new_n9320, n5330, new_n9348);
and_5  g07000(new_n9348, n12341, new_n9349);
xnor_4 g07001(new_n9348, n12341, new_n9350);
and_5  g07002(new_n5343, n20986, new_n9351);
and_5  g07003(new_n5344, new_n5342, new_n9352);
nor_5  g07004(new_n9352, new_n9351, new_n9353);
nor_5  g07005(new_n9353, new_n9350, new_n9354);
nor_5  g07006(new_n9354, new_n9349, new_n9355);
nor_5  g07007(new_n9355, new_n9347, new_n9356);
nor_5  g07008(new_n9356, new_n9346, new_n9357);
and_5  g07009(new_n9357, new_n9344_1, new_n9358);
nor_5  g07010(new_n9358, new_n9343, new_n9359);
xnor_4 g07011(new_n9340, n17959, new_n9360);
nor_5  g07012(new_n9360, new_n9359, new_n9361);
nor_5  g07013(new_n9361, new_n9341, new_n9362);
nor_5  g07014(new_n9362, new_n9339, new_n9363);
nor_5  g07015(new_n9363, new_n9338, new_n9364_1);
nor_5  g07016(new_n9364_1, new_n9336, new_n9365);
nor_5  g07017(new_n9365, new_n9335, new_n9366);
nor_5  g07018(new_n9366, new_n9333, new_n9367);
nor_5  g07019(new_n9367, new_n9332, new_n9368);
and_5  g07020(new_n9329, n23895, new_n9369);
nor_5  g07021(new_n9369, new_n9368, new_n9370);
nor_5  g07022(new_n9370, new_n9330, new_n9371_1);
nor_5  g07023(new_n9371_1, new_n9328, new_n9372_1);
or_5   g07024(new_n9372_1, new_n9319, new_n9373);
xnor_4 g07025(new_n9318_1, n8614, new_n9374);
xor_4  g07026(new_n9329, n23895, new_n9375);
xnor_4 g07027(new_n9375, new_n9368, new_n9376);
nor_5  g07028(new_n9376, new_n9374, new_n9377);
xnor_4 g07029(new_n9316, n15182, new_n9378);
xor_4  g07030(new_n9366, new_n9333, new_n9379);
not_10 g07031(new_n9379, new_n9380_1);
nor_5  g07032(new_n9380_1, new_n9378, new_n9381);
xnor_4 g07033(new_n9380_1, new_n9378, new_n9382_1);
xor_4  g07034(new_n9315, n27037, new_n9383);
xor_4  g07035(new_n9364_1, new_n9336, new_n9384);
not_10 g07036(new_n9384, new_n9385);
nor_5  g07037(new_n9385, new_n9383, new_n9386);
xnor_4 g07038(new_n9385, new_n9383, new_n9387);
xor_4  g07039(new_n9314, n8964, new_n9388);
xor_4  g07040(new_n9362, new_n9339, new_n9389);
not_10 g07041(new_n9389, new_n9390);
nor_5  g07042(new_n9390, new_n9388, new_n9391);
xnor_4 g07043(new_n9390, new_n9388, new_n9392);
xnor_4 g07044(new_n9313, new_n9309, new_n9393);
xor_4  g07045(new_n9360, new_n9359, new_n9394);
and_5  g07046(new_n9394, new_n9393, new_n9395);
xnor_4 g07047(new_n9394, new_n9393, new_n9396_1);
xor_4  g07048(new_n9312, n7693, new_n9397);
xor_4  g07049(new_n9357, new_n9344_1, new_n9398);
not_10 g07050(new_n9398, new_n9399_1);
nor_5  g07051(new_n9399_1, new_n9397, new_n9400);
xnor_4 g07052(new_n9399_1, new_n9397, new_n9401);
xor_4  g07053(new_n9311, n10405, new_n9402);
xor_4  g07054(new_n9345, n7731, new_n9403_1);
xnor_4 g07055(new_n9403_1, new_n9355, new_n9404);
nor_5  g07056(new_n9404, new_n9402, new_n9405);
xnor_4 g07057(new_n9404, new_n9402, new_n9406);
xor_4  g07058(new_n9353, new_n9350, new_n9407);
xnor_4 g07059(new_n5348, n11302, new_n9408);
nor_5  g07060(new_n9408, new_n9407, new_n9409);
xnor_4 g07061(new_n9408, new_n9407, new_n9410);
nor_5  g07062(new_n5352, new_n5345, new_n9411);
nor_5  g07063(new_n9411, new_n5351_1, new_n9412);
nor_5  g07064(new_n9412, new_n9410, new_n9413);
nor_5  g07065(new_n9413, new_n9409, new_n9414);
nor_5  g07066(new_n9414, new_n9406, new_n9415);
nor_5  g07067(new_n9415, new_n9405, new_n9416);
nor_5  g07068(new_n9416, new_n9401, new_n9417);
nor_5  g07069(new_n9417, new_n9400, new_n9418);
nor_5  g07070(new_n9418, new_n9396_1, new_n9419_1);
nor_5  g07071(new_n9419_1, new_n9395, new_n9420);
nor_5  g07072(new_n9420, new_n9392, new_n9421);
nor_5  g07073(new_n9421, new_n9391, new_n9422);
nor_5  g07074(new_n9422, new_n9387, new_n9423_1);
nor_5  g07075(new_n9423_1, new_n9386, new_n9424);
nor_5  g07076(new_n9424, new_n9382_1, new_n9425);
nor_5  g07077(new_n9425, new_n9381, new_n9426);
xor_4  g07078(new_n9376, new_n9374, new_n9427);
and_5  g07079(new_n9427, new_n9426, new_n9428);
or_5   g07080(new_n9428, new_n9377, new_n9429);
nor_5  g07081(new_n9429, new_n9373, new_n9430_1);
xnor_4 g07082(new_n9430_1, new_n9308_1, new_n9431);
xor_4  g07083(new_n9307, new_n5117, new_n9432);
xor_4  g07084(new_n9372_1, new_n9319, new_n9433);
xnor_4 g07085(new_n9433, new_n9429, new_n9434);
nor_5  g07086(new_n9434, new_n9432, new_n9435_1);
xor_4  g07087(new_n9434, new_n9432, new_n9436);
xnor_4 g07088(new_n9305, new_n9271, new_n9437);
xor_4  g07089(new_n9427, new_n9426, new_n9438);
and_5  g07090(new_n9438, new_n9437, new_n9439);
xnor_4 g07091(new_n9438, new_n9437, new_n9440);
xor_4  g07092(new_n9424, new_n9382_1, new_n9441);
xor_4  g07093(new_n9303, new_n9273, new_n9442);
nor_5  g07094(new_n9442, new_n9441, new_n9443);
xnor_4 g07095(new_n9422, new_n9387, new_n9444);
xnor_4 g07096(new_n9301, new_n9275, new_n9445_1);
nor_5  g07097(new_n9445_1, new_n9444, new_n9446);
xor_4  g07098(new_n9445_1, new_n9444, new_n9447);
xor_4  g07099(new_n9420, new_n9392, new_n9448);
xor_4  g07100(new_n9299, new_n9277, new_n9449);
nor_5  g07101(new_n9449, new_n9448, new_n9450);
xnor_4 g07102(new_n9418, new_n9396_1, new_n9451_1);
xnor_4 g07103(new_n9297, new_n9279, new_n9452);
nor_5  g07104(new_n9452, new_n9451_1, new_n9453);
xor_4  g07105(new_n9452, new_n9451_1, new_n9454);
xor_4  g07106(new_n9416, new_n9401, new_n9455);
xor_4  g07107(new_n9295, new_n9281, new_n9456);
nor_5  g07108(new_n9456, new_n9455, new_n9457);
xnor_4 g07109(new_n9456, new_n9455, new_n9458_1);
xor_4  g07110(new_n9414, new_n9406, new_n9459_1);
nor_5  g07111(new_n9292, new_n9285, new_n9460_1);
xnor_4 g07112(new_n9460_1, new_n9283, new_n9461);
and_5  g07113(new_n9461, new_n9459_1, new_n9462);
xnor_4 g07114(new_n9461, new_n9459_1, new_n9463);
xnor_4 g07115(new_n9412, new_n9410, new_n9464);
xnor_4 g07116(new_n5202, n13044, new_n9465);
xnor_4 g07117(new_n9465, new_n9291, new_n9466);
nor_5  g07118(new_n9466, new_n9464, new_n9467);
and_5  g07119(new_n5353_1, new_n5341, new_n9468);
and_5  g07120(new_n5354, new_n5337_1, new_n9469);
or_5   g07121(new_n9469, new_n9468, new_n9470);
xor_4  g07122(new_n9466, new_n9464, new_n9471);
and_5  g07123(new_n9471, new_n9470, new_n9472);
nor_5  g07124(new_n9472, new_n9467, new_n9473);
nor_5  g07125(new_n9473, new_n9463, new_n9474);
or_5   g07126(new_n9474, new_n9462, new_n9475);
nor_5  g07127(new_n9475, new_n9458_1, new_n9476);
nor_5  g07128(new_n9476, new_n9457, new_n9477);
and_5  g07129(new_n9477, new_n9454, new_n9478);
or_5   g07130(new_n9478, new_n9453, new_n9479);
xnor_4 g07131(new_n9449, new_n9448, new_n9480);
nor_5  g07132(new_n9480, new_n9479, new_n9481);
nor_5  g07133(new_n9481, new_n9450, new_n9482);
and_5  g07134(new_n9482, new_n9447, new_n9483);
or_5   g07135(new_n9483, new_n9446, new_n9484);
xnor_4 g07136(new_n9442, new_n9441, new_n9485);
nor_5  g07137(new_n9485, new_n9484, new_n9486);
nor_5  g07138(new_n9486, new_n9443, new_n9487);
nor_5  g07139(new_n9487, new_n9440, new_n9488);
nor_5  g07140(new_n9488, new_n9439, new_n9489);
and_5  g07141(new_n9489, new_n9436, new_n9490);
nor_5  g07142(new_n9490, new_n9435_1, new_n9491);
xnor_4 g07143(new_n9491, new_n9431, n1357);
xnor_4 g07144(new_n7247, n25240, new_n9493_1);
nor_5  g07145(new_n7251, n10125, new_n9494);
xnor_4 g07146(new_n7251, n10125, new_n9495);
nor_5  g07147(new_n7255, n8067, new_n9496);
xnor_4 g07148(new_n7255, n8067, new_n9497);
nor_5  g07149(new_n7259, n20923, new_n9498);
xnor_4 g07150(new_n7259, n20923, new_n9499);
nor_5  g07151(new_n7263, n18157, new_n9500);
nor_5  g07152(new_n7683, new_n7674_1, new_n9501);
nor_5  g07153(new_n9501, new_n9500, new_n9502);
nor_5  g07154(new_n9502, new_n9499, new_n9503);
nor_5  g07155(new_n9503, new_n9498, new_n9504);
nor_5  g07156(new_n9504, new_n9497, new_n9505);
nor_5  g07157(new_n9505, new_n9496, new_n9506);
nor_5  g07158(new_n9506, new_n9495, new_n9507_1);
nor_5  g07159(new_n9507_1, new_n9494, new_n9508_1);
xnor_4 g07160(new_n9508_1, new_n9493_1, new_n9509);
xnor_4 g07161(n6381, n1099, new_n9510);
nor_5  g07162(n14345, n2113, new_n9511);
xnor_4 g07163(n14345, n2113, new_n9512_1);
nor_5  g07164(n21134, n11356, new_n9513);
xnor_4 g07165(n21134, n11356, new_n9514);
and_5  g07166(n6369, n3164, new_n9515);
or_5   g07167(n6369, n3164, new_n9516);
nor_5  g07168(n25797, n10611, new_n9517);
nor_5  g07169(new_n5995, new_n5986, new_n9518);
nor_5  g07170(new_n9518, new_n9517, new_n9519);
and_5  g07171(new_n9519, new_n9516, new_n9520);
or_5   g07172(new_n9520, new_n9515, new_n9521);
nor_5  g07173(new_n9521, new_n9514, new_n9522);
nor_5  g07174(new_n9522, new_n9513, new_n9523);
nor_5  g07175(new_n9523, new_n9512_1, new_n9524);
nor_5  g07176(new_n9524, new_n9511, new_n9525);
xnor_4 g07177(new_n9525, new_n9510, new_n9526);
xnor_4 g07178(new_n9526, n5077, new_n9527);
xnor_4 g07179(new_n9523, new_n9512_1, new_n9528);
nand_5 g07180(new_n9528, n15546, new_n9529);
xnor_4 g07181(new_n9528, n15546, new_n9530);
xnor_4 g07182(new_n9521, new_n9514, new_n9531);
nor_5  g07183(new_n9531, n26452, new_n9532);
xnor_4 g07184(n6369, n3164, new_n9533);
xnor_4 g07185(new_n9533, new_n9519, new_n9534);
and_5  g07186(new_n9534, n19905, new_n9535);
xnor_4 g07187(new_n9534, n19905, new_n9536);
and_5  g07188(new_n5996, n17035, new_n9537);
and_5  g07189(new_n7711, new_n7708_1, new_n9538);
nor_5  g07190(new_n9538, new_n9537, new_n9539);
nor_5  g07191(new_n9539, new_n9536, new_n9540);
or_5   g07192(new_n9540, new_n9535, new_n9541);
xnor_4 g07193(new_n9531, n26452, new_n9542);
nor_5  g07194(new_n9542, new_n9541, new_n9543);
nor_5  g07195(new_n9543, new_n9532, new_n9544);
not_10 g07196(new_n9544, new_n9545);
or_5   g07197(new_n9545, new_n9530, new_n9546);
nand_5 g07198(new_n9546, new_n9529, new_n9547);
xor_4  g07199(new_n9547, new_n9527, new_n9548);
xnor_4 g07200(new_n9548, new_n9509, new_n9549);
xor_4  g07201(new_n9506, new_n9495, new_n9550);
xnor_4 g07202(new_n9544, new_n9530, new_n9551);
and_5  g07203(new_n9551, new_n9550, new_n9552_1);
xnor_4 g07204(new_n9551, new_n9550, new_n9553);
xnor_4 g07205(new_n9504, new_n9497, new_n9554_1);
xor_4  g07206(new_n9542, new_n9541, new_n9555);
nor_5  g07207(new_n9555, new_n9554_1, new_n9556_1);
xnor_4 g07208(new_n9555, new_n9554_1, new_n9557_1);
xnor_4 g07209(new_n9502, new_n9499, new_n9558_1);
xor_4  g07210(new_n9539, new_n9536, new_n9559);
not_10 g07211(new_n9559, new_n9560);
nor_5  g07212(new_n9560, new_n9558_1, new_n9561);
xnor_4 g07213(new_n9559, new_n9558_1, new_n9562);
and_5  g07214(new_n7706, new_n7684, new_n9563);
not_10 g07215(new_n7712, new_n9564);
and_5  g07216(new_n9564, new_n7707, new_n9565);
nor_5  g07217(new_n9565, new_n9563, new_n9566);
and_5  g07218(new_n9566, new_n9562, new_n9567);
nor_5  g07219(new_n9567, new_n9561, new_n9568);
nor_5  g07220(new_n9568, new_n9557_1, new_n9569);
nor_5  g07221(new_n9569, new_n9556_1, new_n9570);
nor_5  g07222(new_n9570, new_n9553, new_n9571);
nor_5  g07223(new_n9571, new_n9552_1, new_n9572);
xnor_4 g07224(new_n9572, new_n9549, n1371);
xor_4  g07225(n17250, n15241, new_n9574);
nor_5  g07226(new_n6983_1, n7678, new_n9575);
nor_5  g07227(new_n6986, n3785, new_n9576);
xor_4  g07228(n16524, n3785, new_n9577);
nor_5  g07229(new_n4073, n11056, new_n9578);
nor_5  g07230(n15271, new_n4075, new_n9579);
xor_4  g07231(n15271, n5822, new_n9580);
nor_5  g07232(new_n4080, n25877, new_n9581);
and_5  g07233(new_n5317, new_n5316, new_n9582);
nor_5  g07234(new_n9582, new_n9581, new_n9583);
nor_5  g07235(new_n9583, new_n9580, new_n9584);
nor_5  g07236(new_n9584, new_n9579, new_n9585);
xor_4  g07237(n20250, n11056, new_n9586);
nor_5  g07238(new_n9586, new_n9585, new_n9587);
or_5   g07239(new_n9587, new_n9578, new_n9588);
nor_5  g07240(new_n9588, new_n9577, new_n9589);
nor_5  g07241(new_n9589, new_n9576, new_n9590);
xor_4  g07242(n23160, n7678, new_n9591);
nor_5  g07243(new_n9591, new_n9590, new_n9592);
nor_5  g07244(new_n9592, new_n9575, new_n9593);
xor_4  g07245(new_n9593, new_n9574, new_n9594);
xnor_4 g07246(new_n8753, n13783, new_n9595);
nor_5  g07247(new_n8756, n26660, new_n9596);
xor_4  g07248(new_n8756, n26660, new_n9597);
and_5  g07249(new_n8759, n3018, new_n9598_1);
nor_5  g07250(new_n8759, n3018, new_n9599);
and_5  g07251(new_n8573, n3480, new_n9600);
nor_5  g07252(new_n8581_1, new_n8574, new_n9601);
nor_5  g07253(new_n9601, new_n9600, new_n9602);
nor_5  g07254(new_n9602, new_n9599, new_n9603);
nor_5  g07255(new_n9603, new_n9598_1, new_n9604);
and_5  g07256(new_n9604, new_n9597, new_n9605);
nor_5  g07257(new_n9605, new_n9596, new_n9606);
xor_4  g07258(new_n9606, new_n9595, new_n9607);
xor_4  g07259(new_n9607, new_n9594, new_n9608);
xnor_4 g07260(new_n9604, new_n9597, new_n9609);
xor_4  g07261(new_n9591, new_n9590, new_n9610);
and_5  g07262(new_n9610, new_n9609, new_n9611);
xnor_4 g07263(new_n9610, new_n9609, new_n9612);
xor_4  g07264(new_n9588, new_n9577, new_n9613);
xor_4  g07265(new_n8759, n3018, new_n9614);
xnor_4 g07266(new_n9614, new_n9602, new_n9615);
nor_5  g07267(new_n9615, new_n9613, new_n9616_1);
xnor_4 g07268(new_n9615, new_n9613, new_n9617);
xnor_4 g07269(new_n9586, new_n9585, new_n9618);
nor_5  g07270(new_n9618, new_n8582, new_n9619);
xor_4  g07271(new_n9618, new_n8582, new_n9620);
xor_4  g07272(new_n9583, new_n9580, new_n9621);
nor_5  g07273(new_n9621, new_n8584, new_n9622_1);
xnor_4 g07274(new_n9621, new_n8584, new_n9623);
nor_5  g07275(new_n5318, new_n5315, new_n9624);
nor_5  g07276(new_n5326, new_n5319, new_n9625);
nor_5  g07277(new_n9625, new_n9624, new_n9626_1);
nor_5  g07278(new_n9626_1, new_n9623, new_n9627);
nor_5  g07279(new_n9627, new_n9622_1, new_n9628);
and_5  g07280(new_n9628, new_n9620, new_n9629);
nor_5  g07281(new_n9629, new_n9619, new_n9630);
nor_5  g07282(new_n9630, new_n9617, new_n9631);
or_5   g07283(new_n9631, new_n9616_1, new_n9632);
nor_5  g07284(new_n9632, new_n9612, new_n9633_1);
nor_5  g07285(new_n9633_1, new_n9611, new_n9634);
xnor_4 g07286(new_n9634, new_n9608, new_n9635_1);
xnor_4 g07287(new_n9635_1, new_n5183, new_n9636);
xor_4  g07288(new_n9632, new_n9612, new_n9637);
nor_5  g07289(new_n9637, new_n5187, new_n9638);
xor_4  g07290(new_n9637, new_n5187, new_n9639);
xor_4  g07291(new_n9630, new_n9617, new_n9640);
nor_5  g07292(new_n9640, new_n5192, new_n9641);
xor_4  g07293(new_n9628, new_n9620, new_n9642);
not_10 g07294(new_n9642, new_n9643);
nor_5  g07295(new_n9643, new_n5196, new_n9644);
xnor_4 g07296(new_n9642, new_n5196, new_n9645);
xnor_4 g07297(new_n9626_1, new_n9623, new_n9646_1);
nor_5  g07298(new_n9646_1, new_n5202, new_n9647);
nand_5 g07299(new_n5313, new_n9287_1, new_n9648_1);
not_10 g07300(new_n5327, new_n9649);
or_5   g07301(new_n9649, new_n5314, new_n9650);
and_5  g07302(new_n9650, new_n9648_1, new_n9651);
xnor_4 g07303(new_n9646_1, new_n5202, new_n9652);
nor_5  g07304(new_n9652, new_n9651, new_n9653);
nor_5  g07305(new_n9653, new_n9647, new_n9654);
and_5  g07306(new_n9654, new_n9645, new_n9655_1);
or_5   g07307(new_n9655_1, new_n9644, new_n9656);
xor_4  g07308(new_n9640, new_n5191, new_n9657);
nor_5  g07309(new_n9657, new_n9656, new_n9658);
nor_5  g07310(new_n9658, new_n9641, new_n9659);
and_5  g07311(new_n9659, new_n9639, new_n9660);
or_5   g07312(new_n9660, new_n9638, new_n9661);
xor_4  g07313(new_n9661, new_n9636, n1385);
xor_4  g07314(new_n8309_1, new_n8267_1, new_n9663);
xor_4  g07315(n26808, n24732, new_n9664);
and_5  g07316(n26808, n24732, new_n9665);
xnor_4 g07317(n7339, n6631, new_n9666);
xnor_4 g07318(new_n9666, new_n9665, new_n9667);
nor_5  g07319(new_n9667, new_n9664, new_n9668);
xnor_4 g07320(n14684, n1667, new_n9669);
nor_5  g07321(n7339, n6631, new_n9670);
nor_5  g07322(new_n9666, new_n9665, new_n9671);
nor_5  g07323(new_n9671, new_n9670, new_n9672);
xor_4  g07324(new_n9672, new_n9669, new_n9673);
nand_5 g07325(new_n9673, new_n9668, new_n9674);
xnor_4 g07326(n17035, n2680, new_n9675);
nor_5  g07327(n14684, n1667, new_n9676);
nor_5  g07328(new_n9672, new_n9669, new_n9677);
nor_5  g07329(new_n9677, new_n9676, new_n9678);
xor_4  g07330(new_n9678, new_n9675, new_n9679);
not_10 g07331(new_n9679, new_n9680);
or_5   g07332(new_n9680, new_n9674, new_n9681);
xnor_4 g07333(n19905, n2547, new_n9682);
nor_5  g07334(n17035, n2680, new_n9683);
nor_5  g07335(new_n9678, new_n9675, new_n9684);
nor_5  g07336(new_n9684, new_n9683, new_n9685);
xor_4  g07337(new_n9685, new_n9682, new_n9686);
not_10 g07338(new_n9686, new_n9687);
or_5   g07339(new_n9687, new_n9681, new_n9688);
xnor_4 g07340(n26452, n2999, new_n9689_1);
nor_5  g07341(n19905, n2547, new_n9690);
nor_5  g07342(new_n9685, new_n9682, new_n9691);
nor_5  g07343(new_n9691, new_n9690, new_n9692);
xor_4  g07344(new_n9692, new_n9689_1, new_n9693);
not_10 g07345(new_n9693, new_n9694);
or_5   g07346(new_n9694, new_n9688, new_n9695_1);
xnor_4 g07347(n15546, n14702, new_n9696);
nor_5  g07348(n26452, n2999, new_n9697);
nor_5  g07349(new_n9692, new_n9689_1, new_n9698);
nor_5  g07350(new_n9698, new_n9697, new_n9699_1);
xor_4  g07351(new_n9699_1, new_n9696, new_n9700);
not_10 g07352(new_n9700, new_n9701);
or_5   g07353(new_n9701, new_n9695_1, new_n9702);
xnor_4 g07354(n13914, n5077, new_n9703);
nor_5  g07355(n15546, n14702, new_n9704);
nor_5  g07356(new_n9699_1, new_n9696, new_n9705);
nor_5  g07357(new_n9705, new_n9704, new_n9706);
xor_4  g07358(new_n9706, new_n9703, new_n9707);
not_10 g07359(new_n9707, new_n9708);
or_5   g07360(new_n9708, new_n9702, new_n9709);
xnor_4 g07361(n18035, n3279, new_n9710);
nor_5  g07362(n13914, n5077, new_n9711);
nor_5  g07363(new_n9706, new_n9703, new_n9712);
nor_5  g07364(new_n9712, new_n9711, new_n9713);
xor_4  g07365(new_n9713, new_n9710, new_n9714);
not_10 g07366(new_n9714, new_n9715);
or_5   g07367(new_n9715, new_n9709, new_n9716);
xnor_4 g07368(n8827, n4306, new_n9717);
nor_5  g07369(n18035, n3279, new_n9718);
nor_5  g07370(new_n9713, new_n9710, new_n9719);
nor_5  g07371(new_n9719, new_n9718, new_n9720);
xor_4  g07372(new_n9720, new_n9717, new_n9721);
xnor_4 g07373(new_n9721, new_n9716, new_n9722);
xnor_4 g07374(new_n9722, new_n7239, new_n9723);
xnor_4 g07375(new_n9714, new_n9709, new_n9724);
nor_5  g07376(new_n9724, new_n7243, new_n9725);
xnor_4 g07377(new_n9724, new_n7243, new_n9726_1);
xnor_4 g07378(new_n9707, new_n9702, new_n9727);
nor_5  g07379(new_n9727, new_n7247, new_n9728);
xnor_4 g07380(new_n9727, new_n7247, new_n9729);
xnor_4 g07381(new_n9700, new_n9695_1, new_n9730);
nor_5  g07382(new_n9730, new_n7251, new_n9731);
xnor_4 g07383(new_n9730, new_n7251, new_n9732);
xnor_4 g07384(new_n9693, new_n9688, new_n9733);
nor_5  g07385(new_n9733, new_n7255, new_n9734);
xnor_4 g07386(new_n9733, new_n7255, new_n9735);
xnor_4 g07387(new_n9686, new_n9681, new_n9736);
nor_5  g07388(new_n9736, new_n7259, new_n9737);
xnor_4 g07389(new_n9736, new_n7259, new_n9738);
xnor_4 g07390(new_n9679, new_n9674, new_n9739);
nor_5  g07391(new_n9739, new_n7263, new_n9740);
xnor_4 g07392(new_n9739, new_n7263, new_n9741);
xor_4  g07393(new_n9673, new_n9668, new_n9742);
nor_5  g07394(new_n9742, new_n7267, new_n9743);
xnor_4 g07395(new_n9742, new_n7267, new_n9744);
not_10 g07396(new_n9664, new_n9745);
or_5   g07397(new_n9745, new_n2523, new_n9746);
and_5  g07398(new_n9746, new_n7273, new_n9747);
nor_5  g07399(new_n9666, new_n9745, new_n9748);
or_5   g07400(new_n9748, new_n9668, new_n9749);
nor_5  g07401(new_n9746, new_n7222, new_n9750);
nor_5  g07402(new_n9750, new_n9747, new_n9751);
and_5  g07403(new_n9751, new_n9749, new_n9752);
nor_5  g07404(new_n9752, new_n9747, new_n9753_1);
nor_5  g07405(new_n9753_1, new_n9744, new_n9754);
nor_5  g07406(new_n9754, new_n9743, new_n9755);
nor_5  g07407(new_n9755, new_n9741, new_n9756);
nor_5  g07408(new_n9756, new_n9740, new_n9757);
nor_5  g07409(new_n9757, new_n9738, new_n9758);
nor_5  g07410(new_n9758, new_n9737, new_n9759);
nor_5  g07411(new_n9759, new_n9735, new_n9760);
nor_5  g07412(new_n9760, new_n9734, new_n9761_1);
nor_5  g07413(new_n9761_1, new_n9732, new_n9762);
nor_5  g07414(new_n9762, new_n9731, new_n9763_1);
nor_5  g07415(new_n9763_1, new_n9729, new_n9764);
nor_5  g07416(new_n9764, new_n9728, new_n9765);
nor_5  g07417(new_n9765, new_n9726_1, new_n9766);
nor_5  g07418(new_n9766, new_n9725, new_n9767_1);
xor_4  g07419(new_n9767_1, new_n9723, new_n9768);
xnor_4 g07420(new_n9768, new_n9663, new_n9769);
xor_4  g07421(new_n9765, new_n9726_1, new_n9770);
and_5  g07422(new_n9770, new_n8313, new_n9771_1);
xnor_4 g07423(new_n9770, new_n8313, new_n9772);
xor_4  g07424(new_n9763_1, new_n9729, new_n9773);
and_5  g07425(new_n9773, new_n8317, new_n9774);
xnor_4 g07426(new_n9773, new_n8317, new_n9775);
xor_4  g07427(new_n9761_1, new_n9732, new_n9776);
and_5  g07428(new_n9776, new_n8321_1, new_n9777);
xnor_4 g07429(new_n9776, new_n8321_1, new_n9778_1);
xor_4  g07430(new_n9759, new_n9735, new_n9779);
and_5  g07431(new_n9779, new_n8325, new_n9780);
xnor_4 g07432(new_n9779, new_n8325, new_n9781);
xor_4  g07433(new_n9757, new_n9738, new_n9782);
and_5  g07434(new_n9782, new_n8328, new_n9783_1);
xnor_4 g07435(new_n9782, new_n8328, new_n9784);
xor_4  g07436(new_n9755, new_n9741, new_n9785);
and_5  g07437(new_n9785, new_n8332, new_n9786);
not_10 g07438(new_n8336, new_n9787);
xor_4  g07439(new_n9753_1, new_n9744, new_n9788);
and_5  g07440(new_n9788, new_n9787, new_n9789);
xnor_4 g07441(new_n9788, new_n9787, new_n9790);
xnor_4 g07442(new_n9664, new_n2523, new_n9791);
or_5   g07443(new_n9791, new_n8344, new_n9792);
nor_5  g07444(new_n9792, new_n8341, new_n9793);
xor_4  g07445(new_n9792, new_n8341, new_n9794);
xor_4  g07446(new_n9751, new_n9749, new_n9795);
and_5  g07447(new_n9795, new_n9794, new_n9796);
nor_5  g07448(new_n9796, new_n9793, new_n9797);
nor_5  g07449(new_n9797, new_n9790, new_n9798);
nor_5  g07450(new_n9798, new_n9789, new_n9799);
xnor_4 g07451(new_n9785, new_n8332, new_n9800);
nor_5  g07452(new_n9800, new_n9799, new_n9801);
nor_5  g07453(new_n9801, new_n9786, new_n9802);
nor_5  g07454(new_n9802, new_n9784, new_n9803_1);
nor_5  g07455(new_n9803_1, new_n9783_1, new_n9804);
nor_5  g07456(new_n9804, new_n9781, new_n9805);
nor_5  g07457(new_n9805, new_n9780, new_n9806);
nor_5  g07458(new_n9806, new_n9778_1, new_n9807);
nor_5  g07459(new_n9807, new_n9777, new_n9808);
nor_5  g07460(new_n9808, new_n9775, new_n9809);
nor_5  g07461(new_n9809, new_n9774, new_n9810);
nor_5  g07462(new_n9810, new_n9772, new_n9811);
nor_5  g07463(new_n9811, new_n9771_1, new_n9812);
xnor_4 g07464(new_n9812, new_n9769, n1498);
xor_4  g07465(n20658, n9090, new_n9814);
xnor_4 g07466(new_n9814, new_n5465, new_n9815);
xor_4  g07467(new_n9815, new_n4626, n1501);
or_5   g07468(n15506, n11473, new_n9817);
nor_5  g07469(new_n9817, n5131, new_n9818);
not_10 g07470(new_n9818, new_n9819);
or_5   g07471(new_n9819, n21538, new_n9820);
or_5   g07472(new_n9820, n25094, new_n9821);
nor_5  g07473(new_n9821, n1611, new_n9822);
xnor_4 g07474(new_n9822, n752, new_n9823);
xnor_4 g07475(new_n9823, new_n8792, new_n9824);
xnor_4 g07476(new_n8734, new_n8716_1, new_n9825);
xor_4  g07477(new_n9821, n1611, new_n9826);
nor_5  g07478(new_n9826, new_n9825, new_n9827);
xor_4  g07479(new_n9826, new_n8794, new_n9828);
xnor_4 g07480(new_n9820, n25094, new_n9829);
and_5  g07481(new_n9829, new_n8798, new_n9830);
xor_4  g07482(new_n9820, n25094, new_n9831);
xnor_4 g07483(new_n9831, new_n8798, new_n9832_1);
xnor_4 g07484(new_n9818, n21538, new_n9833_1);
not_10 g07485(new_n9833_1, new_n9834);
nor_5  g07486(new_n9834, new_n8803_1, new_n9835);
xor_4  g07487(new_n9817, n5131, new_n9836);
nor_5  g07488(new_n9836, new_n8807, new_n9837);
xnor_4 g07489(new_n9836, new_n8807, new_n9838_1);
nand_5 g07490(new_n8814, n15506, new_n9839);
xnor_4 g07491(n15506, n11473, new_n9840);
and_5  g07492(new_n9840, new_n9839, new_n9841);
nor_5  g07493(new_n9839, n11473, new_n9842);
nor_5  g07494(new_n9842, new_n9841, new_n9843);
and_5  g07495(new_n9843, new_n8811, new_n9844);
nor_5  g07496(new_n9844, new_n9841, new_n9845);
nor_5  g07497(new_n9845, new_n9838_1, new_n9846);
or_5   g07498(new_n9846, new_n9837, new_n9847);
xnor_4 g07499(new_n9834, new_n8803_1, new_n9848);
nor_5  g07500(new_n9848, new_n9847, new_n9849);
nor_5  g07501(new_n9849, new_n9835, new_n9850);
and_5  g07502(new_n9850, new_n9832_1, new_n9851);
nor_5  g07503(new_n9851, new_n9830, new_n9852);
nor_5  g07504(new_n9852, new_n9828, new_n9853);
or_5   g07505(new_n9853, new_n9827, new_n9854);
xor_4  g07506(new_n9854, new_n9824, new_n9855);
xnor_4 g07507(n20470, n3366, new_n9856);
and_5  g07508(n26565, n21222, new_n9857);
or_5   g07509(n26565, n21222, new_n9858);
nor_5  g07510(n9832, n3959, new_n9859);
nor_5  g07511(new_n8646, new_n8633, new_n9860);
nor_5  g07512(new_n9860, new_n9859, new_n9861);
and_5  g07513(new_n9861, new_n9858, new_n9862);
or_5   g07514(new_n9862, new_n9857, new_n9863);
xor_4  g07515(new_n9863, new_n9856, new_n9864);
xnor_4 g07516(new_n9864, new_n9855, new_n9865);
xor_4  g07517(new_n9852, new_n9828, new_n9866);
xnor_4 g07518(n26565, n21222, new_n9867_1);
xnor_4 g07519(new_n9867_1, new_n9861, new_n9868);
and_5  g07520(new_n9868, new_n9866, new_n9869);
xnor_4 g07521(new_n9868, new_n9866, new_n9870);
xor_4  g07522(new_n9850, new_n9832_1, new_n9871);
and_5  g07523(new_n9871, new_n8647, new_n9872_1);
xnor_4 g07524(new_n9871, new_n8647, new_n9873);
xor_4  g07525(new_n9848, new_n9847, new_n9874);
nor_5  g07526(new_n9874, new_n8691, new_n9875);
xor_4  g07527(new_n9874, new_n8691, new_n9876);
not_10 g07528(new_n8695, new_n9877);
xor_4  g07529(new_n9845, new_n9838_1, new_n9878);
nor_5  g07530(new_n9878, new_n9877, new_n9879);
xnor_4 g07531(new_n9843, new_n8811, new_n9880);
nor_5  g07532(new_n9880, new_n8700, new_n9881);
xor_4  g07533(new_n8814, n15506, new_n9882);
nor_5  g07534(new_n9882, new_n6522, new_n9883);
xor_4  g07535(new_n9880, new_n8700, new_n9884);
and_5  g07536(new_n9884, new_n9883, new_n9885);
or_5   g07537(new_n9885, new_n9881, new_n9886);
xnor_4 g07538(new_n9878, new_n9877, new_n9887);
nor_5  g07539(new_n9887, new_n9886, new_n9888);
nor_5  g07540(new_n9888, new_n9879, new_n9889);
and_5  g07541(new_n9889, new_n9876, new_n9890_1);
nor_5  g07542(new_n9890_1, new_n9875, new_n9891);
nor_5  g07543(new_n9891, new_n9873, new_n9892);
nor_5  g07544(new_n9892, new_n9872_1, new_n9893);
nor_5  g07545(new_n9893, new_n9870, new_n9894);
nor_5  g07546(new_n9894, new_n9869, new_n9895);
xnor_4 g07547(new_n9895, new_n9865, n1518);
nor_5  g07548(new_n6526, n14826, new_n9897);
xor_4  g07549(n17458, n14826, new_n9898);
nor_5  g07550(n23493, new_n6529, new_n9899);
xor_4  g07551(n23493, n1222, new_n9900);
nor_5  g07552(new_n6532, n10275, new_n9901);
xor_4  g07553(n25240, n10275, new_n9902);
nor_5  g07554(n15146, new_n6535, new_n9903);
xor_4  g07555(n15146, n10125, new_n9904);
nor_5  g07556(n11579, new_n6538, new_n9905);
xor_4  g07557(n11579, n8067, new_n9906);
nor_5  g07558(new_n6541, n21, new_n9907);
xor_4  g07559(n20923, n21, new_n9908);
nor_5  g07560(new_n6544, n1682, new_n9909);
xor_4  g07561(n18157, n1682, new_n9910);
not_10 g07562(n7963, new_n9911);
nor_5  g07563(n12161, new_n9911, new_n9912);
nor_5  g07564(new_n6547, n7963, new_n9913);
not_10 g07565(n10017, new_n9914);
nor_5  g07566(new_n9914, n5026, new_n9915);
or_5   g07567(n10017, new_n6550, new_n9916);
not_10 g07568(n3618, new_n9917_1);
nor_5  g07569(n8581, new_n9917_1, new_n9918);
and_5  g07570(new_n9918, new_n9916, new_n9919_1);
nor_5  g07571(new_n9919_1, new_n9915, new_n9920);
nor_5  g07572(new_n9920, new_n9913, new_n9921);
or_5   g07573(new_n9921, new_n9912, new_n9922);
nor_5  g07574(new_n9922, new_n9910, new_n9923);
nor_5  g07575(new_n9923, new_n9909, new_n9924);
nor_5  g07576(new_n9924, new_n9908, new_n9925);
nor_5  g07577(new_n9925, new_n9907, new_n9926_1);
nor_5  g07578(new_n9926_1, new_n9906, new_n9927);
nor_5  g07579(new_n9927, new_n9905, new_n9928);
nor_5  g07580(new_n9928, new_n9904, new_n9929);
nor_5  g07581(new_n9929, new_n9903, new_n9930);
nor_5  g07582(new_n9930, new_n9902, new_n9931);
nor_5  g07583(new_n9931, new_n9901, new_n9932);
nor_5  g07584(new_n9932, new_n9900, new_n9933);
nor_5  g07585(new_n9933, new_n9899, new_n9934_1);
nor_5  g07586(new_n9934_1, new_n9898, new_n9935);
nor_5  g07587(new_n9935, new_n9897, new_n9936);
or_5   g07588(new_n3915, n3468, new_n9937);
or_5   g07589(new_n9937, n12821, new_n9938_1);
or_5   g07590(new_n9938_1, n22492, new_n9939);
or_5   g07591(new_n9939, n7330, new_n9940);
or_5   g07592(new_n9940, n767, new_n9941);
xor_4  g07593(new_n9941, n2944, new_n9942_1);
and_5  g07594(new_n9942_1, n19282, new_n9943);
nor_5  g07595(new_n9941, n2944, new_n9944);
xor_4  g07596(new_n9940, n767, new_n9945);
nor_5  g07597(new_n9945, n12657, new_n9946_1);
xnor_4 g07598(new_n9945, n12657, new_n9947);
xor_4  g07599(new_n9939, n7330, new_n9948);
and_5  g07600(new_n9948, n17077, new_n9949);
xnor_4 g07601(new_n9948, n17077, new_n9950);
xor_4  g07602(new_n9938_1, n22492, new_n9951);
and_5  g07603(new_n9951, n26510, new_n9952);
xnor_4 g07604(new_n9951, n26510, new_n9953);
xor_4  g07605(new_n9937, n12821, new_n9954);
and_5  g07606(new_n9954, n23068, new_n9955);
nor_5  g07607(new_n9954, n23068, new_n9956);
and_5  g07608(new_n3916, n19514, new_n9957);
nor_5  g07609(new_n3933, new_n3917, new_n9958);
nor_5  g07610(new_n9958, new_n9957, new_n9959);
nor_5  g07611(new_n9959, new_n9956, new_n9960);
nor_5  g07612(new_n9960, new_n9955, new_n9961);
nor_5  g07613(new_n9961, new_n9953, new_n9962);
nor_5  g07614(new_n9962, new_n9952, new_n9963);
nor_5  g07615(new_n9963, new_n9950, new_n9964);
or_5   g07616(new_n9964, new_n9949, new_n9965);
nor_5  g07617(new_n9965, new_n9947, new_n9966);
nor_5  g07618(new_n9966, new_n9946_1, new_n9967_1);
or_5   g07619(new_n9942_1, n19282, new_n9968_1);
and_5  g07620(new_n9968_1, new_n9967_1, new_n9969);
or_5   g07621(new_n9969, new_n9944, new_n9970);
nor_5  g07622(new_n9970, new_n9943, new_n9971);
nor_5  g07623(new_n9971, new_n9936, new_n9972);
xor_4  g07624(new_n9934_1, new_n9898, new_n9973);
xnor_4 g07625(new_n9942_1, n19282, new_n9974);
xnor_4 g07626(new_n9974, new_n9967_1, new_n9975);
nor_5  g07627(new_n9975, new_n9973, new_n9976);
xnor_4 g07628(new_n9975, new_n9973, new_n9977);
xor_4  g07629(new_n9932, new_n9900, new_n9978);
xnor_4 g07630(new_n9965, new_n9947, new_n9979);
nor_5  g07631(new_n9979, new_n9978, new_n9980);
xnor_4 g07632(new_n9979, new_n9978, new_n9981);
xor_4  g07633(new_n9930, new_n9902, new_n9982);
xor_4  g07634(new_n9963, new_n9950, new_n9983);
nor_5  g07635(new_n9983, new_n9982, new_n9984);
xnor_4 g07636(new_n9983, new_n9982, new_n9985);
xor_4  g07637(new_n9928, new_n9904, new_n9986);
xor_4  g07638(new_n9961, new_n9953, new_n9987);
nor_5  g07639(new_n9987, new_n9986, new_n9988);
xnor_4 g07640(new_n9987, new_n9986, new_n9989);
xor_4  g07641(new_n9926_1, new_n9906, new_n9990);
xor_4  g07642(new_n9954, n23068, new_n9991);
xnor_4 g07643(new_n9991, new_n9959, new_n9992);
nor_5  g07644(new_n9992, new_n9990, new_n9993);
xnor_4 g07645(new_n9992, new_n9990, new_n9994);
xor_4  g07646(new_n9924, new_n9908, new_n9995);
nor_5  g07647(new_n9995, new_n3934_1, new_n9996);
xor_4  g07648(new_n9922, new_n9910, new_n9997);
nor_5  g07649(new_n9997, new_n3958, new_n9998);
xnor_4 g07650(new_n9997, new_n3958, new_n9999);
not_10 g07651(new_n3974, new_n10000);
xnor_4 g07652(n12161, n7963, new_n10001);
xnor_4 g07653(new_n10001, new_n9920, new_n10002);
and_5  g07654(new_n10002, new_n10000, new_n10003);
xnor_4 g07655(new_n10002, new_n10000, new_n10004);
xnor_4 g07656(n8581, n3618, new_n10005);
nor_5  g07657(new_n10005, new_n3968, new_n10006);
xor_4  g07658(n10017, n5026, new_n10007);
xnor_4 g07659(new_n10007, new_n9918, new_n10008);
not_10 g07660(new_n10008, new_n10009_1);
nor_5  g07661(new_n10009_1, new_n10006, new_n10010_1);
xnor_4 g07662(new_n10008, new_n10006, new_n10011);
and_5  g07663(new_n10011, new_n3964, new_n10012);
nor_5  g07664(new_n10012, new_n10010_1, new_n10013);
nor_5  g07665(new_n10013, new_n10004, new_n10014);
nor_5  g07666(new_n10014, new_n10003, new_n10015);
nor_5  g07667(new_n10015, new_n9999, new_n10016);
nor_5  g07668(new_n10016, new_n9998, new_n10017_1);
xnor_4 g07669(new_n9995, new_n3934_1, new_n10018_1);
nor_5  g07670(new_n10018_1, new_n10017_1, new_n10019_1);
nor_5  g07671(new_n10019_1, new_n9996, new_n10020);
nor_5  g07672(new_n10020, new_n9994, new_n10021_1);
nor_5  g07673(new_n10021_1, new_n9993, new_n10022);
nor_5  g07674(new_n10022, new_n9989, new_n10023);
nor_5  g07675(new_n10023, new_n9988, new_n10024);
nor_5  g07676(new_n10024, new_n9985, new_n10025);
nor_5  g07677(new_n10025, new_n9984, new_n10026);
nor_5  g07678(new_n10026, new_n9981, new_n10027);
nor_5  g07679(new_n10027, new_n9980, new_n10028);
nor_5  g07680(new_n10028, new_n9977, new_n10029);
or_5   g07681(new_n10029, new_n9976, new_n10030);
xnor_4 g07682(new_n9971, new_n9936, new_n10031);
nor_5  g07683(new_n10031, new_n10030, new_n10032);
nor_5  g07684(new_n10032, new_n9972, new_n10033);
nor_5  g07685(n20040, new_n6744, new_n10034);
nor_5  g07686(new_n7936, new_n7901, new_n10035);
nor_5  g07687(new_n10035, new_n10034, new_n10036);
xnor_4 g07688(new_n10036, new_n10033, new_n10037);
xor_4  g07689(new_n10031, new_n10030, new_n10038);
nor_5  g07690(new_n10038, new_n10036, new_n10039);
xnor_4 g07691(new_n10028, new_n9977, new_n10040);
nor_5  g07692(new_n10040, new_n7937_1, new_n10041);
xnor_4 g07693(new_n10040, new_n7937_1, new_n10042);
xnor_4 g07694(new_n10026, new_n9981, new_n10043);
nor_5  g07695(new_n10043, new_n7992_1, new_n10044);
xnor_4 g07696(new_n10043, new_n7992_1, new_n10045);
xnor_4 g07697(new_n10024, new_n9985, new_n10046);
nor_5  g07698(new_n10046, new_n7997, new_n10047);
xnor_4 g07699(new_n10046, new_n7997, new_n10048);
xnor_4 g07700(new_n10022, new_n9989, new_n10049);
nor_5  g07701(new_n10049, new_n8002, new_n10050);
xnor_4 g07702(new_n10049, new_n8002, new_n10051);
xor_4  g07703(new_n10020, new_n9994, new_n10052);
and_5  g07704(new_n10052, new_n8006_1, new_n10053_1);
xor_4  g07705(new_n7928, new_n7909, new_n10054);
xnor_4 g07706(new_n10052, new_n10054, new_n10055_1);
xnor_4 g07707(new_n10018_1, new_n10017_1, new_n10056);
and_5  g07708(new_n10056, new_n8013, new_n10057_1);
xnor_4 g07709(new_n10015, new_n9999, new_n10058);
nor_5  g07710(new_n10058, new_n8015, new_n10059);
xnor_4 g07711(new_n10058, new_n8015, new_n10060);
xor_4  g07712(new_n10013, new_n10004, new_n10061);
and_5  g07713(new_n10061, new_n8021, new_n10062);
not_10 g07714(new_n8026, new_n10063);
xnor_4 g07715(new_n10005, new_n3968, new_n10064);
nor_5  g07716(new_n10064, new_n8028, new_n10065);
and_5  g07717(new_n10065, new_n10063, new_n10066);
xnor_4 g07718(new_n10011, new_n3964, new_n10067);
xnor_4 g07719(new_n10065, new_n8026, new_n10068);
and_5  g07720(new_n10068, new_n10067, new_n10069);
nor_5  g07721(new_n10069, new_n10066, new_n10070);
not_10 g07722(new_n8021, new_n10071);
xnor_4 g07723(new_n10061, new_n10071, new_n10072);
and_5  g07724(new_n10072, new_n10070, new_n10073);
nor_5  g07725(new_n10073, new_n10062, new_n10074);
nor_5  g07726(new_n10074, new_n10060, new_n10075);
or_5   g07727(new_n10075, new_n10059, new_n10076);
xnor_4 g07728(new_n10056, new_n8013, new_n10077);
nor_5  g07729(new_n10077, new_n10076, new_n10078);
nor_5  g07730(new_n10078, new_n10057_1, new_n10079);
and_5  g07731(new_n10079, new_n10055_1, new_n10080);
nor_5  g07732(new_n10080, new_n10053_1, new_n10081);
nor_5  g07733(new_n10081, new_n10051, new_n10082);
nor_5  g07734(new_n10082, new_n10050, new_n10083);
nor_5  g07735(new_n10083, new_n10048, new_n10084);
nor_5  g07736(new_n10084, new_n10047, new_n10085);
nor_5  g07737(new_n10085, new_n10045, new_n10086);
nor_5  g07738(new_n10086, new_n10044, new_n10087);
nor_5  g07739(new_n10087, new_n10042, new_n10088);
nor_5  g07740(new_n10088, new_n10041, new_n10089);
xnor_4 g07741(new_n10038, new_n10036, new_n10090);
nor_5  g07742(new_n10090, new_n10089, new_n10091);
or_5   g07743(new_n10091, new_n10039, new_n10092);
xor_4  g07744(new_n10092, new_n10037, n1527);
xor_4  g07745(n25345, n23463, new_n10094);
not_10 g07746(n13074, new_n10095);
nor_5  g07747(new_n10095, n9655, new_n10096_1);
xor_4  g07748(n13074, n9655, new_n10097);
not_10 g07749(n10739, new_n10098);
nor_5  g07750(n13490, new_n10098, new_n10099);
xor_4  g07751(n13490, n10739, new_n10100);
nor_5  g07752(n22660, new_n2350, new_n10101_1);
xor_4  g07753(n22660, n21753, new_n10102);
nor_5  g07754(new_n2353, n1777, new_n10103);
xor_4  g07755(n21832, n1777, new_n10104);
nor_5  g07756(new_n2356, n8745, new_n10105);
nor_5  g07757(n16223, new_n5092, new_n10106);
nor_5  g07758(new_n8845, new_n8840, new_n10107);
or_5   g07759(new_n10107, new_n10106, new_n10108);
xor_4  g07760(n26913, n8745, new_n10109);
nor_5  g07761(new_n10109, new_n10108, new_n10110);
nor_5  g07762(new_n10110, new_n10105, new_n10111_1);
nor_5  g07763(new_n10111_1, new_n10104, new_n10112);
nor_5  g07764(new_n10112, new_n10103, new_n10113);
nor_5  g07765(new_n10113, new_n10102, new_n10114);
nor_5  g07766(new_n10114, new_n10101_1, new_n10115);
nor_5  g07767(new_n10115, new_n10100, new_n10116);
nor_5  g07768(new_n10116, new_n10099, new_n10117_1);
nor_5  g07769(new_n10117_1, new_n10097, new_n10118);
nor_5  g07770(new_n10118, new_n10096_1, new_n10119);
xor_4  g07771(new_n10119, new_n10094, new_n10120);
xnor_4 g07772(new_n10120, new_n7144, new_n10121);
xor_4  g07773(new_n10117_1, new_n10097, new_n10122);
nor_5  g07774(new_n10122, new_n7149_1, new_n10123);
xnor_4 g07775(new_n10122, new_n7149_1, new_n10124);
xor_4  g07776(new_n10115, new_n10100, new_n10125_1);
nor_5  g07777(new_n10125_1, new_n7154, new_n10126);
xnor_4 g07778(new_n10125_1, new_n7154, new_n10127);
xor_4  g07779(new_n10113, new_n10102, new_n10128);
nor_5  g07780(new_n10128, new_n7158, new_n10129);
xnor_4 g07781(new_n10128, new_n7158, new_n10130);
xor_4  g07782(new_n10111_1, new_n10104, new_n10131);
nor_5  g07783(new_n10131, new_n7165, new_n10132);
xnor_4 g07784(new_n10131, new_n7165, new_n10133);
xor_4  g07785(new_n10109, new_n10108, new_n10134);
nor_5  g07786(new_n10134, new_n7168, new_n10135);
and_5  g07787(new_n8846, new_n7173, new_n10136);
nor_5  g07788(new_n8855, new_n8847, new_n10137);
nor_5  g07789(new_n10137, new_n10136, new_n10138);
xnor_4 g07790(new_n10134, new_n7168, new_n10139);
nor_5  g07791(new_n10139, new_n10138, new_n10140);
nor_5  g07792(new_n10140, new_n10135, new_n10141);
nor_5  g07793(new_n10141, new_n10133, new_n10142);
nor_5  g07794(new_n10142, new_n10132, new_n10143);
nor_5  g07795(new_n10143, new_n10130, new_n10144);
nor_5  g07796(new_n10144, new_n10129, new_n10145);
nor_5  g07797(new_n10145, new_n10127, new_n10146);
nor_5  g07798(new_n10146, new_n10126, new_n10147);
nor_5  g07799(new_n10147, new_n10124, new_n10148);
or_5   g07800(new_n10148, new_n10123, new_n10149);
xor_4  g07801(new_n10149, new_n10121, n1580);
xnor_4 g07802(n18962, n12315, new_n10151);
or_5   g07803(new_n10151, new_n6717, new_n10152);
or_5   g07804(new_n7918, n12315, new_n10153);
xor_4  g07805(n10158, n3952, new_n10154);
xor_4  g07806(new_n10154, new_n10153, new_n10155);
xnor_4 g07807(new_n10155, new_n10152, new_n10156);
xor_4  g07808(new_n10156, new_n6722, n1586);
xor_4  g07809(n19539, n1483, new_n10158_1);
not_10 g07810(n8194, new_n10159);
nor_5  g07811(n24093, new_n10159, new_n10160);
xor_4  g07812(n24093, n8194, new_n10161);
not_10 g07813(n23657, new_n10162);
nor_5  g07814(new_n10162, n23035, new_n10163);
xor_4  g07815(n23657, n23035, new_n10164);
not_10 g07816(n16911, new_n10165_1);
nor_5  g07817(new_n10165_1, n7773, new_n10166);
nor_5  g07818(new_n5874, new_n5846, new_n10167);
nor_5  g07819(new_n10167, new_n10166, new_n10168);
nor_5  g07820(new_n10168, new_n10164, new_n10169);
nor_5  g07821(new_n10169, new_n10163, new_n10170);
nor_5  g07822(new_n10170, new_n10161, new_n10171);
nor_5  g07823(new_n10171, new_n10160, new_n10172);
xnor_4 g07824(new_n10172, new_n10158_1, new_n10173);
xor_4  g07825(n25494, n1314, new_n10174);
not_10 g07826(n3306, new_n10175);
nor_5  g07827(n10117, new_n10175, new_n10176);
xor_4  g07828(n10117, n3306, new_n10177);
not_10 g07829(n22335, new_n10178);
nor_5  g07830(new_n10178, n13460, new_n10179);
xor_4  g07831(n22335, n13460, new_n10180);
not_10 g07832(n24048, new_n10181);
nor_5  g07833(new_n10181, n6104, new_n10182);
not_10 g07834(n1525, new_n10183);
nor_5  g07835(n4119, new_n10183, new_n10184);
nor_5  g07836(new_n4313, new_n4292, new_n10185);
nor_5  g07837(new_n10185, new_n10184, new_n10186);
xor_4  g07838(n24048, n6104, new_n10187);
nor_5  g07839(new_n10187, new_n10186, new_n10188);
nor_5  g07840(new_n10188, new_n10182, new_n10189);
nor_5  g07841(new_n10189, new_n10180, new_n10190);
nor_5  g07842(new_n10190, new_n10179, new_n10191);
nor_5  g07843(new_n10191, new_n10177, new_n10192);
nor_5  g07844(new_n10192, new_n10176, new_n10193);
xor_4  g07845(new_n10193, new_n10174, new_n10194);
xor_4  g07846(n25296, n23717, new_n10195);
not_10 g07847(n7788, new_n10196);
nor_5  g07848(n20013, new_n10196, new_n10197);
xor_4  g07849(n20013, n7788, new_n10198);
not_10 g07850(n5443, new_n10199);
nor_5  g07851(new_n10199, n1320, new_n10200);
xor_4  g07852(n5443, n1320, new_n10201_1);
not_10 g07853(n18584, new_n10202);
nor_5  g07854(n19803, new_n10202, new_n10203);
nor_5  g07855(new_n5844, new_n5840_1, new_n10204);
nor_5  g07856(new_n10204, new_n10203, new_n10205);
nor_5  g07857(new_n10205, new_n10201_1, new_n10206);
nor_5  g07858(new_n10206, new_n10200, new_n10207);
nor_5  g07859(new_n10207, new_n10198, new_n10208);
nor_5  g07860(new_n10208, new_n10197, new_n10209);
xor_4  g07861(new_n10209, new_n10195, new_n10210);
xnor_4 g07862(new_n10210, new_n10194, new_n10211);
xor_4  g07863(new_n10191, new_n10177, new_n10212);
xor_4  g07864(new_n10207, new_n10198, new_n10213);
and_5  g07865(new_n10213, new_n10212, new_n10214);
xnor_4 g07866(new_n10213, new_n10212, new_n10215);
xor_4  g07867(new_n10189, new_n10180, new_n10216);
xor_4  g07868(new_n10205, new_n10201_1, new_n10217);
nor_5  g07869(new_n10217, new_n10216, new_n10218);
xnor_4 g07870(new_n10217, new_n10216, new_n10219);
xor_4  g07871(new_n10187, new_n10186, new_n10220);
not_10 g07872(new_n10220, new_n10221);
nor_5  g07873(new_n10221, new_n5845, new_n10222);
xor_4  g07874(new_n10220, new_n5845, new_n10223);
and_5  g07875(new_n4338, new_n4314, new_n10224);
nor_5  g07876(new_n4371, new_n4339, new_n10225);
nor_5  g07877(new_n10225, new_n10224, new_n10226);
nor_5  g07878(new_n10226, new_n10223, new_n10227);
or_5   g07879(new_n10227, new_n10222, new_n10228);
nor_5  g07880(new_n10228, new_n10219, new_n10229);
or_5   g07881(new_n10229, new_n10218, new_n10230);
nor_5  g07882(new_n10230, new_n10215, new_n10231);
nor_5  g07883(new_n10231, new_n10214, new_n10232);
xnor_4 g07884(new_n10232, new_n10211, new_n10233);
xnor_4 g07885(new_n10233, new_n10173, new_n10234);
xor_4  g07886(new_n10170, new_n10161, new_n10235);
xor_4  g07887(new_n10230, new_n10215, new_n10236_1);
nor_5  g07888(new_n10236_1, new_n10235, new_n10237);
xnor_4 g07889(new_n10236_1, new_n10235, new_n10238);
xor_4  g07890(new_n10168, new_n10164, new_n10239_1);
xnor_4 g07891(new_n10228, new_n10219, new_n10240);
nor_5  g07892(new_n10240, new_n10239_1, new_n10241);
xnor_4 g07893(new_n10240, new_n10239_1, new_n10242);
xor_4  g07894(new_n5874, new_n5846, new_n10243);
xor_4  g07895(new_n10226, new_n10223, new_n10244_1);
nor_5  g07896(new_n10244_1, new_n10243, new_n10245);
xnor_4 g07897(new_n10244_1, new_n10243, new_n10246);
xor_4  g07898(new_n5872, new_n5849, new_n10247);
nor_5  g07899(new_n10247, new_n4372, new_n10248);
nor_5  g07900(new_n5919, new_n4375, new_n10249);
xnor_4 g07901(new_n5919, new_n4375, new_n10250_1);
nor_5  g07902(new_n5923, new_n4378, new_n10251);
and_5  g07903(new_n5928, new_n4381, new_n10252);
xnor_4 g07904(new_n5928, new_n4381, new_n10253);
nor_5  g07905(new_n5932, new_n4387, new_n10254);
nor_5  g07906(new_n10254, new_n5936_1, new_n10255);
xnor_4 g07907(new_n10254, new_n5935, new_n10256);
and_5  g07908(new_n10256, new_n4392, new_n10257);
nor_5  g07909(new_n10257, new_n10255, new_n10258);
nor_5  g07910(new_n10258, new_n10253, new_n10259);
nor_5  g07911(new_n10259, new_n10252, new_n10260);
xnor_4 g07912(new_n5923, new_n4378, new_n10261_1);
nor_5  g07913(new_n10261_1, new_n10260, new_n10262_1);
nor_5  g07914(new_n10262_1, new_n10251, new_n10263);
nor_5  g07915(new_n10263, new_n10250_1, new_n10264);
nor_5  g07916(new_n10264, new_n10249, new_n10265);
xnor_4 g07917(new_n10247, new_n4372, new_n10266);
nor_5  g07918(new_n10266, new_n10265, new_n10267);
nor_5  g07919(new_n10267, new_n10248, new_n10268);
nor_5  g07920(new_n10268, new_n10246, new_n10269);
nor_5  g07921(new_n10269, new_n10245, new_n10270);
nor_5  g07922(new_n10270, new_n10242, new_n10271);
nor_5  g07923(new_n10271, new_n10241, new_n10272);
nor_5  g07924(new_n10272, new_n10238, new_n10273);
or_5   g07925(new_n10273, new_n10237, new_n10274);
xor_4  g07926(new_n10274, new_n10234, n1590);
xnor_4 g07927(new_n6906, new_n6892, n1602);
xor_4  g07928(new_n2763, new_n2715, n1634);
xnor_4 g07929(new_n10272, new_n10238, n1636);
nor_5  g07930(n10514, n4514, new_n10279);
xnor_4 g07931(n10514, n4514, new_n10280);
nor_5  g07932(n18649, n3984, new_n10281);
xnor_4 g07933(n18649, n3984, new_n10282);
and_5  g07934(n19652, n6218, new_n10283);
or_5   g07935(n19652, n6218, new_n10284);
nor_5  g07936(n20470, n3366, new_n10285);
nor_5  g07937(new_n9863, new_n9856, new_n10286);
nor_5  g07938(new_n10286, new_n10285, new_n10287_1);
and_5  g07939(new_n10287_1, new_n10284, new_n10288);
or_5   g07940(new_n10288, new_n10283, new_n10289);
nor_5  g07941(new_n10289, new_n10282, new_n10290);
nor_5  g07942(new_n10290, new_n10281, new_n10291);
nor_5  g07943(new_n10291, new_n10280, new_n10292);
or_5   g07944(new_n10292, new_n10279, new_n10293);
xnor_4 g07945(n18880, n2978, new_n10294);
nor_5  g07946(n25475, n23697, new_n10295_1);
nor_5  g07947(new_n6155, new_n6126, new_n10296);
nor_5  g07948(new_n10296, new_n10295_1, new_n10297);
xnor_4 g07949(new_n10297, new_n10294, new_n10298);
and_5  g07950(new_n10298, n20040, new_n10299);
xnor_4 g07951(new_n10298, n20040, new_n10300);
nand_5 g07952(new_n6156, n19531, new_n10301);
xnor_4 g07953(new_n6156, n19531, new_n10302);
nor_5  g07954(new_n6158, n18345, new_n10303);
xnor_4 g07955(new_n6158, n18345, new_n10304);
or_5   g07956(new_n6161, n13190, new_n10305);
xnor_4 g07957(new_n6161, n13190, new_n10306);
and_5  g07958(new_n6164, n3460, new_n10307);
and_5  g07959(new_n6166, n5226, new_n10308);
nor_5  g07960(new_n8665, new_n8652, new_n10309);
nor_5  g07961(new_n10309, new_n10308, new_n10310);
xnor_4 g07962(new_n6164, n3460, new_n10311);
nor_5  g07963(new_n10311, new_n10310, new_n10312);
nor_5  g07964(new_n10312, new_n10307, new_n10313);
not_10 g07965(new_n10313, new_n10314);
or_5   g07966(new_n10314, new_n10306, new_n10315);
and_5  g07967(new_n10315, new_n10305, new_n10316);
nor_5  g07968(new_n10316, new_n10304, new_n10317);
or_5   g07969(new_n10317, new_n10303, new_n10318);
or_5   g07970(new_n10318, new_n10302, new_n10319);
and_5  g07971(new_n10319, new_n10301, new_n10320);
nor_5  g07972(new_n10320, new_n10300, new_n10321_1);
nor_5  g07973(new_n10321_1, new_n10299, new_n10322);
nor_5  g07974(n18880, n2978, new_n10323);
nor_5  g07975(new_n10297, new_n10294, new_n10324);
or_5   g07976(new_n10324, new_n10323, new_n10325);
xnor_4 g07977(new_n10325, new_n10322, new_n10326_1);
nor_5  g07978(new_n8650, n19575, new_n10327_1);
not_10 g07979(new_n10327_1, new_n10328);
or_5   g07980(new_n10328, n26512, new_n10329);
or_5   g07981(new_n10329, n26191, new_n10330_1);
or_5   g07982(new_n10330_1, n5386, new_n10331);
or_5   g07983(new_n10331, n17037, new_n10332);
nor_5  g07984(new_n10332, n7569, new_n10333);
xnor_4 g07985(new_n10333, new_n10326_1, new_n10334);
xor_4  g07986(new_n10320, new_n10300, new_n10335);
xor_4  g07987(new_n10332, n7569, new_n10336);
nor_5  g07988(new_n10336, new_n10335, new_n10337);
xnor_4 g07989(new_n10336, new_n10335, new_n10338);
xor_4  g07990(new_n10318, new_n10302, new_n10339);
xor_4  g07991(new_n10331, n17037, new_n10340_1);
nor_5  g07992(new_n10340_1, new_n10339, new_n10341);
xnor_4 g07993(new_n10340_1, new_n10339, new_n10342);
xnor_4 g07994(new_n10316, new_n10304, new_n10343);
xor_4  g07995(new_n10330_1, n5386, new_n10344);
nor_5  g07996(new_n10344, new_n10343, new_n10345_1);
xor_4  g07997(new_n10316, new_n10304, new_n10346);
xor_4  g07998(new_n10344, new_n10346, new_n10347);
xnor_4 g07999(new_n10313, new_n10306, new_n10348);
not_10 g08000(new_n10348, new_n10349);
xor_4  g08001(new_n10329, n26191, new_n10350);
or_5   g08002(new_n10350, new_n10349, new_n10351);
xnor_4 g08003(new_n10327_1, n26512, new_n10352);
xor_4  g08004(new_n10311, new_n10310, new_n10353);
and_5  g08005(new_n10353, new_n10352, new_n10354);
xor_4  g08006(new_n10353, new_n10352, new_n10355);
nor_5  g08007(new_n8666, new_n8651, new_n10356_1);
nor_5  g08008(new_n8687_1, new_n8667, new_n10357);
nor_5  g08009(new_n10357, new_n10356_1, new_n10358);
and_5  g08010(new_n10358, new_n10355, new_n10359);
nor_5  g08011(new_n10359, new_n10354, new_n10360);
not_10 g08012(new_n10360, new_n10361);
xor_4  g08013(new_n10350, new_n10348, new_n10362);
or_5   g08014(new_n10362, new_n10361, new_n10363);
and_5  g08015(new_n10363, new_n10351, new_n10364);
nor_5  g08016(new_n10364, new_n10347, new_n10365);
nor_5  g08017(new_n10365, new_n10345_1, new_n10366);
nor_5  g08018(new_n10366, new_n10342, new_n10367);
nor_5  g08019(new_n10367, new_n10341, new_n10368);
nor_5  g08020(new_n10368, new_n10338, new_n10369);
nor_5  g08021(new_n10369, new_n10337, new_n10370);
xnor_4 g08022(new_n10370, new_n10334, new_n10371);
xnor_4 g08023(new_n10371, new_n10293, new_n10372_1);
xnor_4 g08024(new_n10368, new_n10338, new_n10373);
xor_4  g08025(new_n10291, new_n10280, new_n10374);
nor_5  g08026(new_n10374, new_n10373, new_n10375);
xnor_4 g08027(new_n10374, new_n10373, new_n10376);
xnor_4 g08028(new_n10366, new_n10342, new_n10377);
xor_4  g08029(new_n10289, new_n10282, new_n10378);
nor_5  g08030(new_n10378, new_n10377, new_n10379);
xnor_4 g08031(new_n10378, new_n10377, new_n10380);
xnor_4 g08032(new_n10364, new_n10347, new_n10381);
xor_4  g08033(n19652, n6218, new_n10382);
xnor_4 g08034(new_n10382, new_n10287_1, new_n10383);
nor_5  g08035(new_n10383, new_n10381, new_n10384);
xnor_4 g08036(new_n10383, new_n10381, new_n10385_1);
xnor_4 g08037(new_n9863, new_n9856, new_n10386);
xnor_4 g08038(new_n10362, new_n10360, new_n10387_1);
and_5  g08039(new_n10387_1, new_n10386, new_n10388_1);
xnor_4 g08040(new_n10387_1, new_n9864, new_n10389);
not_10 g08041(new_n9868, new_n10390_1);
xor_4  g08042(new_n10358, new_n10355, new_n10391);
and_5  g08043(new_n10391, new_n10390_1, new_n10392);
nor_5  g08044(new_n10391, new_n10390_1, new_n10393);
nor_5  g08045(new_n8688, new_n8647, new_n10394);
nor_5  g08046(new_n8709, new_n8689, new_n10395);
nor_5  g08047(new_n10395, new_n10394, new_n10396);
nor_5  g08048(new_n10396, new_n10393, new_n10397);
nor_5  g08049(new_n10397, new_n10392, new_n10398);
and_5  g08050(new_n10398, new_n10389, new_n10399);
nor_5  g08051(new_n10399, new_n10388_1, new_n10400);
nor_5  g08052(new_n10400, new_n10385_1, new_n10401);
nor_5  g08053(new_n10401, new_n10384, new_n10402);
nor_5  g08054(new_n10402, new_n10380, new_n10403);
nor_5  g08055(new_n10403, new_n10379, new_n10404_1);
nor_5  g08056(new_n10404_1, new_n10376, new_n10405_1);
nor_5  g08057(new_n10405_1, new_n10375, new_n10406);
xnor_4 g08058(new_n10406, new_n10372_1, n1684);
xnor_4 g08059(new_n5669, n3984, new_n10408);
nor_5  g08060(new_n5672, n19652, new_n10409_1);
xnor_4 g08061(new_n5672, n19652, new_n10410);
nor_5  g08062(new_n5675, n3366, new_n10411_1);
xnor_4 g08063(new_n5675, n3366, new_n10412);
nor_5  g08064(new_n3763, n26565, new_n10413);
xnor_4 g08065(new_n3763, n26565, new_n10414);
nor_5  g08066(new_n3765, n3959, new_n10415);
xnor_4 g08067(new_n3765, n3959, new_n10416);
nor_5  g08068(new_n3767, n11566, new_n10417);
xnor_4 g08069(new_n3767, n11566, new_n10418);
nor_5  g08070(new_n3770, n26744, new_n10419);
xnor_4 g08071(new_n3770, n26744, new_n10420_1);
nor_5  g08072(new_n3773, n26625, new_n10421);
and_5  g08073(n19922, n14230, new_n10422);
xnor_4 g08074(new_n3773, n26625, new_n10423);
nor_5  g08075(new_n10423, new_n10422, new_n10424);
nor_5  g08076(new_n10424, new_n10421, new_n10425);
nor_5  g08077(new_n10425, new_n10420_1, new_n10426);
nor_5  g08078(new_n10426, new_n10419, new_n10427);
nor_5  g08079(new_n10427, new_n10418, new_n10428);
nor_5  g08080(new_n10428, new_n10417, new_n10429);
nor_5  g08081(new_n10429, new_n10416, new_n10430);
nor_5  g08082(new_n10430, new_n10415, new_n10431);
nor_5  g08083(new_n10431, new_n10414, new_n10432_1);
nor_5  g08084(new_n10432_1, new_n10413, new_n10433);
nor_5  g08085(new_n10433, new_n10412, new_n10434);
nor_5  g08086(new_n10434, new_n10411_1, new_n10435);
nor_5  g08087(new_n10435, new_n10410, new_n10436);
nor_5  g08088(new_n10436, new_n10409_1, new_n10437);
xor_4  g08089(new_n10437, new_n10408, new_n10438);
nor_5  g08090(new_n10438, n13026, new_n10439);
xnor_4 g08091(new_n10438, n13026, new_n10440);
xor_4  g08092(new_n10435, new_n10410, new_n10441);
nor_5  g08093(new_n10441, n2175, new_n10442);
xnor_4 g08094(new_n10441, n2175, new_n10443);
xor_4  g08095(new_n10433, new_n10412, new_n10444);
nor_5  g08096(new_n10444, n752, new_n10445);
xnor_4 g08097(new_n10444, n752, new_n10446);
xor_4  g08098(new_n10431, new_n10414, new_n10447);
nor_5  g08099(new_n10447, n1611, new_n10448);
xor_4  g08100(new_n10429, new_n10416, new_n10449);
nor_5  g08101(new_n10449, n25094, new_n10450);
xnor_4 g08102(new_n10449, n25094, new_n10451);
xor_4  g08103(new_n10427, new_n10418, new_n10452);
nor_5  g08104(new_n10452, n21538, new_n10453);
xnor_4 g08105(new_n10452, n21538, new_n10454);
xor_4  g08106(new_n10425, new_n10420_1, new_n10455);
nor_5  g08107(new_n10455, n5131, new_n10456);
xor_4  g08108(new_n10423, new_n10422, new_n10457);
nor_5  g08109(new_n10457, n11473, new_n10458);
xnor_4 g08110(n19922, n14230, new_n10459);
and_5  g08111(new_n10459, n15506, new_n10460);
xnor_4 g08112(new_n10457, n11473, new_n10461);
nor_5  g08113(new_n10461, new_n10460, new_n10462);
nor_5  g08114(new_n10462, new_n10458, new_n10463);
xnor_4 g08115(new_n10455, n5131, new_n10464);
nor_5  g08116(new_n10464, new_n10463, new_n10465);
nor_5  g08117(new_n10465, new_n10456, new_n10466);
nor_5  g08118(new_n10466, new_n10454, new_n10467);
nor_5  g08119(new_n10467, new_n10453, new_n10468);
nor_5  g08120(new_n10468, new_n10451, new_n10469);
nor_5  g08121(new_n10469, new_n10450, new_n10470);
xnor_4 g08122(new_n10447, n1611, new_n10471);
nor_5  g08123(new_n10471, new_n10470, new_n10472);
nor_5  g08124(new_n10472, new_n10448, new_n10473);
nor_5  g08125(new_n10473, new_n10446, new_n10474);
nor_5  g08126(new_n10474, new_n10445, new_n10475);
nor_5  g08127(new_n10475, new_n10443, new_n10476);
nor_5  g08128(new_n10476, new_n10442, new_n10477);
nor_5  g08129(new_n10477, new_n10440, new_n10478);
nor_5  g08130(new_n10478, new_n10439, new_n10479);
and_5  g08131(new_n10479, n23912, new_n10480);
xnor_4 g08132(new_n10479, n23912, new_n10481);
nor_5  g08133(new_n5669, n3984, new_n10482);
nor_5  g08134(new_n10437, new_n10408, new_n10483);
or_5   g08135(new_n10483, new_n10482, new_n10484_1);
xor_4  g08136(new_n5665, n4514, new_n10485);
xnor_4 g08137(new_n10485, new_n10484_1, new_n10486);
nor_5  g08138(new_n10486, new_n10481, new_n10487);
or_5   g08139(new_n10487, new_n10480, new_n10488);
and_5  g08140(new_n5665, n4514, new_n10489_1);
nor_5  g08141(new_n5665, n4514, new_n10490);
nor_5  g08142(new_n10490, new_n10484_1, new_n10491);
or_5   g08143(new_n10491, new_n5667, new_n10492);
nor_5  g08144(new_n10492, new_n10489_1, new_n10493);
nor_5  g08145(new_n10493, new_n10488, new_n10494);
not_10 g08146(new_n4148, new_n10495);
nor_5  g08147(new_n10495, n15766, new_n10496);
xor_4  g08148(new_n4148, n15766, new_n10497);
nor_5  g08149(new_n4153_1, n25629, new_n10498);
xnor_4 g08150(new_n4153_1, n25629, new_n10499);
nor_5  g08151(new_n4157, n7692, new_n10500);
xnor_4 g08152(new_n4157, n7692, new_n10501);
nor_5  g08153(new_n4161, n23039, new_n10502);
xnor_4 g08154(new_n4161, n23039, new_n10503);
nor_5  g08155(new_n3725_1, n13677, new_n10504);
nor_5  g08156(new_n3750, new_n3726, new_n10505);
nor_5  g08157(new_n10505, new_n10504, new_n10506);
nor_5  g08158(new_n10506, new_n10503, new_n10507);
nor_5  g08159(new_n10507, new_n10502, new_n10508);
nor_5  g08160(new_n10508, new_n10501, new_n10509);
nor_5  g08161(new_n10509, new_n10500, new_n10510);
nor_5  g08162(new_n10510, new_n10499, new_n10511);
nor_5  g08163(new_n10511, new_n10498, new_n10512);
nor_5  g08164(new_n10512, new_n10497, new_n10513);
or_5   g08165(new_n10513, new_n10496, new_n10514_1);
or_5   g08166(new_n10514_1, new_n4136, new_n10515);
xnor_4 g08167(new_n10514_1, new_n4135, new_n10516);
xor_4  g08168(new_n10493, new_n10488, new_n10517);
nor_5  g08169(new_n10517, new_n10516, new_n10518);
xnor_4 g08170(new_n10517, new_n10516, new_n10519);
xor_4  g08171(new_n10512, new_n10497, new_n10520);
xor_4  g08172(new_n10486, new_n10481, new_n10521);
and_5  g08173(new_n10521, new_n10520, new_n10522);
xor_4  g08174(new_n10510, new_n10499, new_n10523);
not_10 g08175(new_n10523, new_n10524);
xor_4  g08176(new_n10477, new_n10440, new_n10525_1);
nor_5  g08177(new_n10525_1, new_n10524, new_n10526);
xor_4  g08178(new_n10525_1, new_n10523, new_n10527);
xor_4  g08179(new_n10508, new_n10501, new_n10528);
not_10 g08180(new_n10528, new_n10529);
xor_4  g08181(new_n10475, new_n10443, new_n10530);
nor_5  g08182(new_n10530, new_n10529, new_n10531);
xor_4  g08183(new_n10530, new_n10528, new_n10532);
xnor_4 g08184(new_n10506, new_n10503, new_n10533);
xor_4  g08185(new_n10473, new_n10446, new_n10534);
nor_5  g08186(new_n10534, new_n10533, new_n10535);
xnor_4 g08187(new_n10534, new_n10533, new_n10536);
xor_4  g08188(new_n10471, new_n10470, new_n10537);
nor_5  g08189(new_n10537, new_n3751, new_n10538);
xnor_4 g08190(new_n10537, new_n3751, new_n10539);
not_10 g08191(new_n3817, new_n10540_1);
xor_4  g08192(new_n10468, new_n10451, new_n10541);
nor_5  g08193(new_n10541, new_n10540_1, new_n10542);
xor_4  g08194(new_n10466, new_n10454, new_n10543);
nor_5  g08195(new_n10543, new_n3821, new_n10544);
xnor_4 g08196(new_n10543, new_n3821, new_n10545);
xor_4  g08197(new_n10464, new_n10463, new_n10546);
nor_5  g08198(new_n10546, new_n3824, new_n10547);
xor_4  g08199(new_n10461, new_n10460, new_n10548);
nor_5  g08200(new_n10548, new_n3829, new_n10549);
xor_4  g08201(new_n10459, n15506, new_n10550);
or_5   g08202(new_n10550, new_n2531, new_n10551);
xor_4  g08203(new_n10548, new_n3829, new_n10552);
and_5  g08204(new_n10552, new_n10551, new_n10553);
nor_5  g08205(new_n10553, new_n10549, new_n10554);
xnor_4 g08206(new_n10546, new_n3824, new_n10555);
nor_5  g08207(new_n10555, new_n10554, new_n10556);
nor_5  g08208(new_n10556, new_n10547, new_n10557);
nor_5  g08209(new_n10557, new_n10545, new_n10558);
or_5   g08210(new_n10558, new_n10544, new_n10559);
xnor_4 g08211(new_n10541, new_n3817, new_n10560);
and_5  g08212(new_n10560, new_n10559, new_n10561_1);
nor_5  g08213(new_n10561_1, new_n10542, new_n10562);
nor_5  g08214(new_n10562, new_n10539, new_n10563);
nor_5  g08215(new_n10563, new_n10538, new_n10564_1);
nor_5  g08216(new_n10564_1, new_n10536, new_n10565);
nor_5  g08217(new_n10565, new_n10535, new_n10566);
nor_5  g08218(new_n10566, new_n10532, new_n10567);
nor_5  g08219(new_n10567, new_n10531, new_n10568);
nor_5  g08220(new_n10568, new_n10527, new_n10569);
or_5   g08221(new_n10569, new_n10526, new_n10570);
xor_4  g08222(new_n10521, new_n10520, new_n10571);
and_5  g08223(new_n10571, new_n10570, new_n10572);
nor_5  g08224(new_n10572, new_n10522, new_n10573);
nor_5  g08225(new_n10573, new_n10519, new_n10574);
nor_5  g08226(new_n10574, new_n10518, new_n10575);
xnor_4 g08227(new_n10575, new_n10515, new_n10576);
xnor_4 g08228(new_n10576, new_n10494, n1701);
xnor_4 g08229(new_n3693, new_n3663, n1703);
xnor_4 g08230(new_n4260, new_n4213, n1721);
nor_5  g08231(new_n7018, new_n4052, new_n10580);
nor_5  g08232(new_n8145, new_n8144, new_n10581);
or_5   g08233(new_n10581, new_n10580, new_n10582);
and_5  g08234(new_n10582, new_n8193, new_n10583);
nor_5  g08235(new_n8193, new_n8146, new_n10584);
nor_5  g08236(new_n8254, new_n8194_1, new_n10585);
nor_5  g08237(new_n10585, new_n10584, new_n10586);
nor_5  g08238(new_n10586, new_n10583, new_n10587);
nor_5  g08239(new_n10582, new_n8193, new_n10588_1);
nor_5  g08240(new_n10588_1, new_n10585, new_n10589);
nor_5  g08241(new_n10589, new_n10587, n1760);
xnor_4 g08242(new_n3834, new_n3827, n1791);
xor_4  g08243(new_n3216, new_n3215, n1808);
and_5  g08244(new_n7018, new_n6970, new_n10593_1);
nor_5  g08245(new_n7080, new_n7019, new_n10594);
nor_5  g08246(new_n10594, new_n10593_1, new_n10595_1);
not_10 g08247(n4319, new_n10596);
nor_5  g08248(n13494, new_n10596, new_n10597);
xor_4  g08249(n13494, n4319, new_n10598);
not_10 g08250(n23463, new_n10599);
nor_5  g08251(n25345, new_n10599, new_n10600);
nor_5  g08252(new_n10119, new_n10094, new_n10601);
nor_5  g08253(new_n10601, new_n10600, new_n10602);
nor_5  g08254(new_n10602, new_n10598, new_n10603);
nor_5  g08255(new_n10603, new_n10597, new_n10604);
and_5  g08256(new_n10604, new_n10595_1, new_n10605);
nor_5  g08257(new_n10604, new_n7081, new_n10606);
xor_4  g08258(new_n10604, new_n7081, new_n10607);
xor_4  g08259(new_n10602, new_n10598, new_n10608);
and_5  g08260(new_n10608, new_n7139_1, new_n10609);
xnor_4 g08261(new_n10608, new_n7139_1, new_n10610);
and_5  g08262(new_n10120, new_n7144, new_n10611_1);
nor_5  g08263(new_n10149, new_n10121, new_n10612);
nor_5  g08264(new_n10612, new_n10611_1, new_n10613);
nor_5  g08265(new_n10613, new_n10610, new_n10614_1);
nor_5  g08266(new_n10614_1, new_n10609, new_n10615);
and_5  g08267(new_n10615, new_n10607, new_n10616);
nor_5  g08268(new_n10616, new_n10606, new_n10617_1);
nor_5  g08269(new_n10617_1, new_n10605, new_n10618);
nor_5  g08270(new_n10604, new_n10595_1, new_n10619);
nor_5  g08271(new_n10619, new_n10616, new_n10620);
nor_5  g08272(new_n10620, new_n10618, n1821);
xor_4  g08273(new_n6290, new_n6288, n1832);
xnor_4 g08274(n9934, n2272, new_n10623);
nor_5  g08275(n25331, n18496, new_n10624);
xnor_4 g08276(n25331, n18496, new_n10625);
nor_5  g08277(n26224, n18483, new_n10626);
xnor_4 g08278(n26224, n18483, new_n10627);
nor_5  g08279(n21934, n19327, new_n10628_1);
xnor_4 g08280(n21934, n19327, new_n10629);
nor_5  g08281(n22597, n18901, new_n10630);
xnor_4 g08282(n22597, n18901, new_n10631);
nor_5  g08283(n26107, n4376, new_n10632);
xnor_4 g08284(n26107, n4376, new_n10633);
nor_5  g08285(n14570, n342, new_n10634);
xnor_4 g08286(n14570, n342, new_n10635);
nor_5  g08287(n26553, n23775, new_n10636);
xnor_4 g08288(n26553, n23775, new_n10637);
nor_5  g08289(n8259, n4964, new_n10638);
and_5  g08290(n11479, n7876, new_n10639);
xnor_4 g08291(n8259, n4964, new_n10640);
nor_5  g08292(new_n10640, new_n10639, new_n10641);
nor_5  g08293(new_n10641, new_n10638, new_n10642);
nor_5  g08294(new_n10642, new_n10637, new_n10643);
nor_5  g08295(new_n10643, new_n10636, new_n10644);
nor_5  g08296(new_n10644, new_n10635, new_n10645);
nor_5  g08297(new_n10645, new_n10634, new_n10646);
nor_5  g08298(new_n10646, new_n10633, new_n10647_1);
nor_5  g08299(new_n10647_1, new_n10632, new_n10648);
nor_5  g08300(new_n10648, new_n10631, new_n10649);
nor_5  g08301(new_n10649, new_n10630, new_n10650_1);
nor_5  g08302(new_n10650_1, new_n10629, new_n10651);
nor_5  g08303(new_n10651, new_n10628_1, new_n10652);
nor_5  g08304(new_n10652, new_n10627, new_n10653_1);
nor_5  g08305(new_n10653_1, new_n10626, new_n10654);
nor_5  g08306(new_n10654, new_n10625, new_n10655);
nor_5  g08307(new_n10655, new_n10624, new_n10656);
xor_4  g08308(new_n10656, new_n10623, new_n10657);
xnor_4 g08309(new_n10657, n2160, new_n10658);
xor_4  g08310(new_n10654, new_n10625, new_n10659);
nor_5  g08311(new_n10659, n10763, new_n10660);
xor_4  g08312(new_n10659, n10763, new_n10661);
xor_4  g08313(new_n10652, new_n10627, new_n10662);
and_5  g08314(new_n10662, n7437, new_n10663);
xnor_4 g08315(new_n10662, n7437, new_n10664);
xor_4  g08316(new_n10650_1, new_n10629, new_n10665);
and_5  g08317(new_n10665, n20700, new_n10666);
xnor_4 g08318(new_n10665, n20700, new_n10667);
xor_4  g08319(new_n10648, new_n10631, new_n10668);
and_5  g08320(new_n10668, n7099, new_n10669);
xnor_4 g08321(new_n10668, n7099, new_n10670);
xor_4  g08322(new_n10646, new_n10633, new_n10671);
and_5  g08323(new_n10671, n12811, new_n10672);
xnor_4 g08324(new_n10671, n12811, new_n10673);
xor_4  g08325(new_n10644, new_n10635, new_n10674);
and_5  g08326(new_n10674, n1118, new_n10675);
xnor_4 g08327(new_n10674, n1118, new_n10676);
xor_4  g08328(new_n10642, new_n10637, new_n10677);
and_5  g08329(new_n10677, n25974, new_n10678);
xor_4  g08330(new_n10677, n25974, new_n10679);
xnor_4 g08331(n11479, n7876, new_n10680);
and_5  g08332(new_n10680, n1451, new_n10681);
nor_5  g08333(new_n10681, n1630, new_n10682);
xor_4  g08334(new_n10640, new_n10639, new_n10683);
xnor_4 g08335(new_n10681, n1630, new_n10684);
nor_5  g08336(new_n10684, new_n10683, new_n10685);
nor_5  g08337(new_n10685, new_n10682, new_n10686);
and_5  g08338(new_n10686, new_n10679, new_n10687);
nor_5  g08339(new_n10687, new_n10678, new_n10688);
nor_5  g08340(new_n10688, new_n10676, new_n10689);
nor_5  g08341(new_n10689, new_n10675, new_n10690);
nor_5  g08342(new_n10690, new_n10673, new_n10691);
nor_5  g08343(new_n10691, new_n10672, new_n10692_1);
nor_5  g08344(new_n10692_1, new_n10670, new_n10693);
nor_5  g08345(new_n10693, new_n10669, new_n10694_1);
nor_5  g08346(new_n10694_1, new_n10667, new_n10695);
nor_5  g08347(new_n10695, new_n10666, new_n10696);
nor_5  g08348(new_n10696, new_n10664, new_n10697);
nor_5  g08349(new_n10697, new_n10663, new_n10698);
and_5  g08350(new_n10698, new_n10661, new_n10699);
nor_5  g08351(new_n10699, new_n10660, new_n10700);
xnor_4 g08352(new_n10700, new_n10658, new_n10701_1);
or_5   g08353(new_n3620, n4325, new_n10702);
or_5   g08354(new_n10702, n11926, new_n10703);
or_5   g08355(new_n10703, n5521, new_n10704);
xor_4  g08356(new_n10704, n21784, new_n10705);
xnor_4 g08357(new_n10705, new_n6591, new_n10706);
xor_4  g08358(new_n10703, n5521, new_n10707);
nor_5  g08359(new_n10707, new_n6595, new_n10708);
xnor_4 g08360(new_n10707, new_n6595, new_n10709);
xor_4  g08361(new_n10702, n11926, new_n10710_1);
nor_5  g08362(new_n10710_1, new_n6599, new_n10711);
xnor_4 g08363(new_n10710_1, new_n6599, new_n10712_1);
nor_5  g08364(new_n3621, new_n3614, new_n10713);
nor_5  g08365(new_n3656, new_n3622, new_n10714);
nor_5  g08366(new_n10714, new_n10713, new_n10715);
nor_5  g08367(new_n10715, new_n10712_1, new_n10716);
nor_5  g08368(new_n10716, new_n10711, new_n10717);
nor_5  g08369(new_n10717, new_n10709, new_n10718);
nor_5  g08370(new_n10718, new_n10708, new_n10719);
xor_4  g08371(new_n10719, new_n10706, new_n10720);
xnor_4 g08372(new_n10720, new_n10701_1, new_n10721);
xnor_4 g08373(new_n10698, new_n10661, new_n10722);
xor_4  g08374(new_n10717, new_n10709, new_n10723);
and_5  g08375(new_n10723, new_n10722, new_n10724);
xnor_4 g08376(new_n10723, new_n10722, new_n10725);
xor_4  g08377(new_n10696, new_n10664, new_n10726);
xor_4  g08378(new_n10715, new_n10712_1, new_n10727);
and_5  g08379(new_n10727, new_n10726, new_n10728);
xnor_4 g08380(new_n10727, new_n10726, new_n10729);
xor_4  g08381(new_n10694_1, new_n10667, new_n10730);
and_5  g08382(new_n10730, new_n3657, new_n10731);
xnor_4 g08383(new_n10730, new_n3657, new_n10732);
xor_4  g08384(new_n10692_1, new_n10670, new_n10733);
and_5  g08385(new_n10733, new_n3659, new_n10734);
xnor_4 g08386(new_n10733, new_n3659, new_n10735);
xor_4  g08387(new_n10690, new_n10673, new_n10736);
and_5  g08388(new_n10736, new_n3664, new_n10737);
xnor_4 g08389(new_n10736, new_n3664, new_n10738);
xor_4  g08390(new_n10688, new_n10676, new_n10739_1);
and_5  g08391(new_n10739_1, new_n3669, new_n10740);
xnor_4 g08392(new_n10739_1, new_n3669, new_n10741);
xnor_4 g08393(new_n10686, new_n10679, new_n10742);
nor_5  g08394(new_n10742, new_n3674, new_n10743);
xor_4  g08395(new_n10742, new_n3674, new_n10744);
xor_4  g08396(new_n10680, n1451, new_n10745);
nor_5  g08397(new_n10745, new_n3683, new_n10746);
xor_4  g08398(new_n10684, new_n10683, new_n10747);
and_5  g08399(new_n10747, new_n10746, new_n10748);
xor_4  g08400(new_n10747, new_n10746, new_n10749);
and_5  g08401(new_n10749, new_n3678, new_n10750);
nor_5  g08402(new_n10750, new_n10748, new_n10751);
and_5  g08403(new_n10751, new_n10744, new_n10752);
nor_5  g08404(new_n10752, new_n10743, new_n10753);
nor_5  g08405(new_n10753, new_n10741, new_n10754);
nor_5  g08406(new_n10754, new_n10740, new_n10755);
nor_5  g08407(new_n10755, new_n10738, new_n10756_1);
nor_5  g08408(new_n10756_1, new_n10737, new_n10757);
nor_5  g08409(new_n10757, new_n10735, new_n10758);
nor_5  g08410(new_n10758, new_n10734, new_n10759);
nor_5  g08411(new_n10759, new_n10732, new_n10760);
nor_5  g08412(new_n10760, new_n10731, new_n10761);
nor_5  g08413(new_n10761, new_n10729, new_n10762);
nor_5  g08414(new_n10762, new_n10728, new_n10763_1);
nor_5  g08415(new_n10763_1, new_n10725, new_n10764);
nor_5  g08416(new_n10764, new_n10724, new_n10765);
xnor_4 g08417(new_n10765, new_n10721, n1859);
xnor_4 g08418(new_n4815, new_n4792, n1860);
or_5   g08419(new_n10325, new_n10322, new_n10768);
nor_5  g08420(n21915, n15182, new_n10769);
nor_5  g08421(new_n6221, new_n6198, new_n10770);
nor_5  g08422(new_n10770, new_n10769, new_n10771);
xnor_4 g08423(n25972, n8614, new_n10772);
xnor_4 g08424(new_n10772, new_n10771, new_n10773);
and_5  g08425(new_n10773, n10250, new_n10774);
xnor_4 g08426(new_n10773, n10250, new_n10775_1);
and_5  g08427(new_n6222, n7674, new_n10776);
xnor_4 g08428(new_n6222, n7674, new_n10777);
and_5  g08429(new_n6224, n6397, new_n10778);
xnor_4 g08430(new_n6224, n6397, new_n10779);
and_5  g08431(new_n6227, n19196, new_n10780_1);
xnor_4 g08432(new_n6227, n19196, new_n10781);
nand_5 g08433(new_n6230, n23586, new_n10782);
or_5   g08434(new_n6233_1, n21226, new_n10783);
xnor_4 g08435(new_n6233_1, n21226, new_n10784);
and_5  g08436(new_n6237, n4426, new_n10785);
xnor_4 g08437(new_n6237, n4426, new_n10786);
and_5  g08438(new_n3848, new_n7878, new_n10787);
nor_5  g08439(new_n3860, new_n3851, new_n10788);
nand_5 g08440(new_n3864, n9380, new_n10789);
xor_4  g08441(new_n3860, n11192, new_n10790);
nor_5  g08442(new_n10790, new_n10789, new_n10791);
nor_5  g08443(new_n10791, new_n10788, new_n10792_1);
xnor_4 g08444(new_n3848, n20036, new_n10793);
and_5  g08445(new_n10793, new_n10792_1, new_n10794);
or_5   g08446(new_n10794, new_n10787, new_n10795);
nor_5  g08447(new_n10795, new_n10786, new_n10796);
nor_5  g08448(new_n10796, new_n10785, new_n10797);
not_10 g08449(new_n10797, new_n10798);
or_5   g08450(new_n10798, new_n10784, new_n10799);
nand_5 g08451(new_n10799, new_n10783, new_n10800);
xnor_4 g08452(new_n6230, n23586, new_n10801);
or_5   g08453(new_n10801, new_n10800, new_n10802);
and_5  g08454(new_n10802, new_n10782, new_n10803);
nor_5  g08455(new_n10803, new_n10781, new_n10804);
nor_5  g08456(new_n10804, new_n10780_1, new_n10805);
nor_5  g08457(new_n10805, new_n10779, new_n10806);
nor_5  g08458(new_n10806, new_n10778, new_n10807);
nor_5  g08459(new_n10807, new_n10777, new_n10808);
nor_5  g08460(new_n10808, new_n10776, new_n10809);
nor_5  g08461(new_n10809, new_n10775_1, new_n10810);
nor_5  g08462(new_n10810, new_n10774, new_n10811);
and_5  g08463(n25972, n8614, new_n10812);
or_5   g08464(n25972, n8614, new_n10813);
and_5  g08465(new_n10813, new_n10771, new_n10814);
nor_5  g08466(new_n10814, new_n10812, new_n10815);
nor_5  g08467(new_n10815, new_n10811, new_n10816);
nor_5  g08468(new_n10816, new_n10768, new_n10817_1);
xnor_4 g08469(new_n10816, new_n10768, new_n10818);
not_10 g08470(new_n10815, new_n10819);
xnor_4 g08471(new_n10819, new_n10811, new_n10820);
nor_5  g08472(new_n10820, new_n10326_1, new_n10821);
xnor_4 g08473(new_n10820, new_n10326_1, new_n10822);
xnor_4 g08474(new_n10320, new_n10300, new_n10823);
xor_4  g08475(new_n10809, new_n10775_1, new_n10824);
nor_5  g08476(new_n10824, new_n10823, new_n10825);
xnor_4 g08477(new_n10824, new_n10823, new_n10826);
xnor_4 g08478(new_n10318, new_n10302, new_n10827);
xor_4  g08479(new_n10807, new_n10777, new_n10828);
nor_5  g08480(new_n10828, new_n10827, new_n10829);
xnor_4 g08481(new_n10828, new_n10827, new_n10830);
xor_4  g08482(new_n10805, new_n10779, new_n10831);
nor_5  g08483(new_n10831, new_n10346, new_n10832);
xnor_4 g08484(new_n10831, new_n10346, new_n10833);
xor_4  g08485(new_n10803, new_n10781, new_n10834_1);
nor_5  g08486(new_n10834_1, new_n10348, new_n10835);
xnor_4 g08487(new_n10834_1, new_n10348, new_n10836);
not_10 g08488(new_n10353, new_n10837);
xor_4  g08489(new_n10801, new_n10800, new_n10838);
nor_5  g08490(new_n10838, new_n10837, new_n10839);
xor_4  g08491(new_n10838, new_n10353, new_n10840);
xnor_4 g08492(new_n10797, new_n10784, new_n10841);
and_5  g08493(new_n10841, new_n8666, new_n10842);
xnor_4 g08494(new_n10841, new_n8666, new_n10843);
not_10 g08495(new_n8668, new_n10844);
xor_4  g08496(new_n10795, new_n10786, new_n10845);
nor_5  g08497(new_n10845, new_n10844, new_n10846);
xor_4  g08498(new_n10845, new_n8668, new_n10847);
xor_4  g08499(new_n10793, new_n10792_1, new_n10848);
and_5  g08500(new_n10848, new_n8672, new_n10849);
xnor_4 g08501(new_n10848, new_n8672, new_n10850);
xor_4  g08502(new_n10790, new_n10789, new_n10851_1);
nor_5  g08503(new_n10851_1, new_n8676, new_n10852);
not_10 g08504(new_n6523, new_n10853);
xor_4  g08505(new_n3864, n9380, new_n10854);
nor_5  g08506(new_n10854, new_n10853, new_n10855);
xor_4  g08507(new_n10851_1, new_n8676, new_n10856);
and_5  g08508(new_n10856, new_n10855, new_n10857);
nor_5  g08509(new_n10857, new_n10852, new_n10858);
nor_5  g08510(new_n10858, new_n10850, new_n10859);
nor_5  g08511(new_n10859, new_n10849, new_n10860);
nor_5  g08512(new_n10860, new_n10847, new_n10861);
nor_5  g08513(new_n10861, new_n10846, new_n10862);
nor_5  g08514(new_n10862, new_n10843, new_n10863);
nor_5  g08515(new_n10863, new_n10842, new_n10864);
nor_5  g08516(new_n10864, new_n10840, new_n10865);
nor_5  g08517(new_n10865, new_n10839, new_n10866);
nor_5  g08518(new_n10866, new_n10836, new_n10867);
nor_5  g08519(new_n10867, new_n10835, new_n10868);
nor_5  g08520(new_n10868, new_n10833, new_n10869);
nor_5  g08521(new_n10869, new_n10832, new_n10870);
nor_5  g08522(new_n10870, new_n10830, new_n10871);
nor_5  g08523(new_n10871, new_n10829, new_n10872);
nor_5  g08524(new_n10872, new_n10826, new_n10873);
nor_5  g08525(new_n10873, new_n10825, new_n10874_1);
nor_5  g08526(new_n10874_1, new_n10822, new_n10875);
nor_5  g08527(new_n10875, new_n10821, new_n10876);
nor_5  g08528(new_n10876, new_n10818, new_n10877);
or_5   g08529(new_n10877, new_n10817_1, n1861);
or_5   g08530(n13714, n12593, new_n10879);
or_5   g08531(new_n10879, n19144, new_n10880);
or_5   g08532(new_n10880, n8309, new_n10881);
or_5   g08533(new_n10881, n19081, new_n10882);
or_5   g08534(new_n10882, n26054, new_n10883);
xor_4  g08535(new_n10883, n26318, new_n10884);
xor_4  g08536(new_n10884, new_n4933, new_n10885);
not_10 g08537(new_n4937, new_n10886);
xor_4  g08538(new_n10882, n26054, new_n10887);
nor_5  g08539(new_n10887, new_n10886, new_n10888);
xor_4  g08540(new_n10881, n19081, new_n10889);
nor_5  g08541(new_n10889, new_n4964_1, new_n10890);
xnor_4 g08542(new_n10889, new_n4964_1, new_n10891);
not_10 g08543(new_n4940, new_n10892);
xor_4  g08544(new_n10880, n8309, new_n10893);
nor_5  g08545(new_n10893, new_n10892, new_n10894);
not_10 g08546(new_n4944, new_n10895);
xor_4  g08547(new_n10879, n19144, new_n10896);
or_5   g08548(new_n10896, new_n10895, new_n10897);
xor_4  g08549(new_n10896, new_n4944, new_n10898);
and_5  g08550(new_n4950, n13714, new_n10899);
xnor_4 g08551(new_n10899, n12593, new_n10900);
nor_5  g08552(new_n10900, new_n4946, new_n10901);
not_10 g08553(n13714, new_n10902);
or_5   g08554(new_n4950, new_n10902, new_n10903);
nor_5  g08555(new_n10903, n12593, new_n10904);
nor_5  g08556(new_n10904, new_n10901, new_n10905);
not_10 g08557(new_n10905, new_n10906);
or_5   g08558(new_n10906, new_n10898, new_n10907);
and_5  g08559(new_n10907, new_n10897, new_n10908);
xor_4  g08560(new_n10893, new_n4940, new_n10909);
nor_5  g08561(new_n10909, new_n10908, new_n10910);
nor_5  g08562(new_n10910, new_n10894, new_n10911);
nor_5  g08563(new_n10911, new_n10891, new_n10912);
nor_5  g08564(new_n10912, new_n10890, new_n10913);
xor_4  g08565(new_n10887, new_n4937, new_n10914);
nor_5  g08566(new_n10914, new_n10913, new_n10915);
nor_5  g08567(new_n10915, new_n10888, new_n10916);
xnor_4 g08568(new_n10916, new_n10885, new_n10917);
or_5   g08569(new_n7799, n19228, new_n10918);
or_5   g08570(new_n10918, n20179, new_n10919);
xnor_4 g08571(new_n10919, new_n6753, new_n10920);
xnor_4 g08572(new_n10920, new_n6602, new_n10921);
xnor_4 g08573(new_n10918, new_n6756, new_n10922);
and_5  g08574(new_n10922, new_n6605, new_n10923);
xnor_4 g08575(new_n10922, new_n6605, new_n10924_1);
nor_5  g08576(new_n7800, new_n6608, new_n10925);
xnor_4 g08577(new_n7800, new_n6608, new_n10926);
nor_5  g08578(new_n7802, new_n6611_1, new_n10927);
xnor_4 g08579(new_n7802, new_n6611_1, new_n10928);
not_10 g08580(new_n6615, new_n10929);
and_5  g08581(new_n7805, new_n10929, new_n10930);
nor_5  g08582(new_n7805, new_n10929, new_n10931);
not_10 g08583(new_n7808, new_n10932);
and_5  g08584(new_n10932, new_n6619, new_n10933);
or_5   g08585(new_n6621, new_n7918, new_n10934);
xnor_4 g08586(new_n7808, new_n6619, new_n10935);
and_5  g08587(new_n10935, new_n10934, new_n10936);
or_5   g08588(new_n10936, new_n10933, new_n10937);
nor_5  g08589(new_n10937, new_n10931, new_n10938);
or_5   g08590(new_n10938, new_n10930, new_n10939);
nor_5  g08591(new_n10939, new_n10928, new_n10940);
nor_5  g08592(new_n10940, new_n10927, new_n10941);
nor_5  g08593(new_n10941, new_n10926, new_n10942);
or_5   g08594(new_n10942, new_n10925, new_n10943_1);
nor_5  g08595(new_n10943_1, new_n10924_1, new_n10944);
nor_5  g08596(new_n10944, new_n10923, new_n10945);
xor_4  g08597(new_n10945, new_n10921, new_n10946);
xnor_4 g08598(new_n10946, new_n10917, new_n10947);
xnor_4 g08599(new_n10943_1, new_n10924_1, new_n10948);
xor_4  g08600(new_n10914, new_n10913, new_n10949);
and_5  g08601(new_n10949, new_n10948, new_n10950);
xnor_4 g08602(new_n10949, new_n10948, new_n10951);
xor_4  g08603(new_n10911, new_n10891, new_n10952);
xor_4  g08604(new_n10941, new_n10926, new_n10953);
and_5  g08605(new_n10953, new_n10952, new_n10954);
xnor_4 g08606(new_n10953, new_n10952, new_n10955);
xor_4  g08607(new_n10909, new_n10908, new_n10956);
xor_4  g08608(new_n10939, new_n10928, new_n10957);
and_5  g08609(new_n10957, new_n10956, new_n10958);
xnor_4 g08610(new_n10957, new_n10956, new_n10959);
xnor_4 g08611(new_n10905, new_n10898, new_n10960);
not_10 g08612(new_n10960, new_n10961_1);
xnor_4 g08613(new_n7805, new_n6615, new_n10962);
xnor_4 g08614(new_n10962, new_n10937, new_n10963);
nor_5  g08615(new_n10963, new_n10961_1, new_n10964);
xnor_4 g08616(new_n10963, new_n10961_1, new_n10965);
xnor_4 g08617(new_n10935, new_n10934, new_n10966);
xor_4  g08618(new_n10900, new_n4946, new_n10967);
nor_5  g08619(new_n10967, new_n10966, new_n10968);
xor_4  g08620(new_n6621, n18962, new_n10969);
xor_4  g08621(new_n4950, n13714, new_n10970);
or_5   g08622(new_n10970, new_n10969, new_n10971);
xor_4  g08623(new_n10967, new_n10966, new_n10972);
and_5  g08624(new_n10972, new_n10971, new_n10973);
nor_5  g08625(new_n10973, new_n10968, new_n10974);
nor_5  g08626(new_n10974, new_n10965, new_n10975);
nor_5  g08627(new_n10975, new_n10964, new_n10976);
nor_5  g08628(new_n10976, new_n10959, new_n10977);
nor_5  g08629(new_n10977, new_n10958, new_n10978);
nor_5  g08630(new_n10978, new_n10955, new_n10979);
nor_5  g08631(new_n10979, new_n10954, new_n10980);
nor_5  g08632(new_n10980, new_n10951, new_n10981);
nor_5  g08633(new_n10981, new_n10950, new_n10982);
xnor_4 g08634(new_n10982, new_n10947, n1891);
xor_4  g08635(new_n5944, new_n5960, new_n10984);
xor_4  g08636(n20169, n1949, new_n10985);
and_5  g08637(n9323, new_n3753, new_n10986);
nor_5  g08638(n9323, new_n3753, new_n10987);
not_10 g08639(n6729, new_n10988);
and_5  g08640(n10792, new_n10988, new_n10989);
or_5   g08641(n10792, new_n10988, new_n10990);
not_10 g08642(n19922, new_n10991);
nor_5  g08643(n21687, new_n10991, new_n10992);
and_5  g08644(new_n10992, new_n10990, new_n10993);
nor_5  g08645(new_n10993, new_n10989, new_n10994);
nor_5  g08646(new_n10994, new_n10987, new_n10995);
nor_5  g08647(new_n10995, new_n10986, new_n10996);
xor_4  g08648(new_n10996, new_n10985, new_n10997);
xnor_4 g08649(new_n10997, new_n10984, new_n10998);
xor_4  g08650(new_n5941, new_n5930, new_n10999);
xnor_4 g08651(n9323, n8285, new_n11000);
xnor_4 g08652(new_n11000, new_n10994, new_n11001);
and_5  g08653(new_n11001, new_n10999, new_n11002);
xnor_4 g08654(new_n11001, new_n10999, new_n11003);
xnor_4 g08655(n21687, n19922, new_n11004);
or_5   g08656(new_n11004, new_n5967, new_n11005_1);
xor_4  g08657(n10792, n6729, new_n11006);
xnor_4 g08658(new_n11006, new_n10992, new_n11007);
and_5  g08659(new_n11007, new_n11005_1, new_n11008);
xor_4  g08660(new_n11007, new_n11005_1, new_n11009);
and_5  g08661(new_n11009, new_n5970, new_n11010);
nor_5  g08662(new_n11010, new_n11008, new_n11011_1);
nor_5  g08663(new_n11011_1, new_n11003, new_n11012);
nor_5  g08664(new_n11012, new_n11002, new_n11013);
xnor_4 g08665(new_n11013, new_n10998, n1925);
xnor_4 g08666(new_n6910, new_n6884, n1942);
xnor_4 g08667(new_n5834_1, new_n5785, n1972);
and_5  g08668(new_n7990, new_n7937_1, new_n11017);
nor_5  g08669(new_n8047, new_n7991, new_n11018);
nor_5  g08670(new_n11018, new_n11017, new_n11019);
and_5  g08671(new_n7945, new_n7204, new_n11020);
and_5  g08672(new_n7946, n12507, new_n11021);
nor_5  g08673(new_n7946, n12507, new_n11022);
nor_5  g08674(new_n7989, new_n11022, new_n11023_1);
or_5   g08675(new_n11023_1, new_n11021, new_n11024);
nor_5  g08676(new_n11024, new_n11020, new_n11025_1);
not_10 g08677(new_n11025_1, new_n11026);
nor_5  g08678(new_n11026, new_n10036, new_n11027);
and_5  g08679(new_n11027, new_n11019, new_n11028);
nand_5 g08680(new_n11026, new_n10036, new_n11029);
nor_5  g08681(new_n11029, new_n11019, new_n11030);
or_5   g08682(new_n11030, new_n11028, new_n11031);
nor_5  g08683(new_n11031, new_n9936, new_n11032);
nor_5  g08684(new_n11030, new_n11028, new_n11033);
xor_4  g08685(new_n11033, new_n9936, new_n11034);
xor_4  g08686(new_n11025_1, new_n10036, new_n11035);
xnor_4 g08687(new_n11035, new_n11019, new_n11036);
nor_5  g08688(new_n11036, new_n9936, new_n11037);
xnor_4 g08689(new_n11036, new_n9936, new_n11038);
nor_5  g08690(new_n9973, new_n8048, new_n11039);
nor_5  g08691(new_n9978, new_n8051, new_n11040);
xnor_4 g08692(new_n9978, new_n8051, new_n11041);
xnor_4 g08693(new_n8043, new_n8001, new_n11042);
nor_5  g08694(new_n9982, new_n11042, new_n11043);
xnor_4 g08695(new_n9982, new_n11042, new_n11044_1);
xnor_4 g08696(new_n8041, new_n8005, new_n11045);
nor_5  g08697(new_n9986, new_n11045, new_n11046);
xnor_4 g08698(new_n9986, new_n11045, new_n11047);
xnor_4 g08699(new_n8039, new_n8009, new_n11048);
nor_5  g08700(new_n9990, new_n11048, new_n11049);
xnor_4 g08701(new_n9990, new_n11048, new_n11050);
xnor_4 g08702(new_n8037, new_n8014, new_n11051);
nor_5  g08703(new_n9995, new_n11051, new_n11052);
xnor_4 g08704(new_n9995, new_n11051, new_n11053);
nor_5  g08705(new_n9997, new_n8070, new_n11054);
xnor_4 g08706(new_n9997, new_n8070, new_n11055);
and_5  g08707(new_n10002, new_n8074, new_n11056_1);
xnor_4 g08708(new_n10002, new_n8074, new_n11057);
nor_5  g08709(new_n10005, new_n8080, new_n11058);
nor_5  g08710(new_n11058, new_n10009_1, new_n11059);
xnor_4 g08711(new_n11058, new_n10008, new_n11060);
and_5  g08712(new_n11060, new_n8085, new_n11061);
nor_5  g08713(new_n11061, new_n11059, new_n11062);
nor_5  g08714(new_n11062, new_n11057, new_n11063_1);
nor_5  g08715(new_n11063_1, new_n11056_1, new_n11064);
nor_5  g08716(new_n11064, new_n11055, new_n11065);
nor_5  g08717(new_n11065, new_n11054, new_n11066);
nor_5  g08718(new_n11066, new_n11053, new_n11067);
nor_5  g08719(new_n11067, new_n11052, new_n11068);
nor_5  g08720(new_n11068, new_n11050, new_n11069);
nor_5  g08721(new_n11069, new_n11049, new_n11070);
nor_5  g08722(new_n11070, new_n11047, new_n11071);
nor_5  g08723(new_n11071, new_n11046, new_n11072);
nor_5  g08724(new_n11072, new_n11044_1, new_n11073);
nor_5  g08725(new_n11073, new_n11043, new_n11074);
nor_5  g08726(new_n11074, new_n11041, new_n11075);
or_5   g08727(new_n11075, new_n11040, new_n11076);
xor_4  g08728(new_n9973, new_n8048, new_n11077);
and_5  g08729(new_n11077, new_n11076, new_n11078_1);
nor_5  g08730(new_n11078_1, new_n11039, new_n11079);
nor_5  g08731(new_n11079, new_n11038, new_n11080_1);
or_5   g08732(new_n11080_1, new_n11037, new_n11081);
nor_5  g08733(new_n11081, new_n11034, new_n11082);
nor_5  g08734(new_n11082, new_n11032, n1981);
xnor_4 g08735(new_n11077, new_n11076, n2004);
not_10 g08736(n5140, new_n11085);
nor_5  g08737(n6105, new_n11085, new_n11086);
xor_4  g08738(n6105, n5140, new_n11087);
not_10 g08739(n6204, new_n11088);
nor_5  g08740(new_n11088, n3795, new_n11089);
xor_4  g08741(n6204, n3795, new_n11090);
not_10 g08742(n3349, new_n11091);
nor_5  g08743(n25464, new_n11091, new_n11092);
xor_4  g08744(n25464, n3349, new_n11093);
not_10 g08745(n1742, new_n11094_1);
nor_5  g08746(n4590, new_n11094_1, new_n11095);
xor_4  g08747(n4590, n1742, new_n11096);
not_10 g08748(n4858, new_n11097);
nor_5  g08749(n26752, new_n11097, new_n11098);
xor_4  g08750(n26752, n4858, new_n11099);
not_10 g08751(n8244, new_n11100);
or_5   g08752(new_n11100, n6513, new_n11101_1);
xor_4  g08753(n8244, n6513, new_n11102);
not_10 g08754(n9493, new_n11103_1);
or_5   g08755(new_n11103_1, n3918, new_n11104);
xor_4  g08756(n9493, n3918, new_n11105);
not_10 g08757(n15167, new_n11106);
and_5  g08758(new_n11106, n919, new_n11107);
nor_5  g08759(new_n11106, n919, new_n11108);
not_10 g08760(n21095, new_n11109);
and_5  g08761(n25316, new_n11109, new_n11110);
or_5   g08762(n25316, new_n11109, new_n11111);
not_10 g08763(n20385, new_n11112);
nor_5  g08764(new_n11112, n8656, new_n11113);
and_5  g08765(new_n11113, new_n11111, new_n11114);
nor_5  g08766(new_n11114, new_n11110, new_n11115);
nor_5  g08767(new_n11115, new_n11108, new_n11116);
nor_5  g08768(new_n11116, new_n11107, new_n11117);
not_10 g08769(new_n11117, new_n11118);
or_5   g08770(new_n11118, new_n11105, new_n11119);
and_5  g08771(new_n11119, new_n11104, new_n11120_1);
or_5   g08772(new_n11120_1, new_n11102, new_n11121_1);
and_5  g08773(new_n11121_1, new_n11101_1, new_n11122);
nor_5  g08774(new_n11122, new_n11099, new_n11123);
nor_5  g08775(new_n11123, new_n11098, new_n11124);
nor_5  g08776(new_n11124, new_n11096, new_n11125);
nor_5  g08777(new_n11125, new_n11095, new_n11126);
nor_5  g08778(new_n11126, new_n11093, new_n11127_1);
nor_5  g08779(new_n11127_1, new_n11092, new_n11128);
nor_5  g08780(new_n11128, new_n11090, new_n11129);
nor_5  g08781(new_n11129, new_n11089, new_n11130);
nor_5  g08782(new_n11130, new_n11087, new_n11131);
nor_5  g08783(new_n11131, new_n11086, new_n11132_1);
not_10 g08784(n10018, new_n11133);
and_5  g08785(new_n5665, new_n11133, new_n11134_1);
nor_5  g08786(new_n5665, new_n11133, new_n11135);
xnor_4 g08787(new_n5663, n1288, new_n11136);
nor_5  g08788(new_n11136, n2184, new_n11137);
xnor_4 g08789(new_n11136, n2184, new_n11138_1);
xnor_4 g08790(new_n5662, n1752, new_n11139);
nor_5  g08791(new_n11139, n3541, new_n11140);
xnor_4 g08792(new_n11139, n3541, new_n11141);
not_10 g08793(n16818, new_n11142);
and_5  g08794(new_n5675, new_n11142, new_n11143);
xor_4  g08795(new_n5675, n16818, new_n11144);
and_5  g08796(new_n3763, new_n5876, new_n11145);
xor_4  g08797(new_n3763, n1269, new_n11146);
and_5  g08798(new_n3765, new_n5877, new_n11147);
xor_4  g08799(new_n3765, n14576, new_n11148);
or_5   g08800(new_n3767, new_n5892, new_n11149);
xor_4  g08801(new_n3767, n2985, new_n11150);
and_5  g08802(new_n3770, new_n5878, new_n11151);
not_10 g08803(new_n3773, new_n11152);
and_5  g08804(new_n11152, n15652, new_n11153);
not_10 g08805(n4939, new_n11154);
or_5   g08806(n19922, new_n11154, new_n11155);
xor_4  g08807(new_n3773, n15652, new_n11156);
nor_5  g08808(new_n11156, new_n11155, new_n11157);
nor_5  g08809(new_n11157, new_n11153, new_n11158);
xnor_4 g08810(new_n3770, n5605, new_n11159);
and_5  g08811(new_n11159, new_n11158, new_n11160);
nor_5  g08812(new_n11160, new_n11151, new_n11161);
not_10 g08813(new_n11161, new_n11162);
or_5   g08814(new_n11162, new_n11150, new_n11163);
nand_5 g08815(new_n11163, new_n11149, new_n11164);
nor_5  g08816(new_n11164, new_n11148, new_n11165);
nor_5  g08817(new_n11165, new_n11147, new_n11166);
nor_5  g08818(new_n11166, new_n11146, new_n11167);
nor_5  g08819(new_n11167, new_n11145, new_n11168);
nor_5  g08820(new_n11168, new_n11144, new_n11169);
nor_5  g08821(new_n11169, new_n11143, new_n11170);
nor_5  g08822(new_n11170, new_n11141, new_n11171);
nor_5  g08823(new_n11171, new_n11140, new_n11172);
nor_5  g08824(new_n11172, new_n11138_1, new_n11173);
nor_5  g08825(new_n11173, new_n11137, new_n11174);
nor_5  g08826(new_n11174, new_n11135, new_n11175);
xor_4  g08827(new_n11175, new_n5667, new_n11176);
nor_5  g08828(new_n11176, new_n11134_1, new_n11177);
xnor_4 g08829(new_n11177, new_n5660, new_n11178);
xnor_4 g08830(new_n5665, n10018, new_n11179);
xnor_4 g08831(new_n11179, new_n11174, new_n11180);
nor_5  g08832(new_n11180, new_n5692, new_n11181);
xnor_4 g08833(new_n11180, new_n5692, new_n11182_1);
xor_4  g08834(new_n11172, new_n11138_1, new_n11183);
nor_5  g08835(new_n11183, new_n5697, new_n11184_1);
xnor_4 g08836(new_n11183, new_n5697, new_n11185);
xor_4  g08837(new_n11170, new_n11141, new_n11186);
nor_5  g08838(new_n11186, new_n5701, new_n11187);
xnor_4 g08839(new_n11186, new_n5701, new_n11188);
xor_4  g08840(new_n11168, new_n11144, new_n11189);
nor_5  g08841(new_n11189, new_n5704_1, new_n11190);
xor_4  g08842(new_n11166, new_n11146, new_n11191);
nor_5  g08843(new_n11191, new_n5707, new_n11192_1);
xnor_4 g08844(new_n11191, new_n5707, new_n11193);
xor_4  g08845(new_n11164, new_n11148, new_n11194);
nor_5  g08846(new_n11194, new_n5710, new_n11195);
xnor_4 g08847(new_n11194, new_n5710, new_n11196);
xor_4  g08848(new_n5646, new_n5637, new_n11197);
xnor_4 g08849(new_n11161, new_n11150, new_n11198);
and_5  g08850(new_n11198, new_n11197, new_n11199);
not_10 g08851(new_n5713, new_n11200);
xor_4  g08852(new_n11159, new_n11158, new_n11201_1);
and_5  g08853(new_n11201_1, new_n11200, new_n11202);
xnor_4 g08854(new_n11201_1, new_n11200, new_n11203);
xor_4  g08855(new_n11156, new_n11155, new_n11204);
nor_5  g08856(new_n11204, new_n5716, new_n11205);
not_10 g08857(new_n5718, new_n11206);
xnor_4 g08858(n19922, n4939, new_n11207);
or_5   g08859(new_n11207, new_n11206, new_n11208);
xnor_4 g08860(new_n11204, new_n5716, new_n11209);
nor_5  g08861(new_n11209, new_n11208, new_n11210);
nor_5  g08862(new_n11210, new_n11205, new_n11211);
nor_5  g08863(new_n11211, new_n11203, new_n11212);
or_5   g08864(new_n11212, new_n11202, new_n11213);
xnor_4 g08865(new_n11198, new_n11197, new_n11214);
nor_5  g08866(new_n11214, new_n11213, new_n11215);
nor_5  g08867(new_n11215, new_n11199, new_n11216);
nor_5  g08868(new_n11216, new_n11196, new_n11217);
nor_5  g08869(new_n11217, new_n11195, new_n11218);
nor_5  g08870(new_n11218, new_n11193, new_n11219);
nor_5  g08871(new_n11219, new_n11192_1, new_n11220_1);
xnor_4 g08872(new_n11189, new_n5704_1, new_n11221);
nor_5  g08873(new_n11221, new_n11220_1, new_n11222);
nor_5  g08874(new_n11222, new_n11190, new_n11223_1);
nor_5  g08875(new_n11223_1, new_n11188, new_n11224);
nor_5  g08876(new_n11224, new_n11187, new_n11225);
nor_5  g08877(new_n11225, new_n11185, new_n11226);
nor_5  g08878(new_n11226, new_n11184_1, new_n11227);
nor_5  g08879(new_n11227, new_n11182_1, new_n11228);
or_5   g08880(new_n11228, new_n11181, new_n11229);
xnor_4 g08881(new_n11229, new_n11178, new_n11230);
nor_5  g08882(new_n11230, new_n11132_1, new_n11231);
xnor_4 g08883(new_n11230, new_n11132_1, new_n11232);
xnor_4 g08884(new_n11130, new_n11087, new_n11233);
xor_4  g08885(new_n11227, new_n11182_1, new_n11234_1);
and_5  g08886(new_n11234_1, new_n11233, new_n11235);
xnor_4 g08887(new_n11234_1, new_n11233, new_n11236);
xnor_4 g08888(new_n11128, new_n11090, new_n11237);
xor_4  g08889(new_n11225, new_n11185, new_n11238);
and_5  g08890(new_n11238, new_n11237, new_n11239);
xnor_4 g08891(new_n11238, new_n11237, new_n11240);
xnor_4 g08892(new_n11126, new_n11093, new_n11241);
xor_4  g08893(new_n11223_1, new_n11188, new_n11242);
and_5  g08894(new_n11242, new_n11241, new_n11243);
xnor_4 g08895(new_n11242, new_n11241, new_n11244);
xnor_4 g08896(new_n11124, new_n11096, new_n11245_1);
xor_4  g08897(new_n11221, new_n11220_1, new_n11246);
and_5  g08898(new_n11246, new_n11245_1, new_n11247);
xnor_4 g08899(new_n11246, new_n11245_1, new_n11248);
xnor_4 g08900(new_n11122, new_n11099, new_n11249);
xor_4  g08901(new_n11218, new_n11193, new_n11250);
and_5  g08902(new_n11250, new_n11249, new_n11251);
xnor_4 g08903(new_n11250, new_n11249, new_n11252);
xnor_4 g08904(new_n11120_1, new_n11102, new_n11253);
xor_4  g08905(new_n11216, new_n11196, new_n11254);
and_5  g08906(new_n11254, new_n11253, new_n11255);
xnor_4 g08907(new_n11254, new_n11253, new_n11256);
xor_4  g08908(new_n11117, new_n11105, new_n11257);
xor_4  g08909(new_n11214, new_n11213, new_n11258);
and_5  g08910(new_n11258, new_n11257, new_n11259);
xnor_4 g08911(new_n11258, new_n11257, new_n11260);
xnor_4 g08912(new_n11211, new_n11203, new_n11261_1);
xnor_4 g08913(n15167, n919, new_n11262);
xnor_4 g08914(new_n11262, new_n11115, new_n11263);
and_5  g08915(new_n11263, new_n11261_1, new_n11264);
xnor_4 g08916(new_n11263, new_n11261_1, new_n11265);
xor_4  g08917(new_n11207, new_n5718, new_n11266_1);
xnor_4 g08918(n20385, n8656, new_n11267);
nor_5  g08919(new_n11267, new_n11266_1, new_n11268);
xor_4  g08920(n25316, n21095, new_n11269);
xnor_4 g08921(new_n11269, new_n11113, new_n11270);
not_10 g08922(new_n11270, new_n11271);
nor_5  g08923(new_n11271, new_n11268, new_n11272);
xnor_4 g08924(new_n11209, new_n11208, new_n11273_1);
xnor_4 g08925(new_n11270, new_n11268, new_n11274);
and_5  g08926(new_n11274, new_n11273_1, new_n11275_1);
nor_5  g08927(new_n11275_1, new_n11272, new_n11276);
nor_5  g08928(new_n11276, new_n11265, new_n11277);
nor_5  g08929(new_n11277, new_n11264, new_n11278);
nor_5  g08930(new_n11278, new_n11260, new_n11279);
nor_5  g08931(new_n11279, new_n11259, new_n11280);
nor_5  g08932(new_n11280, new_n11256, new_n11281);
nor_5  g08933(new_n11281, new_n11255, new_n11282);
nor_5  g08934(new_n11282, new_n11252, new_n11283);
nor_5  g08935(new_n11283, new_n11251, new_n11284);
nor_5  g08936(new_n11284, new_n11248, new_n11285);
nor_5  g08937(new_n11285, new_n11247, new_n11286);
nor_5  g08938(new_n11286, new_n11244, new_n11287);
nor_5  g08939(new_n11287, new_n11243, new_n11288);
nor_5  g08940(new_n11288, new_n11240, new_n11289);
nor_5  g08941(new_n11289, new_n11239, new_n11290_1);
nor_5  g08942(new_n11290_1, new_n11236, new_n11291);
nor_5  g08943(new_n11291, new_n11235, new_n11292);
nor_5  g08944(new_n11292, new_n11232, new_n11293);
or_5   g08945(new_n11293, new_n11231, new_n11294);
not_10 g08946(new_n5660, new_n11295);
nor_5  g08947(new_n11177, new_n11295, new_n11296);
and_5  g08948(new_n11175, new_n5667, new_n11297);
and_5  g08949(new_n11177, new_n11295, new_n11298);
nor_5  g08950(new_n11229, new_n11298, new_n11299);
or_5   g08951(new_n11299, new_n11297, new_n11300);
nor_5  g08952(new_n11300, new_n11296, new_n11301);
and_5  g08953(new_n11301, new_n11294, n2007);
xnor_4 g08954(new_n8088, new_n8078, n2061);
not_10 g08955(new_n6450, new_n11304);
xnor_4 g08956(new_n10212, new_n11304, new_n11305);
not_10 g08957(new_n6454, new_n11306);
nor_5  g08958(new_n10216, new_n11306, new_n11307);
xnor_4 g08959(new_n10216, new_n11306, new_n11308);
and_5  g08960(new_n10221, new_n6458, new_n11309);
not_10 g08961(new_n4314, new_n11310);
and_5  g08962(new_n6462, new_n11310, new_n11311);
xor_4  g08963(new_n6462, new_n4314, new_n11312);
and_5  g08964(new_n6466, new_n4340_1, new_n11313_1);
xnor_4 g08965(new_n6466, new_n4340_1, new_n11314);
nor_5  g08966(new_n6469, new_n4344, new_n11315);
nor_5  g08967(new_n6476_1, new_n4349, new_n11316);
xnor_4 g08968(new_n6472, new_n4349, new_n11317);
not_10 g08969(new_n4356, new_n11318);
nor_5  g08970(new_n6478, new_n4360, new_n11319);
and_5  g08971(new_n11319, new_n11318, new_n11320);
xor_4  g08972(new_n11319, new_n4356, new_n11321);
nor_5  g08973(new_n11321, new_n6484, new_n11322);
nor_5  g08974(new_n11322, new_n11320, new_n11323);
and_5  g08975(new_n11323, new_n11317, new_n11324);
nor_5  g08976(new_n11324, new_n11316, new_n11325_1);
xnor_4 g08977(new_n6469, new_n4344, new_n11326_1);
nor_5  g08978(new_n11326_1, new_n11325_1, new_n11327);
nor_5  g08979(new_n11327, new_n11315, new_n11328);
nor_5  g08980(new_n11328, new_n11314, new_n11329);
nor_5  g08981(new_n11329, new_n11313_1, new_n11330_1);
nor_5  g08982(new_n11330_1, new_n11312, new_n11331);
nor_5  g08983(new_n11331, new_n11311, new_n11332);
xor_4  g08984(new_n10220, new_n6458, new_n11333);
nor_5  g08985(new_n11333, new_n11332, new_n11334);
nor_5  g08986(new_n11334, new_n11309, new_n11335);
nor_5  g08987(new_n11335, new_n11308, new_n11336);
nor_5  g08988(new_n11336, new_n11307, new_n11337);
xnor_4 g08989(new_n11337, new_n11305, n2092);
xnor_4 g08990(n22253, n10650, new_n11339);
nor_5  g08991(n12900, n1255, new_n11340);
xnor_4 g08992(n12900, n1255, new_n11341);
nor_5  g08993(n20411, n9512, new_n11342);
xnor_4 g08994(n20411, n9512, new_n11343);
nor_5  g08995(n17069, n16608, new_n11344);
xnor_4 g08996(n17069, n16608, new_n11345);
nor_5  g08997(n21735, n15918, new_n11346);
xnor_4 g08998(n21735, n15918, new_n11347_1);
nor_5  g08999(n24085, n17784, new_n11348_1);
xnor_4 g09000(n24085, n17784, new_n11349);
nor_5  g09001(n14323, n14071, new_n11350);
xnor_4 g09002(n14323, n14071, new_n11351);
nor_5  g09003(n2886, n1738, new_n11352_1);
xnor_4 g09004(n2886, n1738, new_n11353);
nor_5  g09005(n12152, n1040, new_n11354);
and_5  g09006(n19107, n9090, new_n11355);
xnor_4 g09007(n12152, n1040, new_n11356_1);
nor_5  g09008(new_n11356_1, new_n11355, new_n11357);
nor_5  g09009(new_n11357, new_n11354, new_n11358);
nor_5  g09010(new_n11358, new_n11353, new_n11359);
nor_5  g09011(new_n11359, new_n11352_1, new_n11360);
nor_5  g09012(new_n11360, new_n11351, new_n11361);
nor_5  g09013(new_n11361, new_n11350, new_n11362);
nor_5  g09014(new_n11362, new_n11349, new_n11363);
nor_5  g09015(new_n11363, new_n11348_1, new_n11364);
nor_5  g09016(new_n11364, new_n11347_1, new_n11365);
nor_5  g09017(new_n11365, new_n11346, new_n11366);
nor_5  g09018(new_n11366, new_n11345, new_n11367);
nor_5  g09019(new_n11367, new_n11344, new_n11368);
nor_5  g09020(new_n11368, new_n11343, new_n11369);
nor_5  g09021(new_n11369, new_n11342, new_n11370);
nor_5  g09022(new_n11370, new_n11341, new_n11371);
nor_5  g09023(new_n11371, new_n11340, new_n11372);
xor_4  g09024(new_n11372, new_n11339, new_n11373);
and_5  g09025(new_n11373, n2272, new_n11374);
xnor_4 g09026(new_n11373, n2272, new_n11375_1);
xor_4  g09027(new_n11370, new_n11341, new_n11376);
and_5  g09028(new_n11376, n25331, new_n11377);
xnor_4 g09029(new_n11376, n25331, new_n11378);
xor_4  g09030(new_n11368, new_n11343, new_n11379_1);
and_5  g09031(new_n11379_1, n18483, new_n11380);
xnor_4 g09032(new_n11379_1, n18483, new_n11381);
xor_4  g09033(new_n11366, new_n11345, new_n11382);
and_5  g09034(new_n11382, n21934, new_n11383);
xnor_4 g09035(new_n11382, n21934, new_n11384);
xor_4  g09036(new_n11364, new_n11347_1, new_n11385);
and_5  g09037(new_n11385, n18901, new_n11386_1);
xnor_4 g09038(new_n11385, n18901, new_n11387);
xor_4  g09039(new_n11362, new_n11349, new_n11388);
and_5  g09040(new_n11388, n4376, new_n11389);
xnor_4 g09041(new_n11388, n4376, new_n11390);
xor_4  g09042(new_n11360, new_n11351, new_n11391_1);
and_5  g09043(new_n11391_1, n14570, new_n11392);
xnor_4 g09044(new_n11391_1, n14570, new_n11393);
xor_4  g09045(new_n11358, new_n11353, new_n11394);
and_5  g09046(new_n11394, n23775, new_n11395);
xnor_4 g09047(new_n11394, n23775, new_n11396);
xnor_4 g09048(n19107, n9090, new_n11397);
and_5  g09049(new_n11397, n11479, new_n11398_1);
nor_5  g09050(new_n11398_1, n8259, new_n11399);
xor_4  g09051(new_n11356_1, new_n11355, new_n11400);
xnor_4 g09052(new_n11398_1, n8259, new_n11401);
nor_5  g09053(new_n11401, new_n11400, new_n11402);
or_5   g09054(new_n11402, new_n11399, new_n11403_1);
nor_5  g09055(new_n11403_1, new_n11396, new_n11404);
nor_5  g09056(new_n11404, new_n11395, new_n11405);
nor_5  g09057(new_n11405, new_n11393, new_n11406);
nor_5  g09058(new_n11406, new_n11392, new_n11407);
nor_5  g09059(new_n11407, new_n11390, new_n11408);
nor_5  g09060(new_n11408, new_n11389, new_n11409);
nor_5  g09061(new_n11409, new_n11387, new_n11410);
nor_5  g09062(new_n11410, new_n11386_1, new_n11411);
nor_5  g09063(new_n11411, new_n11384, new_n11412);
nor_5  g09064(new_n11412, new_n11383, new_n11413);
nor_5  g09065(new_n11413, new_n11381, new_n11414);
nor_5  g09066(new_n11414, new_n11380, new_n11415);
nor_5  g09067(new_n11415, new_n11378, new_n11416);
nor_5  g09068(new_n11416, new_n11377, new_n11417);
nor_5  g09069(new_n11417, new_n11375_1, new_n11418);
nor_5  g09070(new_n11418, new_n11374, new_n11419_1);
nor_5  g09071(n22253, n10650, new_n11420);
nor_5  g09072(new_n11372, new_n11339, new_n11421);
nor_5  g09073(new_n11421, new_n11420, new_n11422);
nor_5  g09074(new_n11422, new_n11419_1, new_n11423);
nor_5  g09075(n7876, n4964, new_n11424_1);
not_10 g09076(new_n11424_1, new_n11425);
or_5   g09077(new_n11425, n26553, new_n11426);
or_5   g09078(new_n11426, n342, new_n11427);
or_5   g09079(new_n11427, n26107, new_n11428);
or_5   g09080(new_n11428, n22597, new_n11429);
or_5   g09081(new_n11429, n19327, new_n11430);
or_5   g09082(new_n11430, n26224, new_n11431);
or_5   g09083(new_n11431, n18496, new_n11432);
nor_5  g09084(new_n11432, n9934, new_n11433);
xnor_4 g09085(new_n11432, n9934, new_n11434);
or_5   g09086(n18409, n5704, new_n11435);
or_5   g09087(new_n11435, n13708, new_n11436);
or_5   g09088(new_n11436, n19911, new_n11437);
or_5   g09089(new_n11437, n2731, new_n11438);
or_5   g09090(new_n11438, n18907, new_n11439_1);
or_5   g09091(new_n11439_1, n22332, new_n11440);
or_5   g09092(new_n11440, n4256, new_n11441);
xor_4  g09093(new_n11441, n21287, new_n11442);
nor_5  g09094(new_n11442, n12861, new_n11443);
xnor_4 g09095(new_n11442, n12861, new_n11444);
xor_4  g09096(new_n11440, n4256, new_n11445);
nor_5  g09097(new_n11445, n13333, new_n11446);
xnor_4 g09098(new_n11445, n13333, new_n11447);
xor_4  g09099(new_n11439_1, n22332, new_n11448);
nor_5  g09100(new_n11448, n2210, new_n11449);
xnor_4 g09101(new_n11448, n2210, new_n11450);
xor_4  g09102(new_n11438, n18907, new_n11451);
nor_5  g09103(new_n11451, n20604, new_n11452);
xnor_4 g09104(new_n11451, n20604, new_n11453);
xor_4  g09105(new_n11437, n2731, new_n11454);
nor_5  g09106(new_n11454, n16158, new_n11455_1);
xnor_4 g09107(new_n11454, n16158, new_n11456);
xor_4  g09108(new_n11436, n19911, new_n11457);
nor_5  g09109(new_n11457, n5752, new_n11458);
xor_4  g09110(new_n11435, n13708, new_n11459);
nor_5  g09111(new_n11459, n18171, new_n11460);
xnor_4 g09112(new_n11459, n18171, new_n11461);
xor_4  g09113(n18409, n5704, new_n11462_1);
nor_5  g09114(new_n11462_1, n25073, new_n11463);
nand_5 g09115(n22309, n5704, new_n11464);
xor_4  g09116(new_n11462_1, n25073, new_n11465);
and_5  g09117(new_n11465, new_n11464, new_n11466);
nor_5  g09118(new_n11466, new_n11463, new_n11467);
nor_5  g09119(new_n11467, new_n11461, new_n11468);
nor_5  g09120(new_n11468, new_n11460, new_n11469);
xnor_4 g09121(new_n11457, n5752, new_n11470_1);
nor_5  g09122(new_n11470_1, new_n11469, new_n11471);
nor_5  g09123(new_n11471, new_n11458, new_n11472_1);
nor_5  g09124(new_n11472_1, new_n11456, new_n11473_1);
nor_5  g09125(new_n11473_1, new_n11455_1, new_n11474);
nor_5  g09126(new_n11474, new_n11453, new_n11475);
nor_5  g09127(new_n11475, new_n11452, new_n11476);
nor_5  g09128(new_n11476, new_n11450, new_n11477);
nor_5  g09129(new_n11477, new_n11449, new_n11478);
nor_5  g09130(new_n11478, new_n11447, new_n11479_1);
nor_5  g09131(new_n11479_1, new_n11446, new_n11480);
nor_5  g09132(new_n11480, new_n11444, new_n11481_1);
nor_5  g09133(new_n11481_1, new_n11443, new_n11482);
nor_5  g09134(new_n11441, n21287, new_n11483);
xnor_4 g09135(new_n11483, n26986, new_n11484);
xor_4  g09136(new_n11484, n8305, new_n11485);
xnor_4 g09137(new_n11485, new_n11482, new_n11486_1);
nor_5  g09138(new_n11486_1, new_n11434, new_n11487);
xnor_4 g09139(new_n11486_1, new_n11434, new_n11488);
xnor_4 g09140(new_n11431, n18496, new_n11489);
xor_4  g09141(new_n11480, new_n11444, new_n11490);
nor_5  g09142(new_n11490, new_n11489, new_n11491);
xnor_4 g09143(new_n11490, new_n11489, new_n11492);
xnor_4 g09144(new_n11430, n26224, new_n11493);
xor_4  g09145(new_n11478, new_n11447, new_n11494);
nor_5  g09146(new_n11494, new_n11493, new_n11495);
xnor_4 g09147(new_n11494, new_n11493, new_n11496_1);
xnor_4 g09148(new_n11429, n19327, new_n11497);
xor_4  g09149(new_n11476, new_n11450, new_n11498);
nor_5  g09150(new_n11498, new_n11497, new_n11499);
xnor_4 g09151(new_n11498, new_n11497, new_n11500);
xnor_4 g09152(new_n11428, n22597, new_n11501);
xor_4  g09153(new_n11474, new_n11453, new_n11502);
nor_5  g09154(new_n11502, new_n11501, new_n11503_1);
xnor_4 g09155(new_n11502, new_n11501, new_n11504);
xnor_4 g09156(new_n11427, n26107, new_n11505);
xor_4  g09157(new_n11472_1, new_n11456, new_n11506_1);
nor_5  g09158(new_n11506_1, new_n11505, new_n11507);
xnor_4 g09159(new_n11506_1, new_n11505, new_n11508);
xnor_4 g09160(new_n11426, n342, new_n11509);
xor_4  g09161(new_n11470_1, new_n11469, new_n11510);
nor_5  g09162(new_n11510, new_n11509, new_n11511);
xnor_4 g09163(new_n11510, new_n11509, new_n11512);
xor_4  g09164(new_n11467, new_n11461, new_n11513);
xor_4  g09165(new_n11424_1, n26553, new_n11514);
nor_5  g09166(new_n11514, new_n11513, new_n11515_1);
xnor_4 g09167(new_n11514, new_n11513, new_n11516);
xnor_4 g09168(n7876, n4964, new_n11517);
xor_4  g09169(new_n11465, new_n11464, new_n11518);
nor_5  g09170(new_n11518, new_n11517, new_n11519);
xor_4  g09171(n22309, n5704, new_n11520);
and_5  g09172(new_n11520, n7876, new_n11521);
xor_4  g09173(new_n11518, new_n11517, new_n11522);
and_5  g09174(new_n11522, new_n11521, new_n11523);
nor_5  g09175(new_n11523, new_n11519, new_n11524);
nor_5  g09176(new_n11524, new_n11516, new_n11525);
nor_5  g09177(new_n11525, new_n11515_1, new_n11526);
nor_5  g09178(new_n11526, new_n11512, new_n11527);
nor_5  g09179(new_n11527, new_n11511, new_n11528);
nor_5  g09180(new_n11528, new_n11508, new_n11529);
nor_5  g09181(new_n11529, new_n11507, new_n11530);
nor_5  g09182(new_n11530, new_n11504, new_n11531);
nor_5  g09183(new_n11531, new_n11503_1, new_n11532);
nor_5  g09184(new_n11532, new_n11500, new_n11533);
nor_5  g09185(new_n11533, new_n11499, new_n11534);
nor_5  g09186(new_n11534, new_n11496_1, new_n11535);
nor_5  g09187(new_n11535, new_n11495, new_n11536);
nor_5  g09188(new_n11536, new_n11492, new_n11537);
nor_5  g09189(new_n11537, new_n11491, new_n11538_1);
nor_5  g09190(new_n11538_1, new_n11488, new_n11539);
or_5   g09191(new_n11539, new_n11487, new_n11540);
nor_5  g09192(new_n11540, new_n11433, new_n11541);
not_10 g09193(new_n11541, new_n11542);
and_5  g09194(new_n11483, new_n6505, new_n11543);
nor_5  g09195(new_n11484, n8305, new_n11544);
and_5  g09196(new_n11484, n8305, new_n11545);
nor_5  g09197(new_n11545, new_n11482, new_n11546);
nor_5  g09198(new_n11546, new_n11544, new_n11547);
nor_5  g09199(new_n11547, new_n11543, new_n11548_1);
or_5   g09200(new_n11548_1, new_n11542, new_n11549);
xor_4  g09201(new_n11549, new_n11423, new_n11550);
xor_4  g09202(new_n11422, new_n11419_1, new_n11551);
xnor_4 g09203(new_n11548_1, new_n11541, new_n11552);
and_5  g09204(new_n11552, new_n11551, new_n11553);
xnor_4 g09205(new_n11552, new_n11551, new_n11554);
xnor_4 g09206(new_n11417, new_n11375_1, new_n11555);
xor_4  g09207(new_n11538_1, new_n11488, new_n11556);
nor_5  g09208(new_n11556, new_n11555, new_n11557);
xnor_4 g09209(new_n11556, new_n11555, new_n11558);
xnor_4 g09210(new_n11415, new_n11378, new_n11559);
xor_4  g09211(new_n11536, new_n11492, new_n11560);
nor_5  g09212(new_n11560, new_n11559, new_n11561);
xnor_4 g09213(new_n11560, new_n11559, new_n11562);
xnor_4 g09214(new_n11413, new_n11381, new_n11563);
xor_4  g09215(new_n11534, new_n11496_1, new_n11564_1);
nor_5  g09216(new_n11564_1, new_n11563, new_n11565);
xnor_4 g09217(new_n11564_1, new_n11563, new_n11566_1);
xnor_4 g09218(new_n11411, new_n11384, new_n11567);
xor_4  g09219(new_n11532, new_n11500, new_n11568);
nor_5  g09220(new_n11568, new_n11567, new_n11569);
xnor_4 g09221(new_n11568, new_n11567, new_n11570);
xnor_4 g09222(new_n11409, new_n11387, new_n11571);
xor_4  g09223(new_n11530, new_n11504, new_n11572);
nor_5  g09224(new_n11572, new_n11571, new_n11573);
xnor_4 g09225(new_n11572, new_n11571, new_n11574);
xnor_4 g09226(new_n11407, new_n11390, new_n11575);
xor_4  g09227(new_n11528, new_n11508, new_n11576);
nor_5  g09228(new_n11576, new_n11575, new_n11577);
xnor_4 g09229(new_n11576, new_n11575, new_n11578);
xnor_4 g09230(new_n11405, new_n11393, new_n11579_1);
xor_4  g09231(new_n11526, new_n11512, new_n11580_1);
nor_5  g09232(new_n11580_1, new_n11579_1, new_n11581);
xnor_4 g09233(new_n11580_1, new_n11579_1, new_n11582);
xnor_4 g09234(new_n11403_1, new_n11396, new_n11583);
xor_4  g09235(new_n11524, new_n11516, new_n11584);
nor_5  g09236(new_n11584, new_n11583, new_n11585);
xor_4  g09237(new_n11584, new_n11583, new_n11586);
xnor_4 g09238(new_n11522, new_n11521, new_n11587);
xnor_4 g09239(new_n11401, new_n11400, new_n11588);
nor_5  g09240(new_n11588, new_n11587, new_n11589);
xnor_4 g09241(new_n11397, n11479, new_n11590);
xnor_4 g09242(n22309, n5704, new_n11591_1);
xnor_4 g09243(new_n11591_1, n7876, new_n11592);
nand_5 g09244(new_n11592, new_n11590, new_n11593);
xnor_4 g09245(new_n11588, new_n11587, new_n11594);
nor_5  g09246(new_n11594, new_n11593, new_n11595);
nor_5  g09247(new_n11595, new_n11589, new_n11596);
and_5  g09248(new_n11596, new_n11586, new_n11597);
nor_5  g09249(new_n11597, new_n11585, new_n11598);
nor_5  g09250(new_n11598, new_n11582, new_n11599);
nor_5  g09251(new_n11599, new_n11581, new_n11600);
nor_5  g09252(new_n11600, new_n11578, new_n11601);
nor_5  g09253(new_n11601, new_n11577, new_n11602);
nor_5  g09254(new_n11602, new_n11574, new_n11603);
nor_5  g09255(new_n11603, new_n11573, new_n11604);
nor_5  g09256(new_n11604, new_n11570, new_n11605);
nor_5  g09257(new_n11605, new_n11569, new_n11606);
nor_5  g09258(new_n11606, new_n11566_1, new_n11607_1);
nor_5  g09259(new_n11607_1, new_n11565, new_n11608);
nor_5  g09260(new_n11608, new_n11562, new_n11609);
nor_5  g09261(new_n11609, new_n11561, new_n11610);
nor_5  g09262(new_n11610, new_n11558, new_n11611);
nor_5  g09263(new_n11611, new_n11557, new_n11612);
nor_5  g09264(new_n11612, new_n11554, new_n11613);
nor_5  g09265(new_n11613, new_n11553, new_n11614);
xnor_4 g09266(new_n11614, new_n11550, n2095);
xnor_4 g09267(new_n10266, new_n10265, n2105);
xnor_4 g09268(n23166, n11898, new_n11617);
and_5  g09269(n19941, n10577, new_n11618);
or_5   g09270(n19941, n10577, new_n11619);
nor_5  g09271(n6381, n1099, new_n11620);
nor_5  g09272(new_n9525, new_n9510, new_n11621);
nor_5  g09273(new_n11621, new_n11620, new_n11622);
and_5  g09274(new_n11622, new_n11619, new_n11623);
or_5   g09275(new_n11623, new_n11618, new_n11624);
xnor_4 g09276(new_n11624, new_n11617, new_n11625);
xnor_4 g09277(new_n11625, n8827, new_n11626);
xnor_4 g09278(n19941, n10577, new_n11627);
xnor_4 g09279(new_n11627, new_n11622, new_n11628);
nand_5 g09280(new_n11628, n18035, new_n11629);
xnor_4 g09281(new_n11628, n18035, new_n11630_1);
nor_5  g09282(new_n9526, n5077, new_n11631);
nor_5  g09283(new_n9547, new_n9527, new_n11632);
or_5   g09284(new_n11632, new_n11631, new_n11633);
or_5   g09285(new_n11633, new_n11630_1, new_n11634);
and_5  g09286(new_n11634, new_n11629, new_n11635);
xor_4  g09287(new_n11635, new_n11626, new_n11636);
xor_4  g09288(new_n11636, new_n5570, new_n11637);
not_10 g09289(new_n5572, new_n11638);
xor_4  g09290(new_n11633, new_n11630_1, new_n11639);
and_5  g09291(new_n11639, new_n11638, new_n11640);
xor_4  g09292(new_n11639, new_n5572, new_n11641);
nor_5  g09293(new_n9548, new_n5577, new_n11642);
xnor_4 g09294(new_n9548, new_n5577, new_n11643);
not_10 g09295(new_n5581, new_n11644);
and_5  g09296(new_n9551, new_n11644, new_n11645);
xor_4  g09297(new_n9551, new_n5581, new_n11646);
nor_5  g09298(new_n9555, new_n5585, new_n11647_1);
xnor_4 g09299(new_n9555, new_n5585, new_n11648);
nor_5  g09300(new_n9560, new_n5589, new_n11649);
xor_4  g09301(new_n9559, new_n5589, new_n11650);
nor_5  g09302(new_n9564, new_n5593_1, new_n11651);
xor_4  g09303(new_n7712, new_n5593_1, new_n11652);
nor_5  g09304(new_n7693_1, new_n5597, new_n11653);
xnor_4 g09305(new_n7693_1, new_n5597, new_n11654);
not_10 g09306(new_n5601, new_n11655);
nor_5  g09307(new_n7696, new_n11655, new_n11656);
nor_5  g09308(new_n7699, new_n5330_1, new_n11657);
xnor_4 g09309(new_n7696, new_n5601, new_n11658);
and_5  g09310(new_n11658, new_n11657, new_n11659);
nor_5  g09311(new_n11659, new_n11656, new_n11660);
nor_5  g09312(new_n11660, new_n11654, new_n11661);
nor_5  g09313(new_n11661, new_n11653, new_n11662);
nor_5  g09314(new_n11662, new_n11652, new_n11663);
nor_5  g09315(new_n11663, new_n11651, new_n11664);
nor_5  g09316(new_n11664, new_n11650, new_n11665);
nor_5  g09317(new_n11665, new_n11649, new_n11666);
nor_5  g09318(new_n11666, new_n11648, new_n11667_1);
nor_5  g09319(new_n11667_1, new_n11647_1, new_n11668);
nor_5  g09320(new_n11668, new_n11646, new_n11669);
nor_5  g09321(new_n11669, new_n11645, new_n11670);
nor_5  g09322(new_n11670, new_n11643, new_n11671);
nor_5  g09323(new_n11671, new_n11642, new_n11672);
nor_5  g09324(new_n11672, new_n11641, new_n11673);
nor_5  g09325(new_n11673, new_n11640, new_n11674_1);
xnor_4 g09326(new_n11674_1, new_n11637, n2122);
xnor_4 g09327(new_n2755, new_n2733, n2147);
xnor_4 g09328(new_n9482, new_n9447, n2209);
xor_4  g09329(new_n5312, new_n5209, n2214);
not_10 g09330(new_n3912, new_n11679);
xnor_4 g09331(new_n10056, new_n11679, new_n11680);
nor_5  g09332(new_n10058, new_n3982, new_n11681);
xor_4  g09333(new_n10058, new_n3982, new_n11682_1);
nor_5  g09334(new_n10061, new_n3987, new_n11683);
xnor_4 g09335(new_n10061, new_n3987, new_n11684);
not_10 g09336(new_n3994, new_n11685);
nor_5  g09337(new_n10067, new_n11685, new_n11686);
or_5   g09338(new_n10064, new_n3996, new_n11687);
xnor_4 g09339(new_n10067, new_n3994, new_n11688);
and_5  g09340(new_n11688, new_n11687, new_n11689);
or_5   g09341(new_n11689, new_n11686, new_n11690);
nor_5  g09342(new_n11690, new_n11684, new_n11691);
nor_5  g09343(new_n11691, new_n11683, new_n11692);
and_5  g09344(new_n11692, new_n11682_1, new_n11693);
nor_5  g09345(new_n11693, new_n11681, new_n11694);
xnor_4 g09346(new_n11694, new_n11680, n2238);
xor_4  g09347(new_n10077, new_n10076, n2327);
xnor_4 g09348(new_n5296, new_n5267, n2343);
xnor_4 g09349(new_n9534, n13453, new_n11698);
and_5  g09350(new_n5996, n7421, new_n11699);
nor_5  g09351(new_n6010, new_n5997, new_n11700);
nor_5  g09352(new_n11700, new_n11699, new_n11701);
xnor_4 g09353(new_n11701, new_n11698, new_n11702);
xnor_4 g09354(n20923, n16524, new_n11703);
nor_5  g09355(n18157, n11056, new_n11704);
nor_5  g09356(new_n6021, new_n6012_1, new_n11705);
nor_5  g09357(new_n11705, new_n11704, new_n11706);
xnor_4 g09358(new_n11706, new_n11703, new_n11707);
xnor_4 g09359(new_n11707, n3785, new_n11708);
nor_5  g09360(new_n6022_1, n20250, new_n11709);
nor_5  g09361(new_n6035, new_n6023, new_n11710_1);
nor_5  g09362(new_n11710_1, new_n11709, new_n11711);
xnor_4 g09363(new_n11711, new_n11708, new_n11712_1);
xnor_4 g09364(new_n11712_1, new_n11702, new_n11713);
not_10 g09365(new_n6036, new_n11714);
nor_5  g09366(new_n11714, new_n6011, new_n11715);
and_5  g09367(new_n6053, new_n6037, new_n11716);
nor_5  g09368(new_n11716, new_n11715, new_n11717);
xnor_4 g09369(new_n11717, new_n11713, n2361);
xor_4  g09370(new_n3498, new_n3497, n2363);
xnor_4 g09371(new_n4254, new_n4225, n2374);
xnor_4 g09372(n7305, n1204, new_n11721);
nor_5  g09373(n25872, n19618, new_n11722);
nor_5  g09374(new_n5361, new_n5356, new_n11723);
nor_5  g09375(new_n11723, new_n11722, new_n11724_1);
xor_4  g09376(new_n11724_1, new_n11721, new_n11725);
and_5  g09377(new_n11725, new_n4500, new_n11726);
xor_4  g09378(new_n11725, new_n4499, new_n11727);
nor_5  g09379(new_n5362, new_n4504, new_n11728);
nor_5  g09380(new_n5370, new_n5363, new_n11729);
or_5   g09381(new_n11729, new_n11728, new_n11730);
nor_5  g09382(new_n11730, new_n11727, new_n11731);
or_5   g09383(new_n11731, new_n11726, new_n11732);
xnor_4 g09384(n20826, n626, new_n11733);
nor_5  g09385(n7305, n1204, new_n11734);
nor_5  g09386(new_n11724_1, new_n11721, new_n11735);
nor_5  g09387(new_n11735, new_n11734, new_n11736_1);
xor_4  g09388(new_n11736_1, new_n11733, new_n11737);
xor_4  g09389(new_n11737, new_n11732, new_n11738);
xnor_4 g09390(new_n11738, new_n4496, new_n11739);
xnor_4 g09391(new_n11739, new_n3557, new_n11740);
xor_4  g09392(new_n11730, new_n11727, new_n11741_1);
nor_5  g09393(new_n11741_1, new_n3561_1, new_n11742);
and_5  g09394(new_n5371, new_n3564, new_n11743);
nor_5  g09395(new_n5380, new_n5372, new_n11744);
nor_5  g09396(new_n11744, new_n11743, new_n11745);
xnor_4 g09397(new_n11741_1, new_n3561_1, new_n11746);
nor_5  g09398(new_n11746, new_n11745, new_n11747);
nor_5  g09399(new_n11747, new_n11742, new_n11748);
xor_4  g09400(new_n11748, new_n11740, n2388);
xnor_4 g09401(n7335, n2160, new_n11750);
nor_5  g09402(n10763, n5696, new_n11751);
nor_5  g09403(new_n4925_1, new_n4896, new_n11752);
nor_5  g09404(new_n11752, new_n11751, new_n11753);
xor_4  g09405(new_n11753, new_n11750, new_n11754);
xnor_4 g09406(n11220, n3425, new_n11755);
nor_5  g09407(n22379, n9967, new_n11756);
nor_5  g09408(new_n4894, new_n4865, new_n11757);
nor_5  g09409(new_n11757, new_n11756, new_n11758);
xnor_4 g09410(new_n11758, new_n11755, new_n11759);
xnor_4 g09411(new_n11759, new_n11754, new_n11760);
nor_5  g09412(new_n4926, new_n4895, new_n11761);
nor_5  g09413(new_n4974, new_n4927, new_n11762);
nor_5  g09414(new_n11762, new_n11761, new_n11763);
xnor_4 g09415(new_n11763, new_n11760, new_n11764);
or_5   g09416(new_n4825, n337, new_n11765);
xor_4  g09417(new_n11765, n7593, new_n11766);
xor_4  g09418(new_n11766, n5025, new_n11767);
nor_5  g09419(new_n4826, n6485, new_n11768);
nor_5  g09420(new_n4863, new_n4827, new_n11769);
nor_5  g09421(new_n11769, new_n11768, new_n11770_1);
xnor_4 g09422(new_n11770_1, new_n11767, new_n11771_1);
xnor_4 g09423(new_n11771_1, new_n11764, new_n11772);
and_5  g09424(new_n4975, new_n4864, new_n11773);
nor_5  g09425(new_n5022, new_n4976, new_n11774);
nor_5  g09426(new_n11774, new_n11773, new_n11775_1);
xor_4  g09427(new_n11775_1, new_n11772, n2440);
xnor_4 g09428(new_n10400, new_n10385_1, n2444);
xor_4  g09429(new_n4697, new_n3112, n2513);
xnor_4 g09430(new_n5456, n14323, new_n11779);
and_5  g09431(new_n5461, n2886, new_n11780);
xnor_4 g09432(new_n5461, n2886, new_n11781);
and_5  g09433(new_n5471, n1040, new_n11782);
and_5  g09434(n20658, n9090, new_n11783);
xor_4  g09435(new_n5471, n1040, new_n11784);
and_5  g09436(new_n11784, new_n11783, new_n11785);
nor_5  g09437(new_n11785, new_n11782, new_n11786);
nor_5  g09438(new_n11786, new_n11781, new_n11787);
nor_5  g09439(new_n11787, new_n11780, new_n11788);
xor_4  g09440(new_n11788, new_n11779, new_n11789);
xnor_4 g09441(new_n11789, n12562, new_n11790);
xor_4  g09442(new_n11786, new_n11781, new_n11791);
nor_5  g09443(new_n11791, n7949, new_n11792);
xnor_4 g09444(new_n11791, n7949, new_n11793);
and_5  g09445(new_n9814, n14575, new_n11794);
nor_5  g09446(new_n11794, n24374, new_n11795);
xor_4  g09447(new_n11784, new_n11783, new_n11796);
xnor_4 g09448(new_n11794, n24374, new_n11797);
nor_5  g09449(new_n11797, new_n11796, new_n11798);
nor_5  g09450(new_n11798, new_n11795, new_n11799);
nor_5  g09451(new_n11799, new_n11793, new_n11800);
or_5   g09452(new_n11800, new_n11792, new_n11801);
xor_4  g09453(new_n11801, new_n11790, new_n11802);
xnor_4 g09454(new_n11802, new_n11580_1, new_n11803);
not_10 g09455(new_n11584, new_n11804);
xor_4  g09456(new_n11799, new_n11793, new_n11805);
and_5  g09457(new_n11805, new_n11804, new_n11806);
xor_4  g09458(new_n11805, new_n11584, new_n11807);
xor_4  g09459(new_n11797, new_n11796, new_n11808);
and_5  g09460(new_n11808, new_n11587, new_n11809);
xor_4  g09461(new_n9814, n14575, new_n11810);
nand_5 g09462(new_n11810, new_n11592, new_n11811);
xor_4  g09463(new_n11808, new_n11587, new_n11812);
and_5  g09464(new_n11812, new_n11811, new_n11813);
nor_5  g09465(new_n11813, new_n11809, new_n11814);
nor_5  g09466(new_n11814, new_n11807, new_n11815);
nor_5  g09467(new_n11815, new_n11806, new_n11816);
xnor_4 g09468(new_n11816, new_n11803, n2515);
xnor_4 g09469(new_n9806, new_n9778_1, n2533);
nor_5  g09470(n26986, new_n3073, new_n11819);
xor_4  g09471(n26986, n3425, new_n11820);
nor_5  g09472(n21287, new_n3054, new_n11821);
xor_4  g09473(n21287, n9967, new_n11822);
nor_5  g09474(new_n3055, n4256, new_n11823);
xor_4  g09475(n20946, n4256, new_n11824);
nor_5  g09476(n22332, new_n3056, new_n11825);
xor_4  g09477(n22332, n7751, new_n11826);
nor_5  g09478(new_n3057, n18907, new_n11827);
xor_4  g09479(n26823, n18907, new_n11828);
nor_5  g09480(new_n3058, n2731, new_n11829);
nor_5  g09481(new_n7651, new_n7637, new_n11830);
nor_5  g09482(new_n11830, new_n11829, new_n11831);
nor_5  g09483(new_n11831, new_n11828, new_n11832);
nor_5  g09484(new_n11832, new_n11827, new_n11833);
nor_5  g09485(new_n11833, new_n11826, new_n11834);
nor_5  g09486(new_n11834, new_n11825, new_n11835);
nor_5  g09487(new_n11835, new_n11824, new_n11836);
nor_5  g09488(new_n11836, new_n11823, new_n11837_1);
nor_5  g09489(new_n11837_1, new_n11822, new_n11838);
nor_5  g09490(new_n11838, new_n11821, new_n11839);
nor_5  g09491(new_n11839, new_n11820, new_n11840);
nor_5  g09492(new_n11840, new_n11819, new_n11841_1);
not_10 g09493(new_n6444, new_n11842_1);
not_10 g09494(new_n6390, new_n11843_1);
not_10 g09495(new_n6394, new_n11844);
or_5   g09496(new_n6401, new_n4729, new_n11845);
or_5   g09497(new_n6397_1, new_n11845, new_n11846);
or_5   g09498(new_n11846, new_n11844, new_n11847);
or_5   g09499(new_n11847, new_n11843_1, new_n11848);
nor_5  g09500(new_n11848, new_n11842_1, new_n11849);
and_5  g09501(new_n11849, new_n6512, new_n11850);
nor_5  g09502(new_n11849, new_n6514_1, new_n11851);
nor_5  g09503(new_n11851, new_n11850, new_n11852);
nor_5  g09504(new_n11852, new_n3051, new_n11853);
not_10 g09505(new_n3001, new_n11854);
xnor_4 g09506(new_n11848, new_n6444, new_n11855);
nor_5  g09507(new_n11855, new_n11854, new_n11856);
xnor_4 g09508(new_n11855, new_n11854, new_n11857);
not_10 g09509(new_n3004, new_n11858);
xnor_4 g09510(new_n11847, new_n6390, new_n11859);
nor_5  g09511(new_n11859, new_n11858, new_n11860);
xnor_4 g09512(new_n11859, new_n11858, new_n11861);
not_10 g09513(new_n3007, new_n11862);
xnor_4 g09514(new_n11846, new_n6394, new_n11863);
nor_5  g09515(new_n11863, new_n11862, new_n11864);
xnor_4 g09516(new_n11863, new_n11862, new_n11865);
not_10 g09517(new_n3010_1, new_n11866);
xor_4  g09518(new_n6397_1, new_n11845, new_n11867);
nor_5  g09519(new_n11867, new_n11866, new_n11868);
xnor_4 g09520(new_n11867, new_n11866, new_n11869);
nor_5  g09521(new_n4735, new_n4703, new_n11870);
nor_5  g09522(new_n4765, new_n4736, new_n11871);
nor_5  g09523(new_n11871, new_n11870, new_n11872);
nor_5  g09524(new_n11872, new_n11869, new_n11873);
nor_5  g09525(new_n11873, new_n11868, new_n11874);
nor_5  g09526(new_n11874, new_n11865, new_n11875);
nor_5  g09527(new_n11875, new_n11864, new_n11876);
nor_5  g09528(new_n11876, new_n11861, new_n11877);
nor_5  g09529(new_n11877, new_n11860, new_n11878);
nor_5  g09530(new_n11878, new_n11857, new_n11879);
nor_5  g09531(new_n11879, new_n11856, new_n11880);
and_5  g09532(new_n11852, new_n3051, new_n11881);
nor_5  g09533(new_n11881, new_n11880, new_n11882);
nor_5  g09534(new_n11882, new_n11853, new_n11883);
nor_5  g09535(new_n11883, new_n11850, new_n11884);
xnor_4 g09536(new_n11884, new_n11841_1, new_n11885);
xnor_4 g09537(new_n11852, new_n3051, new_n11886);
xnor_4 g09538(new_n11886, new_n11880, new_n11887);
nor_5  g09539(new_n11887, new_n11841_1, new_n11888);
xnor_4 g09540(new_n11887, new_n11841_1, new_n11889);
xnor_4 g09541(new_n11839, new_n11820, new_n11890);
xor_4  g09542(new_n11878, new_n11857, new_n11891);
and_5  g09543(new_n11891, new_n11890, new_n11892);
xnor_4 g09544(new_n11891, new_n11890, new_n11893);
xnor_4 g09545(new_n11837_1, new_n11822, new_n11894);
xor_4  g09546(new_n11876, new_n11861, new_n11895);
and_5  g09547(new_n11895, new_n11894, new_n11896);
xnor_4 g09548(new_n11895, new_n11894, new_n11897);
xnor_4 g09549(new_n11835, new_n11824, new_n11898_1);
xor_4  g09550(new_n11874, new_n11865, new_n11899);
and_5  g09551(new_n11899, new_n11898_1, new_n11900);
xnor_4 g09552(new_n11899, new_n11898_1, new_n11901);
xor_4  g09553(new_n11833, new_n11826, new_n11902);
xnor_4 g09554(new_n11872, new_n11869, new_n11903);
nor_5  g09555(new_n11903, new_n11902, new_n11904);
xor_4  g09556(new_n11903, new_n11902, new_n11905_1);
xor_4  g09557(new_n11831, new_n11828, new_n11906);
and_5  g09558(new_n11906, new_n4766_1, new_n11907);
xnor_4 g09559(new_n11906, new_n4766_1, new_n11908);
and_5  g09560(new_n7652, new_n7636, new_n11909);
nor_5  g09561(new_n7672, new_n7653, new_n11910);
nor_5  g09562(new_n11910, new_n11909, new_n11911);
nor_5  g09563(new_n11911, new_n11908, new_n11912);
nor_5  g09564(new_n11912, new_n11907, new_n11913);
and_5  g09565(new_n11913, new_n11905_1, new_n11914);
nor_5  g09566(new_n11914, new_n11904, new_n11915);
nor_5  g09567(new_n11915, new_n11901, new_n11916);
nor_5  g09568(new_n11916, new_n11900, new_n11917);
nor_5  g09569(new_n11917, new_n11897, new_n11918);
nor_5  g09570(new_n11918, new_n11896, new_n11919);
nor_5  g09571(new_n11919, new_n11893, new_n11920);
nor_5  g09572(new_n11920, new_n11892, new_n11921);
nor_5  g09573(new_n11921, new_n11889, new_n11922);
nor_5  g09574(new_n11922, new_n11888, new_n11923);
xnor_4 g09575(new_n11923, new_n11885, n2535);
or_5   g09576(n20259, n3925, new_n11925);
or_5   g09577(new_n11925, n25872, new_n11926_1);
or_5   g09578(new_n11926_1, n7305, new_n11927);
or_5   g09579(new_n11927, n20826, new_n11928);
xor_4  g09580(new_n11928, n22198, new_n11929);
xnor_4 g09581(new_n11929, n21674, new_n11930);
xor_4  g09582(new_n11927, n20826, new_n11931);
nor_5  g09583(new_n11931, n17251, new_n11932);
xnor_4 g09584(new_n11931, n17251, new_n11933);
xor_4  g09585(new_n11926_1, n7305, new_n11934);
nor_5  g09586(new_n11934, n14790, new_n11935);
xor_4  g09587(new_n11925, n25872, new_n11936);
nor_5  g09588(new_n11936, n10096, new_n11937);
xnor_4 g09589(new_n11936, n10096, new_n11938);
xor_4  g09590(n20259, n3925, new_n11939);
nor_5  g09591(new_n11939, n16994, new_n11940);
and_5  g09592(n9246, n3925, new_n11941);
xnor_4 g09593(new_n11939, n16994, new_n11942);
nor_5  g09594(new_n11942, new_n11941, new_n11943);
nor_5  g09595(new_n11943, new_n11940, new_n11944);
nor_5  g09596(new_n11944, new_n11938, new_n11945);
nor_5  g09597(new_n11945, new_n11937, new_n11946);
xnor_4 g09598(new_n11934, n14790, new_n11947);
nor_5  g09599(new_n11947, new_n11946, new_n11948);
nor_5  g09600(new_n11948, new_n11935, new_n11949);
nor_5  g09601(new_n11949, new_n11933, new_n11950);
nor_5  g09602(new_n11950, new_n11932, new_n11951);
xnor_4 g09603(new_n11951, new_n11930, new_n11952);
xnor_4 g09604(new_n11952, new_n7037, new_n11953);
xnor_4 g09605(new_n11949, new_n11933, new_n11954);
nor_5  g09606(new_n11954, new_n7041, new_n11955);
xnor_4 g09607(new_n11954, new_n7041, new_n11956);
xnor_4 g09608(new_n11947, new_n11946, new_n11957);
nor_5  g09609(new_n11957, new_n7045, new_n11958);
xnor_4 g09610(new_n11957, new_n7045, new_n11959);
xor_4  g09611(new_n11944, new_n11938, new_n11960);
nor_5  g09612(new_n11960, new_n7051, new_n11961);
xnor_4 g09613(new_n11960, new_n7051, new_n11962);
xor_4  g09614(new_n11942, new_n11941, new_n11963);
nor_5  g09615(new_n11963, new_n7057_1, new_n11964);
or_5   g09616(new_n8836, new_n7060, new_n11965_1);
xnor_4 g09617(new_n11963, new_n7057_1, new_n11966);
nor_5  g09618(new_n11966, new_n11965_1, new_n11967);
nor_5  g09619(new_n11967, new_n11964, new_n11968);
nor_5  g09620(new_n11968, new_n11962, new_n11969);
or_5   g09621(new_n11969, new_n11961, new_n11970);
nor_5  g09622(new_n11970, new_n11959, new_n11971);
nor_5  g09623(new_n11971, new_n11958, new_n11972);
nor_5  g09624(new_n11972, new_n11956, new_n11973);
nor_5  g09625(new_n11973, new_n11955, new_n11974);
xor_4  g09626(new_n11974, new_n11953, new_n11975);
xor_4  g09627(n1163, n329, new_n11976);
not_10 g09628(n24170, new_n11977);
nor_5  g09629(new_n11977, n18537, new_n11978);
xor_4  g09630(n24170, n18537, new_n11979);
not_10 g09631(n2409, new_n11980_1);
nor_5  g09632(n7057, new_n11980_1, new_n11981);
xor_4  g09633(n7057, n2409, new_n11982);
nor_5  g09634(n8869, new_n8602, new_n11983);
and_5  g09635(n8869, new_n8602, new_n11984);
nor_5  g09636(new_n4660, n10372, new_n11985);
nor_5  g09637(new_n8606, n7428, new_n11986);
nand_5 g09638(new_n4660, n10372, new_n11987);
and_5  g09639(new_n11987, new_n11986, new_n11988);
nor_5  g09640(new_n11988, new_n11985, new_n11989);
nor_5  g09641(new_n11989, new_n11984, new_n11990);
or_5   g09642(new_n11990, new_n11983, new_n11991);
nor_5  g09643(new_n11991, new_n11982, new_n11992);
nor_5  g09644(new_n11992, new_n11981, new_n11993);
nor_5  g09645(new_n11993, new_n11979, new_n11994);
nor_5  g09646(new_n11994, new_n11978, new_n11995);
xor_4  g09647(new_n11995, new_n11976, new_n11996);
xor_4  g09648(new_n11996, new_n11975, new_n11997);
xnor_4 g09649(new_n11993, new_n11979, new_n11998);
xor_4  g09650(new_n11972, new_n11956, new_n11999);
and_5  g09651(new_n11999, new_n11998, new_n12000_1);
xnor_4 g09652(new_n11999, new_n11998, new_n12001);
xnor_4 g09653(new_n11970, new_n11959, new_n12002);
xor_4  g09654(new_n11991, new_n11982, new_n12003_1);
nor_5  g09655(new_n12003_1, new_n12002, new_n12004);
xnor_4 g09656(new_n12003_1, new_n12002, new_n12005);
xor_4  g09657(new_n11968, new_n11962, new_n12006);
not_10 g09658(new_n12006, new_n12007);
xnor_4 g09659(n8869, n8381, new_n12008);
xnor_4 g09660(new_n12008, new_n11989, new_n12009);
and_5  g09661(new_n12009, new_n12007, new_n12010);
xor_4  g09662(new_n12009, new_n12006, new_n12011_1);
or_5   g09663(new_n8838, new_n8837, new_n12012);
xor_4  g09664(n20235, n10372, new_n12013);
xnor_4 g09665(new_n12013, new_n11986, new_n12014);
and_5  g09666(new_n12014, new_n12012, new_n12015);
xnor_4 g09667(new_n11966, new_n11965_1, new_n12016);
xor_4  g09668(new_n12014, new_n12012, new_n12017);
and_5  g09669(new_n12017, new_n12016, new_n12018);
nor_5  g09670(new_n12018, new_n12015, new_n12019);
nor_5  g09671(new_n12019, new_n12011_1, new_n12020);
nor_5  g09672(new_n12020, new_n12010, new_n12021);
nor_5  g09673(new_n12021, new_n12005, new_n12022);
nor_5  g09674(new_n12022, new_n12004, new_n12023);
nor_5  g09675(new_n12023, new_n12001, new_n12024);
nor_5  g09676(new_n12024, new_n12000_1, new_n12025);
xnor_4 g09677(new_n12025, new_n11997, n2537);
xnor_4 g09678(new_n9954, new_n2880, new_n12027);
and_5  g09679(new_n3916, new_n2884, new_n12028);
xnor_4 g09680(new_n3916, new_n2884, new_n12029);
nor_5  g09681(new_n3918_1, new_n2888, new_n12030);
xnor_4 g09682(new_n3918_1, new_n2888, new_n12031);
and_5  g09683(new_n3921, new_n2892, new_n12032);
xor_4  g09684(new_n3921, new_n2892, new_n12033);
nor_5  g09685(new_n3924, new_n2896, new_n12034);
nor_5  g09686(new_n2899, n1152, new_n12035);
xor_4  g09687(new_n3924, new_n2896, new_n12036);
and_5  g09688(new_n12036, new_n12035, new_n12037);
nor_5  g09689(new_n12037, new_n12034, new_n12038);
and_5  g09690(new_n12038, new_n12033, new_n12039);
or_5   g09691(new_n12039, new_n12032, new_n12040);
nor_5  g09692(new_n12040, new_n12031, new_n12041);
or_5   g09693(new_n12041, new_n12030, new_n12042);
nor_5  g09694(new_n12042, new_n12029, new_n12043);
nor_5  g09695(new_n12043, new_n12028, new_n12044);
xor_4  g09696(new_n12044, new_n12027, new_n12045);
xnor_4 g09697(new_n12045, new_n10353, new_n12046);
xor_4  g09698(new_n12042, new_n12029, new_n12047);
nor_5  g09699(new_n12047, new_n8666, new_n12048);
xnor_4 g09700(new_n12047, new_n8666, new_n12049);
xor_4  g09701(new_n12040, new_n12031, new_n12050);
and_5  g09702(new_n12050, new_n10844, new_n12051);
xnor_4 g09703(new_n12050, new_n8668, new_n12052);
xor_4  g09704(new_n12038, new_n12033, new_n12053);
and_5  g09705(new_n12053, new_n8672, new_n12054);
xnor_4 g09706(new_n12053, new_n8672, new_n12055);
xor_4  g09707(new_n12036, new_n12035, new_n12056);
and_5  g09708(new_n12056, new_n8676, new_n12057);
xor_4  g09709(new_n2899, n1152, new_n12058);
or_5   g09710(new_n12058, new_n10853, new_n12059);
xor_4  g09711(new_n12056, new_n8676, new_n12060);
and_5  g09712(new_n12060, new_n12059, new_n12061);
or_5   g09713(new_n12061, new_n12057, new_n12062);
nor_5  g09714(new_n12062, new_n12055, new_n12063);
nor_5  g09715(new_n12063, new_n12054, new_n12064);
and_5  g09716(new_n12064, new_n12052, new_n12065);
nor_5  g09717(new_n12065, new_n12051, new_n12066);
nor_5  g09718(new_n12066, new_n12049, new_n12067);
nor_5  g09719(new_n12067, new_n12048, new_n12068);
xnor_4 g09720(new_n12068, new_n12046, n2553);
xnor_4 g09721(new_n10755, new_n10738, n2555);
xnor_4 g09722(new_n9664, n12892, new_n12071);
nor_5  g09723(new_n12071, new_n9073, new_n12072_1);
nand_5 g09724(new_n9664, n12892, new_n12073);
xor_4  g09725(new_n9667, n12209, new_n12074);
xor_4  g09726(new_n12074, new_n12073, new_n12075);
xnor_4 g09727(new_n12075, new_n9070, new_n12076);
xnor_4 g09728(new_n12076, new_n12072_1, n2560);
nor_5  g09729(n26180, n10650, new_n12078);
xnor_4 g09730(n26180, n10650, new_n12079);
nor_5  g09731(n24004, n12900, new_n12080);
xnor_4 g09732(n24004, n12900, new_n12081);
nor_5  g09733(n20411, n12871, new_n12082);
xnor_4 g09734(n20411, n12871, new_n12083);
nor_5  g09735(n23304, n17069, new_n12084);
xnor_4 g09736(n23304, n17069, new_n12085);
nor_5  g09737(n19361, n15918, new_n12086);
xnor_4 g09738(n19361, n15918, new_n12087);
nor_5  g09739(n17784, n1437, new_n12088);
xnor_4 g09740(n17784, n1437, new_n12089);
nor_5  g09741(n14323, n4722, new_n12090);
xnor_4 g09742(n14323, n4722, new_n12091);
nor_5  g09743(n14633, n2886, new_n12092);
xnor_4 g09744(n14633, n2886, new_n12093);
nor_5  g09745(n8721, n1040, new_n12094);
and_5  g09746(n18578, n9090, new_n12095);
xnor_4 g09747(n8721, n1040, new_n12096);
nor_5  g09748(new_n12096, new_n12095, new_n12097);
nor_5  g09749(new_n12097, new_n12094, new_n12098);
nor_5  g09750(new_n12098, new_n12093, new_n12099);
nor_5  g09751(new_n12099, new_n12092, new_n12100);
nor_5  g09752(new_n12100, new_n12091, new_n12101);
nor_5  g09753(new_n12101, new_n12090, new_n12102);
nor_5  g09754(new_n12102, new_n12089, new_n12103);
nor_5  g09755(new_n12103, new_n12088, new_n12104);
nor_5  g09756(new_n12104, new_n12087, new_n12105);
nor_5  g09757(new_n12105, new_n12086, new_n12106);
nor_5  g09758(new_n12106, new_n12085, new_n12107);
nor_5  g09759(new_n12107, new_n12084, new_n12108);
nor_5  g09760(new_n12108, new_n12083, new_n12109);
nor_5  g09761(new_n12109, new_n12082, new_n12110);
nor_5  g09762(new_n12110, new_n12081, new_n12111);
nor_5  g09763(new_n12111, new_n12080, new_n12112);
nor_5  g09764(new_n12112, new_n12079, new_n12113_1);
nor_5  g09765(new_n12113_1, new_n12078, new_n12114);
nor_5  g09766(n9259, n6456, new_n12115);
nor_5  g09767(new_n5429, new_n5396, new_n12116);
nor_5  g09768(new_n12116, new_n12115, new_n12117);
not_10 g09769(new_n12117, new_n12118);
nor_5  g09770(new_n12118, new_n12114, new_n12119);
xor_4  g09771(new_n12117, new_n12114, new_n12120);
not_10 g09772(new_n5430_1, new_n12121_1);
xor_4  g09773(new_n12112, new_n12079, new_n12122);
and_5  g09774(new_n12122, new_n12121_1, new_n12123);
xor_4  g09775(new_n12122, new_n5430_1, new_n12124);
xor_4  g09776(new_n12110, new_n12081, new_n12125);
and_5  g09777(new_n12125, new_n5434, new_n12126);
xnor_4 g09778(new_n12125, new_n5434, new_n12127);
not_10 g09779(new_n5439_1, new_n12128);
xor_4  g09780(new_n12108, new_n12083, new_n12129);
and_5  g09781(new_n12129, new_n12128, new_n12130);
xor_4  g09782(new_n12129, new_n5439_1, new_n12131_1);
not_10 g09783(new_n5444, new_n12132);
xor_4  g09784(new_n12106, new_n12085, new_n12133);
and_5  g09785(new_n12133, new_n12132, new_n12134);
xor_4  g09786(new_n12133, new_n5444, new_n12135);
not_10 g09787(new_n5448, new_n12136);
xor_4  g09788(new_n12104, new_n12087, new_n12137);
nand_5 g09789(new_n12137, new_n12136, new_n12138);
xor_4  g09790(new_n12137, new_n5448, new_n12139);
not_10 g09791(new_n5453, new_n12140);
xor_4  g09792(new_n12102, new_n12089, new_n12141);
nor_5  g09793(new_n12141, new_n12140, new_n12142);
xor_4  g09794(new_n12141, new_n5453, new_n12143);
xor_4  g09795(new_n12100, new_n12091, new_n12144);
nor_5  g09796(new_n12144, new_n5459, new_n12145);
xor_4  g09797(new_n12144, new_n5457, new_n12146_1);
not_10 g09798(new_n5462, new_n12147);
xor_4  g09799(new_n12098, new_n12093, new_n12148);
nor_5  g09800(new_n12148, new_n12147, new_n12149);
xor_4  g09801(new_n12148, new_n5462, new_n12150);
xor_4  g09802(n18578, n9090, new_n12151);
or_5   g09803(new_n12151, new_n5466, new_n12152_1);
and_5  g09804(new_n12152_1, new_n5469, new_n12153_1);
xor_4  g09805(new_n12096, new_n12095, new_n12154);
nor_5  g09806(new_n12152_1, new_n5413, new_n12155);
or_5   g09807(new_n12155, new_n12153_1, new_n12156);
nor_5  g09808(new_n12156, new_n12154, new_n12157_1);
nor_5  g09809(new_n12157_1, new_n12153_1, new_n12158_1);
nor_5  g09810(new_n12158_1, new_n12150, new_n12159);
nor_5  g09811(new_n12159, new_n12149, new_n12160);
nor_5  g09812(new_n12160, new_n12146_1, new_n12161_1);
nor_5  g09813(new_n12161_1, new_n12145, new_n12162);
nor_5  g09814(new_n12162, new_n12143, new_n12163);
nor_5  g09815(new_n12163, new_n12142, new_n12164);
not_10 g09816(new_n12164, new_n12165);
or_5   g09817(new_n12165, new_n12139, new_n12166);
and_5  g09818(new_n12166, new_n12138, new_n12167);
nor_5  g09819(new_n12167, new_n12135, new_n12168);
nor_5  g09820(new_n12168, new_n12134, new_n12169);
nor_5  g09821(new_n12169, new_n12131_1, new_n12170);
nor_5  g09822(new_n12170, new_n12130, new_n12171);
nor_5  g09823(new_n12171, new_n12127, new_n12172);
nor_5  g09824(new_n12172, new_n12126, new_n12173);
nor_5  g09825(new_n12173, new_n12124, new_n12174);
nor_5  g09826(new_n12174, new_n12123, new_n12175);
nor_5  g09827(new_n12175, new_n12120, new_n12176);
or_5   g09828(new_n12176, new_n12119, new_n12177);
xor_4  g09829(new_n12175, new_n12120, new_n12178);
not_10 g09830(n2743, new_n12179_1);
nor_5  g09831(n3506, new_n12179_1, new_n12180);
nor_5  g09832(new_n3395, new_n3352, new_n12181);
nor_5  g09833(new_n12181, new_n12180, new_n12182);
and_5  g09834(new_n12182, new_n12178, new_n12183);
xnor_4 g09835(new_n12182, new_n12178, new_n12184);
xor_4  g09836(new_n12173, new_n12124, new_n12185);
and_5  g09837(new_n12185, new_n3396, new_n12186);
xnor_4 g09838(new_n12185, new_n3396, new_n12187);
xor_4  g09839(new_n12171, new_n12127, new_n12188);
and_5  g09840(new_n12188, new_n3408, new_n12189);
xnor_4 g09841(new_n12188, new_n3408, new_n12190);
xor_4  g09842(new_n12169, new_n12131_1, new_n12191);
and_5  g09843(new_n12191, new_n3412, new_n12192_1);
xnor_4 g09844(new_n12191, new_n3412, new_n12193);
xor_4  g09845(new_n12167, new_n12135, new_n12194);
and_5  g09846(new_n12194, new_n3416, new_n12195);
xnor_4 g09847(new_n12194, new_n3416, new_n12196);
xnor_4 g09848(new_n12164, new_n12139, new_n12197);
and_5  g09849(new_n12197, new_n3420, new_n12198);
xnor_4 g09850(new_n12197, new_n3420, new_n12199);
xnor_4 g09851(new_n3385, new_n3367, new_n12200);
xor_4  g09852(new_n12162, new_n12143, new_n12201);
nor_5  g09853(new_n12201, new_n12200, new_n12202);
xnor_4 g09854(new_n12201, new_n12200, new_n12203);
not_10 g09855(new_n3429, new_n12204);
xor_4  g09856(new_n12160, new_n12146_1, new_n12205);
nor_5  g09857(new_n12205, new_n12204, new_n12206);
xnor_4 g09858(new_n12205, new_n12204, new_n12207);
xor_4  g09859(new_n12158_1, new_n12150, new_n12208);
nor_5  g09860(new_n12208, new_n3433, new_n12209_1);
xnor_4 g09861(new_n12208, new_n3433, new_n12210);
xor_4  g09862(new_n12156, new_n12154, new_n12211);
nor_5  g09863(new_n12211, new_n3439, new_n12212);
xor_4  g09864(new_n12151, new_n5465, new_n12213);
nor_5  g09865(new_n12213, new_n3442, new_n12214);
xor_4  g09866(new_n12211, new_n3439, new_n12215);
and_5  g09867(new_n12215, new_n12214, new_n12216);
nor_5  g09868(new_n12216, new_n12212, new_n12217);
nor_5  g09869(new_n12217, new_n12210, new_n12218);
nor_5  g09870(new_n12218, new_n12209_1, new_n12219);
nor_5  g09871(new_n12219, new_n12207, new_n12220);
nor_5  g09872(new_n12220, new_n12206, new_n12221);
nor_5  g09873(new_n12221, new_n12203, new_n12222);
nor_5  g09874(new_n12222, new_n12202, new_n12223_1);
nor_5  g09875(new_n12223_1, new_n12199, new_n12224);
nor_5  g09876(new_n12224, new_n12198, new_n12225_1);
nor_5  g09877(new_n12225_1, new_n12196, new_n12226);
nor_5  g09878(new_n12226, new_n12195, new_n12227);
nor_5  g09879(new_n12227, new_n12193, new_n12228_1);
nor_5  g09880(new_n12228_1, new_n12192_1, new_n12229);
nor_5  g09881(new_n12229, new_n12190, new_n12230);
nor_5  g09882(new_n12230, new_n12189, new_n12231);
nor_5  g09883(new_n12231, new_n12187, new_n12232);
nor_5  g09884(new_n12232, new_n12186, new_n12233);
nor_5  g09885(new_n12233, new_n12184, new_n12234);
or_5   g09886(new_n12234, new_n12183, new_n12235_1);
xor_4  g09887(new_n12235_1, new_n12177, n2561);
xor_4  g09888(new_n7665, new_n7663, n2573);
xor_4  g09889(n18558, n10411, new_n12238);
nor_5  g09890(new_n9119, n7149, new_n12239);
nor_5  g09891(n16971, new_n2783_1, new_n12240);
nor_5  g09892(n14148, new_n9123, new_n12241);
or_5   g09893(new_n2787, n11503, new_n12242);
nor_5  g09894(new_n9126, n1152, new_n12243);
and_5  g09895(new_n12243, new_n12242, new_n12244);
nor_5  g09896(new_n12244, new_n12241, new_n12245);
nor_5  g09897(new_n12245, new_n12240, new_n12246);
nor_5  g09898(new_n12246, new_n12239, new_n12247);
xor_4  g09899(new_n12247, new_n12238, new_n12248);
and_5  g09900(new_n9911, n6590, new_n12249);
nor_5  g09901(new_n9911, n6590, new_n12250);
and_5  g09902(n20349, new_n9914, new_n12251);
or_5   g09903(n20349, new_n9914, new_n12252);
and_5  g09904(n15936, new_n9917_1, new_n12253);
and_5  g09905(new_n12253, new_n12252, new_n12254);
nor_5  g09906(new_n12254, new_n12251, new_n12255);
nor_5  g09907(new_n12255, new_n12250, new_n12256);
nor_5  g09908(new_n12256, new_n12249, new_n12257);
xnor_4 g09909(new_n12257, new_n8996, new_n12258);
xnor_4 g09910(new_n12258, new_n12248, new_n12259);
xnor_4 g09911(n16971, n7149, new_n12260);
xnor_4 g09912(new_n12260, new_n12245, new_n12261);
xor_4  g09913(new_n12255, new_n9000, new_n12262);
not_10 g09914(new_n12262, new_n12263);
nor_5  g09915(new_n12263, new_n12261, new_n12264);
xor_4  g09916(new_n12262, new_n12261, new_n12265);
xnor_4 g09917(n18151, n1152, new_n12266);
or_5   g09918(new_n12266, new_n9006, new_n12267);
xor_4  g09919(n14148, n11503, new_n12268);
xnor_4 g09920(new_n12268, new_n12243, new_n12269);
and_5  g09921(new_n12269, new_n12267, new_n12270);
xnor_4 g09922(new_n12269, new_n12267, new_n12271);
xnor_4 g09923(new_n12253, new_n9003_1, new_n12272);
nor_5  g09924(new_n12272, new_n12271, new_n12273);
or_5   g09925(new_n12273, new_n12270, new_n12274);
nor_5  g09926(new_n12274, new_n12265, new_n12275);
nor_5  g09927(new_n12275, new_n12264, new_n12276);
xor_4  g09928(new_n12276, new_n12259, new_n12277);
xor_4  g09929(n19515, n17035, new_n12278);
not_10 g09930(n14684, new_n12279);
and_5  g09931(n22588, new_n12279, new_n12280);
nor_5  g09932(n22588, new_n12279, new_n12281);
and_5  g09933(n12209, new_n7687, new_n12282);
or_5   g09934(n12209, new_n7687, new_n12283);
not_10 g09935(n12892, new_n12284);
nor_5  g09936(n24732, new_n12284, new_n12285);
and_5  g09937(new_n12285, new_n12283, new_n12286);
nor_5  g09938(new_n12286, new_n12282, new_n12287);
nor_5  g09939(new_n12287, new_n12281, new_n12288);
nor_5  g09940(new_n12288, new_n12280, new_n12289);
xnor_4 g09941(new_n12289, new_n12278, new_n12290);
xnor_4 g09942(new_n12290, new_n12277, new_n12291);
xor_4  g09943(new_n12274, new_n12265, new_n12292);
xor_4  g09944(n22588, n14684, new_n12293);
xnor_4 g09945(new_n12293, new_n12287, new_n12294);
nor_5  g09946(new_n12294, new_n12292, new_n12295);
xnor_4 g09947(n24732, n12892, new_n12296);
xnor_4 g09948(new_n12266, new_n9006, new_n12297);
nor_5  g09949(new_n12297, new_n12296, new_n12298);
xor_4  g09950(n12209, n6631, new_n12299);
xnor_4 g09951(new_n12299, new_n12285, new_n12300);
not_10 g09952(new_n12300, new_n12301);
nor_5  g09953(new_n12301, new_n12298, new_n12302_1);
xnor_4 g09954(new_n12300, new_n12298, new_n12303);
xor_4  g09955(new_n12272, new_n12271, new_n12304_1);
and_5  g09956(new_n12304_1, new_n12303, new_n12305);
or_5   g09957(new_n12305, new_n12302_1, new_n12306);
xor_4  g09958(new_n12294, new_n12292, new_n12307);
and_5  g09959(new_n12307, new_n12306, new_n12308);
nor_5  g09960(new_n12308, new_n12295, new_n12309);
xnor_4 g09961(new_n12309, new_n12291, n2578);
not_10 g09962(new_n7137, new_n12311);
and_5  g09963(new_n10595_1, new_n12311, new_n12312);
xnor_4 g09964(new_n10595_1, new_n12311, new_n12313);
and_5  g09965(new_n7137, new_n7081, new_n12314);
nor_5  g09966(new_n7202, new_n7138, new_n12315_1);
nor_5  g09967(new_n12315_1, new_n12314, new_n12316);
nor_5  g09968(new_n12316, new_n12313, new_n12317);
nor_5  g09969(new_n12317, new_n12312, n2582);
xor_4  g09970(new_n4000_1, new_n3989, n2602);
nor_5  g09971(n22201, n2420, new_n12320);
not_10 g09972(new_n12320, new_n12321);
or_5   g09973(new_n12321, n24485, new_n12322);
or_5   g09974(new_n12322, n21078, new_n12323);
or_5   g09975(new_n12323, n12546, new_n12324_1);
xor_4  g09976(new_n12324_1, n8324, new_n12325_1);
xnor_4 g09977(new_n12325_1, new_n3725_1, new_n12326);
xor_4  g09978(new_n12323, n12546, new_n12327);
nor_5  g09979(new_n12327, new_n3727, new_n12328);
xor_4  g09980(new_n12322, n21078, new_n12329_1);
nor_5  g09981(new_n12329_1, new_n3729, new_n12330_1);
xnor_4 g09982(new_n12329_1, new_n3729, new_n12331);
xor_4  g09983(new_n12320, n24485, new_n12332);
nor_5  g09984(new_n12332, new_n3733_1, new_n12333);
xnor_4 g09985(new_n12332, new_n3733_1, new_n12334);
xor_4  g09986(n22201, n2420, new_n12335);
nor_5  g09987(new_n12335, new_n3738, new_n12336);
nand_5 g09988(new_n2530, n22201, new_n12337);
xnor_4 g09989(new_n12335, new_n3737, new_n12338);
and_5  g09990(new_n12338, new_n12337, new_n12339);
or_5   g09991(new_n12339, new_n12336, new_n12340);
nor_5  g09992(new_n12340, new_n12334, new_n12341_1);
or_5   g09993(new_n12341_1, new_n12333, new_n12342);
nor_5  g09994(new_n12342, new_n12331, new_n12343);
nor_5  g09995(new_n12343, new_n12330_1, new_n12344);
xnor_4 g09996(new_n12327, new_n3727, new_n12345);
nor_5  g09997(new_n12345, new_n12344, new_n12346_1);
nor_5  g09998(new_n12346_1, new_n12328, new_n12347);
xor_4  g09999(new_n12347, new_n12326, new_n12348);
not_10 g10000(new_n12348, new_n12349_1);
xnor_4 g10001(new_n7357, n7678, new_n12350);
nor_5  g10002(new_n7360, n3785, new_n12351);
xnor_4 g10003(new_n7360, n3785, new_n12352);
nor_5  g10004(new_n7363_1, n20250, new_n12353);
xnor_4 g10005(new_n7363_1, n20250, new_n12354);
nor_5  g10006(new_n7367, new_n4075, new_n12355);
and_5  g10007(new_n7367, new_n4075, new_n12356);
and_5  g10008(new_n7372, new_n4080, new_n12357);
or_5   g10009(new_n2525, new_n4084, new_n12358);
xnor_4 g10010(new_n7372, n26443, new_n12359);
and_5  g10011(new_n12359, new_n12358, new_n12360);
or_5   g10012(new_n12360, new_n12357, new_n12361);
nor_5  g10013(new_n12361, new_n12356, new_n12362);
or_5   g10014(new_n12362, new_n12355, new_n12363);
nor_5  g10015(new_n12363, new_n12354, new_n12364_1);
nor_5  g10016(new_n12364_1, new_n12353, new_n12365);
nor_5  g10017(new_n12365, new_n12352, new_n12366);
or_5   g10018(new_n12366, new_n12351, new_n12367);
xor_4  g10019(new_n12367, new_n12350, new_n12368);
xnor_4 g10020(new_n12368, new_n12349_1, new_n12369);
xor_4  g10021(new_n12365, new_n12352, new_n12370);
xor_4  g10022(new_n12345, new_n12344, new_n12371);
and_5  g10023(new_n12371, new_n12370, new_n12372);
xnor_4 g10024(new_n12371, new_n12370, new_n12373);
xor_4  g10025(new_n12342, new_n12331, new_n12374);
xor_4  g10026(new_n12363, new_n12354, new_n12375);
and_5  g10027(new_n12375, new_n12374, new_n12376);
not_10 g10028(new_n12374, new_n12377);
xnor_4 g10029(new_n12375, new_n12377, new_n12378);
xor_4  g10030(new_n12340, new_n12334, new_n12379);
xnor_4 g10031(new_n7367, n5822, new_n12380_1);
xnor_4 g10032(new_n12380_1, new_n12361, new_n12381);
and_5  g10033(new_n12381, new_n12379, new_n12382);
xor_4  g10034(new_n12338, new_n12337, new_n12383_1);
xor_4  g10035(new_n12359, new_n12358, new_n12384_1);
and_5  g10036(new_n12384_1, new_n12383_1, new_n12385);
xor_4  g10037(new_n2525, n1681, new_n12386);
xnor_4 g10038(new_n2530, n22201, new_n12387);
or_5   g10039(new_n12387, new_n12386, new_n12388);
not_10 g10040(new_n12383_1, new_n12389);
xnor_4 g10041(new_n12384_1, new_n12389, new_n12390);
and_5  g10042(new_n12390, new_n12388, new_n12391);
or_5   g10043(new_n12391, new_n12385, new_n12392);
xnor_4 g10044(new_n12381, new_n12379, new_n12393);
nor_5  g10045(new_n12393, new_n12392, new_n12394);
nor_5  g10046(new_n12394, new_n12382, new_n12395);
and_5  g10047(new_n12395, new_n12378, new_n12396);
nor_5  g10048(new_n12396, new_n12376, new_n12397_1);
nor_5  g10049(new_n12397_1, new_n12373, new_n12398_1);
nor_5  g10050(new_n12398_1, new_n12372, new_n12399);
xnor_4 g10051(new_n12399, new_n12369, n2619);
nor_5  g10052(new_n11548_1, new_n11542, new_n12401);
nor_5  g10053(new_n5432, n12900, new_n12402);
xnor_4 g10054(new_n5432, n12900, new_n12403);
nor_5  g10055(new_n5438_1, n20411, new_n12404);
xnor_4 g10056(new_n5438_1, n20411, new_n12405);
nor_5  g10057(new_n5443_1, n17069, new_n12406);
xnor_4 g10058(new_n5443_1, n17069, new_n12407);
nor_5  g10059(new_n5447, n15918, new_n12408_1);
nor_5  g10060(new_n5452, n17784, new_n12409);
xnor_4 g10061(new_n5452, n17784, new_n12410);
and_5  g10062(new_n5456, n14323, new_n12411);
nor_5  g10063(new_n11788, new_n11779, new_n12412);
or_5   g10064(new_n12412, new_n12411, new_n12413);
nor_5  g10065(new_n12413, new_n12410, new_n12414);
nor_5  g10066(new_n12414, new_n12409, new_n12415);
xnor_4 g10067(new_n5447, n15918, new_n12416);
nor_5  g10068(new_n12416, new_n12415, new_n12417);
nor_5  g10069(new_n12417, new_n12408_1, new_n12418);
nor_5  g10070(new_n12418, new_n12407, new_n12419);
nor_5  g10071(new_n12419, new_n12406, new_n12420);
nor_5  g10072(new_n12420, new_n12405, new_n12421);
nor_5  g10073(new_n12421, new_n12404, new_n12422);
nor_5  g10074(new_n12422, new_n12403, new_n12423);
or_5   g10075(new_n12423, new_n12402, new_n12424);
xor_4  g10076(new_n5395, n10650, new_n12425);
xnor_4 g10077(new_n12425, new_n12424, new_n12426);
nor_5  g10078(new_n12426, n6456, new_n12427);
xnor_4 g10079(new_n12426, n6456, new_n12428);
xnor_4 g10080(new_n12422, new_n12403, new_n12429);
nor_5  g10081(new_n12429, n4085, new_n12430);
xnor_4 g10082(new_n12429, n4085, new_n12431);
xnor_4 g10083(new_n12420, new_n12405, new_n12432);
nor_5  g10084(new_n12432, n26725, new_n12433);
xnor_4 g10085(new_n12432, n26725, new_n12434);
xnor_4 g10086(new_n12418, new_n12407, new_n12435);
nor_5  g10087(new_n12435, n11980, new_n12436);
xnor_4 g10088(new_n12435, n11980, new_n12437);
xnor_4 g10089(new_n12416, new_n12415, new_n12438);
nor_5  g10090(new_n12438, n3253, new_n12439);
xor_4  g10091(new_n12438, n3253, new_n12440);
xnor_4 g10092(new_n12413, new_n12410, new_n12441);
and_5  g10093(new_n12441, n7759, new_n12442);
xnor_4 g10094(new_n12441, n7759, new_n12443);
and_5  g10095(new_n11789, n12562, new_n12444);
nor_5  g10096(new_n11801, new_n11790, new_n12445);
nor_5  g10097(new_n12445, new_n12444, new_n12446_1);
nor_5  g10098(new_n12446_1, new_n12443, new_n12447);
nor_5  g10099(new_n12447, new_n12442, new_n12448);
and_5  g10100(new_n12448, new_n12440, new_n12449_1);
nor_5  g10101(new_n12449_1, new_n12439, new_n12450);
nor_5  g10102(new_n12450, new_n12437, new_n12451);
nor_5  g10103(new_n12451, new_n12436, new_n12452);
nor_5  g10104(new_n12452, new_n12434, new_n12453);
nor_5  g10105(new_n12453, new_n12433, new_n12454);
nor_5  g10106(new_n12454, new_n12431, new_n12455);
nor_5  g10107(new_n12455, new_n12430, new_n12456);
nor_5  g10108(new_n12456, new_n12428, new_n12457);
nor_5  g10109(new_n12457, new_n12427, new_n12458);
nor_5  g10110(new_n5395, n10650, new_n12459);
nor_5  g10111(new_n12459, new_n12424, new_n12460);
nor_5  g10112(new_n5394, n2979, new_n12461_1);
and_5  g10113(new_n5395, n10650, new_n12462_1);
or_5   g10114(new_n12462_1, new_n12461_1, new_n12463);
nor_5  g10115(new_n12463, new_n12460, new_n12464);
and_5  g10116(new_n12464, new_n12458, new_n12465);
nor_5  g10117(new_n12465, new_n12401, new_n12466);
xnor_4 g10118(new_n12465, new_n12401, new_n12467_1);
not_10 g10119(new_n11552, new_n12468);
xor_4  g10120(new_n12464, new_n12458, new_n12469_1);
nor_5  g10121(new_n12469_1, new_n12468, new_n12470);
xnor_4 g10122(new_n12469_1, new_n12468, new_n12471);
not_10 g10123(new_n11556, new_n12472);
xor_4  g10124(new_n12456, new_n12428, new_n12473);
and_5  g10125(new_n12473, new_n12472, new_n12474);
xnor_4 g10126(new_n12473, new_n12472, new_n12475);
not_10 g10127(new_n11560, new_n12476);
xor_4  g10128(new_n12454, new_n12431, new_n12477);
and_5  g10129(new_n12477, new_n12476, new_n12478);
xnor_4 g10130(new_n12477, new_n12476, new_n12479);
not_10 g10131(new_n11564_1, new_n12480);
xor_4  g10132(new_n12452, new_n12434, new_n12481);
and_5  g10133(new_n12481, new_n12480, new_n12482);
xnor_4 g10134(new_n12481, new_n12480, new_n12483);
not_10 g10135(new_n11568, new_n12484);
xor_4  g10136(new_n12450, new_n12437, new_n12485);
and_5  g10137(new_n12485, new_n12484, new_n12486);
xnor_4 g10138(new_n12485, new_n12484, new_n12487);
not_10 g10139(new_n11572, new_n12488);
xor_4  g10140(new_n12448, new_n12440, new_n12489);
and_5  g10141(new_n12489, new_n12488, new_n12490);
xnor_4 g10142(new_n12489, new_n12488, new_n12491);
xor_4  g10143(new_n12446_1, new_n12443, new_n12492);
nor_5  g10144(new_n12492, new_n11576, new_n12493);
xnor_4 g10145(new_n12492, new_n11576, new_n12494);
nor_5  g10146(new_n11802, new_n11580_1, new_n12495_1);
nor_5  g10147(new_n11816, new_n11803, new_n12496);
nor_5  g10148(new_n12496, new_n12495_1, new_n12497);
nor_5  g10149(new_n12497, new_n12494, new_n12498);
nor_5  g10150(new_n12498, new_n12493, new_n12499);
nor_5  g10151(new_n12499, new_n12491, new_n12500);
nor_5  g10152(new_n12500, new_n12490, new_n12501);
nor_5  g10153(new_n12501, new_n12487, new_n12502);
nor_5  g10154(new_n12502, new_n12486, new_n12503);
nor_5  g10155(new_n12503, new_n12483, new_n12504);
nor_5  g10156(new_n12504, new_n12482, new_n12505);
nor_5  g10157(new_n12505, new_n12479, new_n12506);
nor_5  g10158(new_n12506, new_n12478, new_n12507_1);
nor_5  g10159(new_n12507_1, new_n12475, new_n12508);
nor_5  g10160(new_n12508, new_n12474, new_n12509);
nor_5  g10161(new_n12509, new_n12471, new_n12510);
nor_5  g10162(new_n12510, new_n12470, new_n12511);
nor_5  g10163(new_n12511, new_n12467_1, new_n12512);
nor_5  g10164(new_n12512, new_n12466, n2661);
xnor_4 g10165(new_n10072, new_n10070, n2693);
xor_4  g10166(new_n12248, new_n6611_1, new_n12515_1);
nor_5  g10167(new_n12261, new_n6615, new_n12516_1);
xnor_4 g10168(new_n12261, new_n6615, new_n12517);
nor_5  g10169(new_n12269, new_n6619, new_n12518);
nor_5  g10170(new_n12266, new_n6621, new_n12519);
xor_4  g10171(new_n12269, new_n6619, new_n12520);
and_5  g10172(new_n12520, new_n12519, new_n12521);
nor_5  g10173(new_n12521, new_n12518, new_n12522);
nor_5  g10174(new_n12522, new_n12517, new_n12523);
nor_5  g10175(new_n12523, new_n12516_1, new_n12524);
xor_4  g10176(new_n12524, new_n12515_1, new_n12525);
xor_4  g10177(n8309, n4665, new_n12526);
nor_5  g10178(new_n9121, n19005, new_n12527);
nor_5  g10179(n19144, new_n2785, new_n12528);
nor_5  g10180(new_n7968_1, n4326, new_n12529);
or_5   g10181(n12593, new_n2789, new_n12530);
nor_5  g10182(new_n10902, n5438, new_n12531);
and_5  g10183(new_n12531, new_n12530, new_n12532);
nor_5  g10184(new_n12532, new_n12529, new_n12533);
nor_5  g10185(new_n12533, new_n12528, new_n12534);
nor_5  g10186(new_n12534, new_n12527, new_n12535);
xor_4  g10187(new_n12535, new_n12526, new_n12536);
xor_4  g10188(new_n12536, new_n12525, new_n12537);
xor_4  g10189(new_n12522, new_n12517, new_n12538);
not_10 g10190(new_n12538, new_n12539);
xnor_4 g10191(n19144, n19005, new_n12540_1);
xnor_4 g10192(new_n12540_1, new_n12533, new_n12541);
and_5  g10193(new_n12541, new_n12539, new_n12542);
xor_4  g10194(new_n12541, new_n12538, new_n12543);
xnor_4 g10195(n13714, n5438, new_n12544);
xnor_4 g10196(new_n12266, new_n6621, new_n12545_1);
or_5   g10197(new_n12545_1, new_n12544, new_n12546_1);
xor_4  g10198(n12593, n4326, new_n12547);
xnor_4 g10199(new_n12547, new_n12531, new_n12548);
and_5  g10200(new_n12548, new_n12546_1, new_n12549);
xnor_4 g10201(new_n12520, new_n12519, new_n12550);
xor_4  g10202(new_n12548, new_n12546_1, new_n12551);
and_5  g10203(new_n12551, new_n12550, new_n12552_1);
nor_5  g10204(new_n12552_1, new_n12549, new_n12553);
nor_5  g10205(new_n12553, new_n12543, new_n12554);
nor_5  g10206(new_n12554, new_n12542, new_n12555);
xnor_4 g10207(new_n12555, new_n12537, n2703);
xnor_4 g10208(new_n11662, new_n11652, n2706);
not_10 g10209(n1831, new_n12558);
nor_5  g10210(n3320, new_n12558, new_n12559);
xor_4  g10211(n3320, n1831, new_n12560);
not_10 g10212(n13137, new_n12561);
nor_5  g10213(new_n12561, n1288, new_n12562_1);
xor_4  g10214(n13137, n1288, new_n12563);
not_10 g10215(n18452, new_n12564);
nor_5  g10216(new_n12564, n1752, new_n12565);
xor_4  g10217(n18452, n1752, new_n12566_1);
not_10 g10218(n21317, new_n12567);
nor_5  g10219(new_n12567, n13110, new_n12568);
xor_4  g10220(n21317, n13110, new_n12569_1);
not_10 g10221(n12398, new_n12570);
nor_5  g10222(n25694, new_n12570, new_n12571);
xor_4  g10223(n25694, n12398, new_n12572);
nor_5  g10224(new_n3752, n15424, new_n12573);
xor_4  g10225(n19789, n15424, new_n12574);
not_10 g10226(n1949, new_n12575);
nor_5  g10227(n20169, new_n12575, new_n12576);
nor_5  g10228(new_n10996, new_n10985, new_n12577);
or_5   g10229(new_n12577, new_n12576, new_n12578);
nor_5  g10230(new_n12578, new_n12574, new_n12579);
nor_5  g10231(new_n12579, new_n12573, new_n12580);
nor_5  g10232(new_n12580, new_n12572, new_n12581);
nor_5  g10233(new_n12581, new_n12571, new_n12582);
nor_5  g10234(new_n12582, new_n12569_1, new_n12583);
nor_5  g10235(new_n12583, new_n12568, new_n12584);
nor_5  g10236(new_n12584, new_n12566_1, new_n12585);
nor_5  g10237(new_n12585, new_n12565, new_n12586);
nor_5  g10238(new_n12586, new_n12563, new_n12587_1);
nor_5  g10239(new_n12587_1, new_n12562_1, new_n12588);
nor_5  g10240(new_n12588, new_n12560, new_n12589);
nor_5  g10241(new_n12589, new_n12559, new_n12590);
not_10 g10242(n1483, new_n12591);
nor_5  g10243(n19539, new_n12591, new_n12592);
nor_5  g10244(new_n10172, new_n10158_1, new_n12593_1);
nor_5  g10245(new_n12593_1, new_n12592, new_n12594);
and_5  g10246(new_n5883, new_n11142, new_n12595);
not_10 g10247(new_n12595, new_n12596);
or_5   g10248(new_n12596, n3541, new_n12597);
xnor_4 g10249(new_n12597, n2184, new_n12598);
and_5  g10250(new_n12598, new_n11088, new_n12599);
xor_4  g10251(new_n12597, n2184, new_n12600);
xnor_4 g10252(new_n12600, n6204, new_n12601);
xnor_4 g10253(new_n12595, n3541, new_n12602);
and_5  g10254(new_n12602, n3349, new_n12603);
nor_5  g10255(new_n12602, n3349, new_n12604);
and_5  g10256(new_n5884, n1742, new_n12605);
nor_5  g10257(new_n5884, n1742, new_n12606);
nor_5  g10258(new_n5912, new_n12606, new_n12607_1);
nor_5  g10259(new_n12607_1, new_n12605, new_n12608);
nor_5  g10260(new_n12608, new_n12604, new_n12609);
or_5   g10261(new_n12609, new_n12603, new_n12610);
nor_5  g10262(new_n12610, new_n12601, new_n12611);
nor_5  g10263(new_n12611, new_n12599, new_n12612);
nor_5  g10264(new_n12597, n2184, new_n12613);
xnor_4 g10265(new_n12613, n10018, new_n12614);
xor_4  g10266(new_n12614, n5140, new_n12615);
xnor_4 g10267(new_n12615, new_n12612, new_n12616);
and_5  g10268(new_n12616, new_n10173, new_n12617);
xnor_4 g10269(new_n12616, new_n10173, new_n12618);
xnor_4 g10270(new_n10170, new_n10161, new_n12619);
xor_4  g10271(new_n12610, new_n12601, new_n12620_1);
and_5  g10272(new_n12620_1, new_n12619, new_n12621_1);
xnor_4 g10273(new_n12620_1, new_n12619, new_n12622);
xnor_4 g10274(new_n12602, new_n11091, new_n12623);
xnor_4 g10275(new_n12623, new_n12608, new_n12624);
and_5  g10276(new_n12624, new_n10239_1, new_n12625);
xnor_4 g10277(new_n12624, new_n10239_1, new_n12626_1);
nor_5  g10278(new_n5913, new_n5875, new_n12627);
nor_5  g10279(new_n5950, new_n5914, new_n12628);
nor_5  g10280(new_n12628, new_n12627, new_n12629);
nor_5  g10281(new_n12629, new_n12626_1, new_n12630);
or_5   g10282(new_n12630, new_n12625, new_n12631);
nor_5  g10283(new_n12631, new_n12622, new_n12632);
nor_5  g10284(new_n12632, new_n12621_1, new_n12633);
nor_5  g10285(new_n12633, new_n12618, new_n12634);
or_5   g10286(new_n12634, new_n12617, new_n12635);
and_5  g10287(new_n12613, new_n11133, new_n12636);
nor_5  g10288(new_n12614, n5140, new_n12637);
and_5  g10289(new_n12614, n5140, new_n12638);
nor_5  g10290(new_n12638, new_n12612, new_n12639);
nor_5  g10291(new_n12639, new_n12637, new_n12640);
nor_5  g10292(new_n12640, new_n12636, new_n12641);
nor_5  g10293(new_n12641, new_n12635, new_n12642);
and_5  g10294(new_n12642, new_n12594, new_n12643);
nand_5 g10295(new_n12641, new_n12635, new_n12644);
nor_5  g10296(new_n12644, new_n12594, new_n12645);
nor_5  g10297(new_n12645, new_n12643, new_n12646);
xnor_4 g10298(new_n12646, new_n12590, new_n12647);
xor_4  g10299(new_n12641, new_n12635, new_n12648);
xnor_4 g10300(new_n12648, new_n12594, new_n12649);
and_5  g10301(new_n12649, new_n12590, new_n12650_1);
nor_5  g10302(new_n12649, new_n12590, new_n12651);
xnor_4 g10303(new_n12588, new_n12560, new_n12652);
xor_4  g10304(new_n12633, new_n12618, new_n12653);
and_5  g10305(new_n12653, new_n12652, new_n12654_1);
xnor_4 g10306(new_n12653, new_n12652, new_n12655);
xnor_4 g10307(new_n12586, new_n12563, new_n12656);
xor_4  g10308(new_n12631, new_n12622, new_n12657_1);
and_5  g10309(new_n12657_1, new_n12656, new_n12658);
xnor_4 g10310(new_n12657_1, new_n12656, new_n12659);
xor_4  g10311(new_n12584, new_n12566_1, new_n12660);
xor_4  g10312(new_n12629, new_n12626_1, new_n12661);
nor_5  g10313(new_n12661, new_n12660, new_n12662);
xnor_4 g10314(new_n12661, new_n12660, new_n12663);
xor_4  g10315(new_n5950, new_n5914, new_n12664);
xor_4  g10316(new_n12582, new_n12569_1, new_n12665_1);
nor_5  g10317(new_n12665_1, new_n12664, new_n12666);
xor_4  g10318(new_n12580, new_n12572, new_n12667);
nor_5  g10319(new_n12667, new_n5953, new_n12668);
xnor_4 g10320(new_n12667, new_n5953, new_n12669);
xor_4  g10321(new_n5956, new_n5922, new_n12670_1);
xor_4  g10322(new_n12578, new_n12574, new_n12671);
nor_5  g10323(new_n12671, new_n12670_1, new_n12672);
xnor_4 g10324(new_n12671, new_n12670_1, new_n12673);
and_5  g10325(new_n10997, new_n10984, new_n12674);
nor_5  g10326(new_n11013, new_n10998, new_n12675);
nor_5  g10327(new_n12675, new_n12674, new_n12676);
nor_5  g10328(new_n12676, new_n12673, new_n12677);
nor_5  g10329(new_n12677, new_n12672, new_n12678);
nor_5  g10330(new_n12678, new_n12669, new_n12679);
or_5   g10331(new_n12679, new_n12668, new_n12680);
xnor_4 g10332(new_n12665_1, new_n5951, new_n12681);
and_5  g10333(new_n12681, new_n12680, new_n12682);
nor_5  g10334(new_n12682, new_n12666, new_n12683);
nor_5  g10335(new_n12683, new_n12663, new_n12684);
nor_5  g10336(new_n12684, new_n12662, new_n12685);
nor_5  g10337(new_n12685, new_n12659, new_n12686);
nor_5  g10338(new_n12686, new_n12658, new_n12687);
nor_5  g10339(new_n12687, new_n12655, new_n12688);
or_5   g10340(new_n12688, new_n12654_1, new_n12689);
nor_5  g10341(new_n12689, new_n12651, new_n12690);
nor_5  g10342(new_n12690, new_n12650_1, new_n12691);
xnor_4 g10343(new_n12691, new_n12647, n2711);
xor_4  g10344(n10611, n2680, new_n12693);
and_5  g10345(new_n8287, n1667, new_n12694);
nor_5  g10346(new_n8287, n1667, new_n12695);
and_5  g10347(new_n8290, n7339, new_n12696);
or_5   g10348(new_n8290, n7339, new_n12697);
nor_5  g10349(new_n8343, n18, new_n12698);
and_5  g10350(new_n12698, new_n12697, new_n12699);
nor_5  g10351(new_n12699, new_n12696, new_n12700);
nor_5  g10352(new_n12700, new_n12695, new_n12701);
nor_5  g10353(new_n12701, new_n12694, new_n12702_1);
xor_4  g10354(new_n12702_1, new_n12693, new_n12703);
xnor_4 g10355(new_n12703, new_n8219, new_n12704);
xnor_4 g10356(n2783, n1667, new_n12705);
xnor_4 g10357(new_n12705, new_n12700, new_n12706);
and_5  g10358(new_n12706, new_n8223, new_n12707_1);
xnor_4 g10359(new_n12706, new_n8223, new_n12708);
xnor_4 g10360(n26808, n18, new_n12709);
or_5   g10361(new_n12709, new_n8229, new_n12710);
xor_4  g10362(n15490, n7339, new_n12711);
xnor_4 g10363(new_n12711, new_n12698, new_n12712);
and_5  g10364(new_n12712, new_n12710, new_n12713);
xor_4  g10365(new_n12712, new_n12710, new_n12714);
and_5  g10366(new_n12714, new_n8234, new_n12715);
nor_5  g10367(new_n12715, new_n12713, new_n12716);
nor_5  g10368(new_n12716, new_n12708, new_n12717);
nor_5  g10369(new_n12717, new_n12707_1, new_n12718);
xnor_4 g10370(new_n12718, new_n12704, n2761);
xnor_4 g10371(n25120, n8526, new_n12720);
nor_5  g10372(n8363, n2816, new_n12721);
xnor_4 g10373(n8363, n2816, new_n12722);
nor_5  g10374(n20359, n14680, new_n12723);
xnor_4 g10375(n20359, n14680, new_n12724);
nor_5  g10376(n17250, n4409, new_n12725_1);
nor_5  g10377(new_n8488, new_n8467, new_n12726);
nor_5  g10378(new_n12726, new_n12725_1, new_n12727_1);
nor_5  g10379(new_n12727_1, new_n12724, new_n12728);
nor_5  g10380(new_n12728, new_n12723, new_n12729);
nor_5  g10381(new_n12729, new_n12722, new_n12730);
nor_5  g10382(new_n12730, new_n12721, new_n12731);
xnor_4 g10383(new_n12731, new_n12720, new_n12732);
nor_5  g10384(new_n12732, n17458, new_n12733);
xor_4  g10385(new_n12732, n17458, new_n12734);
xnor_4 g10386(new_n12729, new_n12722, new_n12735);
and_5  g10387(new_n12735, n1222, new_n12736);
xnor_4 g10388(new_n12727_1, new_n12724, new_n12737);
nor_5  g10389(new_n12737, n25240, new_n12738);
xor_4  g10390(new_n12737, n25240, new_n12739);
and_5  g10391(new_n8489_1, n10125, new_n12740_1);
xnor_4 g10392(new_n8489_1, n10125, new_n12741);
and_5  g10393(new_n8491, n8067, new_n12742_1);
xnor_4 g10394(new_n8491, n8067, new_n12743);
and_5  g10395(new_n8494, n20923, new_n12744);
xnor_4 g10396(new_n8494, n20923, new_n12745);
and_5  g10397(new_n8497, n18157, new_n12746_1);
xnor_4 g10398(new_n8497, n18157, new_n12747);
and_5  g10399(new_n8500, n12161, new_n12748);
nor_5  g10400(new_n8502, n5026, new_n12749);
nand_5 g10401(new_n8504, n8581, new_n12750);
xor_4  g10402(new_n8502, n5026, new_n12751);
and_5  g10403(new_n12751, new_n12750, new_n12752);
nor_5  g10404(new_n12752, new_n12749, new_n12753);
xor_4  g10405(new_n8500, n12161, new_n12754);
and_5  g10406(new_n12754, new_n12753, new_n12755);
nor_5  g10407(new_n12755, new_n12748, new_n12756_1);
nor_5  g10408(new_n12756_1, new_n12747, new_n12757);
nor_5  g10409(new_n12757, new_n12746_1, new_n12758);
nor_5  g10410(new_n12758, new_n12745, new_n12759);
nor_5  g10411(new_n12759, new_n12744, new_n12760);
nor_5  g10412(new_n12760, new_n12743, new_n12761);
nor_5  g10413(new_n12761, new_n12742_1, new_n12762);
nor_5  g10414(new_n12762, new_n12741, new_n12763);
nor_5  g10415(new_n12763, new_n12740_1, new_n12764);
and_5  g10416(new_n12764, new_n12739, new_n12765);
or_5   g10417(new_n12765, new_n12738, new_n12766);
xnor_4 g10418(new_n12735, n1222, new_n12767);
nor_5  g10419(new_n12767, new_n12766, new_n12768);
nor_5  g10420(new_n12768, new_n12736, new_n12769);
and_5  g10421(new_n12769, new_n12734, new_n12770);
nor_5  g10422(new_n12770, new_n12733, new_n12771);
or_5   g10423(n25120, n8526, new_n12772);
or_5   g10424(new_n12731, new_n12720, new_n12773);
and_5  g10425(new_n12773, new_n12772, new_n12774);
and_5  g10426(new_n12774, new_n12771, new_n12775);
or_5   g10427(new_n3522, n2113, new_n12776);
or_5   g10428(new_n12776, n1099, new_n12777);
or_5   g10429(new_n12777, n19941, new_n12778);
xor_4  g10430(new_n12778, n11898, new_n12779);
nor_5  g10431(new_n12779, new_n4476_1, new_n12780);
xnor_4 g10432(new_n12779, new_n4476_1, new_n12781);
xor_4  g10433(new_n12777, n19941, new_n12782);
nor_5  g10434(new_n12782, new_n4479, new_n12783_1);
xnor_4 g10435(new_n12782, new_n4479, new_n12784);
xor_4  g10436(new_n12776, n1099, new_n12785);
nor_5  g10437(new_n12785, new_n4483, new_n12786);
xnor_4 g10438(new_n12785, new_n4483, new_n12787);
nor_5  g10439(new_n4487, new_n3523, new_n12788);
xnor_4 g10440(new_n4487, new_n3523, new_n12789);
nor_5  g10441(new_n4491, new_n3525, new_n12790);
xnor_4 g10442(new_n4491, new_n3525, new_n12791);
nor_5  g10443(new_n4495, new_n3528_1, new_n12792);
xnor_4 g10444(new_n4495, new_n3528_1, new_n12793);
nor_5  g10445(new_n4499, new_n3531, new_n12794);
xnor_4 g10446(new_n4499, new_n3531, new_n12795);
nor_5  g10447(new_n4503, new_n3533, new_n12796);
xnor_4 g10448(new_n4503, new_n3533, new_n12797);
nor_5  g10449(new_n4508, n25435, new_n12798);
and_5  g10450(new_n12798, new_n3901, new_n12799);
or_5   g10451(new_n4508, n25435, new_n12800);
and_5  g10452(new_n12800, new_n3536, new_n12801_1);
nor_5  g10453(new_n12801_1, new_n12799, new_n12802);
and_5  g10454(new_n12802, new_n4506, new_n12803);
nor_5  g10455(new_n12803, new_n12799, new_n12804);
nor_5  g10456(new_n12804, new_n12797, new_n12805);
nor_5  g10457(new_n12805, new_n12796, new_n12806);
nor_5  g10458(new_n12806, new_n12795, new_n12807);
nor_5  g10459(new_n12807, new_n12794, new_n12808);
nor_5  g10460(new_n12808, new_n12793, new_n12809);
nor_5  g10461(new_n12809, new_n12792, new_n12810);
nor_5  g10462(new_n12810, new_n12791, new_n12811_1);
nor_5  g10463(new_n12811_1, new_n12790, new_n12812_1);
nor_5  g10464(new_n12812_1, new_n12789, new_n12813);
nor_5  g10465(new_n12813, new_n12788, new_n12814);
nor_5  g10466(new_n12814, new_n12787, new_n12815);
nor_5  g10467(new_n12815, new_n12786, new_n12816_1);
nor_5  g10468(new_n12816_1, new_n12784, new_n12817);
nor_5  g10469(new_n12817, new_n12783_1, new_n12818);
nor_5  g10470(new_n12818, new_n12781, new_n12819);
nor_5  g10471(new_n12819, new_n12780, new_n12820);
nor_5  g10472(new_n12778, n11898, new_n12821_1);
and_5  g10473(new_n12821_1, new_n4533, new_n12822);
and_5  g10474(new_n12822, new_n12820, new_n12823);
or_5   g10475(new_n12821_1, new_n4533, new_n12824);
nor_5  g10476(new_n12824, new_n12820, new_n12825);
nor_5  g10477(new_n12825, new_n12823, new_n12826);
and_5  g10478(new_n12826, new_n12775, new_n12827);
or_5   g10479(new_n12826, new_n12775, new_n12828);
not_10 g10480(new_n12774, new_n12829);
xnor_4 g10481(new_n12829, new_n12771, new_n12830);
xor_4  g10482(new_n12821_1, new_n4533, new_n12831);
xnor_4 g10483(new_n12831, new_n12820, new_n12832);
nor_5  g10484(new_n12832, new_n12830, new_n12833);
xnor_4 g10485(new_n12832, new_n12830, new_n12834);
xor_4  g10486(new_n12769, new_n12734, new_n12835);
xor_4  g10487(new_n12818, new_n12781, new_n12836);
and_5  g10488(new_n12836, new_n12835, new_n12837);
xnor_4 g10489(new_n12836, new_n12835, new_n12838);
xnor_4 g10490(new_n12816_1, new_n12784, new_n12839);
xor_4  g10491(new_n12767, new_n12766, new_n12840);
nor_5  g10492(new_n12840, new_n12839, new_n12841);
xnor_4 g10493(new_n12840, new_n12839, new_n12842);
xor_4  g10494(new_n12764, new_n12739, new_n12843_1);
xor_4  g10495(new_n12814, new_n12787, new_n12844);
and_5  g10496(new_n12844, new_n12843_1, new_n12845);
xnor_4 g10497(new_n12844, new_n12843_1, new_n12846);
xnor_4 g10498(new_n12812_1, new_n12789, new_n12847);
xor_4  g10499(new_n12762, new_n12741, new_n12848);
nor_5  g10500(new_n12848, new_n12847, new_n12849);
xnor_4 g10501(new_n12848, new_n12847, new_n12850);
xnor_4 g10502(new_n12810, new_n12791, new_n12851);
xor_4  g10503(new_n12760, new_n12743, new_n12852);
nor_5  g10504(new_n12852, new_n12851, new_n12853);
xnor_4 g10505(new_n12852, new_n12851, new_n12854);
xnor_4 g10506(new_n12808, new_n12793, new_n12855);
xor_4  g10507(new_n12758, new_n12745, new_n12856);
nor_5  g10508(new_n12856, new_n12855, new_n12857);
xnor_4 g10509(new_n12856, new_n12855, new_n12858);
xnor_4 g10510(new_n12806, new_n12795, new_n12859);
xor_4  g10511(new_n12756_1, new_n12747, new_n12860);
nor_5  g10512(new_n12860, new_n12859, new_n12861_1);
xor_4  g10513(new_n12860, new_n12859, new_n12862);
xnor_4 g10514(new_n12804, new_n12797, new_n12863);
xor_4  g10515(new_n12754, new_n12753, new_n12864_1);
and_5  g10516(new_n12864_1, new_n12863, new_n12865_1);
xnor_4 g10517(new_n12864_1, new_n12863, new_n12866);
xor_4  g10518(new_n12751, new_n12750, new_n12867);
xor_4  g10519(new_n12802, new_n4506, new_n12868);
and_5  g10520(new_n12868, new_n12867, new_n12869);
xor_4  g10521(new_n8504, n8581, new_n12870_1);
xnor_4 g10522(new_n4508, n25435, new_n12871_1);
nand_5 g10523(new_n12871_1, new_n12870_1, new_n12872);
not_10 g10524(new_n12867, new_n12873_1);
xnor_4 g10525(new_n12868, new_n12873_1, new_n12874);
and_5  g10526(new_n12874, new_n12872, new_n12875_1);
or_5   g10527(new_n12875_1, new_n12869, new_n12876);
nor_5  g10528(new_n12876, new_n12866, new_n12877);
nor_5  g10529(new_n12877, new_n12865_1, new_n12878);
and_5  g10530(new_n12878, new_n12862, new_n12879);
nor_5  g10531(new_n12879, new_n12861_1, new_n12880);
nor_5  g10532(new_n12880, new_n12858, new_n12881);
nor_5  g10533(new_n12881, new_n12857, new_n12882);
nor_5  g10534(new_n12882, new_n12854, new_n12883);
nor_5  g10535(new_n12883, new_n12853, new_n12884);
nor_5  g10536(new_n12884, new_n12850, new_n12885);
nor_5  g10537(new_n12885, new_n12849, new_n12886);
nor_5  g10538(new_n12886, new_n12846, new_n12887);
nor_5  g10539(new_n12887, new_n12845, new_n12888);
nor_5  g10540(new_n12888, new_n12842, new_n12889);
nor_5  g10541(new_n12889, new_n12841, new_n12890);
nor_5  g10542(new_n12890, new_n12838, new_n12891);
nor_5  g10543(new_n12891, new_n12837, new_n12892_1);
nor_5  g10544(new_n12892_1, new_n12834, new_n12893);
nor_5  g10545(new_n12893, new_n12833, new_n12894);
and_5  g10546(new_n12894, new_n12828, new_n12895);
or_5   g10547(new_n12895, new_n12823, new_n12896);
nor_5  g10548(new_n12896, new_n12827, n2774);
or_5   g10549(new_n8556, n20478, new_n12898);
or_5   g10550(new_n12898, n987, new_n12899);
or_5   g10551(new_n12899, n2421, new_n12900_1);
or_5   g10552(new_n12900_1, n11044, new_n12901);
or_5   g10553(new_n12901, n5031, new_n12902);
xor_4  g10554(new_n12902, n2145, new_n12903);
xor_4  g10555(new_n12903, n2858, new_n12904_1);
xor_4  g10556(new_n12901, n5031, new_n12905);
nor_5  g10557(new_n12905, n2659, new_n12906);
xnor_4 g10558(new_n12905, n2659, new_n12907);
xor_4  g10559(new_n12900_1, n11044, new_n12908);
nor_5  g10560(new_n12908, n24327, new_n12909);
xnor_4 g10561(new_n12908, n24327, new_n12910);
xor_4  g10562(new_n12899, n2421, new_n12911);
nor_5  g10563(new_n12911, n22198, new_n12912);
xor_4  g10564(new_n12898, n987, new_n12913);
and_5  g10565(new_n12913, n20826, new_n12914);
xnor_4 g10566(new_n12913, n20826, new_n12915);
and_5  g10567(new_n8557, n7305, new_n12916);
nor_5  g10568(new_n8569, new_n8558, new_n12917_1);
nor_5  g10569(new_n12917_1, new_n12916, new_n12918);
nor_5  g10570(new_n12918, new_n12915, new_n12919);
nor_5  g10571(new_n12919, new_n12914, new_n12920);
xor_4  g10572(new_n12911, n22198, new_n12921);
and_5  g10573(new_n12921, new_n12920, new_n12922);
nor_5  g10574(new_n12922, new_n12912, new_n12923);
nor_5  g10575(new_n12923, new_n12910, new_n12924);
nor_5  g10576(new_n12924, new_n12909, new_n12925);
nor_5  g10577(new_n12925, new_n12907, new_n12926);
nor_5  g10578(new_n12926, new_n12906, new_n12927);
xnor_4 g10579(new_n12927, new_n12904_1, new_n12928);
xnor_4 g10580(new_n12928, new_n3306_1, new_n12929);
xor_4  g10581(new_n12925, new_n12907, new_n12930);
nor_5  g10582(new_n12930, new_n3309, new_n12931);
xor_4  g10583(new_n12923, new_n12910, new_n12932);
not_10 g10584(new_n12932, new_n12933);
nor_5  g10585(new_n12933, new_n3313, new_n12934);
xnor_4 g10586(new_n12933, new_n3313, new_n12935);
xnor_4 g10587(new_n12921, new_n12920, new_n12936);
nor_5  g10588(new_n12936, new_n3316_1, new_n12937);
xnor_4 g10589(new_n12936, new_n3316_1, new_n12938);
xor_4  g10590(new_n12918, new_n12915, new_n12939);
nor_5  g10591(new_n12939, new_n3319, new_n12940);
xnor_4 g10592(new_n12939, new_n3319, new_n12941_1);
and_5  g10593(new_n8570, new_n3322, new_n12942_1);
xnor_4 g10594(new_n8570, new_n3322, new_n12943);
and_5  g10595(new_n8585, new_n3325, new_n12944);
xnor_4 g10596(new_n8585, new_n3325, new_n12945);
nor_5  g10597(new_n8590, new_n3330, new_n12946);
not_10 g10598(new_n3332_1, new_n12947);
or_5   g10599(new_n8592, new_n12947, new_n12948);
xor_4  g10600(new_n8589, new_n3330, new_n12949);
nor_5  g10601(new_n12949, new_n12948, new_n12950);
nor_5  g10602(new_n12950, new_n12946, new_n12951);
nor_5  g10603(new_n12951, new_n12945, new_n12952);
nor_5  g10604(new_n12952, new_n12944, new_n12953);
nor_5  g10605(new_n12953, new_n12943, new_n12954);
or_5   g10606(new_n12954, new_n12942_1, new_n12955);
nor_5  g10607(new_n12955, new_n12941_1, new_n12956_1);
nor_5  g10608(new_n12956_1, new_n12940, new_n12957);
nor_5  g10609(new_n12957, new_n12938, new_n12958);
nor_5  g10610(new_n12958, new_n12937, new_n12959);
nor_5  g10611(new_n12959, new_n12935, new_n12960);
nor_5  g10612(new_n12960, new_n12934, new_n12961);
xor_4  g10613(new_n12930, new_n3309, new_n12962);
and_5  g10614(new_n12962, new_n12961, new_n12963);
nor_5  g10615(new_n12963, new_n12931, new_n12964);
xor_4  g10616(new_n12964, new_n12929, new_n12965);
xor_4  g10617(new_n3409, n7026, new_n12966);
and_5  g10618(new_n3413, n13719, new_n12967);
or_5   g10619(new_n3413, n13719, new_n12968);
nor_5  g10620(new_n3417, n442, new_n12969);
xnor_4 g10621(new_n3417, n442, new_n12970);
nor_5  g10622(new_n3421, n9172, new_n12971);
xnor_4 g10623(new_n3421, n9172, new_n12972);
nor_5  g10624(new_n3424, n4913, new_n12973);
xnor_4 g10625(new_n3424, n4913, new_n12974);
nor_5  g10626(new_n3428, n604, new_n12975);
xor_4  g10627(new_n3397, n11273, new_n12976);
nor_5  g10628(new_n12976, n16824, new_n12977);
xnor_4 g10629(new_n12976, n16824, new_n12978_1);
nor_5  g10630(new_n3436, n16521, new_n12979);
nand_5 g10631(n21993, n7139, new_n12980_1);
xor_4  g10632(new_n3436, n16521, new_n12981);
and_5  g10633(new_n12981, new_n12980_1, new_n12982);
nor_5  g10634(new_n12982, new_n12979, new_n12983);
nor_5  g10635(new_n12983, new_n12978_1, new_n12984);
nor_5  g10636(new_n12984, new_n12977, new_n12985_1);
xnor_4 g10637(new_n3428, n604, new_n12986);
nor_5  g10638(new_n12986, new_n12985_1, new_n12987_1);
nor_5  g10639(new_n12987_1, new_n12975, new_n12988);
nor_5  g10640(new_n12988, new_n12974, new_n12989);
nor_5  g10641(new_n12989, new_n12973, new_n12990);
nor_5  g10642(new_n12990, new_n12972, new_n12991);
nor_5  g10643(new_n12991, new_n12971, new_n12992_1);
nor_5  g10644(new_n12992_1, new_n12970, new_n12993);
nor_5  g10645(new_n12993, new_n12969, new_n12994);
and_5  g10646(new_n12994, new_n12968, new_n12995);
nor_5  g10647(new_n12995, new_n12967, new_n12996);
xor_4  g10648(new_n12996, new_n12966, new_n12997);
xor_4  g10649(new_n12997, new_n12965, new_n12998);
xor_4  g10650(new_n12962, new_n12961, new_n12999);
xnor_4 g10651(new_n3413, n13719, new_n13000);
xnor_4 g10652(new_n13000, new_n12994, new_n13001);
and_5  g10653(new_n13001, new_n12999, new_n13002);
xnor_4 g10654(new_n13001, new_n12999, new_n13003);
xor_4  g10655(new_n12992_1, new_n12970, new_n13004);
xor_4  g10656(new_n12959, new_n12935, new_n13005_1);
and_5  g10657(new_n13005_1, new_n13004, new_n13006);
xnor_4 g10658(new_n13005_1, new_n13004, new_n13007);
xor_4  g10659(new_n12990, new_n12972, new_n13008);
xor_4  g10660(new_n12957, new_n12938, new_n13009);
and_5  g10661(new_n13009, new_n13008, new_n13010);
xor_4  g10662(new_n13009, new_n13008, new_n13011);
xor_4  g10663(new_n12988, new_n12974, new_n13012);
xor_4  g10664(new_n12955, new_n12941_1, new_n13013);
nor_5  g10665(new_n13013, new_n13012, new_n13014);
xor_4  g10666(new_n12986, new_n12985_1, new_n13015);
xnor_4 g10667(new_n12953, new_n12943, new_n13016);
nor_5  g10668(new_n13016, new_n13015, new_n13017);
xnor_4 g10669(new_n13016, new_n13015, new_n13018);
xnor_4 g10670(new_n12983, new_n12978_1, new_n13019);
xor_4  g10671(new_n12951, new_n12945, new_n13020);
and_5  g10672(new_n13020, new_n13019, new_n13021);
xnor_4 g10673(new_n13020, new_n13019, new_n13022);
xor_4  g10674(new_n12949, new_n12948, new_n13023);
nor_5  g10675(new_n13023, new_n12981, new_n13024);
not_10 g10676(new_n13023, new_n13025);
xor_4  g10677(new_n12981, new_n12980_1, new_n13026_1);
or_5   g10678(new_n13026_1, new_n13025, new_n13027);
xnor_4 g10679(n21993, n7139, new_n13028);
xor_4  g10680(new_n8592, new_n3332_1, new_n13029);
or_5   g10681(new_n13029, new_n13028, new_n13030);
and_5  g10682(new_n13030, new_n13027, new_n13031);
or_5   g10683(new_n13031, new_n13024, new_n13032);
nor_5  g10684(new_n13032, new_n13022, new_n13033);
nor_5  g10685(new_n13033, new_n13021, new_n13034);
nor_5  g10686(new_n13034, new_n13018, new_n13035);
nor_5  g10687(new_n13035, new_n13017, new_n13036);
xnor_4 g10688(new_n13013, new_n13012, new_n13037);
nor_5  g10689(new_n13037, new_n13036, new_n13038);
nor_5  g10690(new_n13038, new_n13014, new_n13039);
and_5  g10691(new_n13039, new_n13011, new_n13040);
nor_5  g10692(new_n13040, new_n13010, new_n13041);
nor_5  g10693(new_n13041, new_n13007, new_n13042);
or_5   g10694(new_n13042, new_n13006, new_n13043_1);
nor_5  g10695(new_n13043_1, new_n13003, new_n13044_1);
nor_5  g10696(new_n13044_1, new_n13002, new_n13045);
xnor_4 g10697(new_n13045, new_n12998, n2779);
xor_4  g10698(new_n9305, new_n9271, new_n13047);
nor_5  g10699(new_n9331, n25751, new_n13048_1);
xnor_4 g10700(new_n9331, n25751, new_n13049);
nor_5  g10701(new_n9334, n26053, new_n13050);
xnor_4 g10702(new_n9334, n26053, new_n13051);
nor_5  g10703(new_n9337, n7917, new_n13052);
xnor_4 g10704(new_n9337, n7917, new_n13053);
nor_5  g10705(new_n9340, n17302, new_n13054_1);
xnor_4 g10706(new_n9340, n17302, new_n13055);
nor_5  g10707(new_n9342, n2013, new_n13056);
xnor_4 g10708(new_n9342, n2013, new_n13057);
nor_5  g10709(new_n9345, n23755, new_n13058);
nor_5  g10710(new_n9348, n19163, new_n13059);
xnor_4 g10711(new_n9348, n19163, new_n13060);
nor_5  g10712(new_n5343, n22358, new_n13061);
and_5  g10713(n25926, n9646, new_n13062);
xnor_4 g10714(new_n5343, n22358, new_n13063);
nor_5  g10715(new_n13063, new_n13062, new_n13064);
nor_5  g10716(new_n13064, new_n13061, new_n13065);
nor_5  g10717(new_n13065, new_n13060, new_n13066);
nor_5  g10718(new_n13066, new_n13059, new_n13067);
xnor_4 g10719(new_n9345, n23755, new_n13068);
nor_5  g10720(new_n13068, new_n13067, new_n13069);
nor_5  g10721(new_n13069, new_n13058, new_n13070);
nor_5  g10722(new_n13070, new_n13057, new_n13071);
nor_5  g10723(new_n13071, new_n13056, new_n13072);
nor_5  g10724(new_n13072, new_n13055, new_n13073);
nor_5  g10725(new_n13073, new_n13054_1, new_n13074_1);
nor_5  g10726(new_n13074_1, new_n13053, new_n13075);
nor_5  g10727(new_n13075, new_n13052, new_n13076);
nor_5  g10728(new_n13076, new_n13051, new_n13077);
nor_5  g10729(new_n13077, new_n13050, new_n13078);
nor_5  g10730(new_n13078, new_n13049, new_n13079);
or_5   g10731(new_n13079, new_n13048_1, new_n13080);
xnor_4 g10732(new_n9329, n25586, new_n13081);
xnor_4 g10733(new_n13081, new_n13080, new_n13082_1);
xor_4  g10734(new_n13082_1, n4514, new_n13083);
xor_4  g10735(new_n13078, new_n13049, new_n13084);
nor_5  g10736(new_n13084, n3984, new_n13085);
xnor_4 g10737(new_n13084, n3984, new_n13086);
xor_4  g10738(new_n13076, new_n13051, new_n13087);
nor_5  g10739(new_n13087, n19652, new_n13088);
xnor_4 g10740(new_n13087, n19652, new_n13089);
xor_4  g10741(new_n13074_1, new_n13053, new_n13090);
nor_5  g10742(new_n13090, n3366, new_n13091);
xor_4  g10743(new_n13072, new_n13055, new_n13092);
nor_5  g10744(new_n13092, n26565, new_n13093);
xnor_4 g10745(new_n13092, n26565, new_n13094);
xor_4  g10746(new_n13070, new_n13057, new_n13095);
nor_5  g10747(new_n13095, n3959, new_n13096_1);
xnor_4 g10748(new_n13095, n3959, new_n13097);
xor_4  g10749(new_n13068, new_n13067, new_n13098);
nor_5  g10750(new_n13098, n11566, new_n13099);
xnor_4 g10751(new_n13098, n11566, new_n13100);
xor_4  g10752(new_n13065, new_n13060, new_n13101);
nor_5  g10753(new_n13101, n26744, new_n13102);
xor_4  g10754(new_n13063, new_n13062, new_n13103);
nor_5  g10755(new_n13103, n26625, new_n13104);
and_5  g10756(new_n5983, n14230, new_n13105);
xnor_4 g10757(new_n13103, n26625, new_n13106);
nor_5  g10758(new_n13106, new_n13105, new_n13107);
nor_5  g10759(new_n13107, new_n13104, new_n13108);
xnor_4 g10760(new_n13101, n26744, new_n13109);
nor_5  g10761(new_n13109, new_n13108, new_n13110_1);
nor_5  g10762(new_n13110_1, new_n13102, new_n13111);
nor_5  g10763(new_n13111, new_n13100, new_n13112);
nor_5  g10764(new_n13112, new_n13099, new_n13113);
nor_5  g10765(new_n13113, new_n13097, new_n13114);
nor_5  g10766(new_n13114, new_n13096_1, new_n13115);
nor_5  g10767(new_n13115, new_n13094, new_n13116_1);
nor_5  g10768(new_n13116_1, new_n13093, new_n13117);
xnor_4 g10769(new_n13090, n3366, new_n13118);
nor_5  g10770(new_n13118, new_n13117, new_n13119);
nor_5  g10771(new_n13119, new_n13091, new_n13120);
nor_5  g10772(new_n13120, new_n13089, new_n13121);
nor_5  g10773(new_n13121, new_n13088, new_n13122_1);
nor_5  g10774(new_n13122_1, new_n13086, new_n13123);
nor_5  g10775(new_n13123, new_n13085, new_n13124);
xor_4  g10776(new_n13124, new_n13083, new_n13125);
and_5  g10777(new_n13125, new_n13047, new_n13126);
xnor_4 g10778(new_n13125, new_n13047, new_n13127);
xnor_4 g10779(new_n9303, new_n9273, new_n13128);
xor_4  g10780(new_n13122_1, new_n13086, new_n13129);
nor_5  g10781(new_n13129, new_n13128, new_n13130);
xnor_4 g10782(new_n13129, new_n13128, new_n13131);
xor_4  g10783(new_n13120, new_n13089, new_n13132);
nor_5  g10784(new_n13132, new_n9445_1, new_n13133);
xnor_4 g10785(new_n13132, new_n9445_1, new_n13134);
xnor_4 g10786(new_n9299, new_n9277, new_n13135);
xor_4  g10787(new_n13118, new_n13117, new_n13136);
nor_5  g10788(new_n13136, new_n13135, new_n13137_1);
xnor_4 g10789(new_n13136, new_n13135, new_n13138);
xor_4  g10790(new_n13115, new_n13094, new_n13139);
nor_5  g10791(new_n13139, new_n9452, new_n13140);
xnor_4 g10792(new_n13139, new_n9452, new_n13141_1);
xnor_4 g10793(new_n9295, new_n9281, new_n13142);
xor_4  g10794(new_n13113, new_n13097, new_n13143);
nor_5  g10795(new_n13143, new_n13142, new_n13144_1);
xnor_4 g10796(new_n13143, new_n13142, new_n13145);
xor_4  g10797(new_n9460_1, new_n9283, new_n13146);
xor_4  g10798(new_n13111, new_n13100, new_n13147);
nor_5  g10799(new_n13147, new_n13146, new_n13148);
xnor_4 g10800(new_n13147, new_n13146, new_n13149);
xor_4  g10801(new_n13109, new_n13108, new_n13150);
nor_5  g10802(new_n13150, new_n9466, new_n13151);
xnor_4 g10803(new_n13150, new_n9466, new_n13152);
xor_4  g10804(new_n13106, new_n13105, new_n13153);
nor_5  g10805(new_n13153, new_n5340, new_n13154);
or_5   g10806(new_n5984, new_n5336, new_n13155);
not_10 g10807(new_n13153, new_n13156);
or_5   g10808(new_n13156, new_n5341, new_n13157);
and_5  g10809(new_n13157, new_n13155, new_n13158);
nor_5  g10810(new_n13158, new_n13154, new_n13159);
nor_5  g10811(new_n13159, new_n13152, new_n13160);
nor_5  g10812(new_n13160, new_n13151, new_n13161);
nor_5  g10813(new_n13161, new_n13149, new_n13162);
nor_5  g10814(new_n13162, new_n13148, new_n13163);
nor_5  g10815(new_n13163, new_n13145, new_n13164);
nor_5  g10816(new_n13164, new_n13144_1, new_n13165);
nor_5  g10817(new_n13165, new_n13141_1, new_n13166);
nor_5  g10818(new_n13166, new_n13140, new_n13167);
nor_5  g10819(new_n13167, new_n13138, new_n13168_1);
nor_5  g10820(new_n13168_1, new_n13137_1, new_n13169);
nor_5  g10821(new_n13169, new_n13134, new_n13170);
nor_5  g10822(new_n13170, new_n13133, new_n13171);
nor_5  g10823(new_n13171, new_n13131, new_n13172);
nor_5  g10824(new_n13172, new_n13130, new_n13173);
nor_5  g10825(new_n13173, new_n13127, new_n13174);
nor_5  g10826(new_n13174, new_n13126, new_n13175);
xnor_4 g10827(new_n13175, new_n9432, new_n13176);
and_5  g10828(new_n13082_1, n4514, new_n13177);
and_5  g10829(new_n13124, new_n13083, new_n13178);
nor_5  g10830(new_n13178, new_n13177, new_n13179);
nor_5  g10831(new_n9329, n25586, new_n13180);
nor_5  g10832(new_n13180, new_n13080, new_n13181);
and_5  g10833(new_n9329, n25586, new_n13182);
or_5   g10834(new_n13182, new_n9328, new_n13183);
or_5   g10835(new_n13183, new_n13181, new_n13184);
xnor_4 g10836(new_n13184, new_n13179, new_n13185);
xor_4  g10837(new_n13185, new_n13176, n2826);
and_5  g10838(new_n5692, n5140, new_n13187);
xnor_4 g10839(new_n5692, n5140, new_n13188);
and_5  g10840(new_n5697, n6204, new_n13189);
xnor_4 g10841(new_n5697, n6204, new_n13190_1);
and_5  g10842(new_n5701, n3349, new_n13191);
xnor_4 g10843(new_n5701, n3349, new_n13192);
and_5  g10844(new_n5704_1, n1742, new_n13193);
xnor_4 g10845(new_n5704_1, n1742, new_n13194);
nand_5 g10846(new_n5707, n4858, new_n13195);
or_5   g10847(new_n5710, n8244, new_n13196);
xnor_4 g10848(new_n5710, n8244, new_n13197);
and_5  g10849(new_n5711, n9493, new_n13198_1);
xnor_4 g10850(new_n5711, n9493, new_n13199_1);
and_5  g10851(new_n5713, new_n11106, new_n13200);
nor_5  g10852(new_n5716, new_n11109, new_n13201);
nand_5 g10853(new_n5718, n8656, new_n13202);
xor_4  g10854(new_n5716, n21095, new_n13203);
nor_5  g10855(new_n13203, new_n13202, new_n13204_1);
nor_5  g10856(new_n13204_1, new_n13201, new_n13205);
xnor_4 g10857(new_n5713, n15167, new_n13206);
and_5  g10858(new_n13206, new_n13205, new_n13207);
or_5   g10859(new_n13207, new_n13200, new_n13208);
nor_5  g10860(new_n13208, new_n13199_1, new_n13209_1);
nor_5  g10861(new_n13209_1, new_n13198_1, new_n13210);
not_10 g10862(new_n13210, new_n13211);
or_5   g10863(new_n13211, new_n13197, new_n13212);
nand_5 g10864(new_n13212, new_n13196, new_n13213);
xnor_4 g10865(new_n5707, n4858, new_n13214);
or_5   g10866(new_n13214, new_n13213, new_n13215);
and_5  g10867(new_n13215, new_n13195, new_n13216);
nor_5  g10868(new_n13216, new_n13194, new_n13217);
nor_5  g10869(new_n13217, new_n13193, new_n13218);
nor_5  g10870(new_n13218, new_n13192, new_n13219);
nor_5  g10871(new_n13219, new_n13191, new_n13220);
nor_5  g10872(new_n13220, new_n13190_1, new_n13221);
nor_5  g10873(new_n13221, new_n13189, new_n13222);
nor_5  g10874(new_n13222, new_n13188, new_n13223);
nor_5  g10875(new_n13223, new_n13187, new_n13224);
or_5   g10876(new_n13224, new_n11295, new_n13225);
and_5  g10877(new_n2567, n25365, new_n13226);
nor_5  g10878(new_n2612, new_n2568, new_n13227);
nor_5  g10879(new_n13227, new_n13226, new_n13228);
nor_5  g10880(n20040, n9396, new_n13229);
nor_5  g10881(new_n2566, new_n2533_1, new_n13230);
or_5   g10882(new_n13230, new_n13229, new_n13231);
nor_5  g10883(new_n13231, new_n13228, new_n13232);
xnor_4 g10884(new_n13232, new_n13225, new_n13233);
xnor_4 g10885(new_n13224, new_n11295, new_n13234);
xor_4  g10886(new_n13231, new_n13228, new_n13235);
and_5  g10887(new_n13235, new_n13234, new_n13236);
xnor_4 g10888(new_n13235, new_n13234, new_n13237);
xor_4  g10889(new_n13222, new_n13188, new_n13238);
nor_5  g10890(new_n13238, new_n2613, new_n13239);
xnor_4 g10891(new_n13238, new_n2613, new_n13240);
xnor_4 g10892(new_n2610, new_n2571, new_n13241);
xor_4  g10893(new_n13220, new_n13190_1, new_n13242);
nor_5  g10894(new_n13242, new_n13241, new_n13243);
xnor_4 g10895(new_n13242, new_n13241, new_n13244);
xor_4  g10896(new_n13218, new_n13192, new_n13245);
nor_5  g10897(new_n13245, new_n2716, new_n13246);
xnor_4 g10898(new_n13245, new_n2716, new_n13247);
xor_4  g10899(new_n13216, new_n13194, new_n13248);
nor_5  g10900(new_n13248, new_n2721, new_n13249);
xnor_4 g10901(new_n13248, new_n2721, new_n13250);
xor_4  g10902(new_n13214, new_n13213, new_n13251);
nor_5  g10903(new_n13251, new_n2726, new_n13252);
xnor_4 g10904(new_n13251, new_n2726, new_n13253);
not_10 g10905(new_n2730, new_n13254);
xnor_4 g10906(new_n13210, new_n13197, new_n13255);
and_5  g10907(new_n13255, new_n13254, new_n13256);
xor_4  g10908(new_n13255, new_n2730, new_n13257);
not_10 g10909(new_n2735, new_n13258);
xor_4  g10910(new_n13208, new_n13199_1, new_n13259);
nor_5  g10911(new_n13259, new_n13258, new_n13260);
xor_4  g10912(new_n13259, new_n2735, new_n13261);
xor_4  g10913(new_n13206, new_n13205, new_n13262);
and_5  g10914(new_n13262, new_n2739, new_n13263_1);
xnor_4 g10915(new_n13262, new_n2739, new_n13264);
xor_4  g10916(new_n13203, new_n13202, new_n13265);
nor_5  g10917(new_n13265, new_n2743_1, new_n13266);
xor_4  g10918(new_n5718, n8656, new_n13267);
nor_5  g10919(new_n13267, new_n2746, new_n13268);
xor_4  g10920(new_n13265, new_n2743_1, new_n13269);
and_5  g10921(new_n13269, new_n13268, new_n13270_1);
nor_5  g10922(new_n13270_1, new_n13266, new_n13271);
nor_5  g10923(new_n13271, new_n13264, new_n13272);
nor_5  g10924(new_n13272, new_n13263_1, new_n13273_1);
nor_5  g10925(new_n13273_1, new_n13261, new_n13274);
nor_5  g10926(new_n13274, new_n13260, new_n13275);
nor_5  g10927(new_n13275, new_n13257, new_n13276);
nor_5  g10928(new_n13276, new_n13256, new_n13277);
nor_5  g10929(new_n13277, new_n13253, new_n13278);
nor_5  g10930(new_n13278, new_n13252, new_n13279);
nor_5  g10931(new_n13279, new_n13250, new_n13280);
nor_5  g10932(new_n13280, new_n13249, new_n13281);
nor_5  g10933(new_n13281, new_n13247, new_n13282);
nor_5  g10934(new_n13282, new_n13246, new_n13283);
nor_5  g10935(new_n13283, new_n13244, new_n13284);
nor_5  g10936(new_n13284, new_n13243, new_n13285_1);
nor_5  g10937(new_n13285_1, new_n13240, new_n13286);
nor_5  g10938(new_n13286, new_n13239, new_n13287);
nor_5  g10939(new_n13287, new_n13237, new_n13288);
nor_5  g10940(new_n13288, new_n13236, new_n13289);
xnor_4 g10941(new_n13289, new_n13233, n2853);
xor_4  g10942(n7099, n2035, new_n13291);
not_10 g10943(n12811, new_n13292);
nor_5  g10944(new_n13292, n5213, new_n13293);
xor_4  g10945(n12811, n5213, new_n13294);
not_10 g10946(n1118, new_n13295);
nor_5  g10947(n4665, new_n13295, new_n13296);
xor_4  g10948(n4665, n1118, new_n13297);
nor_5  g10949(n25974, new_n2785, new_n13298);
not_10 g10950(n25974, new_n13299);
nor_5  g10951(new_n13299, n19005, new_n13300);
nor_5  g10952(new_n2789, n1630, new_n13301);
not_10 g10953(n1630, new_n13302);
or_5   g10954(n4326, new_n13302, new_n13303);
nor_5  g10955(new_n2791, n1451, new_n13304);
and_5  g10956(new_n13304, new_n13303, new_n13305);
nor_5  g10957(new_n13305, new_n13301, new_n13306);
nor_5  g10958(new_n13306, new_n13300, new_n13307);
or_5   g10959(new_n13307, new_n13298, new_n13308);
nor_5  g10960(new_n13308, new_n13297, new_n13309);
nor_5  g10961(new_n13309, new_n13296, new_n13310);
nor_5  g10962(new_n13310, new_n13294, new_n13311);
nor_5  g10963(new_n13311, new_n13293, new_n13312);
xor_4  g10964(new_n13312, new_n13291, new_n13313);
or_5   g10965(new_n3937, n13668, new_n13314);
xor_4  g10966(new_n13314, n3570, new_n13315);
xnor_4 g10967(new_n13315, n5337, new_n13316);
and_5  g10968(new_n3938, n626, new_n13317);
nor_5  g10969(new_n3955, new_n3939, new_n13318);
nor_5  g10970(new_n13318, new_n13317, new_n13319_1);
xnor_4 g10971(new_n13319_1, new_n13316, new_n13320);
xor_4  g10972(new_n13320, new_n9992, new_n13321);
and_5  g10973(new_n3956, new_n3934_1, new_n13322);
nor_5  g10974(new_n3979, new_n3957, new_n13323);
nor_5  g10975(new_n13323, new_n13322, new_n13324);
xor_4  g10976(new_n13324, new_n13321, new_n13325);
xnor_4 g10977(new_n13325, new_n13313, new_n13326);
xor_4  g10978(new_n13310, new_n13294, new_n13327);
nor_5  g10979(new_n13327, new_n3980, new_n13328);
xor_4  g10980(new_n13308, new_n13297, new_n13329);
nor_5  g10981(new_n13329, new_n3983_1, new_n13330);
xnor_4 g10982(new_n13329, new_n3983_1, new_n13331);
xnor_4 g10983(n25974, n19005, new_n13332);
xnor_4 g10984(new_n13332, new_n13306, new_n13333_1);
and_5  g10985(new_n13333_1, new_n3986, new_n13334);
xor_4  g10986(new_n13333_1, new_n3986, new_n13335);
xnor_4 g10987(n5438, n1451, new_n13336);
or_5   g10988(new_n13336, new_n3997, new_n13337);
xor_4  g10989(n4326, n1630, new_n13338_1);
xnor_4 g10990(new_n13338_1, new_n13304, new_n13339);
nor_5  g10991(new_n13339, new_n13337, new_n13340);
xor_4  g10992(new_n13339, new_n13337, new_n13341);
and_5  g10993(new_n13341, new_n3990, new_n13342);
nor_5  g10994(new_n13342, new_n13340, new_n13343);
and_5  g10995(new_n13343, new_n13335, new_n13344);
nor_5  g10996(new_n13344, new_n13334, new_n13345);
nor_5  g10997(new_n13345, new_n13331, new_n13346);
or_5   g10998(new_n13346, new_n13330, new_n13347);
xor_4  g10999(new_n13327, new_n3980, new_n13348);
and_5  g11000(new_n13348, new_n13347, new_n13349);
or_5   g11001(new_n13349, new_n13328, new_n13350);
xor_4  g11002(new_n13350, new_n13326, n2860);
xnor_4 g11003(new_n12503, new_n12483, n2887);
or_5   g11004(new_n13314, n3570, new_n13353);
or_5   g11005(new_n13353, n4409, new_n13354);
or_5   g11006(new_n13354, n20359, new_n13355);
or_5   g11007(new_n13355, n2816, new_n13356);
xor_4  g11008(new_n13356, n8526, new_n13357);
nor_5  g11009(new_n13357, n21784, new_n13358);
xor_4  g11010(new_n13355, n2816, new_n13359);
and_5  g11011(new_n13359, n5521, new_n13360);
or_5   g11012(new_n13359, n5521, new_n13361);
xor_4  g11013(new_n13354, n20359, new_n13362);
nor_5  g11014(new_n13362, n11926, new_n13363);
xor_4  g11015(new_n13362, n11926, new_n13364);
xor_4  g11016(new_n13353, n4409, new_n13365);
and_5  g11017(new_n13365, n4325, new_n13366);
nor_5  g11018(new_n13365, n4325, new_n13367_1);
and_5  g11019(new_n13315, n5337, new_n13368);
nor_5  g11020(new_n13315, n5337, new_n13369);
nor_5  g11021(new_n13319_1, new_n13369, new_n13370);
nor_5  g11022(new_n13370, new_n13368, new_n13371);
nor_5  g11023(new_n13371, new_n13367_1, new_n13372);
nor_5  g11024(new_n13372, new_n13366, new_n13373);
and_5  g11025(new_n13373, new_n13364, new_n13374);
nor_5  g11026(new_n13374, new_n13363, new_n13375);
and_5  g11027(new_n13375, new_n13361, new_n13376);
nor_5  g11028(new_n13376, new_n13360, new_n13377);
nor_5  g11029(new_n13377, new_n13358, new_n13378);
nor_5  g11030(new_n13356, n8526, new_n13379);
and_5  g11031(new_n13357, n21784, new_n13380);
or_5   g11032(new_n13380, new_n13379, new_n13381);
nor_5  g11033(new_n13381, new_n13378, new_n13382);
xor_4  g11034(new_n13382, new_n9971, new_n13383);
xor_4  g11035(new_n13357, n21784, new_n13384);
xnor_4 g11036(new_n13384, new_n13377, new_n13385);
and_5  g11037(new_n13385, new_n9975, new_n13386);
xor_4  g11038(new_n13385, new_n9975, new_n13387);
xnor_4 g11039(new_n13359, n5521, new_n13388);
xnor_4 g11040(new_n13388, new_n13375, new_n13389);
nor_5  g11041(new_n13389, new_n9979, new_n13390);
xnor_4 g11042(new_n13389, new_n9979, new_n13391);
xor_4  g11043(new_n13373, new_n13364, new_n13392);
not_10 g11044(new_n13392, new_n13393);
nor_5  g11045(new_n13393, new_n9983, new_n13394);
xor_4  g11046(new_n13365, n4325, new_n13395);
xnor_4 g11047(new_n13395, new_n13371, new_n13396);
and_5  g11048(new_n13396, new_n9987, new_n13397);
xnor_4 g11049(new_n13396, new_n9987, new_n13398);
not_10 g11050(new_n13320, new_n13399);
and_5  g11051(new_n13399, new_n9992, new_n13400);
nor_5  g11052(new_n13324, new_n13321, new_n13401);
nor_5  g11053(new_n13401, new_n13400, new_n13402);
nor_5  g11054(new_n13402, new_n13398, new_n13403);
or_5   g11055(new_n13403, new_n13397, new_n13404);
xor_4  g11056(new_n13392, new_n9983, new_n13405);
nor_5  g11057(new_n13405, new_n13404, new_n13406);
nor_5  g11058(new_n13406, new_n13394, new_n13407_1);
nor_5  g11059(new_n13407_1, new_n13391, new_n13408);
nor_5  g11060(new_n13408, new_n13390, new_n13409_1);
and_5  g11061(new_n13409_1, new_n13387, new_n13410);
nor_5  g11062(new_n13410, new_n13386, new_n13411);
xnor_4 g11063(new_n13411, new_n13383, new_n13412);
not_10 g11064(n8827, new_n13413);
or_5   g11065(new_n3892, n19905, new_n13414);
or_5   g11066(new_n13414, n26452, new_n13415);
or_5   g11067(new_n13415, n15546, new_n13416);
or_5   g11068(new_n13416, n5077, new_n13417);
nor_5  g11069(new_n13417, n18035, new_n13418);
and_5  g11070(new_n13418, new_n13413, new_n13419_1);
xnor_4 g11071(new_n13418, n8827, new_n13420);
nor_5  g11072(new_n13420, n11898, new_n13421);
xor_4  g11073(new_n13417, n18035, new_n13422);
nor_5  g11074(new_n13422, n19941, new_n13423);
xnor_4 g11075(new_n13422, n19941, new_n13424_1);
xor_4  g11076(new_n13416, n5077, new_n13425);
nor_5  g11077(new_n13425, n1099, new_n13426);
xnor_4 g11078(new_n13425, n1099, new_n13427);
xor_4  g11079(new_n13415, n15546, new_n13428);
nor_5  g11080(new_n13428, n2113, new_n13429);
xor_4  g11081(new_n13414, n26452, new_n13430);
nor_5  g11082(new_n13430, n21134, new_n13431);
xnor_4 g11083(new_n13430, n21134, new_n13432);
nor_5  g11084(new_n3893, n6369, new_n13433);
and_5  g11085(new_n3911, new_n3894, new_n13434);
nor_5  g11086(new_n13434, new_n13433, new_n13435);
nor_5  g11087(new_n13435, new_n13432, new_n13436);
nor_5  g11088(new_n13436, new_n13431, new_n13437);
xnor_4 g11089(new_n13428, n2113, new_n13438);
nor_5  g11090(new_n13438, new_n13437, new_n13439);
nor_5  g11091(new_n13439, new_n13429, new_n13440);
nor_5  g11092(new_n13440, new_n13427, new_n13441);
nor_5  g11093(new_n13441, new_n13426, new_n13442);
nor_5  g11094(new_n13442, new_n13424_1, new_n13443);
nor_5  g11095(new_n13443, new_n13423, new_n13444);
and_5  g11096(new_n13420, n11898, new_n13445);
nor_5  g11097(new_n13445, new_n13444, new_n13446);
nor_5  g11098(new_n13446, new_n13421, new_n13447);
nor_5  g11099(new_n13447, new_n13419_1, new_n13448);
xnor_4 g11100(new_n13448, new_n13412, new_n13449);
xor_4  g11101(new_n13409_1, new_n13387, new_n13450);
xor_4  g11102(new_n13420, n11898, new_n13451);
xnor_4 g11103(new_n13451, new_n13444, new_n13452);
not_10 g11104(new_n13452, new_n13453_1);
or_5   g11105(new_n13453_1, new_n13450, new_n13454);
xor_4  g11106(new_n13452, new_n13450, new_n13455);
xnor_4 g11107(new_n13442, new_n13424_1, new_n13456_1);
xnor_4 g11108(new_n13407_1, new_n13391, new_n13457_1);
nor_5  g11109(new_n13457_1, new_n13456_1, new_n13458);
xnor_4 g11110(new_n13457_1, new_n13456_1, new_n13459);
xor_4  g11111(new_n13440, new_n13427, new_n13460_1);
not_10 g11112(new_n13460_1, new_n13461);
xnor_4 g11113(new_n13405, new_n13404, new_n13462);
nor_5  g11114(new_n13462, new_n13461, new_n13463);
xor_4  g11115(new_n13462, new_n13460_1, new_n13464);
xnor_4 g11116(new_n13402, new_n13398, new_n13465);
xor_4  g11117(new_n13438, new_n13437, new_n13466);
and_5  g11118(new_n13466, new_n13465, new_n13467);
xnor_4 g11119(new_n13466, new_n13465, new_n13468);
not_10 g11120(new_n13325, new_n13469);
xor_4  g11121(new_n13435, new_n13432, new_n13470);
and_5  g11122(new_n13470, new_n13469, new_n13471);
xnor_4 g11123(new_n13470, new_n13469, new_n13472);
nor_5  g11124(new_n3980, new_n11679, new_n13473);
and_5  g11125(new_n4004, new_n3981, new_n13474);
nor_5  g11126(new_n13474, new_n13473, new_n13475);
nor_5  g11127(new_n13475, new_n13472, new_n13476);
nor_5  g11128(new_n13476, new_n13471, new_n13477_1);
nor_5  g11129(new_n13477_1, new_n13468, new_n13478);
nor_5  g11130(new_n13478, new_n13467, new_n13479);
nor_5  g11131(new_n13479, new_n13464, new_n13480);
nor_5  g11132(new_n13480, new_n13463, new_n13481);
nor_5  g11133(new_n13481, new_n13459, new_n13482);
nor_5  g11134(new_n13482, new_n13458, new_n13483);
or_5   g11135(new_n13483, new_n13455, new_n13484_1);
nand_5 g11136(new_n13484_1, new_n13454, new_n13485);
xor_4  g11137(new_n13485, new_n13449, n2929);
xor_4  g11138(n22793, n767, new_n13487_1);
not_10 g11139(n7330, new_n13488);
nor_5  g11140(n8439, new_n13488, new_n13489);
xor_4  g11141(n8439, n7330, new_n13490_1);
not_10 g11142(n22492, new_n13491);
nor_5  g11143(n25523, new_n13491, new_n13492);
xor_4  g11144(n25523, n22492, new_n13493);
not_10 g11145(n12821, new_n13494_1);
nor_5  g11146(new_n13494_1, n5579, new_n13495);
xor_4  g11147(n12821, n5579, new_n13496);
not_10 g11148(n3468, new_n13497);
nor_5  g11149(n23430, new_n13497, new_n13498);
xor_4  g11150(n23430, n3468, new_n13499);
not_10 g11151(n10411, new_n13500_1);
nor_5  g11152(n18558, new_n13500_1, new_n13501_1);
nor_5  g11153(new_n12247, new_n12238, new_n13502);
or_5   g11154(new_n13502, new_n13501_1, new_n13503);
nor_5  g11155(new_n13503, new_n13499, new_n13504);
nor_5  g11156(new_n13504, new_n13498, new_n13505);
nor_5  g11157(new_n13505, new_n13496, new_n13506_1);
nor_5  g11158(new_n13506_1, new_n13495, new_n13507);
nor_5  g11159(new_n13507, new_n13493, new_n13508);
nor_5  g11160(new_n13508, new_n13492, new_n13509);
nor_5  g11161(new_n13509, new_n13490_1, new_n13510);
nor_5  g11162(new_n13510, new_n13489, new_n13511);
xor_4  g11163(new_n13511, new_n13487_1, new_n13512);
xnor_4 g11164(new_n13512, new_n6594, new_n13513);
xor_4  g11165(new_n13509, new_n13490_1, new_n13514);
and_5  g11166(new_n13514, new_n6598, new_n13515);
xnor_4 g11167(new_n13514, new_n6598, new_n13516);
xor_4  g11168(new_n13507, new_n13493, new_n13517);
nor_5  g11169(new_n13517, new_n6602, new_n13518);
xnor_4 g11170(new_n13517, new_n6602, new_n13519);
xor_4  g11171(new_n13505, new_n13496, new_n13520);
nor_5  g11172(new_n13520, new_n6605, new_n13521);
xnor_4 g11173(new_n13520, new_n6605, new_n13522);
xor_4  g11174(new_n13503, new_n13499, new_n13523);
and_5  g11175(new_n13523, new_n6608, new_n13524);
xnor_4 g11176(new_n13523, new_n6608, new_n13525);
not_10 g11177(new_n6611_1, new_n13526);
nor_5  g11178(new_n12248, new_n13526, new_n13527);
nor_5  g11179(new_n12524, new_n12515_1, new_n13528);
nor_5  g11180(new_n13528, new_n13527, new_n13529);
nor_5  g11181(new_n13529, new_n13525, new_n13530);
or_5   g11182(new_n13530, new_n13524, new_n13531);
nor_5  g11183(new_n13531, new_n13522, new_n13532);
nor_5  g11184(new_n13532, new_n13521, new_n13533);
nor_5  g11185(new_n13533, new_n13519, new_n13534);
or_5   g11186(new_n13534, new_n13518, new_n13535);
nor_5  g11187(new_n13535, new_n13516, new_n13536);
nor_5  g11188(new_n13536, new_n13515, new_n13537);
xor_4  g11189(new_n13537, new_n13513, new_n13538);
xor_4  g11190(n22379, n15077, new_n13539);
nor_5  g11191(n3710, new_n2768, new_n13540);
xor_4  g11192(n3710, n1662, new_n13541);
nor_5  g11193(n26318, new_n2771, new_n13542);
xor_4  g11194(n26318, n12875, new_n13543);
nor_5  g11195(n26054, new_n2774_1, new_n13544);
xor_4  g11196(n26054, n2035, new_n13545);
nor_5  g11197(n19081, new_n2777, new_n13546);
or_5   g11198(new_n9113, n5213, new_n13547);
nor_5  g11199(new_n9116, n4665, new_n13548_1);
nor_5  g11200(new_n12535, new_n12526, new_n13549_1);
nor_5  g11201(new_n13549_1, new_n13548_1, new_n13550);
and_5  g11202(new_n13550, new_n13547, new_n13551_1);
nor_5  g11203(new_n13551_1, new_n13546, new_n13552);
nor_5  g11204(new_n13552, new_n13545, new_n13553);
nor_5  g11205(new_n13553, new_n13544, new_n13554);
nor_5  g11206(new_n13554, new_n13543, new_n13555);
nor_5  g11207(new_n13555, new_n13542, new_n13556);
nor_5  g11208(new_n13556, new_n13541, new_n13557);
nor_5  g11209(new_n13557, new_n13540, new_n13558);
xor_4  g11210(new_n13558, new_n13539, new_n13559);
xnor_4 g11211(new_n13559, new_n13538, new_n13560);
xor_4  g11212(new_n13556, new_n13541, new_n13561);
xor_4  g11213(new_n13535, new_n13516, new_n13562);
nor_5  g11214(new_n13562, new_n13561, new_n13563);
xnor_4 g11215(new_n13562, new_n13561, new_n13564);
xnor_4 g11216(new_n13554, new_n13543, new_n13565);
xor_4  g11217(new_n13533, new_n13519, new_n13566);
and_5  g11218(new_n13566, new_n13565, new_n13567);
xnor_4 g11219(new_n13566, new_n13565, new_n13568);
xnor_4 g11220(new_n13552, new_n13545, new_n13569);
nor_5  g11221(new_n13530, new_n13524, new_n13570);
xnor_4 g11222(new_n13570, new_n13522, new_n13571);
and_5  g11223(new_n13571, new_n13569, new_n13572);
xor_4  g11224(new_n13529, new_n13525, new_n13573);
xor_4  g11225(n19081, n5213, new_n13574);
xnor_4 g11226(new_n13574, new_n13550, new_n13575);
nor_5  g11227(new_n13575, new_n13573, new_n13576);
xnor_4 g11228(new_n13575, new_n13573, new_n13577);
not_10 g11229(new_n12525, new_n13578);
and_5  g11230(new_n12536, new_n13578, new_n13579);
nor_5  g11231(new_n12555, new_n12537, new_n13580);
nor_5  g11232(new_n13580, new_n13579, new_n13581);
nor_5  g11233(new_n13581, new_n13577, new_n13582);
nor_5  g11234(new_n13582, new_n13576, new_n13583);
xnor_4 g11235(new_n13571, new_n13569, new_n13584);
nor_5  g11236(new_n13584, new_n13583, new_n13585);
nor_5  g11237(new_n13585, new_n13572, new_n13586);
nor_5  g11238(new_n13586, new_n13568, new_n13587);
nor_5  g11239(new_n13587, new_n13567, new_n13588);
nor_5  g11240(new_n13588, new_n13564, new_n13589);
nor_5  g11241(new_n13589, new_n13563, new_n13590);
xnor_4 g11242(new_n13590, new_n13560, n2948);
xor_4  g11243(new_n13034, new_n13018, n2961);
xnor_4 g11244(new_n10268, new_n10246, n2971);
xnor_4 g11245(new_n2515_1, new_n2498, n3010);
xor_4  g11246(new_n6119, new_n6111, n3017);
xor_4  g11247(new_n10582, new_n8193, new_n13596);
xnor_4 g11248(new_n13596, new_n10586, n3020);
xnor_4 g11249(new_n5612, new_n5591, n3067);
xnor_4 g11250(n23541, n19234, new_n13599);
xnor_4 g11251(n27134, n4588, new_n13600);
xnor_4 g11252(new_n13600, new_n13599, new_n13601);
xor_4  g11253(new_n13601, new_n9006, n3076);
nor_5  g11254(n15490, n18, new_n13603);
nand_5 g11255(new_n13603, new_n8287, new_n13604);
xnor_4 g11256(new_n13604, new_n8283, new_n13605);
xnor_4 g11257(new_n13605, n7421, new_n13606);
xnor_4 g11258(new_n13603, n2783, new_n13607);
and_5  g11259(new_n13607, n19680, new_n13608);
xor_4  g11260(new_n13607, n19680, new_n13609);
xor_4  g11261(n15490, n18, new_n13610);
nor_5  g11262(new_n13610, n2809, new_n13611);
nand_5 g11263(n15508, n18, new_n13612);
xor_4  g11264(new_n13610, n2809, new_n13613);
and_5  g11265(new_n13613, new_n13612, new_n13614);
nor_5  g11266(new_n13614, new_n13611, new_n13615);
and_5  g11267(new_n13615, new_n13609, new_n13616);
nor_5  g11268(new_n13616, new_n13608, new_n13617);
xor_4  g11269(new_n13617, new_n13606, new_n13618);
xor_4  g11270(new_n13618, new_n9642, new_n13619);
xnor_4 g11271(new_n13615, new_n13609, new_n13620);
nor_5  g11272(new_n13620, new_n9646_1, new_n13621);
xnor_4 g11273(new_n13620, new_n9646_1, new_n13622);
nor_5  g11274(new_n13613, new_n5327, new_n13623);
xor_4  g11275(new_n13613, new_n13612, new_n13624);
or_5   g11276(new_n13624, new_n9649, new_n13625);
xnor_4 g11277(n15508, n18, new_n13626_1);
or_5   g11278(new_n13626_1, new_n5312, new_n13627);
and_5  g11279(new_n13627, new_n13625, new_n13628);
or_5   g11280(new_n13628, new_n13623, new_n13629);
nor_5  g11281(new_n13629, new_n13622, new_n13630);
nor_5  g11282(new_n13630, new_n13621, new_n13631);
xor_4  g11283(new_n13631, new_n13619, n3089);
xor_4  g11284(new_n4803, new_n4802, n3125);
nor_5  g11285(new_n10325, new_n10322, new_n13634);
xnor_4 g11286(n21839, n19282, new_n13635);
nor_5  g11287(n27089, n12657, new_n13636);
nor_5  g11288(new_n2868, new_n2839, new_n13637);
nor_5  g11289(new_n13637, new_n13636, new_n13638);
xor_4  g11290(new_n13638, new_n13635, new_n13639);
nor_5  g11291(new_n13639, new_n9942_1, new_n13640);
xnor_4 g11292(new_n13639, new_n9942_1, new_n13641);
nor_5  g11293(new_n9945, new_n2869, new_n13642);
nor_5  g11294(new_n9948, new_n2872, new_n13643);
xor_4  g11295(new_n9948, new_n2872, new_n13644);
and_5  g11296(new_n9951, new_n2876, new_n13645);
xnor_4 g11297(new_n9951, new_n2876, new_n13646);
and_5  g11298(new_n9954, new_n2880, new_n13647);
nor_5  g11299(new_n12044, new_n12027, new_n13648);
nor_5  g11300(new_n13648, new_n13647, new_n13649);
nor_5  g11301(new_n13649, new_n13646, new_n13650);
nor_5  g11302(new_n13650, new_n13645, new_n13651);
and_5  g11303(new_n13651, new_n13644, new_n13652);
nor_5  g11304(new_n13652, new_n13643, new_n13653);
xnor_4 g11305(new_n9945, new_n2869, new_n13654);
nor_5  g11306(new_n13654, new_n13653, new_n13655);
nor_5  g11307(new_n13655, new_n13642, new_n13656);
nor_5  g11308(new_n13656, new_n13641, new_n13657);
nor_5  g11309(new_n13657, new_n13640, new_n13658);
nor_5  g11310(n21839, n19282, new_n13659);
nor_5  g11311(new_n13638, new_n13635, new_n13660);
nor_5  g11312(new_n13660, new_n13659, new_n13661);
not_10 g11313(new_n13661, new_n13662);
and_5  g11314(new_n13662, new_n9944, new_n13663);
and_5  g11315(new_n13663, new_n13658, new_n13664);
or_5   g11316(new_n13662, new_n9944, new_n13665);
nor_5  g11317(new_n13665, new_n13658, new_n13666);
nor_5  g11318(new_n13666, new_n13664, new_n13667);
xor_4  g11319(new_n13667, new_n13634, new_n13668_1);
xor_4  g11320(new_n10325, new_n10322, new_n13669);
xnor_4 g11321(new_n13661, new_n9944, new_n13670);
xnor_4 g11322(new_n13670, new_n13658, new_n13671);
nor_5  g11323(new_n13671, new_n13669, new_n13672);
xnor_4 g11324(new_n13671, new_n13669, new_n13673);
xor_4  g11325(new_n13656, new_n13641, new_n13674);
and_5  g11326(new_n13674, new_n10823, new_n13675);
xnor_4 g11327(new_n13674, new_n10823, new_n13676);
xor_4  g11328(new_n13654, new_n13653, new_n13677_1);
and_5  g11329(new_n13677_1, new_n10827, new_n13678);
xor_4  g11330(new_n13677_1, new_n10339, new_n13679);
xor_4  g11331(new_n13651, new_n13644, new_n13680);
and_5  g11332(new_n13680, new_n10346, new_n13681);
xnor_4 g11333(new_n13680, new_n10346, new_n13682);
xor_4  g11334(new_n13649, new_n13646, new_n13683_1);
nor_5  g11335(new_n13683_1, new_n10349, new_n13684);
xor_4  g11336(new_n13683_1, new_n10348, new_n13685);
nor_5  g11337(new_n12045, new_n10353, new_n13686);
nor_5  g11338(new_n12068, new_n12046, new_n13687);
nor_5  g11339(new_n13687, new_n13686, new_n13688);
nor_5  g11340(new_n13688, new_n13685, new_n13689);
nor_5  g11341(new_n13689, new_n13684, new_n13690);
nor_5  g11342(new_n13690, new_n13682, new_n13691);
nor_5  g11343(new_n13691, new_n13681, new_n13692);
nor_5  g11344(new_n13692, new_n13679, new_n13693);
nor_5  g11345(new_n13693, new_n13678, new_n13694);
nor_5  g11346(new_n13694, new_n13676, new_n13695);
nor_5  g11347(new_n13695, new_n13675, new_n13696);
nor_5  g11348(new_n13696, new_n13673, new_n13697);
or_5   g11349(new_n13697, new_n13672, new_n13698);
xnor_4 g11350(new_n13698, new_n13668_1, n3126);
xnor_4 g11351(new_n10868, new_n10833, n3208);
xnor_4 g11352(new_n12874, new_n12872, n3219);
xnor_4 g11353(new_n13271, new_n13264, n3235);
xnor_4 g11354(new_n10143, new_n10130, n3244);
not_10 g11355(n15146, new_n13704);
nor_5  g11356(new_n13704, n5532, new_n13705);
not_10 g11357(new_n8968, new_n13706);
not_10 g11358(n11579, new_n13707);
nor_5  g11359(new_n13707, n3962, new_n13708_1);
not_10 g11360(new_n8965, new_n13709);
not_10 g11361(n21, new_n13710_1);
nor_5  g11362(n23513, new_n13710_1, new_n13711);
not_10 g11363(new_n8949, new_n13712);
and_5  g11364(new_n12257, new_n8996, new_n13713);
not_10 g11365(n1682, new_n13714_1);
nor_5  g11366(n6427, new_n13714_1, new_n13715);
nor_5  g11367(new_n13715, new_n13713, new_n13716);
nor_5  g11368(new_n13716, new_n13712, new_n13717);
nor_5  g11369(new_n13717, new_n13711, new_n13718);
nor_5  g11370(new_n13718, new_n13709, new_n13719_1);
nor_5  g11371(new_n13719_1, new_n13708_1, new_n13720);
nor_5  g11372(new_n13720, new_n13706, new_n13721);
nor_5  g11373(new_n13721, new_n13705, new_n13722_1);
xnor_4 g11374(new_n13722_1, new_n8971_1, new_n13723);
xnor_4 g11375(new_n13723, new_n13514, new_n13724);
xnor_4 g11376(new_n13720, new_n8968, new_n13725);
nor_5  g11377(new_n13725, new_n13517, new_n13726);
xnor_4 g11378(new_n13725, new_n13517, new_n13727);
xnor_4 g11379(new_n13718, new_n8965, new_n13728);
nor_5  g11380(new_n13728, new_n13520, new_n13729);
xnor_4 g11381(new_n13728, new_n13520, new_n13730);
xnor_4 g11382(new_n13716, new_n8949, new_n13731);
nor_5  g11383(new_n13731, new_n13523, new_n13732);
xnor_4 g11384(new_n13731, new_n13523, new_n13733);
nor_5  g11385(new_n12258, new_n12248, new_n13734);
nor_5  g11386(new_n12276, new_n12259, new_n13735);
or_5   g11387(new_n13735, new_n13734, new_n13736);
nor_5  g11388(new_n13736, new_n13733, new_n13737);
nor_5  g11389(new_n13737, new_n13732, new_n13738);
nor_5  g11390(new_n13738, new_n13730, new_n13739);
nor_5  g11391(new_n13739, new_n13729, new_n13740);
nor_5  g11392(new_n13740, new_n13727, new_n13741);
nor_5  g11393(new_n13741, new_n13726, new_n13742);
xnor_4 g11394(new_n13742, new_n13724, new_n13743);
or_5   g11395(n23541, n16247, new_n13744);
or_5   g11396(new_n13744, n8638, new_n13745);
or_5   g11397(new_n13745, n15979, new_n13746);
or_5   g11398(new_n13746, n26483, new_n13747);
or_5   g11399(new_n13747, n24768, new_n13748);
or_5   g11400(new_n13748, n8687, new_n13749);
xor_4  g11401(new_n13749, n19270, new_n13750);
xnor_4 g11402(new_n13750, n18345, new_n13751);
xor_4  g11403(new_n13748, n8687, new_n13752);
nor_5  g11404(new_n13752, n13190, new_n13753);
xnor_4 g11405(new_n13752, n13190, new_n13754_1);
xor_4  g11406(new_n13747, n24768, new_n13755);
nor_5  g11407(new_n13755, n3460, new_n13756);
xnor_4 g11408(new_n13755, n3460, new_n13757);
xor_4  g11409(new_n13746, n26483, new_n13758);
nor_5  g11410(new_n13758, n5226, new_n13759);
xnor_4 g11411(new_n13758, n5226, new_n13760);
xor_4  g11412(new_n13745, n15979, new_n13761);
nor_5  g11413(new_n13761, n17664, new_n13762);
xor_4  g11414(new_n13744, n8638, new_n13763);
nor_5  g11415(new_n13763, n23369, new_n13764_1);
xnor_4 g11416(new_n13763, n23369, new_n13765);
xor_4  g11417(n23541, n16247, new_n13766);
nor_5  g11418(new_n13766, n1136, new_n13767);
nand_5 g11419(n23541, n19234, new_n13768);
xor_4  g11420(new_n13766, n1136, new_n13769);
and_5  g11421(new_n13769, new_n13768, new_n13770);
nor_5  g11422(new_n13770, new_n13767, new_n13771);
nor_5  g11423(new_n13771, new_n13765, new_n13772);
nor_5  g11424(new_n13772, new_n13764_1, new_n13773);
xnor_4 g11425(new_n13761, n17664, new_n13774);
nor_5  g11426(new_n13774, new_n13773, new_n13775_1);
nor_5  g11427(new_n13775_1, new_n13762, new_n13776);
nor_5  g11428(new_n13776, new_n13760, new_n13777);
nor_5  g11429(new_n13777, new_n13759, new_n13778);
nor_5  g11430(new_n13778, new_n13757, new_n13779);
nor_5  g11431(new_n13779, new_n13756, new_n13780);
nor_5  g11432(new_n13780, new_n13754_1, new_n13781_1);
nor_5  g11433(new_n13781_1, new_n13753, new_n13782);
xnor_4 g11434(new_n13782, new_n13751, new_n13783_1);
xnor_4 g11435(new_n13783_1, new_n13743, new_n13784);
xnor_4 g11436(new_n13780, new_n13754_1, new_n13785);
xnor_4 g11437(new_n13740, new_n13727, new_n13786);
nor_5  g11438(new_n13786, new_n13785, new_n13787);
xnor_4 g11439(new_n13778, new_n13757, new_n13788);
xnor_4 g11440(new_n13738, new_n13730, new_n13789);
nor_5  g11441(new_n13789, new_n13788, new_n13790);
xnor_4 g11442(new_n13789, new_n13788, new_n13791);
xnor_4 g11443(new_n13776, new_n13760, new_n13792);
xnor_4 g11444(new_n13736, new_n13733, new_n13793);
nor_5  g11445(new_n13793, new_n13792, new_n13794);
xor_4  g11446(new_n13774, new_n13773, new_n13795);
not_10 g11447(new_n13795, new_n13796);
nor_5  g11448(new_n13796, new_n12277, new_n13797);
xnor_4 g11449(new_n13795, new_n12277, new_n13798_1);
not_10 g11450(new_n12292, new_n13799);
xor_4  g11451(new_n13771, new_n13765, new_n13800);
nor_5  g11452(new_n13800, new_n13799, new_n13801);
xor_4  g11453(new_n13800, new_n12292, new_n13802);
and_5  g11454(n23541, n19234, new_n13803);
xnor_4 g11455(new_n13769, new_n13803, new_n13804);
and_5  g11456(new_n13804, new_n12304_1, new_n13805);
or_5   g11457(new_n13599, new_n12297, new_n13806);
not_10 g11458(new_n13804, new_n13807);
xnor_4 g11459(new_n13807, new_n12304_1, new_n13808);
and_5  g11460(new_n13808, new_n13806, new_n13809);
or_5   g11461(new_n13809, new_n13805, new_n13810);
nor_5  g11462(new_n13810, new_n13802, new_n13811);
nor_5  g11463(new_n13811, new_n13801, new_n13812);
and_5  g11464(new_n13812, new_n13798_1, new_n13813);
nor_5  g11465(new_n13813, new_n13797, new_n13814);
xnor_4 g11466(new_n13793, new_n13792, new_n13815);
nor_5  g11467(new_n13815, new_n13814, new_n13816);
nor_5  g11468(new_n13816, new_n13794, new_n13817);
nor_5  g11469(new_n13817, new_n13791, new_n13818);
nor_5  g11470(new_n13818, new_n13790, new_n13819);
xnor_4 g11471(new_n13786, new_n13785, new_n13820);
nor_5  g11472(new_n13820, new_n13819, new_n13821);
nor_5  g11473(new_n13821, new_n13787, new_n13822);
xnor_4 g11474(new_n13822, new_n13784, n3263);
xnor_4 g11475(new_n11066, new_n11053, n3289);
xnor_4 g11476(n21832, n5211, new_n13825);
and_5  g11477(n26913, n12956, new_n13826);
or_5   g11478(n26913, n12956, new_n13827);
nor_5  g11479(n18295, n16223, new_n13828);
nor_5  g11480(new_n4657, new_n4652, new_n13829);
nor_5  g11481(new_n13829, new_n13828, new_n13830);
and_5  g11482(new_n13830, new_n13827, new_n13831);
or_5   g11483(new_n13831, new_n13826, new_n13832);
xor_4  g11484(new_n13832, new_n13825, new_n13833);
xnor_4 g11485(new_n13833, n18537, new_n13834);
xor_4  g11486(n26913, n12956, new_n13835_1);
xnor_4 g11487(new_n13835_1, new_n13830, new_n13836);
nor_5  g11488(new_n13836, n7057, new_n13837);
xnor_4 g11489(new_n13836, n7057, new_n13838);
nor_5  g11490(new_n4658, n8381, new_n13839);
nor_5  g11491(new_n4668, new_n4659, new_n13840);
nor_5  g11492(new_n13840, new_n13839, new_n13841);
nor_5  g11493(new_n13841, new_n13838, new_n13842);
nor_5  g11494(new_n13842, new_n13837, new_n13843);
xor_4  g11495(new_n13843, new_n13834, new_n13844);
xnor_4 g11496(new_n12939, n21649, new_n13845);
nor_5  g11497(new_n8570, n18274, new_n13846);
xnor_4 g11498(new_n8570, n18274, new_n13847);
nor_5  g11499(new_n8585, n3828, new_n13848);
nor_5  g11500(new_n8589, n23842, new_n13849);
not_10 g11501(n21654, new_n13850_1);
nor_5  g11502(new_n8592, new_n13850_1, new_n13851_1);
xnor_4 g11503(new_n8589, n23842, new_n13852);
nor_5  g11504(new_n13852, new_n13851_1, new_n13853);
nor_5  g11505(new_n13853, new_n13849, new_n13854);
xnor_4 g11506(new_n8585, n3828, new_n13855);
nor_5  g11507(new_n13855, new_n13854, new_n13856);
nor_5  g11508(new_n13856, new_n13848, new_n13857);
nor_5  g11509(new_n13857, new_n13847, new_n13858);
or_5   g11510(new_n13858, new_n13846, new_n13859);
xor_4  g11511(new_n13859, new_n13845, new_n13860);
xor_4  g11512(new_n13860, new_n13844, new_n13861);
xor_4  g11513(new_n13841, new_n13838, new_n13862);
xor_4  g11514(new_n13857, new_n13847, new_n13863);
and_5  g11515(new_n13863, new_n13862, new_n13864);
xnor_4 g11516(new_n13863, new_n13862, new_n13865);
xnor_4 g11517(new_n13855, new_n13854, new_n13866);
nor_5  g11518(new_n13866, new_n4669, new_n13867);
xor_4  g11519(new_n13852, new_n13851_1, new_n13868);
and_5  g11520(new_n13868, new_n4692, new_n13869);
xor_4  g11521(new_n8592, n21654, new_n13870);
or_5   g11522(new_n13870, new_n4695, new_n13871);
xnor_4 g11523(new_n13868, new_n4693_1, new_n13872);
and_5  g11524(new_n13872, new_n13871, new_n13873);
or_5   g11525(new_n13873, new_n13869, new_n13874);
xor_4  g11526(new_n13866, new_n4669, new_n13875);
and_5  g11527(new_n13875, new_n13874, new_n13876);
nor_5  g11528(new_n13876, new_n13867, new_n13877);
nor_5  g11529(new_n13877, new_n13865, new_n13878);
nor_5  g11530(new_n13878, new_n13864, new_n13879);
xnor_4 g11531(new_n13879, new_n13861, n3301);
xor_4  g11532(new_n9686, n3030, new_n13881);
not_10 g11533(n19515, new_n13882);
nor_5  g11534(new_n9679, new_n13882, new_n13883);
xor_4  g11535(new_n9679, n19515, new_n13884);
not_10 g11536(n22588, new_n13885);
nor_5  g11537(new_n9673, new_n13885, new_n13886);
xnor_4 g11538(new_n9673, n22588, new_n13887);
nor_5  g11539(new_n9667, n12209, new_n13888);
and_5  g11540(new_n12074, new_n12073, new_n13889);
nor_5  g11541(new_n13889, new_n13888, new_n13890);
and_5  g11542(new_n13890, new_n13887, new_n13891);
nor_5  g11543(new_n13891, new_n13886, new_n13892);
nor_5  g11544(new_n13892, new_n13884, new_n13893);
nor_5  g11545(new_n13893, new_n13883, new_n13894);
xor_4  g11546(new_n13894, new_n13881, new_n13895);
xnor_4 g11547(new_n13895, new_n9058, new_n13896);
xor_4  g11548(new_n13892, new_n13884, new_n13897);
and_5  g11549(new_n13897, new_n9062, new_n13898);
xnor_4 g11550(new_n13897, new_n9062, new_n13899);
xor_4  g11551(new_n13890, new_n13887, new_n13900);
and_5  g11552(new_n13900, new_n9066, new_n13901);
xnor_4 g11553(new_n13900, new_n9066, new_n13902);
not_10 g11554(new_n12075, new_n13903);
and_5  g11555(new_n13903, new_n9070, new_n13904);
and_5  g11556(new_n12076, new_n12072_1, new_n13905);
nor_5  g11557(new_n13905, new_n13904, new_n13906);
nor_5  g11558(new_n13906, new_n13902, new_n13907);
nor_5  g11559(new_n13907, new_n13901, new_n13908);
nor_5  g11560(new_n13908, new_n13899, new_n13909);
or_5   g11561(new_n13909, new_n13898, new_n13910);
xor_4  g11562(new_n13910, new_n13896, n3316);
xnor_4 g11563(new_n12064, new_n12052, n3332);
nor_5  g11564(new_n7239, n17458, new_n13913);
xnor_4 g11565(new_n7239, n17458, new_n13914_1);
nor_5  g11566(new_n7243, n1222, new_n13915);
xnor_4 g11567(new_n7243, n1222, new_n13916);
nor_5  g11568(new_n7247, n25240, new_n13917);
nor_5  g11569(new_n9508_1, new_n9493_1, new_n13918);
nor_5  g11570(new_n13918, new_n13917, new_n13919);
nor_5  g11571(new_n13919, new_n13916, new_n13920);
nor_5  g11572(new_n13920, new_n13915, new_n13921);
nor_5  g11573(new_n13921, new_n13914_1, new_n13922_1);
or_5   g11574(new_n13922_1, new_n13913, new_n13923_1);
or_5   g11575(new_n13923_1, new_n7298_1, new_n13924);
and_5  g11576(new_n11625, n8827, new_n13925);
nor_5  g11577(new_n11635, new_n11626, new_n13926);
nor_5  g11578(new_n13926, new_n13925, new_n13927);
nor_5  g11579(n23166, n11898, new_n13928);
nor_5  g11580(new_n11624, new_n11617, new_n13929);
or_5   g11581(new_n13929, new_n13928, new_n13930);
nor_5  g11582(new_n13930, new_n13927, new_n13931);
xnor_4 g11583(new_n13931, new_n13924, new_n13932);
xnor_4 g11584(new_n13923_1, new_n7297, new_n13933);
xnor_4 g11585(new_n13930, new_n13927, new_n13934);
nor_5  g11586(new_n13934, new_n13933, new_n13935);
xor_4  g11587(new_n13934, new_n13933, new_n13936);
xor_4  g11588(new_n13921, new_n13914_1, new_n13937);
nor_5  g11589(new_n13937, new_n11636, new_n13938);
xnor_4 g11590(new_n13937, new_n11636, new_n13939);
xor_4  g11591(new_n13919, new_n13916, new_n13940);
and_5  g11592(new_n13940, new_n11639, new_n13941);
nor_5  g11593(new_n9548, new_n9509, new_n13942);
nor_5  g11594(new_n9572, new_n9549, new_n13943);
nor_5  g11595(new_n13943, new_n13942, new_n13944);
xnor_4 g11596(new_n13940, new_n11639, new_n13945);
nor_5  g11597(new_n13945, new_n13944, new_n13946);
or_5   g11598(new_n13946, new_n13941, new_n13947);
nor_5  g11599(new_n13947, new_n13939, new_n13948);
nor_5  g11600(new_n13948, new_n13938, new_n13949);
and_5  g11601(new_n13949, new_n13936, new_n13950);
nor_5  g11602(new_n13950, new_n13935, new_n13951_1);
xnor_4 g11603(new_n13951_1, new_n13932, n3340);
xor_4  g11604(n13851, n5077, new_n13953);
not_10 g11605(n15546, new_n13954);
nor_5  g11606(n24937, new_n13954, new_n13955);
xor_4  g11607(n24937, n15546, new_n13956);
not_10 g11608(n26452, new_n13957);
or_5   g11609(new_n13957, n5098, new_n13958);
xor_4  g11610(n26452, n5098, new_n13959);
not_10 g11611(n19905, new_n13960);
or_5   g11612(new_n13960, n3030, new_n13961);
xor_4  g11613(n19905, n3030, new_n13962);
nor_5  g11614(new_n13882, n17035, new_n13963);
nor_5  g11615(new_n12289, new_n12278, new_n13964);
nor_5  g11616(new_n13964, new_n13963, new_n13965);
not_10 g11617(new_n13965, new_n13966);
or_5   g11618(new_n13966, new_n13962, new_n13967);
and_5  g11619(new_n13967, new_n13961, new_n13968);
or_5   g11620(new_n13968, new_n13959, new_n13969);
and_5  g11621(new_n13969, new_n13958, new_n13970);
nor_5  g11622(new_n13970, new_n13956, new_n13971);
nor_5  g11623(new_n13971, new_n13955, new_n13972);
xor_4  g11624(new_n13972, new_n13953, new_n13973);
xnor_4 g11625(new_n13973, new_n13743, new_n13974);
xor_4  g11626(new_n13970, new_n13956, new_n13975);
nor_5  g11627(new_n13975, new_n13786, new_n13976);
xnor_4 g11628(new_n13975, new_n13786, new_n13977);
xor_4  g11629(new_n13968, new_n13959, new_n13978);
nor_5  g11630(new_n13978, new_n13789, new_n13979);
xor_4  g11631(new_n13978, new_n13789, new_n13980);
xnor_4 g11632(new_n13965, new_n13962, new_n13981);
and_5  g11633(new_n13981, new_n13793, new_n13982);
xnor_4 g11634(new_n13981, new_n13793, new_n13983);
nor_5  g11635(new_n12290, new_n12277, new_n13984);
nor_5  g11636(new_n12309, new_n12291, new_n13985);
or_5   g11637(new_n13985, new_n13984, new_n13986);
nor_5  g11638(new_n13986, new_n13983, new_n13987);
nor_5  g11639(new_n13987, new_n13982, new_n13988);
and_5  g11640(new_n13988, new_n13980, new_n13989);
nor_5  g11641(new_n13989, new_n13979, new_n13990);
nor_5  g11642(new_n13990, new_n13977, new_n13991);
or_5   g11643(new_n13991, new_n13976, new_n13992);
xor_4  g11644(new_n13992, new_n13974, n3343);
or_5   g11645(new_n13749, n19270, new_n13994);
or_5   g11646(new_n13994, n14704, new_n13995);
nor_5  g11647(new_n13995, n25365, new_n13996);
xor_4  g11648(new_n13995, n25365, new_n13997);
nor_5  g11649(new_n13997, n20040, new_n13998);
xor_4  g11650(new_n13994, n14704, new_n13999);
nor_5  g11651(new_n13999, n19531, new_n14000);
xnor_4 g11652(new_n13999, n19531, new_n14001);
nor_5  g11653(new_n13750, n18345, new_n14002);
nor_5  g11654(new_n13782, new_n13751, new_n14003);
nor_5  g11655(new_n14003, new_n14002, new_n14004_1);
nor_5  g11656(new_n14004_1, new_n14001, new_n14005);
nor_5  g11657(new_n14005, new_n14000, new_n14006);
and_5  g11658(new_n13997, n20040, new_n14007);
nor_5  g11659(new_n14007, new_n14006, new_n14008);
nor_5  g11660(new_n14008, new_n13998, new_n14009);
nor_5  g11661(new_n14009, new_n13996, new_n14010);
xor_4  g11662(new_n13997, n20040, new_n14011);
xnor_4 g11663(new_n14011, new_n14006, new_n14012);
not_10 g11664(new_n14012, new_n14013);
and_5  g11665(new_n14013, new_n12614, new_n14014);
nor_5  g11666(new_n14013, new_n12614, new_n14015);
xor_4  g11667(new_n14004_1, new_n14001, new_n14016);
not_10 g11668(new_n14016, new_n14017);
and_5  g11669(new_n14017, new_n12600, new_n14018);
xnor_4 g11670(new_n14017, new_n12600, new_n14019);
and_5  g11671(new_n13783_1, new_n12602, new_n14020);
xnor_4 g11672(new_n13783_1, new_n12602, new_n14021);
and_5  g11673(new_n13785, new_n5884, new_n14022);
xnor_4 g11674(new_n13785, new_n5884, new_n14023);
and_5  g11675(new_n13788, new_n5886, new_n14024);
and_5  g11676(new_n13792, new_n5889, new_n14025);
xor_4  g11677(new_n13792, new_n5889, new_n14026);
nor_5  g11678(new_n13796, new_n5893, new_n14027);
xnor_4 g11679(new_n13795, new_n5893, new_n14028);
not_10 g11680(new_n5895, new_n14029);
nor_5  g11681(new_n13800, new_n14029, new_n14030);
xnor_4 g11682(new_n13800, new_n5895, new_n14031);
nor_5  g11683(new_n13807, new_n5898, new_n14032);
nor_5  g11684(new_n13599, new_n11154, new_n14033);
xor_4  g11685(new_n13804, new_n5898, new_n14034);
nor_5  g11686(new_n14034, new_n14033, new_n14035);
nor_5  g11687(new_n14035, new_n14032, new_n14036_1);
and_5  g11688(new_n14036_1, new_n14031, new_n14037);
nor_5  g11689(new_n14037, new_n14030, new_n14038);
and_5  g11690(new_n14038, new_n14028, new_n14039);
nor_5  g11691(new_n14039, new_n14027, new_n14040);
and_5  g11692(new_n14040, new_n14026, new_n14041);
nor_5  g11693(new_n14041, new_n14025, new_n14042);
xnor_4 g11694(new_n13788, new_n5886, new_n14043);
nor_5  g11695(new_n14043, new_n14042, new_n14044);
nor_5  g11696(new_n14044, new_n14024, new_n14045);
nor_5  g11697(new_n14045, new_n14023, new_n14046);
nor_5  g11698(new_n14046, new_n14022, new_n14047);
nor_5  g11699(new_n14047, new_n14021, new_n14048);
nor_5  g11700(new_n14048, new_n14020, new_n14049);
nor_5  g11701(new_n14049, new_n14019, new_n14050);
nor_5  g11702(new_n14050, new_n14018, new_n14051);
nor_5  g11703(new_n14051, new_n14015, new_n14052);
or_5   g11704(new_n14052, new_n12636, new_n14053);
or_5   g11705(new_n14053, new_n14014, new_n14054);
xnor_4 g11706(new_n14054, new_n14010, new_n14055);
nor_5  g11707(new_n11233, n10250, new_n14056);
xnor_4 g11708(new_n11233, n10250, new_n14057);
nor_5  g11709(new_n11237, n7674, new_n14058);
xnor_4 g11710(new_n11237, n7674, new_n14059_1);
nor_5  g11711(new_n11241, n6397, new_n14060);
xnor_4 g11712(new_n11241, n6397, new_n14061);
nor_5  g11713(new_n11245_1, n19196, new_n14062);
xnor_4 g11714(new_n11245_1, n19196, new_n14063);
nor_5  g11715(new_n11249, n23586, new_n14064);
xnor_4 g11716(new_n11249, n23586, new_n14065);
nor_5  g11717(new_n11253, n21226, new_n14066);
xnor_4 g11718(new_n11253, n21226, new_n14067);
nor_5  g11719(new_n11257, n4426, new_n14068);
xnor_4 g11720(new_n11257, n4426, new_n14069);
nor_5  g11721(new_n11263, n20036, new_n14070);
xnor_4 g11722(new_n11263, new_n7878, new_n14071_1);
and_5  g11723(new_n11270, n11192, new_n14072);
or_5   g11724(new_n11267, n9380, new_n14073);
xnor_4 g11725(new_n11270, new_n3851, new_n14074);
and_5  g11726(new_n14074, new_n14073, new_n14075);
nor_5  g11727(new_n14075, new_n14072, new_n14076);
and_5  g11728(new_n14076, new_n14071_1, new_n14077);
nor_5  g11729(new_n14077, new_n14070, new_n14078);
nor_5  g11730(new_n14078, new_n14069, new_n14079);
nor_5  g11731(new_n14079, new_n14068, new_n14080);
nor_5  g11732(new_n14080, new_n14067, new_n14081_1);
nor_5  g11733(new_n14081_1, new_n14066, new_n14082);
nor_5  g11734(new_n14082, new_n14065, new_n14083);
nor_5  g11735(new_n14083, new_n14064, new_n14084);
nor_5  g11736(new_n14084, new_n14063, new_n14085);
nor_5  g11737(new_n14085, new_n14062, new_n14086);
nor_5  g11738(new_n14086, new_n14061, new_n14087);
nor_5  g11739(new_n14087, new_n14060, new_n14088);
nor_5  g11740(new_n14088, new_n14059_1, new_n14089);
nor_5  g11741(new_n14089, new_n14058, new_n14090_1);
nor_5  g11742(new_n14090_1, new_n14057, new_n14091);
or_5   g11743(new_n14091, new_n14056, new_n14092);
xor_4  g11744(new_n14092, new_n11132_1, new_n14093);
nor_5  g11745(new_n14093, new_n14055, new_n14094);
xnor_4 g11746(new_n14090_1, new_n14057, new_n14095_1);
xnor_4 g11747(new_n14012, new_n12614, new_n14096);
xnor_4 g11748(new_n14096, new_n14051, new_n14097);
nor_5  g11749(new_n14097, new_n14095_1, new_n14098);
xnor_4 g11750(new_n14097, new_n14095_1, new_n14099);
xnor_4 g11751(new_n14088, new_n14059_1, new_n14100);
xor_4  g11752(new_n14049, new_n14019, new_n14101);
nor_5  g11753(new_n14101, new_n14100, new_n14102);
xnor_4 g11754(new_n14101, new_n14100, new_n14103);
xnor_4 g11755(new_n14086, new_n14061, new_n14104);
xor_4  g11756(new_n14047, new_n14021, new_n14105);
nor_5  g11757(new_n14105, new_n14104, new_n14106);
xnor_4 g11758(new_n14105, new_n14104, new_n14107_1);
xnor_4 g11759(new_n14084, new_n14063, new_n14108);
xor_4  g11760(new_n14045, new_n14023, new_n14109);
nor_5  g11761(new_n14109, new_n14108, new_n14110);
xnor_4 g11762(new_n14109, new_n14108, new_n14111);
xnor_4 g11763(new_n14082, new_n14065, new_n14112);
xor_4  g11764(new_n14043, new_n14042, new_n14113);
nor_5  g11765(new_n14113, new_n14112, new_n14114);
xnor_4 g11766(new_n14113, new_n14112, new_n14115);
xnor_4 g11767(new_n14080, new_n14067, new_n14116);
xor_4  g11768(new_n14040, new_n14026, new_n14117);
nor_5  g11769(new_n14117, new_n14116, new_n14118);
xnor_4 g11770(new_n14117, new_n14116, new_n14119);
xor_4  g11771(new_n14078, new_n14069, new_n14120);
xor_4  g11772(new_n14038, new_n14028, new_n14121_1);
and_5  g11773(new_n14121_1, new_n14120, new_n14122);
xnor_4 g11774(new_n14121_1, new_n14120, new_n14123);
xnor_4 g11775(new_n14076, new_n14071_1, new_n14124);
xor_4  g11776(new_n14036_1, new_n14031, new_n14125);
nor_5  g11777(new_n14125, new_n14124, new_n14126_1);
xor_4  g11778(new_n14034, new_n14033, new_n14127);
not_10 g11779(new_n14127, new_n14128);
xor_4  g11780(new_n14074, new_n14073, new_n14129);
and_5  g11781(new_n14129, new_n14128, new_n14130_1);
xnor_4 g11782(new_n13599, n4939, new_n14131);
xnor_4 g11783(new_n11267, n9380, new_n14132);
nand_5 g11784(new_n14132, new_n14131, new_n14133);
xnor_4 g11785(new_n14129, new_n14128, new_n14134);
nor_5  g11786(new_n14134, new_n14133, new_n14135);
nor_5  g11787(new_n14135, new_n14130_1, new_n14136_1);
not_10 g11788(new_n14125, new_n14137);
xnor_4 g11789(new_n14137, new_n14124, new_n14138);
and_5  g11790(new_n14138, new_n14136_1, new_n14139);
nor_5  g11791(new_n14139, new_n14126_1, new_n14140);
nor_5  g11792(new_n14140, new_n14123, new_n14141);
nor_5  g11793(new_n14141, new_n14122, new_n14142);
nor_5  g11794(new_n14142, new_n14119, new_n14143);
nor_5  g11795(new_n14143, new_n14118, new_n14144);
nor_5  g11796(new_n14144, new_n14115, new_n14145);
nor_5  g11797(new_n14145, new_n14114, new_n14146);
nor_5  g11798(new_n14146, new_n14111, new_n14147_1);
nor_5  g11799(new_n14147_1, new_n14110, new_n14148_1);
nor_5  g11800(new_n14148_1, new_n14107_1, new_n14149);
nor_5  g11801(new_n14149, new_n14106, new_n14150);
nor_5  g11802(new_n14150, new_n14103, new_n14151);
nor_5  g11803(new_n14151, new_n14102, new_n14152);
nor_5  g11804(new_n14152, new_n14099, new_n14153);
nor_5  g11805(new_n14153, new_n14098, new_n14154);
xnor_4 g11806(new_n14093, new_n14055, new_n14155);
nor_5  g11807(new_n14155, new_n14154, new_n14156);
nor_5  g11808(new_n14156, new_n14094, new_n14157);
or_5   g11809(new_n14054, new_n14010, new_n14158);
or_5   g11810(new_n14092, new_n11132_1, new_n14159);
xor_4  g11811(new_n14159, new_n14158, new_n14160);
xnor_4 g11812(new_n14160, new_n14157, n3390);
xnor_4 g11813(new_n5971, new_n5970, n3426);
xor_4  g11814(new_n4387, new_n4386, n3451);
xnor_4 g11815(new_n10976, new_n10959, n3459);
xnor_4 g11816(n6773, n583, new_n14165);
xor_4  g11817(new_n14165, n21687, new_n14166);
or_5   g11818(new_n14166, new_n12387, new_n14167);
and_5  g11819(new_n14165, n21687, new_n14168);
nor_5  g11820(new_n14168, n6729, new_n14169);
and_5  g11821(n21687, n6729, new_n14170);
and_5  g11822(new_n14165, new_n14170, new_n14171);
or_5   g11823(new_n14171, new_n14169, new_n14172);
and_5  g11824(n6773, n583, new_n14173);
xnor_4 g11825(n22173, n17090, new_n14174_1);
xnor_4 g11826(new_n14174_1, new_n14173, new_n14175);
xor_4  g11827(new_n14175, new_n14172, new_n14176);
xor_4  g11828(new_n14176, new_n12383_1, new_n14177);
xnor_4 g11829(new_n14177, new_n14167, n3502);
xnor_4 g11830(new_n9808, new_n9775, n3516);
nor_5  g11831(n24129, n22274, new_n14180);
not_10 g11832(new_n14180, new_n14181);
nor_5  g11833(new_n14181, n1689, new_n14182);
not_10 g11834(new_n14182, new_n14183);
or_5   g11835(new_n14183, n19608, new_n14184);
or_5   g11836(new_n14184, n25126, new_n14185);
or_5   g11837(new_n14185, n10712, new_n14186);
xnor_4 g11838(new_n14186, n18145, new_n14187);
xnor_4 g11839(new_n14187, n15761, new_n14188);
xnor_4 g11840(new_n14185, n10712, new_n14189);
and_5  g11841(new_n14189, n11201, new_n14190_1);
xnor_4 g11842(new_n14189, n11201, new_n14191);
xnor_4 g11843(new_n14184, n25126, new_n14192);
and_5  g11844(new_n14192, n18690, new_n14193);
xnor_4 g11845(new_n14192, n18690, new_n14194);
xor_4  g11846(new_n14182, n19608, new_n14195);
and_5  g11847(new_n14195, n12153, new_n14196);
xnor_4 g11848(new_n14195, n12153, new_n14197);
xnor_4 g11849(new_n14180, n1689, new_n14198);
nor_5  g11850(new_n14198, new_n9284, new_n14199);
xor_4  g11851(new_n14198, n13044, new_n14200);
xnor_4 g11852(n24129, n22274, new_n14201);
and_5  g11853(new_n14201, n18745, new_n14202);
or_5   g11854(n24129, new_n5338, new_n14203);
xnor_4 g11855(new_n14201, n18745, new_n14204);
nor_5  g11856(new_n14204, new_n14203, new_n14205);
nor_5  g11857(new_n14205, new_n14202, new_n14206);
nor_5  g11858(new_n14206, new_n14200, new_n14207);
nor_5  g11859(new_n14207, new_n14199, new_n14208);
nor_5  g11860(new_n14208, new_n14197, new_n14209);
nor_5  g11861(new_n14209, new_n14196, new_n14210);
nor_5  g11862(new_n14210, new_n14194, new_n14211_1);
nor_5  g11863(new_n14211_1, new_n14193, new_n14212);
nor_5  g11864(new_n14212, new_n14191, new_n14213);
nor_5  g11865(new_n14213, new_n14190_1, new_n14214);
xnor_4 g11866(new_n14214, new_n14188, new_n14215);
xnor_4 g11867(new_n14215, new_n6227, new_n14216);
xnor_4 g11868(new_n14212, new_n14191, new_n14217);
nor_5  g11869(new_n14217, new_n6230, new_n14218);
xnor_4 g11870(new_n14217, new_n6230, new_n14219);
xnor_4 g11871(new_n14210, new_n14194, new_n14220);
nor_5  g11872(new_n14220, new_n6233_1, new_n14221);
xnor_4 g11873(new_n14220, new_n6233_1, new_n14222_1);
xnor_4 g11874(new_n14208, new_n14197, new_n14223);
nor_5  g11875(new_n14223, new_n6237, new_n14224);
xor_4  g11876(new_n14223, new_n6237, new_n14225);
xor_4  g11877(new_n14206, new_n14200, new_n14226);
nor_5  g11878(new_n14226, new_n3848, new_n14227);
xnor_4 g11879(new_n14226, new_n3848, new_n14228);
xor_4  g11880(new_n14204, new_n14203, new_n14229);
nor_5  g11881(new_n14229, new_n3860, new_n14230_1);
xnor_4 g11882(n24129, n16167, new_n14231);
or_5   g11883(new_n14231, new_n3865, new_n14232);
xnor_4 g11884(new_n14229, new_n3860, new_n14233);
nor_5  g11885(new_n14233, new_n14232, new_n14234);
nor_5  g11886(new_n14234, new_n14230_1, new_n14235);
nor_5  g11887(new_n14235, new_n14228, new_n14236);
nor_5  g11888(new_n14236, new_n14227, new_n14237);
and_5  g11889(new_n14237, new_n14225, new_n14238);
nor_5  g11890(new_n14238, new_n14224, new_n14239);
nor_5  g11891(new_n14239, new_n14222_1, new_n14240);
nor_5  g11892(new_n14240, new_n14221, new_n14241);
nor_5  g11893(new_n14241, new_n14219, new_n14242);
nor_5  g11894(new_n14242, new_n14218, new_n14243);
xor_4  g11895(new_n14243, new_n14216, new_n14244);
xnor_4 g11896(new_n14244, new_n9389, new_n14245);
xor_4  g11897(new_n14241, new_n14219, new_n14246);
and_5  g11898(new_n14246, new_n9394, new_n14247);
xnor_4 g11899(new_n14246, new_n9394, new_n14248);
xor_4  g11900(new_n14239, new_n14222_1, new_n14249);
and_5  g11901(new_n14249, new_n9398, new_n14250);
xnor_4 g11902(new_n14249, new_n9398, new_n14251);
not_10 g11903(new_n9404, new_n14252);
xor_4  g11904(new_n14237, new_n14225, new_n14253);
and_5  g11905(new_n14253, new_n14252, new_n14254);
xor_4  g11906(new_n14235, new_n14228, new_n14255);
nor_5  g11907(new_n14255, new_n9407, new_n14256);
xnor_4 g11908(new_n14255, new_n9407, new_n14257);
xor_4  g11909(new_n14233, new_n14232, new_n14258);
nor_5  g11910(new_n14258, new_n5345, new_n14259);
xor_4  g11911(new_n14231, new_n3864, new_n14260);
or_5   g11912(new_n14260, new_n5334, new_n14261);
xor_4  g11913(new_n14258, new_n5345, new_n14262);
and_5  g11914(new_n14262, new_n14261, new_n14263);
nor_5  g11915(new_n14263, new_n14259, new_n14264);
nor_5  g11916(new_n14264, new_n14257, new_n14265);
nor_5  g11917(new_n14265, new_n14256, new_n14266);
xnor_4 g11918(new_n14253, new_n14252, new_n14267_1);
nor_5  g11919(new_n14267_1, new_n14266, new_n14268);
nor_5  g11920(new_n14268, new_n14254, new_n14269);
nor_5  g11921(new_n14269, new_n14251, new_n14270);
nor_5  g11922(new_n14270, new_n14250, new_n14271_1);
nor_5  g11923(new_n14271_1, new_n14248, new_n14272);
or_5   g11924(new_n14272, new_n14247, new_n14273);
xor_4  g11925(new_n14273, new_n14245, n3528);
xnor_4 g11926(new_n8252, new_n8198, n3555);
nor_5  g11927(new_n9165, new_n2622, new_n14276);
nor_5  g11928(new_n2709, new_n2658, new_n14277_1);
nor_5  g11929(new_n14277_1, new_n14276, new_n14278);
or_5   g11930(new_n2621, n13951, new_n14279);
or_5   g11931(new_n9163, new_n14279, new_n14280);
nor_5  g11932(new_n14280, new_n14278, new_n14281);
and_5  g11933(new_n9163, new_n14279, new_n14282);
and_5  g11934(new_n14282, new_n14278, new_n14283);
nor_5  g11935(new_n14283, new_n14281, new_n14284);
nor_5  g11936(new_n14284, new_n13232, new_n14285);
xnor_4 g11937(new_n14284, new_n13232, new_n14286);
xnor_4 g11938(new_n9163, new_n14279, new_n14287);
xnor_4 g11939(new_n14287, new_n14278, new_n14288);
nor_5  g11940(new_n14288, new_n13235, new_n14289);
xnor_4 g11941(new_n14288, new_n13235, new_n14290);
xor_4  g11942(new_n2612, new_n2568, new_n14291);
nor_5  g11943(new_n2710, new_n14291, new_n14292);
and_5  g11944(new_n2765, new_n2711_1, new_n14293);
nor_5  g11945(new_n14293, new_n14292, new_n14294_1);
nor_5  g11946(new_n14294_1, new_n14290, new_n14295);
nor_5  g11947(new_n14295, new_n14289, new_n14296);
nor_5  g11948(new_n14296, new_n14286, new_n14297);
nor_5  g11949(new_n14297, new_n14285, new_n14298);
nor_5  g11950(new_n14298, new_n14281, n3561);
xor_4  g11951(n16439, n14680, new_n14300);
nor_5  g11952(new_n6980, n15241, new_n14301);
nor_5  g11953(new_n9593, new_n9574, new_n14302);
nor_5  g11954(new_n14302, new_n14301, new_n14303);
xor_4  g11955(new_n14303, new_n14300, new_n14304);
xnor_4 g11956(new_n8750, n1654, new_n14305);
nor_5  g11957(new_n8753, n13783, new_n14306);
nor_5  g11958(new_n9606, new_n9595, new_n14307);
nor_5  g11959(new_n14307, new_n14306, new_n14308);
xor_4  g11960(new_n14308, new_n14305, new_n14309);
xor_4  g11961(new_n14309, new_n14304, new_n14310_1);
not_10 g11962(new_n9594, new_n14311);
nor_5  g11963(new_n9607, new_n14311, new_n14312);
nor_5  g11964(new_n9634, new_n9608, new_n14313);
nor_5  g11965(new_n14313, new_n14312, new_n14314);
xor_4  g11966(new_n14314, new_n14310_1, new_n14315);
xnor_4 g11967(new_n14315, new_n5178, new_n14316);
nor_5  g11968(new_n9635_1, new_n5183, new_n14317);
nor_5  g11969(new_n9661, new_n9636, new_n14318);
nor_5  g11970(new_n14318, new_n14317, new_n14319);
xor_4  g11971(new_n14319, new_n14316, n3563);
xor_4  g11972(new_n5606, new_n5605_1, n3617);
xor_4  g11973(new_n10232, new_n10211, new_n14322);
xor_4  g11974(n22253, n8305, new_n14323_1);
not_10 g11975(n1255, new_n14324);
nor_5  g11976(n12861, new_n14324, new_n14325);
xor_4  g11977(n12861, n1255, new_n14326_1);
not_10 g11978(n9512, new_n14327);
nor_5  g11979(n13333, new_n14327, new_n14328);
xor_4  g11980(n13333, n9512, new_n14329);
not_10 g11981(n16608, new_n14330);
nor_5  g11982(new_n14330, n2210, new_n14331);
not_10 g11983(n21735, new_n14332);
nor_5  g11984(new_n14332, n20604, new_n14333);
nor_5  g11985(new_n4290, new_n4268, new_n14334);
nor_5  g11986(new_n14334, new_n14333, new_n14335);
xor_4  g11987(n16608, n2210, new_n14336);
nor_5  g11988(new_n14336, new_n14335, new_n14337);
nor_5  g11989(new_n14337, new_n14331, new_n14338);
nor_5  g11990(new_n14338, new_n14329, new_n14339);
nor_5  g11991(new_n14339, new_n14328, new_n14340);
nor_5  g11992(new_n14340, new_n14326_1, new_n14341);
nor_5  g11993(new_n14341, new_n14325, new_n14342_1);
xor_4  g11994(new_n14342_1, new_n14323_1, new_n14343);
xnor_4 g11995(new_n14343, new_n14322, new_n14344);
xor_4  g11996(new_n14340, new_n14326_1, new_n14345_1);
nor_5  g11997(new_n14345_1, new_n10236_1, new_n14346);
xnor_4 g11998(new_n14345_1, new_n10236_1, new_n14347);
xor_4  g11999(new_n14338, new_n14329, new_n14348);
nor_5  g12000(new_n14348, new_n10240, new_n14349);
xor_4  g12001(new_n14336, new_n14335, new_n14350);
and_5  g12002(new_n14350, new_n10244_1, new_n14351);
xnor_4 g12003(new_n14350, new_n10244_1, new_n14352);
and_5  g12004(new_n4372, new_n4291, new_n14353_1);
nor_5  g12005(new_n4402, new_n4373, new_n14354);
nor_5  g12006(new_n14354, new_n14353_1, new_n14355);
nor_5  g12007(new_n14355, new_n14352, new_n14356);
nor_5  g12008(new_n14356, new_n14351, new_n14357);
xor_4  g12009(new_n14348, new_n10240, new_n14358);
and_5  g12010(new_n14358, new_n14357, new_n14359);
nor_5  g12011(new_n14359, new_n14349, new_n14360);
nor_5  g12012(new_n14360, new_n14347, new_n14361);
or_5   g12013(new_n14361, new_n14346, new_n14362);
xor_4  g12014(new_n14362, new_n14344, n3642);
xnor_4 g12015(n16544, n4319, new_n14364_1);
nor_5  g12016(n23463, n6814, new_n14365);
xnor_4 g12017(n23463, n6814, new_n14366);
nor_5  g12018(n19701, n13074, new_n14367);
xnor_4 g12019(n19701, n13074, new_n14368);
nor_5  g12020(n23529, n10739, new_n14369);
xnor_4 g12021(n23529, n10739, new_n14370);
nor_5  g12022(n24620, n21753, new_n14371);
xnor_4 g12023(n24620, n21753, new_n14372);
nor_5  g12024(n21832, n5211, new_n14373);
nor_5  g12025(new_n13832, new_n13825, new_n14374);
nor_5  g12026(new_n14374, new_n14373, new_n14375_1);
nor_5  g12027(new_n14375_1, new_n14372, new_n14376);
nor_5  g12028(new_n14376, new_n14371, new_n14377);
nor_5  g12029(new_n14377, new_n14370, new_n14378);
nor_5  g12030(new_n14378, new_n14369, new_n14379);
nor_5  g12031(new_n14379, new_n14368, new_n14380);
nor_5  g12032(new_n14380, new_n14367, new_n14381);
nor_5  g12033(new_n14381, new_n14366, new_n14382);
nor_5  g12034(new_n14382, new_n14365, new_n14383);
xor_4  g12035(new_n14383, new_n14364_1, new_n14384);
xnor_4 g12036(new_n14384, n3324, new_n14385);
xor_4  g12037(new_n14381, new_n14366, new_n14386);
or_5   g12038(new_n14386, n17911, new_n14387);
xnor_4 g12039(new_n14386, n17911, new_n14388);
xor_4  g12040(new_n14379, new_n14368, new_n14389);
or_5   g12041(new_n14389, n21997, new_n14390);
xnor_4 g12042(new_n14389, n21997, new_n14391);
xor_4  g12043(new_n14377, new_n14370, new_n14392);
or_5   g12044(new_n14392, n25119, new_n14393);
xnor_4 g12045(new_n14392, n25119, new_n14394);
xor_4  g12046(new_n14375_1, new_n14372, new_n14395);
and_5  g12047(new_n14395, n1163, new_n14396);
nor_5  g12048(new_n13833, n18537, new_n14397);
nor_5  g12049(new_n13843, new_n13834, new_n14398);
or_5   g12050(new_n14398, new_n14397, new_n14399);
xnor_4 g12051(new_n14395, n1163, new_n14400);
nor_5  g12052(new_n14400, new_n14399, new_n14401);
nor_5  g12053(new_n14401, new_n14396, new_n14402);
not_10 g12054(new_n14402, new_n14403);
or_5   g12055(new_n14403, new_n14394, new_n14404);
and_5  g12056(new_n14404, new_n14393, new_n14405);
or_5   g12057(new_n14405, new_n14391, new_n14406);
and_5  g12058(new_n14406, new_n14390, new_n14407);
or_5   g12059(new_n14407, new_n14388, new_n14408);
and_5  g12060(new_n14408, new_n14387, new_n14409);
xor_4  g12061(new_n14409, new_n14385, new_n14410);
xor_4  g12062(n23250, n16507, new_n14411);
not_10 g12063(n11455, new_n14412_1);
nor_5  g12064(n22470, new_n14412_1, new_n14413);
xor_4  g12065(n22470, n11455, new_n14414_1);
not_10 g12066(n3945, new_n14415);
nor_5  g12067(n19116, new_n14415, new_n14416);
xor_4  g12068(n19116, n3945, new_n14417);
not_10 g12069(n5255, new_n14418);
nor_5  g12070(n6861, new_n14418, new_n14419);
xor_4  g12071(n6861, n5255, new_n14420);
nor_5  g12072(new_n4768, n19357, new_n14421);
xor_4  g12073(n21649, n19357, new_n14422);
nor_5  g12074(new_n4771, n2328, new_n14423);
not_10 g12075(n15053, new_n14424);
nor_5  g12076(new_n14424, n3828, new_n14425);
not_10 g12077(new_n4681, new_n14426);
nor_5  g12078(new_n4686, new_n14426, new_n14427);
nor_5  g12079(new_n14427, new_n14425, new_n14428);
xnor_4 g12080(n18274, n2328, new_n14429);
and_5  g12081(new_n14429, new_n14428, new_n14430);
nor_5  g12082(new_n14430, new_n14423, new_n14431);
nor_5  g12083(new_n14431, new_n14422, new_n14432);
nor_5  g12084(new_n14432, new_n14421, new_n14433);
nor_5  g12085(new_n14433, new_n14420, new_n14434);
nor_5  g12086(new_n14434, new_n14419, new_n14435);
nor_5  g12087(new_n14435, new_n14417, new_n14436);
nor_5  g12088(new_n14436, new_n14416, new_n14437);
nor_5  g12089(new_n14437, new_n14414_1, new_n14438);
nor_5  g12090(new_n14438, new_n14413, new_n14439);
xor_4  g12091(new_n14439, new_n14411, new_n14440_1);
nor_5  g12092(new_n14440_1, n4967, new_n14441);
xnor_4 g12093(new_n14440_1, n4967, new_n14442);
xor_4  g12094(new_n14437, new_n14414_1, new_n14443);
nor_5  g12095(new_n14443, n15602, new_n14444);
xor_4  g12096(new_n14435, new_n14417, new_n14445);
and_5  g12097(new_n14445, n8694, new_n14446);
xor_4  g12098(new_n14433, new_n14420, new_n14447);
nor_5  g12099(new_n14447, n12380, new_n14448);
not_10 g12100(n12380, new_n14449);
xnor_4 g12101(new_n14447, new_n14449, new_n14450);
not_10 g12102(new_n14450, new_n14451);
xor_4  g12103(new_n14431, new_n14422, new_n14452);
nor_5  g12104(new_n14452, n8943, new_n14453);
not_10 g12105(n8943, new_n14454);
xnor_4 g12106(new_n14452, new_n14454, new_n14455);
not_10 g12107(new_n14429, new_n14456);
xnor_4 g12108(new_n14456, new_n14428, new_n14457_1);
and_5  g12109(new_n14457_1, n8255, new_n14458);
not_10 g12110(n11184, new_n14459);
nor_5  g12111(new_n4687, new_n14459, new_n14460);
not_10 g12112(new_n4688, new_n14461);
nor_5  g12113(new_n14461, new_n4680, new_n14462);
nor_5  g12114(new_n14462, new_n14460, new_n14463);
not_10 g12115(n8255, new_n14464_1);
xnor_4 g12116(new_n14457_1, new_n14464_1, new_n14465);
not_10 g12117(new_n14465, new_n14466);
nor_5  g12118(new_n14466, new_n14463, new_n14467);
nor_5  g12119(new_n14467, new_n14458, new_n14468);
and_5  g12120(new_n14468, new_n14455, new_n14469);
nor_5  g12121(new_n14469, new_n14453, new_n14470);
nor_5  g12122(new_n14470, new_n14451, new_n14471_1);
nor_5  g12123(new_n14471_1, new_n14448, new_n14472);
not_10 g12124(n8694, new_n14473);
xnor_4 g12125(new_n14445, new_n14473, new_n14474);
and_5  g12126(new_n14474, new_n14472, new_n14475_1);
nor_5  g12127(new_n14475_1, new_n14446, new_n14476);
not_10 g12128(n15602, new_n14477);
xnor_4 g12129(new_n14443, new_n14477, new_n14478);
and_5  g12130(new_n14478, new_n14476, new_n14479);
nor_5  g12131(new_n14479, new_n14444, new_n14480);
nor_5  g12132(new_n14480, new_n14442, new_n14481);
nor_5  g12133(new_n14481, new_n14441, new_n14482);
xor_4  g12134(n6659, n5101, new_n14483);
not_10 g12135(n23250, new_n14484);
nor_5  g12136(new_n14484, n16507, new_n14485);
nor_5  g12137(new_n14439, new_n14411, new_n14486);
nor_5  g12138(new_n14486, new_n14485, new_n14487);
xor_4  g12139(new_n14487, new_n14483, new_n14488);
xnor_4 g12140(new_n14488, n13419, new_n14489);
xor_4  g12141(new_n14489, new_n14482, new_n14490);
xnor_4 g12142(new_n14490, new_n14410, new_n14491);
xor_4  g12143(new_n14407, new_n14388, new_n14492);
xor_4  g12144(new_n14480, new_n14442, new_n14493);
and_5  g12145(new_n14493, new_n14492, new_n14494);
xnor_4 g12146(new_n14493, new_n14492, new_n14495);
xor_4  g12147(new_n14405, new_n14391, new_n14496);
xor_4  g12148(new_n14478, new_n14476, new_n14497);
and_5  g12149(new_n14497, new_n14496, new_n14498);
xnor_4 g12150(new_n14497, new_n14496, new_n14499);
xnor_4 g12151(new_n14402, new_n14394, new_n14500);
not_10 g12152(new_n14500, new_n14501);
xor_4  g12153(new_n14474, new_n14472, new_n14502);
nor_5  g12154(new_n14502, new_n14501, new_n14503);
xnor_4 g12155(new_n14502, new_n14501, new_n14504);
xor_4  g12156(new_n14470, new_n14450, new_n14505);
xor_4  g12157(new_n14400, new_n14399, new_n14506);
nor_5  g12158(new_n14506, new_n14505, new_n14507);
xnor_4 g12159(new_n14506, new_n14505, new_n14508);
xor_4  g12160(new_n14468, new_n14455, new_n14509);
and_5  g12161(new_n14509, new_n13844, new_n14510_1);
xnor_4 g12162(new_n14509, new_n13844, new_n14511);
not_10 g12163(new_n13862, new_n14512);
xnor_4 g12164(new_n14465, new_n14463, new_n14513);
nor_5  g12165(new_n14513, new_n14512, new_n14514);
xnor_4 g12166(new_n14513, new_n14512, new_n14515);
nor_5  g12167(new_n4689, new_n4669, new_n14516);
nor_5  g12168(new_n4701, new_n4690, new_n14517);
nor_5  g12169(new_n14517, new_n14516, new_n14518);
nor_5  g12170(new_n14518, new_n14515, new_n14519);
nor_5  g12171(new_n14519, new_n14514, new_n14520);
nor_5  g12172(new_n14520, new_n14511, new_n14521);
nor_5  g12173(new_n14521, new_n14510_1, new_n14522);
nor_5  g12174(new_n14522, new_n14508, new_n14523);
nor_5  g12175(new_n14523, new_n14507, new_n14524);
nor_5  g12176(new_n14524, new_n14504, new_n14525);
nor_5  g12177(new_n14525, new_n14503, new_n14526);
nor_5  g12178(new_n14526, new_n14499, new_n14527);
nor_5  g12179(new_n14527, new_n14498, new_n14528);
nor_5  g12180(new_n14528, new_n14495, new_n14529);
or_5   g12181(new_n14529, new_n14494, new_n14530);
xor_4  g12182(new_n14530, new_n14491, n3649);
not_10 g12183(n7917, new_n14532);
nor_5  g12184(n26625, n14230, new_n14533);
not_10 g12185(new_n14533, new_n14534);
nor_5  g12186(new_n14534, n26744, new_n14535);
not_10 g12187(new_n14535, new_n14536);
or_5   g12188(new_n14536, n11566, new_n14537);
or_5   g12189(new_n14537, n3959, new_n14538);
or_5   g12190(new_n14538, n26565, new_n14539);
xnor_4 g12191(new_n14539, n3366, new_n14540);
xnor_4 g12192(new_n14540, n26191, new_n14541_1);
xnor_4 g12193(new_n14538, n26565, new_n14542);
nor_5  g12194(new_n14542, n26512, new_n14543);
xnor_4 g12195(new_n14542, n26512, new_n14544);
nor_5  g12196(new_n14536, n11566, new_n14545);
xor_4  g12197(new_n14545, n3959, new_n14546_1);
nor_5  g12198(new_n14546_1, n19575, new_n14547_1);
xnor_4 g12199(new_n14546_1, n19575, new_n14548);
not_10 g12200(n15378, new_n14549);
xnor_4 g12201(new_n14535, n11566, new_n14550);
and_5  g12202(new_n14550, new_n14549, new_n14551);
xnor_4 g12203(new_n14550, new_n14549, new_n14552);
xor_4  g12204(new_n14533, n26744, new_n14553);
nor_5  g12205(new_n14553, n17095, new_n14554);
xnor_4 g12206(n26625, n14230, new_n14555);
and_5  g12207(new_n14555, n22591, new_n14556);
nor_5  g12208(new_n8677, n14230, new_n14557);
xor_4  g12209(new_n14555, n22591, new_n14558);
and_5  g12210(new_n14558, new_n14557, new_n14559);
or_5   g12211(new_n14559, new_n14556, new_n14560);
xnor_4 g12212(new_n14553, n17095, new_n14561);
nor_5  g12213(new_n14561, new_n14560, new_n14562);
nor_5  g12214(new_n14562, new_n14554, new_n14563);
nor_5  g12215(new_n14563, new_n14552, new_n14564);
nor_5  g12216(new_n14564, new_n14551, new_n14565);
nor_5  g12217(new_n14565, new_n14548, new_n14566);
nor_5  g12218(new_n14566, new_n14547_1, new_n14567);
nor_5  g12219(new_n14567, new_n14544, new_n14568);
nor_5  g12220(new_n14568, new_n14543, new_n14569);
xor_4  g12221(new_n14569, new_n14541_1, new_n14570_1);
xnor_4 g12222(new_n14570_1, new_n14532, new_n14571);
not_10 g12223(n17302, new_n14572);
xor_4  g12224(new_n14567, new_n14544, new_n14573);
and_5  g12225(new_n14573, new_n14572, new_n14574);
xnor_4 g12226(new_n14573, new_n14572, new_n14575_1);
not_10 g12227(n2013, new_n14576_1);
xor_4  g12228(new_n14565, new_n14548, new_n14577);
nor_5  g12229(new_n14577, new_n14576_1, new_n14578);
xnor_4 g12230(new_n14577, new_n14576_1, new_n14579);
not_10 g12231(n23755, new_n14580);
xor_4  g12232(new_n14563, new_n14552, new_n14581);
nor_5  g12233(new_n14581, new_n14580, new_n14582);
xnor_4 g12234(new_n14581, new_n14580, new_n14583);
not_10 g12235(n19163, new_n14584);
xor_4  g12236(new_n14561, new_n14560, new_n14585);
nor_5  g12237(new_n14585, new_n14584, new_n14586);
xnor_4 g12238(new_n14585, new_n14584, new_n14587);
xor_4  g12239(new_n14558, new_n14557, new_n14588);
and_5  g12240(new_n14588, n22358, new_n14589);
nor_5  g12241(new_n14588, n22358, new_n14590);
xnor_4 g12242(n26167, n14230, new_n14591);
nand_5 g12243(new_n14591, n9646, new_n14592);
nor_5  g12244(new_n14592, new_n14590, new_n14593_1);
nor_5  g12245(new_n14593_1, new_n14589, new_n14594);
nor_5  g12246(new_n14594, new_n14587, new_n14595);
nor_5  g12247(new_n14595, new_n14586, new_n14596);
nor_5  g12248(new_n14596, new_n14583, new_n14597);
nor_5  g12249(new_n14597, new_n14582, new_n14598);
nor_5  g12250(new_n14598, new_n14579, new_n14599);
or_5   g12251(new_n14599, new_n14578, new_n14600);
nor_5  g12252(new_n14600, new_n14575_1, new_n14601);
nor_5  g12253(new_n14601, new_n14574, new_n14602);
xor_4  g12254(new_n14602, new_n14571, new_n14603_1);
xnor_4 g12255(new_n14603_1, new_n6266, new_n14604);
xor_4  g12256(new_n14600, new_n14575_1, new_n14605);
nor_5  g12257(new_n14605, new_n6270, new_n14606);
xnor_4 g12258(new_n14605, new_n6270, new_n14607);
xor_4  g12259(new_n14598, new_n14579, new_n14608);
and_5  g12260(new_n14608, new_n6273, new_n14609);
xnor_4 g12261(new_n14608, new_n6273, new_n14610);
xor_4  g12262(new_n14596, new_n14583, new_n14611);
and_5  g12263(new_n14611, new_n6277, new_n14612);
xnor_4 g12264(new_n14611, new_n6277, new_n14613);
not_10 g12265(new_n6282, new_n14614);
xor_4  g12266(new_n14594, new_n14587, new_n14615);
and_5  g12267(new_n14615, new_n14614, new_n14616);
xnor_4 g12268(new_n14615, new_n6282, new_n14617);
xor_4  g12269(new_n14588, n22358, new_n14618);
xnor_4 g12270(new_n14618, new_n14592, new_n14619);
nor_5  g12271(new_n14619, new_n6286, new_n14620);
xnor_4 g12272(new_n14591, n9646, new_n14621);
nand_5 g12273(new_n14621, new_n6288, new_n14622);
xnor_4 g12274(new_n14619, new_n6286, new_n14623);
nor_5  g12275(new_n14623, new_n14622, new_n14624);
nor_5  g12276(new_n14624, new_n14620, new_n14625);
and_5  g12277(new_n14625, new_n14617, new_n14626);
nor_5  g12278(new_n14626, new_n14616, new_n14627);
nor_5  g12279(new_n14627, new_n14613, new_n14628);
nor_5  g12280(new_n14628, new_n14612, new_n14629);
nor_5  g12281(new_n14629, new_n14610, new_n14630);
nor_5  g12282(new_n14630, new_n14609, new_n14631);
nor_5  g12283(new_n14631, new_n14607, new_n14632);
nor_5  g12284(new_n14632, new_n14606, new_n14633_1);
xnor_4 g12285(new_n14633_1, new_n14604, n3665);
xor_4  g12286(new_n5336, new_n5335, n3679);
or_5   g12287(n16521, n7139, new_n14636_1);
or_5   g12288(new_n14636_1, n16824, new_n14637);
or_5   g12289(new_n14637, n604, new_n14638);
or_5   g12290(new_n14638, n4913, new_n14639);
or_5   g12291(new_n14639, n9172, new_n14640);
nor_5  g12292(new_n14640, n442, new_n14641);
and_5  g12293(new_n14641, new_n3356, new_n14642);
xnor_4 g12294(new_n14642, new_n3353, new_n14643);
xnor_4 g12295(new_n14643, new_n5434, new_n14644);
xnor_4 g12296(new_n14641, n13719, new_n14645);
and_5  g12297(new_n14645, new_n5439_1, new_n14646);
xnor_4 g12298(new_n14645, new_n5439_1, new_n14647);
xor_4  g12299(new_n14640, n442, new_n14648);
nor_5  g12300(new_n14648, new_n5444, new_n14649);
xnor_4 g12301(new_n14648, new_n5444, new_n14650);
xor_4  g12302(new_n14639, n9172, new_n14651);
nor_5  g12303(new_n14651, new_n5448, new_n14652);
xnor_4 g12304(new_n14651, new_n5448, new_n14653);
xor_4  g12305(new_n14638, n4913, new_n14654);
nor_5  g12306(new_n14654, new_n5453, new_n14655);
xnor_4 g12307(new_n14654, new_n5453, new_n14656);
xor_4  g12308(new_n14637, n604, new_n14657);
nor_5  g12309(new_n14657, new_n5457, new_n14658);
xnor_4 g12310(new_n14657, new_n5457, new_n14659);
xor_4  g12311(new_n14636_1, n16824, new_n14660);
nor_5  g12312(new_n14660, new_n5462, new_n14661);
xnor_4 g12313(new_n14660, new_n5462, new_n14662);
nor_5  g12314(new_n14636_1, new_n5466, new_n14663);
nor_5  g12315(new_n5465, n7139, new_n14664);
xnor_4 g12316(new_n14664, n16521, new_n14665);
nor_5  g12317(new_n14665, new_n5469, new_n14666);
nor_5  g12318(new_n14666, new_n14663, new_n14667);
nor_5  g12319(new_n14667, new_n14662, new_n14668);
nor_5  g12320(new_n14668, new_n14661, new_n14669);
nor_5  g12321(new_n14669, new_n14659, new_n14670);
nor_5  g12322(new_n14670, new_n14658, new_n14671);
nor_5  g12323(new_n14671, new_n14656, new_n14672);
nor_5  g12324(new_n14672, new_n14655, new_n14673);
nor_5  g12325(new_n14673, new_n14653, new_n14674);
nor_5  g12326(new_n14674, new_n14652, new_n14675);
nor_5  g12327(new_n14675, new_n14650, new_n14676);
or_5   g12328(new_n14676, new_n14649, new_n14677);
nor_5  g12329(new_n14677, new_n14647, new_n14678);
nor_5  g12330(new_n14678, new_n14646, new_n14679);
xnor_4 g12331(new_n14679, new_n14644, new_n14680_1);
xor_4  g12332(new_n5528, n2858, new_n14681);
and_5  g12333(new_n5531, n2659, new_n14682);
xnor_4 g12334(new_n5531, n2659, new_n14683);
and_5  g12335(new_n5534, n24327, new_n14684_1);
nor_5  g12336(new_n7735, new_n7714, new_n14685);
nor_5  g12337(new_n14685, new_n14684_1, new_n14686);
nor_5  g12338(new_n14686, new_n14683, new_n14687);
nor_5  g12339(new_n14687, new_n14682, new_n14688);
xor_4  g12340(new_n14688, new_n14681, new_n14689);
xnor_4 g12341(new_n14689, new_n14680_1, new_n14690);
xor_4  g12342(new_n14686, new_n14683, new_n14691);
xor_4  g12343(new_n14677, new_n14647, new_n14692_1);
nor_5  g12344(new_n14692_1, new_n14691, new_n14693);
xnor_4 g12345(new_n14692_1, new_n14691, new_n14694);
not_10 g12346(new_n7736, new_n14695);
xor_4  g12347(new_n14675, new_n14650, new_n14696);
and_5  g12348(new_n14696, new_n14695, new_n14697);
xor_4  g12349(new_n14696, new_n7736, new_n14698);
xor_4  g12350(new_n14673, new_n14653, new_n14699);
and_5  g12351(new_n14699, new_n7761, new_n14700);
xnor_4 g12352(new_n14699, new_n7761, new_n14701_1);
not_10 g12353(new_n7766, new_n14702_1);
xor_4  g12354(new_n14671, new_n14656, new_n14703);
and_5  g12355(new_n14703, new_n14702_1, new_n14704_1);
xor_4  g12356(new_n14703, new_n7766, new_n14705);
xnor_4 g12357(new_n14669, new_n14659, new_n14706);
nor_5  g12358(new_n14706, new_n7770, new_n14707);
xor_4  g12359(new_n14706, new_n7770, new_n14708);
not_10 g12360(new_n7774, new_n14709);
xor_4  g12361(new_n14667, new_n14662, new_n14710);
nor_5  g12362(new_n14710, new_n14709, new_n14711);
xor_4  g12363(new_n14710, new_n7774, new_n14712);
xor_4  g12364(new_n14665, new_n5469, new_n14713);
and_5  g12365(new_n14713, new_n7777, new_n14714);
xnor_4 g12366(new_n5465, n7139, new_n14715);
or_5   g12367(new_n14715, new_n7782, new_n14716);
xor_4  g12368(new_n14713, new_n7777, new_n14717);
and_5  g12369(new_n14717, new_n14716, new_n14718);
or_5   g12370(new_n14718, new_n14714, new_n14719);
nor_5  g12371(new_n14719, new_n14712, new_n14720);
nor_5  g12372(new_n14720, new_n14711, new_n14721);
and_5  g12373(new_n14721, new_n14708, new_n14722);
nor_5  g12374(new_n14722, new_n14707, new_n14723);
nor_5  g12375(new_n14723, new_n14705, new_n14724);
nor_5  g12376(new_n14724, new_n14704_1, new_n14725);
nor_5  g12377(new_n14725, new_n14701_1, new_n14726);
nor_5  g12378(new_n14726, new_n14700, new_n14727);
nor_5  g12379(new_n14727, new_n14698, new_n14728);
nor_5  g12380(new_n14728, new_n14697, new_n14729);
nor_5  g12381(new_n14729, new_n14694, new_n14730);
nor_5  g12382(new_n14730, new_n14693, new_n14731);
xnor_4 g12383(new_n14731, new_n14690, n3725);
not_10 g12384(new_n13382, new_n14733);
nor_5  g12385(n11220, n3425, new_n14734_1);
nor_5  g12386(new_n11758, new_n11755, new_n14735);
nor_5  g12387(new_n14735, new_n14734_1, new_n14736);
nor_5  g12388(n7335, n2160, new_n14737);
nor_5  g12389(new_n11753, new_n11750, new_n14738);
nor_5  g12390(new_n14738, new_n14737, new_n14739);
xor_4  g12391(new_n14739, new_n14736, new_n14740);
nor_5  g12392(new_n11759, new_n11754, new_n14741);
nor_5  g12393(new_n11763, new_n11760, new_n14742);
nor_5  g12394(new_n14742, new_n14741, new_n14743);
xnor_4 g12395(new_n14743, new_n14740, new_n14744);
xnor_4 g12396(new_n14744, new_n14733, new_n14745);
xor_4  g12397(new_n11763, new_n11760, new_n14746_1);
nor_5  g12398(new_n13385, new_n14746_1, new_n14747);
xnor_4 g12399(new_n13385, new_n11764, new_n14748);
and_5  g12400(new_n13389, new_n4975, new_n14749);
xnor_4 g12401(new_n13389, new_n4975, new_n14750);
and_5  g12402(new_n13393, new_n4978, new_n14751);
xnor_4 g12403(new_n4970, new_n4935, new_n14752);
nor_5  g12404(new_n13396, new_n14752, new_n14753);
xor_4  g12405(new_n13396, new_n4982, new_n14754);
and_5  g12406(new_n13320, new_n4986, new_n14755);
xnor_4 g12407(new_n13320, new_n4986, new_n14756);
nor_5  g12408(new_n4990, new_n3956, new_n14757);
nor_5  g12409(new_n4993, new_n3960, new_n14758);
xnor_4 g12410(new_n4993, new_n3960, new_n14759);
nor_5  g12411(new_n4998, new_n3963, new_n14760);
xnor_4 g12412(new_n4998, new_n3963, new_n14761);
nor_5  g12413(new_n5001, new_n3965, new_n14762);
nor_5  g12414(new_n5002, new_n3949, new_n14763_1);
or_5   g12415(new_n5007, new_n3967, new_n14764);
nor_5  g12416(new_n14764, new_n14763_1, new_n14765);
nor_5  g12417(new_n14765, new_n14762, new_n14766);
nor_5  g12418(new_n14766, new_n14761, new_n14767);
nor_5  g12419(new_n14767, new_n14760, new_n14768);
nor_5  g12420(new_n14768, new_n14759, new_n14769);
nor_5  g12421(new_n14769, new_n14758, new_n14770);
not_10 g12422(new_n3956, new_n14771);
xnor_4 g12423(new_n4990, new_n14771, new_n14772_1);
and_5  g12424(new_n14772_1, new_n14770, new_n14773);
nor_5  g12425(new_n14773, new_n14757, new_n14774);
nor_5  g12426(new_n14774, new_n14756, new_n14775);
nor_5  g12427(new_n14775, new_n14755, new_n14776);
nor_5  g12428(new_n14776, new_n14754, new_n14777);
or_5   g12429(new_n14777, new_n14753, new_n14778);
xnor_4 g12430(new_n13393, new_n4978, new_n14779);
nor_5  g12431(new_n14779, new_n14778, new_n14780);
nor_5  g12432(new_n14780, new_n14751, new_n14781);
nor_5  g12433(new_n14781, new_n14750, new_n14782);
nor_5  g12434(new_n14782, new_n14749, new_n14783);
and_5  g12435(new_n14783, new_n14748, new_n14784);
nor_5  g12436(new_n14784, new_n14747, new_n14785);
xnor_4 g12437(new_n14785, new_n14745, n3733);
xor_4  g12438(new_n9700, n24937, new_n14787);
and_5  g12439(new_n9694, n5098, new_n14788);
xor_4  g12440(new_n9693, n5098, new_n14789);
and_5  g12441(new_n9687, n3030, new_n14790_1);
nor_5  g12442(new_n13894, new_n13881, new_n14791);
nor_5  g12443(new_n14791, new_n14790_1, new_n14792);
nor_5  g12444(new_n14792, new_n14789, new_n14793);
nor_5  g12445(new_n14793, new_n14788, new_n14794);
xor_4  g12446(new_n14794, new_n14787, new_n14795);
xnor_4 g12447(new_n14795, new_n9050, new_n14796);
xor_4  g12448(new_n14792, new_n14789, new_n14797);
nor_5  g12449(new_n14797, new_n9054, new_n14798);
xnor_4 g12450(new_n14797, new_n9054, new_n14799);
nor_5  g12451(new_n13895, new_n9058, new_n14800);
nor_5  g12452(new_n13910, new_n13896, new_n14801_1);
nor_5  g12453(new_n14801_1, new_n14800, new_n14802);
nor_5  g12454(new_n14802, new_n14799, new_n14803);
nor_5  g12455(new_n14803, new_n14798, new_n14804);
xor_4  g12456(new_n14804, new_n14796, n3755);
xnor_4 g12457(new_n8244_1, new_n8214, n3758);
not_10 g12458(new_n10773, new_n14807);
not_10 g12459(n2570, new_n14808);
or_5   g12460(new_n14186, n18145, new_n14809);
or_5   g12461(new_n14809, n655, new_n14810);
nor_5  g12462(new_n14810, n19033, new_n14811);
xnor_4 g12463(new_n14811, new_n14808, new_n14812);
xnor_4 g12464(new_n14812, n14692, new_n14813);
xnor_4 g12465(new_n14810, n19033, new_n14814);
and_5  g12466(new_n14814, n4100, new_n14815);
xnor_4 g12467(new_n14814, n4100, new_n14816);
xnor_4 g12468(new_n14809, n655, new_n14817);
and_5  g12469(new_n14817, n21957, new_n14818);
xnor_4 g12470(new_n14817, n21957, new_n14819_1);
and_5  g12471(new_n14187, n15761, new_n14820);
nor_5  g12472(new_n14214, new_n14188, new_n14821);
nor_5  g12473(new_n14821, new_n14820, new_n14822);
nor_5  g12474(new_n14822, new_n14819_1, new_n14823);
nor_5  g12475(new_n14823, new_n14818, new_n14824);
nor_5  g12476(new_n14824, new_n14816, new_n14825);
nor_5  g12477(new_n14825, new_n14815, new_n14826_1);
xor_4  g12478(new_n14826_1, new_n14813, new_n14827_1);
and_5  g12479(new_n14827_1, new_n14807, new_n14828);
xnor_4 g12480(new_n14827_1, new_n14807, new_n14829);
xnor_4 g12481(new_n14824, new_n14816, new_n14830);
nor_5  g12482(new_n14830, new_n6222, new_n14831);
xnor_4 g12483(new_n14830, new_n6222, new_n14832);
xnor_4 g12484(new_n14822, new_n14819_1, new_n14833);
nor_5  g12485(new_n14833, new_n6224, new_n14834);
xnor_4 g12486(new_n14833, new_n6224, new_n14835);
nor_5  g12487(new_n14215, new_n6227, new_n14836);
nor_5  g12488(new_n14243, new_n14216, new_n14837);
nor_5  g12489(new_n14837, new_n14836, new_n14838);
nor_5  g12490(new_n14838, new_n14835, new_n14839_1);
nor_5  g12491(new_n14839_1, new_n14834, new_n14840);
nor_5  g12492(new_n14840, new_n14832, new_n14841);
nor_5  g12493(new_n14841, new_n14831, new_n14842);
nor_5  g12494(new_n14842, new_n14829, new_n14843);
or_5   g12495(new_n14843, new_n14828, new_n14844);
nand_5 g12496(new_n14811, new_n14808, new_n14845);
and_5  g12497(new_n14812, n14692, new_n14846);
nor_5  g12498(new_n14826_1, new_n14813, new_n14847);
or_5   g12499(new_n14847, new_n14846, new_n14848);
xor_4  g12500(new_n14848, new_n14845, new_n14849_1);
xnor_4 g12501(new_n14849_1, new_n10815, new_n14850);
xnor_4 g12502(new_n14850, new_n14844, new_n14851);
nor_5  g12503(new_n14851, new_n9372_1, new_n14852);
xnor_4 g12504(new_n14851, new_n9372_1, new_n14853);
xor_4  g12505(new_n14842, new_n14829, new_n14854);
and_5  g12506(new_n14854, new_n9376, new_n14855);
xnor_4 g12507(new_n14854, new_n9376, new_n14856);
xor_4  g12508(new_n14840, new_n14832, new_n14857);
and_5  g12509(new_n14857, new_n9379, new_n14858);
xnor_4 g12510(new_n14857, new_n9379, new_n14859);
xor_4  g12511(new_n14838, new_n14835, new_n14860);
and_5  g12512(new_n14860, new_n9384, new_n14861);
xnor_4 g12513(new_n14860, new_n9385, new_n14862);
nor_5  g12514(new_n14244, new_n9389, new_n14863);
nor_5  g12515(new_n14273, new_n14245, new_n14864);
nor_5  g12516(new_n14864, new_n14863, new_n14865);
and_5  g12517(new_n14865, new_n14862, new_n14866);
nor_5  g12518(new_n14866, new_n14861, new_n14867);
nor_5  g12519(new_n14867, new_n14859, new_n14868);
nor_5  g12520(new_n14868, new_n14858, new_n14869);
nor_5  g12521(new_n14869, new_n14856, new_n14870);
nor_5  g12522(new_n14870, new_n14855, new_n14871);
nor_5  g12523(new_n14871, new_n14853, new_n14872);
nor_5  g12524(new_n14872, new_n14852, new_n14873);
and_5  g12525(new_n14849_1, new_n10819, new_n14874);
nor_5  g12526(new_n14848, new_n14845, new_n14875);
nor_5  g12527(new_n14849_1, new_n10819, new_n14876);
nor_5  g12528(new_n14876, new_n14844, new_n14877);
or_5   g12529(new_n14877, new_n14875, new_n14878);
or_5   g12530(new_n14878, new_n14874, new_n14879);
xnor_4 g12531(new_n14879, new_n14873, n3760);
xnor_4 g12532(new_n3691, new_n3668, n3781);
xnor_4 g12533(new_n12223_1, new_n12199, n3794);
nor_5  g12534(new_n9815, new_n4626, new_n14883);
nor_5  g12535(new_n14883, new_n4630, new_n14884);
and_5  g12536(new_n14883, new_n4624_1, new_n14885);
or_5   g12537(new_n14885, new_n14884, new_n14886);
and_5  g12538(new_n9814, new_n5465, new_n14887);
nor_5  g12539(new_n5466, new_n5413, new_n14888);
nor_5  g12540(new_n5470, new_n5465, new_n14889);
nor_5  g12541(new_n14889, new_n14888, new_n14890);
xnor_4 g12542(new_n14890, new_n11796, new_n14891_1);
xor_4  g12543(new_n14891_1, new_n14887, new_n14892);
xor_4  g12544(new_n14892, new_n14886, n3842);
xnor_4 g12545(new_n11060, new_n8085, n3850);
xnor_4 g12546(new_n13341, new_n3992, n3869);
xnor_4 g12547(n21749, n919, new_n14896);
nor_5  g12548(n25316, n7769, new_n14897);
and_5  g12549(n21138, n20385, new_n14898);
xnor_4 g12550(n25316, n7769, new_n14899_1);
nor_5  g12551(new_n14899_1, new_n14898, new_n14900);
nor_5  g12552(new_n14900, new_n14897, new_n14901);
xor_4  g12553(new_n14901, new_n14896, new_n14902);
xor_4  g12554(new_n14902, n19584, new_n14903);
xnor_4 g12555(n21138, n20385, new_n14904);
and_5  g12556(new_n14904, n15332, new_n14905);
nor_5  g12557(new_n14905, n5060, new_n14906);
xor_4  g12558(new_n14899_1, new_n14898, new_n14907);
xnor_4 g12559(new_n14905, n5060, new_n14908);
nor_5  g12560(new_n14908, new_n14907, new_n14909);
nor_5  g12561(new_n14909, new_n14906, new_n14910);
xor_4  g12562(new_n14910, new_n14903, new_n14911);
xor_4  g12563(new_n14911, new_n14125, new_n14912);
xor_4  g12564(new_n14908, new_n14907, new_n14913);
nor_5  g12565(new_n14913, new_n14128, new_n14914);
xnor_4 g12566(new_n14904, n15332, new_n14915);
nand_5 g12567(new_n14915, new_n14131, new_n14916);
xnor_4 g12568(new_n14913, new_n14127, new_n14917);
and_5  g12569(new_n14917, new_n14916, new_n14918);
nor_5  g12570(new_n14918, new_n14914, new_n14919);
xnor_4 g12571(new_n14919, new_n14912, n3871);
xor_4  g12572(new_n14719, new_n14712, n3891);
not_10 g12573(new_n5782_1, new_n14922);
xor_4  g12574(n10250, n2570, new_n14923);
not_10 g12575(n7674, new_n14924);
nor_5  g12576(n19033, new_n14924, new_n14925);
xor_4  g12577(n19033, n7674, new_n14926);
not_10 g12578(n6397, new_n14927);
nor_5  g12579(new_n14927, n655, new_n14928);
xor_4  g12580(n6397, n655, new_n14929);
not_10 g12581(n19196, new_n14930);
nor_5  g12582(new_n14930, n18145, new_n14931_1);
xor_4  g12583(n19196, n18145, new_n14932);
not_10 g12584(n23586, new_n14933);
nor_5  g12585(new_n14933, n10712, new_n14934);
xor_4  g12586(n23586, n10712, new_n14935);
not_10 g12587(n21226, new_n14936);
nor_5  g12588(n25126, new_n14936, new_n14937);
xor_4  g12589(n25126, n21226, new_n14938);
not_10 g12590(n4426, new_n14939);
nor_5  g12591(n19608, new_n14939, new_n14940);
and_5  g12592(new_n7878, n1689, new_n14941);
nor_5  g12593(new_n3857, new_n3850_1, new_n14942);
or_5   g12594(new_n14942, new_n14941, new_n14943);
xor_4  g12595(n19608, n4426, new_n14944_1);
nor_5  g12596(new_n14944_1, new_n14943, new_n14945);
nor_5  g12597(new_n14945, new_n14940, new_n14946);
nor_5  g12598(new_n14946, new_n14938, new_n14947);
nor_5  g12599(new_n14947, new_n14937, new_n14948);
nor_5  g12600(new_n14948, new_n14935, new_n14949);
nor_5  g12601(new_n14949, new_n14934, new_n14950);
nor_5  g12602(new_n14950, new_n14932, new_n14951);
nor_5  g12603(new_n14951, new_n14931_1, new_n14952);
nor_5  g12604(new_n14952, new_n14929, new_n14953);
nor_5  g12605(new_n14953, new_n14928, new_n14954_1);
nor_5  g12606(new_n14954_1, new_n14926, new_n14955);
nor_5  g12607(new_n14955, new_n14925, new_n14956);
xor_4  g12608(new_n14956, new_n14923, new_n14957);
xnor_4 g12609(new_n14957, new_n10773, new_n14958);
xor_4  g12610(new_n14954_1, new_n14926, new_n14959);
nor_5  g12611(new_n14959, new_n6222, new_n14960);
xnor_4 g12612(new_n14959, new_n6222, new_n14961);
xor_4  g12613(new_n14952, new_n14929, new_n14962);
nor_5  g12614(new_n14962, new_n6224, new_n14963);
xnor_4 g12615(new_n14962, new_n6224, new_n14964);
xor_4  g12616(new_n14950, new_n14932, new_n14965);
nor_5  g12617(new_n14965, new_n6227, new_n14966);
xnor_4 g12618(new_n14965, new_n6227, new_n14967);
xor_4  g12619(new_n14948, new_n14935, new_n14968);
nor_5  g12620(new_n14968, new_n6230, new_n14969);
xnor_4 g12621(new_n14968, new_n6230, new_n14970);
xor_4  g12622(new_n14946, new_n14938, new_n14971);
nor_5  g12623(new_n14971, new_n6233_1, new_n14972);
xnor_4 g12624(new_n14971, new_n6233_1, new_n14973);
xor_4  g12625(new_n14944_1, new_n14943, new_n14974);
nor_5  g12626(new_n14974, new_n6237, new_n14975);
xnor_4 g12627(new_n14974, new_n6237, new_n14976);
and_5  g12628(new_n3858, new_n3848, new_n14977_1);
and_5  g12629(new_n3870, new_n3859, new_n14978);
nor_5  g12630(new_n14978, new_n14977_1, new_n14979);
nor_5  g12631(new_n14979, new_n14976, new_n14980);
nor_5  g12632(new_n14980, new_n14975, new_n14981);
nor_5  g12633(new_n14981, new_n14973, new_n14982);
nor_5  g12634(new_n14982, new_n14972, new_n14983);
nor_5  g12635(new_n14983, new_n14970, new_n14984);
nor_5  g12636(new_n14984, new_n14969, new_n14985);
nor_5  g12637(new_n14985, new_n14967, new_n14986);
nor_5  g12638(new_n14986, new_n14966, new_n14987);
nor_5  g12639(new_n14987, new_n14964, new_n14988);
nor_5  g12640(new_n14988, new_n14963, new_n14989_1);
nor_5  g12641(new_n14989_1, new_n14961, new_n14990);
nor_5  g12642(new_n14990, new_n14960, new_n14991);
xor_4  g12643(new_n14991, new_n14958, new_n14992);
xnor_4 g12644(new_n14992, new_n14922, new_n14993);
not_10 g12645(new_n5787, new_n14994);
xor_4  g12646(new_n14989_1, new_n14961, new_n14995);
and_5  g12647(new_n14995, new_n14994, new_n14996);
xnor_4 g12648(new_n14995, new_n14994, new_n14997);
not_10 g12649(new_n5791, new_n14998);
xor_4  g12650(new_n14987, new_n14964, new_n14999);
and_5  g12651(new_n14999, new_n14998, new_n15000);
xnor_4 g12652(new_n14999, new_n14998, new_n15001);
not_10 g12653(new_n5794, new_n15002_1);
xor_4  g12654(new_n14985, new_n14967, new_n15003);
and_5  g12655(new_n15003, new_n15002_1, new_n15004_1);
xnor_4 g12656(new_n15003, new_n15002_1, new_n15005);
not_10 g12657(new_n5799, new_n15006);
xor_4  g12658(new_n14983, new_n14970, new_n15007);
and_5  g12659(new_n15007, new_n15006, new_n15008);
xnor_4 g12660(new_n15007, new_n15006, new_n15009);
not_10 g12661(new_n5803, new_n15010);
xor_4  g12662(new_n14981, new_n14973, new_n15011_1);
and_5  g12663(new_n15011_1, new_n15010, new_n15012);
xnor_4 g12664(new_n15011_1, new_n15010, new_n15013);
xor_4  g12665(new_n14979, new_n14976, new_n15014);
and_5  g12666(new_n15014, new_n5808, new_n15015);
xnor_4 g12667(new_n15014, new_n5808, new_n15016);
nor_5  g12668(new_n3878, new_n3871_1, new_n15017);
nor_5  g12669(new_n3888, new_n3879, new_n15018);
nor_5  g12670(new_n15018, new_n15017, new_n15019_1);
nor_5  g12671(new_n15019_1, new_n15016, new_n15020);
nor_5  g12672(new_n15020, new_n15015, new_n15021);
nor_5  g12673(new_n15021, new_n15013, new_n15022);
nor_5  g12674(new_n15022, new_n15012, new_n15023);
nor_5  g12675(new_n15023, new_n15009, new_n15024);
nor_5  g12676(new_n15024, new_n15008, new_n15025);
nor_5  g12677(new_n15025, new_n15005, new_n15026);
nor_5  g12678(new_n15026, new_n15004_1, new_n15027);
nor_5  g12679(new_n15027, new_n15001, new_n15028);
nor_5  g12680(new_n15028, new_n15000, new_n15029);
nor_5  g12681(new_n15029, new_n14997, new_n15030);
nor_5  g12682(new_n15030, new_n14996, new_n15031_1);
xnor_4 g12683(new_n15031_1, new_n14993, n3932);
xnor_4 g12684(new_n3685, new_n3684, n3934);
xnor_4 g12685(new_n3832, new_n3831, n3971);
or_5   g12686(n8581, n5026, new_n15035);
or_5   g12687(new_n15035, n12161, new_n15036);
or_5   g12688(new_n15036, n18157, new_n15037);
or_5   g12689(new_n15037, n20923, new_n15038);
or_5   g12690(new_n15038, n8067, new_n15039);
or_5   g12691(new_n15039, n10125, new_n15040);
or_5   g12692(new_n15040, n25240, new_n15041);
xor_4  g12693(new_n15041, n1222, new_n15042);
xnor_4 g12694(new_n15042, n15077, new_n15043);
xor_4  g12695(new_n15040, n25240, new_n15044);
or_5   g12696(new_n15044, n3710, new_n15045);
xnor_4 g12697(new_n15044, n3710, new_n15046);
xor_4  g12698(new_n15039, n10125, new_n15047);
and_5  g12699(new_n15047, n26318, new_n15048);
or_5   g12700(new_n15047, n26318, new_n15049);
xor_4  g12701(new_n15038, n8067, new_n15050);
nor_5  g12702(new_n15050, n26054, new_n15051);
xnor_4 g12703(new_n15050, n26054, new_n15052_1);
xor_4  g12704(new_n15037, n20923, new_n15053_1);
nor_5  g12705(new_n15053_1, n19081, new_n15054);
xnor_4 g12706(new_n15053_1, n19081, new_n15055);
xor_4  g12707(new_n15036, n18157, new_n15056);
nor_5  g12708(new_n15056, n8309, new_n15057);
xor_4  g12709(new_n15035, n12161, new_n15058);
nor_5  g12710(new_n15058, n19144, new_n15059);
xnor_4 g12711(new_n15058, n19144, new_n15060);
xnor_4 g12712(n8581, n5026, new_n15061);
and_5  g12713(new_n15061, new_n7968_1, new_n15062);
nand_5 g12714(n13714, n8581, new_n15063);
xnor_4 g12715(new_n15061, n12593, new_n15064);
and_5  g12716(new_n15064, new_n15063, new_n15065);
nor_5  g12717(new_n15065, new_n15062, new_n15066);
nor_5  g12718(new_n15066, new_n15060, new_n15067);
nor_5  g12719(new_n15067, new_n15059, new_n15068);
xnor_4 g12720(new_n15056, n8309, new_n15069);
nor_5  g12721(new_n15069, new_n15068, new_n15070);
nor_5  g12722(new_n15070, new_n15057, new_n15071);
nor_5  g12723(new_n15071, new_n15055, new_n15072);
nor_5  g12724(new_n15072, new_n15054, new_n15073);
nor_5  g12725(new_n15073, new_n15052_1, new_n15074);
nor_5  g12726(new_n15074, new_n15051, new_n15075);
and_5  g12727(new_n15075, new_n15049, new_n15076);
nor_5  g12728(new_n15076, new_n15048, new_n15077_1);
not_10 g12729(new_n15077_1, new_n15078);
or_5   g12730(new_n15078, new_n15046, new_n15079);
and_5  g12731(new_n15079, new_n15045, new_n15080);
xor_4  g12732(new_n15080, new_n15043, new_n15081);
xnor_4 g12733(new_n15081, new_n7302, new_n15082_1);
xnor_4 g12734(new_n15077_1, new_n15046, new_n15083);
nor_5  g12735(new_n15083, new_n7305_1, new_n15084);
xnor_4 g12736(new_n15083, new_n7305_1, new_n15085);
xnor_4 g12737(new_n15047, n26318, new_n15086);
xnor_4 g12738(new_n15086, new_n15075, new_n15087);
and_5  g12739(new_n15087, n22554, new_n15088);
xnor_4 g12740(new_n15087, n22554, new_n15089);
xor_4  g12741(new_n15073, new_n15052_1, new_n15090);
nor_5  g12742(new_n15090, new_n7311, new_n15091);
xnor_4 g12743(new_n15090, new_n7311, new_n15092);
xor_4  g12744(new_n15071, new_n15055, new_n15093);
nor_5  g12745(new_n15093, new_n7314, new_n15094_1);
xnor_4 g12746(new_n15093, new_n7314, new_n15095);
xor_4  g12747(new_n15069, new_n15068, new_n15096);
nor_5  g12748(new_n15096, new_n7317, new_n15097);
xnor_4 g12749(new_n15096, new_n7317, new_n15098);
xor_4  g12750(new_n15066, new_n15060, new_n15099);
not_10 g12751(new_n15099, new_n15100);
and_5  g12752(new_n15100, n2146, new_n15101);
xor_4  g12753(new_n15099, n2146, new_n15102);
not_10 g12754(n22173, new_n15103);
and_5  g12755(n13714, n8581, new_n15104);
xnor_4 g12756(new_n15064, new_n15104, new_n15105);
nor_5  g12757(new_n15105, new_n15103, new_n15106);
xor_4  g12758(n13714, n8581, new_n15107);
nand_5 g12759(new_n15107, n583, new_n15108);
xor_4  g12760(new_n15105, n22173, new_n15109);
nor_5  g12761(new_n15109, new_n15108, new_n15110);
nor_5  g12762(new_n15110, new_n15106, new_n15111);
nor_5  g12763(new_n15111, new_n15102, new_n15112);
nor_5  g12764(new_n15112, new_n15101, new_n15113);
nor_5  g12765(new_n15113, new_n15098, new_n15114);
nor_5  g12766(new_n15114, new_n15097, new_n15115);
nor_5  g12767(new_n15115, new_n15095, new_n15116);
nor_5  g12768(new_n15116, new_n15094_1, new_n15117);
nor_5  g12769(new_n15117, new_n15092, new_n15118_1);
nor_5  g12770(new_n15118_1, new_n15091, new_n15119);
nor_5  g12771(new_n15119, new_n15089, new_n15120);
nor_5  g12772(new_n15120, new_n15088, new_n15121);
nor_5  g12773(new_n15121, new_n15085, new_n15122);
or_5   g12774(new_n15122, new_n15084, new_n15123);
xor_4  g12775(new_n15123, new_n15082_1, new_n15124);
xnor_4 g12776(new_n15124, new_n7405, new_n15125);
xnor_4 g12777(new_n7288, new_n7249, new_n15126);
xor_4  g12778(new_n15121, new_n15085, new_n15127);
nor_5  g12779(new_n15127, new_n15126, new_n15128_1);
xnor_4 g12780(new_n15127, new_n15126, new_n15129);
xnor_4 g12781(new_n7286, new_n7253_1, new_n15130);
xor_4  g12782(new_n15119, new_n15089, new_n15131);
nor_5  g12783(new_n15131, new_n15130, new_n15132);
xnor_4 g12784(new_n15131, new_n15130, new_n15133);
xnor_4 g12785(new_n7284, new_n7257, new_n15134);
xor_4  g12786(new_n15117, new_n15092, new_n15135);
nor_5  g12787(new_n15135, new_n15134, new_n15136);
xnor_4 g12788(new_n15135, new_n15134, new_n15137);
xnor_4 g12789(new_n7282, new_n7261, new_n15138);
xor_4  g12790(new_n15115, new_n15095, new_n15139_1);
nor_5  g12791(new_n15139_1, new_n15138, new_n15140);
xnor_4 g12792(new_n15139_1, new_n15138, new_n15141);
not_10 g12793(new_n7425, new_n15142);
xor_4  g12794(new_n15113, new_n15098, new_n15143);
nor_5  g12795(new_n15143, new_n15142, new_n15144);
xor_4  g12796(new_n15143, new_n7425, new_n15145_1);
xor_4  g12797(new_n15111, new_n15102, new_n15146_1);
nor_5  g12798(new_n15146_1, new_n7429, new_n15147);
xnor_4 g12799(new_n15109, new_n15108, new_n15148);
and_5  g12800(new_n15148, new_n7435, new_n15149);
xnor_4 g12801(new_n15107, n583, new_n15150);
or_5   g12802(new_n15150, new_n2524, new_n15151);
xor_4  g12803(new_n15148, new_n7435, new_n15152);
and_5  g12804(new_n15152, new_n15151, new_n15153);
nor_5  g12805(new_n15153, new_n15149, new_n15154);
xnor_4 g12806(new_n15146_1, new_n7429, new_n15155);
nor_5  g12807(new_n15155, new_n15154, new_n15156);
nor_5  g12808(new_n15156, new_n15147, new_n15157);
nor_5  g12809(new_n15157, new_n15145_1, new_n15158);
nor_5  g12810(new_n15158, new_n15144, new_n15159);
nor_5  g12811(new_n15159, new_n15141, new_n15160);
nor_5  g12812(new_n15160, new_n15140, new_n15161);
nor_5  g12813(new_n15161, new_n15137, new_n15162);
nor_5  g12814(new_n15162, new_n15136, new_n15163);
nor_5  g12815(new_n15163, new_n15133, new_n15164);
nor_5  g12816(new_n15164, new_n15132, new_n15165_1);
nor_5  g12817(new_n15165_1, new_n15129, new_n15166);
nor_5  g12818(new_n15166, new_n15128_1, new_n15167_1);
xnor_4 g12819(new_n15167_1, new_n15125, n3983);
xnor_4 g12820(n13714, n583, new_n15169);
xor_4  g12821(new_n15169, n6611, new_n15170);
and_5  g12822(new_n15170, new_n6047, new_n15171);
nor_5  g12823(new_n15169, new_n8174, new_n15172);
and_5  g12824(n13714, n583, new_n15173);
xnor_4 g12825(n22173, n12593, new_n15174);
xnor_4 g12826(new_n15174, new_n15173, new_n15175);
xnor_4 g12827(new_n15175, n27188, new_n15176_1);
xor_4  g12828(new_n15176_1, new_n15172, new_n15177);
xnor_4 g12829(new_n15177, new_n15171, new_n15178);
xor_4  g12830(new_n15178, new_n6043, n4000);
xnor_4 g12831(new_n6632, new_n6607, new_n15180_1);
xor_4  g12832(n26823, n20179, new_n15181);
nor_5  g12833(n19228, new_n3058, new_n15182_1);
xor_4  g12834(n19228, n4812, new_n15183);
nor_5  g12835(new_n3059, n15539, new_n15184);
xor_4  g12836(n24278, n15539, new_n15185);
nor_5  g12837(new_n7641, n8052, new_n15186);
or_5   g12838(n24618, new_n6766, new_n15187);
nor_5  g12839(new_n6769, n3952, new_n15188);
nor_5  g12840(new_n10154, new_n10153, new_n15189);
nor_5  g12841(new_n15189, new_n15188, new_n15190);
and_5  g12842(new_n15190, new_n15187, new_n15191);
nor_5  g12843(new_n15191, new_n15186, new_n15192);
nor_5  g12844(new_n15192, new_n15185, new_n15193);
nor_5  g12845(new_n15193, new_n15184, new_n15194);
nor_5  g12846(new_n15194, new_n15183, new_n15195);
nor_5  g12847(new_n15195, new_n15182_1, new_n15196);
xor_4  g12848(new_n15196, new_n15181, new_n15197);
xnor_4 g12849(new_n15197, new_n15180_1, new_n15198);
xnor_4 g12850(new_n6630_1, new_n6610, new_n15199);
xor_4  g12851(new_n15194, new_n15183, new_n15200);
nor_5  g12852(new_n15200, new_n15199, new_n15201);
xnor_4 g12853(new_n15200, new_n15199, new_n15202);
xor_4  g12854(new_n15192, new_n15185, new_n15203);
nor_5  g12855(new_n15203, new_n6708, new_n15204);
xor_4  g12856(n24618, n8052, new_n15205_1);
xor_4  g12857(new_n15205_1, new_n15190, new_n15206);
and_5  g12858(new_n15206, new_n6711, new_n15207);
xor_4  g12859(new_n15206, new_n6711, new_n15208);
nor_5  g12860(new_n10155, new_n10152, new_n15209);
nor_5  g12861(new_n10156, new_n6722, new_n15210);
nor_5  g12862(new_n15210, new_n15209, new_n15211);
and_5  g12863(new_n15211, new_n15208, new_n15212);
nor_5  g12864(new_n15212, new_n15207, new_n15213);
xnor_4 g12865(new_n15203, new_n6708, new_n15214);
nor_5  g12866(new_n15214, new_n15213, new_n15215);
nor_5  g12867(new_n15215, new_n15204, new_n15216);
nor_5  g12868(new_n15216, new_n15202, new_n15217);
nor_5  g12869(new_n15217, new_n15201, new_n15218);
xnor_4 g12870(new_n15218, new_n15198, n4010);
xor_4  g12871(n11220, n2160, new_n15220);
not_10 g12872(n10763, new_n15221);
nor_5  g12873(n22379, new_n15221, new_n15222);
xor_4  g12874(n22379, n10763, new_n15223);
not_10 g12875(n7437, new_n15224);
nor_5  g12876(new_n15224, n1662, new_n15225);
xor_4  g12877(n7437, n1662, new_n15226);
not_10 g12878(n20700, new_n15227);
nor_5  g12879(new_n15227, n12875, new_n15228);
not_10 g12880(n7099, new_n15229);
nor_5  g12881(new_n15229, n2035, new_n15230_1);
nor_5  g12882(new_n13312, new_n13291, new_n15231);
nor_5  g12883(new_n15231, new_n15230_1, new_n15232);
xor_4  g12884(n20700, n12875, new_n15233);
nor_5  g12885(new_n15233, new_n15232, new_n15234);
nor_5  g12886(new_n15234, new_n15228, new_n15235);
nor_5  g12887(new_n15235, new_n15226, new_n15236);
nor_5  g12888(new_n15236, new_n15225, new_n15237);
nor_5  g12889(new_n15237, new_n15223, new_n15238);
nor_5  g12890(new_n15238, new_n15222, new_n15239);
xor_4  g12891(new_n15239, new_n15220, new_n15240);
xnor_4 g12892(new_n15240, new_n13450, new_n15241_1);
xor_4  g12893(new_n15237, new_n15223, new_n15242);
nor_5  g12894(new_n15242, new_n13457_1, new_n15243);
xnor_4 g12895(new_n15242, new_n13457_1, new_n15244);
xor_4  g12896(new_n15235, new_n15226, new_n15245);
nor_5  g12897(new_n15245, new_n13462, new_n15246);
xnor_4 g12898(new_n15233, new_n15232, new_n15247);
nor_5  g12899(new_n15247, new_n13465, new_n15248);
xnor_4 g12900(new_n15247, new_n13465, new_n15249);
and_5  g12901(new_n13325, new_n13313, new_n15250);
nor_5  g12902(new_n13350, new_n13326, new_n15251);
nor_5  g12903(new_n15251, new_n15250, new_n15252);
nor_5  g12904(new_n15252, new_n15249, new_n15253);
nor_5  g12905(new_n15253, new_n15248, new_n15254);
xor_4  g12906(new_n15245, new_n13462, new_n15255_1);
and_5  g12907(new_n15255_1, new_n15254, new_n15256);
nor_5  g12908(new_n15256, new_n15246, new_n15257);
nor_5  g12909(new_n15257, new_n15244, new_n15258_1);
or_5   g12910(new_n15258_1, new_n15243, new_n15259);
xor_4  g12911(new_n15259, new_n15241_1, n4014);
xnor_4 g12912(new_n12782, n18496, new_n15261);
nor_5  g12913(new_n12785, n26224, new_n15262);
xnor_4 g12914(new_n12785, n26224, new_n15263);
nor_5  g12915(new_n3523, n19327, new_n15264);
nor_5  g12916(new_n3550, new_n3524, new_n15265);
nor_5  g12917(new_n15265, new_n15264, new_n15266);
nor_5  g12918(new_n15266, new_n15263, new_n15267);
nor_5  g12919(new_n15267, new_n15262, new_n15268);
xor_4  g12920(new_n15268, new_n15261, new_n15269);
xor_4  g12921(new_n15269, n647, new_n15270);
xor_4  g12922(new_n15266, new_n15263, new_n15271_1);
nor_5  g12923(new_n15271_1, new_n5437, new_n15272);
xor_4  g12924(new_n15271_1, n20409, new_n15273);
and_5  g12925(new_n3551, n25749, new_n15274);
nor_5  g12926(new_n3582_1, new_n3552, new_n15275_1);
nor_5  g12927(new_n15275_1, new_n15274, new_n15276);
nor_5  g12928(new_n15276, new_n15273, new_n15277);
nor_5  g12929(new_n15277, new_n15272, new_n15278);
xor_4  g12930(new_n15278, new_n15270, new_n15279);
xor_4  g12931(new_n15279, new_n10723, new_n15280);
not_10 g12932(new_n10727, new_n15281);
xor_4  g12933(new_n15276, new_n15273, new_n15282);
nor_5  g12934(new_n15282, new_n15281, new_n15283);
xor_4  g12935(new_n15282, new_n10727, new_n15284);
and_5  g12936(new_n3657, new_n3583, new_n15285);
nor_5  g12937(new_n3695, new_n3658, new_n15286);
nor_5  g12938(new_n15286, new_n15285, new_n15287);
nor_5  g12939(new_n15287, new_n15284, new_n15288);
nor_5  g12940(new_n15288, new_n15283, new_n15289_1);
xnor_4 g12941(new_n15289_1, new_n15280, n4071);
xnor_4 g12942(new_n11660, new_n11654, n4088);
nor_5  g12943(new_n11765, n7593, new_n15292);
nor_5  g12944(new_n11766, n5025, new_n15293);
and_5  g12945(new_n11766, n5025, new_n15294);
nor_5  g12946(new_n11770_1, new_n15294, new_n15295);
nor_5  g12947(new_n15295, new_n15293, new_n15296);
nor_5  g12948(new_n15296, new_n15292, new_n15297);
not_10 g12949(new_n14736, new_n15298);
nor_5  g12950(new_n14739, new_n15298, new_n15299);
nand_5 g12951(new_n14739, new_n15298, new_n15300_1);
and_5  g12952(new_n14743, new_n15300_1, new_n15301);
nor_5  g12953(new_n15301, new_n15299, new_n15302);
and_5  g12954(new_n15302, new_n15297, new_n15303);
not_10 g12955(new_n15297, new_n15304);
and_5  g12956(new_n15304, new_n14744, new_n15305);
or_5   g12957(new_n15304, new_n14744, new_n15306);
nor_5  g12958(new_n11771_1, new_n11764, new_n15307_1);
nor_5  g12959(new_n11775_1, new_n11772, new_n15308);
nor_5  g12960(new_n15308, new_n15307_1, new_n15309);
and_5  g12961(new_n15309, new_n15306, new_n15310);
nor_5  g12962(new_n15310, new_n15305, new_n15311);
nor_5  g12963(new_n15311, new_n15303, new_n15312);
nor_5  g12964(new_n15302, new_n15297, new_n15313);
nor_5  g12965(new_n15313, new_n15310, new_n15314);
nor_5  g12966(new_n15314, new_n15312, n4089);
or_5   g12967(new_n10919, n1112, new_n15316);
xnor_4 g12968(new_n15316, new_n6750, new_n15317);
xnor_4 g12969(new_n15317, n3228, new_n15318);
nor_5  g12970(new_n10920, n5302, new_n15319);
xnor_4 g12971(new_n10920, n5302, new_n15320);
and_5  g12972(new_n10922, n25738, new_n15321);
or_5   g12973(new_n10922, n25738, new_n15322);
nor_5  g12974(new_n7800, n21471, new_n15323);
and_5  g12975(new_n7817, new_n7801, new_n15324);
nor_5  g12976(new_n15324, new_n15323, new_n15325);
and_5  g12977(new_n15325, new_n15322, new_n15326);
or_5   g12978(new_n15326, new_n15321, new_n15327_1);
nor_5  g12979(new_n15327_1, new_n15320, new_n15328);
nor_5  g12980(new_n15328, new_n15319, new_n15329);
xnor_4 g12981(new_n15329, new_n15318, new_n15330);
xnor_4 g12982(new_n15330, n13775, new_n15331);
xnor_4 g12983(new_n15327_1, new_n15320, new_n15332_1);
nor_5  g12984(new_n15332_1, n1293, new_n15333);
xnor_4 g12985(new_n15332_1, new_n7866, new_n15334);
xnor_4 g12986(new_n10922, n25738, new_n15335);
xnor_4 g12987(new_n15335, new_n15325, new_n15336);
and_5  g12988(new_n15336, n19042, new_n15337);
and_5  g12989(new_n7818, n19472, new_n15338);
nor_5  g12990(new_n7838, new_n7819, new_n15339);
nor_5  g12991(new_n15339, new_n15338, new_n15340);
xnor_4 g12992(new_n15336, n19042, new_n15341);
nor_5  g12993(new_n15341, new_n15340, new_n15342);
nor_5  g12994(new_n15342, new_n15337, new_n15343);
and_5  g12995(new_n15343, new_n15334, new_n15344);
nor_5  g12996(new_n15344, new_n15333, new_n15345_1);
xnor_4 g12997(new_n15345_1, new_n15331, new_n15346);
xor_4  g12998(new_n6845, n11736, new_n15347);
and_5  g12999(new_n2439, n23200, new_n15348);
xnor_4 g13000(new_n2439, n23200, new_n15349);
and_5  g13001(new_n2443, n17959, new_n15350);
xnor_4 g13002(new_n2443, n17959, new_n15351);
and_5  g13003(new_n2447, n7566, new_n15352);
nor_5  g13004(new_n6074, new_n6061, new_n15353_1);
nor_5  g13005(new_n15353_1, new_n15352, new_n15354);
nor_5  g13006(new_n15354, new_n15351, new_n15355);
nor_5  g13007(new_n15355, new_n15350, new_n15356);
nor_5  g13008(new_n15356, new_n15349, new_n15357);
nor_5  g13009(new_n15357, new_n15348, new_n15358);
xor_4  g13010(new_n15358, new_n15347, new_n15359);
xnor_4 g13011(new_n15359, new_n15346, new_n15360);
xnor_4 g13012(new_n15343, new_n15334, new_n15361);
xor_4  g13013(new_n15356, new_n15349, new_n15362);
nor_5  g13014(new_n15362, new_n15361, new_n15363);
xnor_4 g13015(new_n15362, new_n15361, new_n15364);
xor_4  g13016(new_n15354, new_n15351, new_n15365);
xor_4  g13017(new_n15341, new_n15340, new_n15366_1);
nor_5  g13018(new_n15366_1, new_n15365, new_n15367);
nor_5  g13019(new_n7839, new_n6075, new_n15368);
nor_5  g13020(new_n7857, new_n7840, new_n15369);
nor_5  g13021(new_n15369, new_n15368, new_n15370);
xnor_4 g13022(new_n15366_1, new_n15365, new_n15371);
nor_5  g13023(new_n15371, new_n15370, new_n15372);
nor_5  g13024(new_n15372, new_n15367, new_n15373);
nor_5  g13025(new_n15373, new_n15364, new_n15374);
nor_5  g13026(new_n15374, new_n15363, new_n15375);
xnor_4 g13027(new_n15375, new_n15360, n4103);
nor_5  g13028(new_n13382, new_n11548_1, new_n15377);
xnor_4 g13029(new_n13382, new_n11548_1, new_n15378_1);
not_10 g13030(new_n11486_1, new_n15379);
nor_5  g13031(new_n13385, new_n15379, new_n15380);
not_10 g13032(new_n11490, new_n15381);
nor_5  g13033(new_n13389, new_n15381, new_n15382_1);
xor_4  g13034(new_n13389, new_n11490, new_n15383);
and_5  g13035(new_n13392, new_n11494, new_n15384);
xnor_4 g13036(new_n13392, new_n11494, new_n15385);
not_10 g13037(new_n11498, new_n15386);
nor_5  g13038(new_n13396, new_n15386, new_n15387);
xor_4  g13039(new_n13396, new_n11498, new_n15388);
and_5  g13040(new_n13320, new_n11502, new_n15389);
and_5  g13041(new_n11506_1, new_n14771, new_n15390);
xnor_4 g13042(new_n11506_1, new_n3956, new_n15391);
nor_5  g13043(new_n11510, new_n3960, new_n15392);
xnor_4 g13044(new_n11510, new_n3960, new_n15393);
and_5  g13045(new_n11513, new_n3963, new_n15394);
xnor_4 g13046(new_n11513, new_n3963, new_n15395);
and_5  g13047(new_n11518, new_n3965, new_n15396);
nor_5  g13048(new_n11591_1, new_n3967, new_n15397);
xnor_4 g13049(new_n11518, new_n3965, new_n15398);
nor_5  g13050(new_n15398, new_n15397, new_n15399);
nor_5  g13051(new_n15399, new_n15396, new_n15400);
nor_5  g13052(new_n15400, new_n15395, new_n15401);
or_5   g13053(new_n15401, new_n15394, new_n15402);
nor_5  g13054(new_n15402, new_n15393, new_n15403);
nor_5  g13055(new_n15403, new_n15392, new_n15404);
and_5  g13056(new_n15404, new_n15391, new_n15405);
nor_5  g13057(new_n15405, new_n15390, new_n15406);
xnor_4 g13058(new_n13320, new_n11502, new_n15407_1);
nor_5  g13059(new_n15407_1, new_n15406, new_n15408);
nor_5  g13060(new_n15408, new_n15389, new_n15409);
nor_5  g13061(new_n15409, new_n15388, new_n15410);
nor_5  g13062(new_n15410, new_n15387, new_n15411);
nor_5  g13063(new_n15411, new_n15385, new_n15412);
nor_5  g13064(new_n15412, new_n15384, new_n15413);
nor_5  g13065(new_n15413, new_n15383, new_n15414);
nor_5  g13066(new_n15414, new_n15382_1, new_n15415);
xor_4  g13067(new_n13385, new_n11486_1, new_n15416);
nor_5  g13068(new_n15416, new_n15415, new_n15417);
or_5   g13069(new_n15417, new_n15380, new_n15418);
nor_5  g13070(new_n15418, new_n15378_1, new_n15419);
nor_5  g13071(new_n15419, new_n15377, new_n15420);
not_10 g13072(new_n15420, new_n15421);
and_5  g13073(new_n5395, n6456, new_n15422);
or_5   g13074(new_n5395, n6456, new_n15423);
nor_5  g13075(new_n5432, n4085, new_n15424_1);
xnor_4 g13076(new_n5432, n4085, new_n15425);
nor_5  g13077(new_n5438_1, n26725, new_n15426);
xnor_4 g13078(new_n5438_1, n26725, new_n15427);
nor_5  g13079(new_n5443_1, n11980, new_n15428_1);
xnor_4 g13080(new_n5443_1, n11980, new_n15429);
nor_5  g13081(new_n5447, n3253, new_n15430);
xnor_4 g13082(new_n5447, n3253, new_n15431);
nor_5  g13083(new_n5452, n7759, new_n15432);
xnor_4 g13084(new_n5452, n7759, new_n15433);
nor_5  g13085(new_n5456, n12562, new_n15434);
nor_5  g13086(new_n5461, n7949, new_n15435_1);
xnor_4 g13087(new_n5461, n7949, new_n15436);
nor_5  g13088(new_n5471, n24374, new_n15437);
nand_5 g13089(n20658, n14575, new_n15438_1);
xor_4  g13090(new_n5471, n24374, new_n15439);
and_5  g13091(new_n15439, new_n15438_1, new_n15440);
nor_5  g13092(new_n15440, new_n15437, new_n15441);
nor_5  g13093(new_n15441, new_n15436, new_n15442);
nor_5  g13094(new_n15442, new_n15435_1, new_n15443);
xnor_4 g13095(new_n5456, n12562, new_n15444);
nor_5  g13096(new_n15444, new_n15443, new_n15445);
nor_5  g13097(new_n15445, new_n15434, new_n15446);
nor_5  g13098(new_n15446, new_n15433, new_n15447);
nor_5  g13099(new_n15447, new_n15432, new_n15448);
nor_5  g13100(new_n15448, new_n15431, new_n15449);
nor_5  g13101(new_n15449, new_n15430, new_n15450);
nor_5  g13102(new_n15450, new_n15429, new_n15451);
nor_5  g13103(new_n15451, new_n15428_1, new_n15452);
nor_5  g13104(new_n15452, new_n15427, new_n15453);
nor_5  g13105(new_n15453, new_n15426, new_n15454);
nor_5  g13106(new_n15454, new_n15425, new_n15455);
nor_5  g13107(new_n15455, new_n15424_1, new_n15456);
and_5  g13108(new_n15456, new_n15423, new_n15457);
or_5   g13109(new_n15457, new_n12461_1, new_n15458);
nor_5  g13110(new_n15458, new_n15422, new_n15459);
and_5  g13111(new_n15459, new_n15421, new_n15460);
xor_4  g13112(new_n15418, new_n15378_1, new_n15461);
nor_5  g13113(new_n15461, new_n15459, new_n15462);
xnor_4 g13114(new_n15461, new_n15459, new_n15463);
xor_4  g13115(new_n15416, new_n15415, new_n15464);
xor_4  g13116(new_n5395, n6456, new_n15465_1);
xnor_4 g13117(new_n15465_1, new_n15456, new_n15466);
and_5  g13118(new_n15466, new_n15464, new_n15467_1);
xnor_4 g13119(new_n15466, new_n15464, new_n15468);
xor_4  g13120(new_n15454, new_n15425, new_n15469);
xor_4  g13121(new_n15413, new_n15383, new_n15470_1);
and_5  g13122(new_n15470_1, new_n15469, new_n15471);
xnor_4 g13123(new_n15470_1, new_n15469, new_n15472);
xor_4  g13124(new_n15452, new_n15427, new_n15473);
xor_4  g13125(new_n15411, new_n15385, new_n15474);
and_5  g13126(new_n15474, new_n15473, new_n15475);
xnor_4 g13127(new_n15474, new_n15473, new_n15476);
xor_4  g13128(new_n15450, new_n15429, new_n15477_1);
xor_4  g13129(new_n15409, new_n15388, new_n15478);
and_5  g13130(new_n15478, new_n15477_1, new_n15479);
xnor_4 g13131(new_n15478, new_n15477_1, new_n15480);
xor_4  g13132(new_n15448, new_n15431, new_n15481_1);
xor_4  g13133(new_n15407_1, new_n15406, new_n15482);
and_5  g13134(new_n15482, new_n15481_1, new_n15483);
xnor_4 g13135(new_n15482, new_n15481_1, new_n15484);
xor_4  g13136(new_n15446, new_n15433, new_n15485);
xor_4  g13137(new_n15404, new_n15391, new_n15486);
and_5  g13138(new_n15486, new_n15485, new_n15487);
xnor_4 g13139(new_n15486, new_n15485, new_n15488);
xor_4  g13140(new_n15402, new_n15393, new_n15489);
xnor_4 g13141(new_n15444, new_n15443, new_n15490_1);
nor_5  g13142(new_n15490_1, new_n15489, new_n15491);
xor_4  g13143(new_n15490_1, new_n15489, new_n15492);
xor_4  g13144(new_n15441, new_n15436, new_n15493);
xor_4  g13145(new_n15400, new_n15395, new_n15494);
nor_5  g13146(new_n15494, new_n15493, new_n15495);
xnor_4 g13147(new_n15494, new_n15493, new_n15496_1);
xor_4  g13148(new_n15398, new_n15397, new_n15497);
not_10 g13149(new_n15497, new_n15498);
nor_5  g13150(new_n15498, new_n15439, new_n15499);
xor_4  g13151(new_n15439, new_n15438_1, new_n15500);
or_5   g13152(new_n15500, new_n15497, new_n15501_1);
xnor_4 g13153(n20658, n14575, new_n15502);
xnor_4 g13154(new_n11591_1, new_n3967, new_n15503);
or_5   g13155(new_n15503, new_n15502, new_n15504);
and_5  g13156(new_n15504, new_n15501_1, new_n15505);
or_5   g13157(new_n15505, new_n15499, new_n15506_1);
nor_5  g13158(new_n15506_1, new_n15496_1, new_n15507);
nor_5  g13159(new_n15507, new_n15495, new_n15508_1);
and_5  g13160(new_n15508_1, new_n15492, new_n15509);
nor_5  g13161(new_n15509, new_n15491, new_n15510);
nor_5  g13162(new_n15510, new_n15488, new_n15511);
nor_5  g13163(new_n15511, new_n15487, new_n15512);
nor_5  g13164(new_n15512, new_n15484, new_n15513);
nor_5  g13165(new_n15513, new_n15483, new_n15514);
nor_5  g13166(new_n15514, new_n15480, new_n15515);
nor_5  g13167(new_n15515, new_n15479, new_n15516);
nor_5  g13168(new_n15516, new_n15476, new_n15517);
nor_5  g13169(new_n15517, new_n15475, new_n15518);
nor_5  g13170(new_n15518, new_n15472, new_n15519);
nor_5  g13171(new_n15519, new_n15471, new_n15520);
nor_5  g13172(new_n15520, new_n15468, new_n15521);
nor_5  g13173(new_n15521, new_n15467_1, new_n15522);
nor_5  g13174(new_n15522, new_n15463, new_n15523);
nor_5  g13175(new_n15523, new_n15462, new_n15524);
nor_5  g13176(new_n15524, new_n15460, new_n15525);
nor_5  g13177(new_n15459, new_n15421, new_n15526);
nor_5  g13178(new_n15526, new_n15523, new_n15527);
nor_5  g13179(new_n15527, new_n15525, n4123);
xnor_4 g13180(new_n11999, new_n7163, new_n15529);
nor_5  g13181(new_n12002, new_n7170, new_n15530);
xnor_4 g13182(new_n12002, new_n7170, new_n15531);
nor_5  g13183(new_n12006, new_n7185, new_n15532);
xor_4  g13184(new_n12006, new_n7185, new_n15533);
nor_5  g13185(new_n12016, new_n7176, new_n15534);
or_5   g13186(new_n8837, new_n7178, new_n15535);
xnor_4 g13187(new_n12016, new_n7176, new_n15536);
nor_5  g13188(new_n15536, new_n15535, new_n15537);
nor_5  g13189(new_n15537, new_n15534, new_n15538);
and_5  g13190(new_n15538, new_n15533, new_n15539_1);
nor_5  g13191(new_n15539_1, new_n15532, new_n15540);
nor_5  g13192(new_n15540, new_n15531, new_n15541);
nor_5  g13193(new_n15541, new_n15530, new_n15542);
xnor_4 g13194(new_n15542, new_n15529, n4134);
xnor_4 g13195(new_n8250, new_n8202, n4146);
xnor_4 g13196(new_n13897, new_n12860, new_n15545);
not_10 g13197(new_n12864_1, new_n15546_1);
nor_5  g13198(new_n13900, new_n15546_1, new_n15547);
xor_4  g13199(new_n13900, new_n12864_1, new_n15548);
nor_5  g13200(new_n12873_1, new_n12075, new_n15549);
nor_5  g13201(new_n12870_1, new_n12071, new_n15550);
xnor_4 g13202(new_n12867, new_n12075, new_n15551);
and_5  g13203(new_n15551, new_n15550, new_n15552);
or_5   g13204(new_n15552, new_n15549, new_n15553);
nor_5  g13205(new_n15553, new_n15548, new_n15554);
nor_5  g13206(new_n15554, new_n15547, new_n15555_1);
xnor_4 g13207(new_n15555_1, new_n15545, n4150);
xnor_4 g13208(new_n11326_1, new_n11325_1, n4151);
xnor_4 g13209(new_n11610, new_n11558, n4152);
xnor_4 g13210(new_n5616, new_n5583, n4153);
not_10 g13211(n25972, new_n15560);
nor_5  g13212(new_n15560, n10250, new_n15561);
nor_5  g13213(new_n7899, new_n7859, new_n15562);
nor_5  g13214(new_n15562, new_n15561, new_n15563);
xnor_4 g13215(new_n15563, new_n11033, new_n15564);
xor_4  g13216(new_n11035, new_n11019, new_n15565);
not_10 g13217(new_n15563, new_n15566);
nor_5  g13218(new_n15566, new_n15565, new_n15567);
nor_5  g13219(new_n15563, new_n11036, new_n15568);
and_5  g13220(new_n8048, new_n7900, new_n15569);
nor_5  g13221(new_n8102, new_n8049, new_n15570_1);
nor_5  g13222(new_n15570_1, new_n15569, new_n15571);
nor_5  g13223(new_n15571, new_n15568, new_n15572);
nor_5  g13224(new_n15572, new_n15567, new_n15573_1);
xnor_4 g13225(new_n15573_1, new_n15564, n4165);
xnor_4 g13226(new_n10404_1, new_n10376, n4172);
xnor_4 g13227(new_n10256, new_n4392, n4173);
xnor_4 g13228(new_n5977, new_n5959, n4176);
xnor_4 g13229(new_n8235, new_n8234, n4186);
xnor_4 g13230(new_n15161, new_n15137, n4204);
and_5  g13231(new_n10298, n13494, new_n15580);
xnor_4 g13232(new_n10298, n13494, new_n15581);
and_5  g13233(new_n6156, n25345, new_n15582);
nor_5  g13234(new_n6196, new_n6157, new_n15583);
nor_5  g13235(new_n15583, new_n15582, new_n15584);
nor_5  g13236(new_n15584, new_n15581, new_n15585);
nor_5  g13237(new_n15585, new_n15580, new_n15586);
nor_5  g13238(new_n15586, new_n10325, new_n15587);
or_5   g13239(new_n14539, n3366, new_n15588_1);
or_5   g13240(new_n15588_1, n19652, new_n15589);
xnor_4 g13241(new_n15589, n3984, new_n15590_1);
nor_5  g13242(new_n15590_1, n17037, new_n15591);
xnor_4 g13243(new_n15590_1, n17037, new_n15592);
xnor_4 g13244(new_n15588_1, n19652, new_n15593);
and_5  g13245(new_n15593, n5386, new_n15594);
nor_5  g13246(new_n14540, n26191, new_n15595);
nor_5  g13247(new_n14569, new_n14541_1, new_n15596);
or_5   g13248(new_n15596, new_n15595, new_n15597);
xnor_4 g13249(new_n15593, n5386, new_n15598_1);
nor_5  g13250(new_n15598_1, new_n15597, new_n15599);
or_5   g13251(new_n15599, new_n15594, new_n15600);
nor_5  g13252(new_n15600, new_n15592, new_n15601);
nor_5  g13253(new_n15601, new_n15591, new_n15602_1);
nor_5  g13254(new_n15589, n3984, new_n15603);
xor_4  g13255(new_n15603, n4514, new_n15604);
xnor_4 g13256(new_n15604, n7569, new_n15605);
xnor_4 g13257(new_n15605, new_n15602_1, new_n15606);
and_5  g13258(new_n15606, n25586, new_n15607);
xnor_4 g13259(new_n15606, n25586, new_n15608);
not_10 g13260(n25751, new_n15609);
xor_4  g13261(new_n15600, new_n15592, new_n15610);
nor_5  g13262(new_n15610, new_n15609, new_n15611);
xnor_4 g13263(new_n15610, new_n15609, new_n15612);
xor_4  g13264(new_n15598_1, new_n15597, new_n15613);
nor_5  g13265(new_n15613, n26053, new_n15614_1);
xnor_4 g13266(new_n15613, n26053, new_n15615);
and_5  g13267(new_n14570_1, new_n14532, new_n15616);
nor_5  g13268(new_n14602, new_n14571, new_n15617);
nor_5  g13269(new_n15617, new_n15616, new_n15618);
nor_5  g13270(new_n15618, new_n15615, new_n15619);
or_5   g13271(new_n15619, new_n15614_1, new_n15620);
nor_5  g13272(new_n15620, new_n15612, new_n15621);
nor_5  g13273(new_n15621, new_n15611, new_n15622);
nor_5  g13274(new_n15622, new_n15608, new_n15623);
nor_5  g13275(new_n15623, new_n15607, new_n15624);
or_5   g13276(new_n15589, n3984, new_n15625);
or_5   g13277(new_n15625, n4514, new_n15626);
and_5  g13278(new_n15604, n7569, new_n15627);
or_5   g13279(new_n15627, new_n15602_1, new_n15628);
nor_5  g13280(new_n15628, new_n15626, new_n15629);
and_5  g13281(new_n15629, new_n15624, new_n15630);
nor_5  g13282(new_n15604, n7569, new_n15631);
xor_4  g13283(new_n15628, new_n15626, new_n15632);
or_5   g13284(new_n15632, new_n15631, new_n15633);
or_5   g13285(new_n15633, new_n15624, new_n15634);
nor_5  g13286(new_n15634, new_n15629, new_n15635);
nor_5  g13287(new_n15635, new_n15630, new_n15636_1);
nor_5  g13288(new_n15636_1, new_n15587, new_n15637);
xnor_4 g13289(new_n15633, new_n15624, new_n15638);
xor_4  g13290(new_n15586, new_n10325, new_n15639);
nor_5  g13291(new_n15639, new_n15638, new_n15640);
xnor_4 g13292(new_n15639, new_n15638, new_n15641);
xnor_4 g13293(new_n15622, new_n15608, new_n15642);
xor_4  g13294(new_n15584, new_n15581, new_n15643);
nor_5  g13295(new_n15643, new_n15642, new_n15644);
xnor_4 g13296(new_n15643, new_n15642, new_n15645);
xor_4  g13297(new_n15620, new_n15612, new_n15646);
and_5  g13298(new_n15646, new_n6197, new_n15647);
xnor_4 g13299(new_n15646, new_n6197, new_n15648);
xor_4  g13300(new_n15618, new_n15615, new_n15649);
nor_5  g13301(new_n15649, new_n6262, new_n15650);
nor_5  g13302(new_n14603_1, new_n6266, new_n15651);
nor_5  g13303(new_n14633_1, new_n14604, new_n15652_1);
nor_5  g13304(new_n15652_1, new_n15651, new_n15653);
xnor_4 g13305(new_n15649, new_n6262, new_n15654);
nor_5  g13306(new_n15654, new_n15653, new_n15655);
nor_5  g13307(new_n15655, new_n15650, new_n15656);
nor_5  g13308(new_n15656, new_n15648, new_n15657);
nor_5  g13309(new_n15657, new_n15647, new_n15658);
nor_5  g13310(new_n15658, new_n15645, new_n15659);
nor_5  g13311(new_n15659, new_n15644, new_n15660);
nor_5  g13312(new_n15660, new_n15641, new_n15661);
or_5   g13313(new_n15661, new_n15640, new_n15662_1);
nor_5  g13314(new_n15662_1, new_n15637, new_n15663);
and_5  g13315(new_n15636_1, new_n15587, new_n15664);
or_5   g13316(new_n15664, new_n15630, new_n15665);
nor_5  g13317(new_n15665, new_n15663, n4205);
or_5   g13318(new_n11928, n22198, new_n15667);
or_5   g13319(new_n15667, n24327, new_n15668);
xor_4  g13320(new_n15668, n2659, new_n15669);
xnor_4 g13321(new_n15669, n18444, new_n15670);
xor_4  g13322(new_n15667, n24327, new_n15671);
nor_5  g13323(new_n15671, n24638, new_n15672);
xnor_4 g13324(new_n15671, n24638, new_n15673);
nor_5  g13325(new_n11929, n21674, new_n15674);
nor_5  g13326(new_n11951, new_n11930, new_n15675);
nor_5  g13327(new_n15675, new_n15674, new_n15676);
nor_5  g13328(new_n15676, new_n15673, new_n15677);
nor_5  g13329(new_n15677, new_n15672, new_n15678);
xor_4  g13330(new_n15678, new_n15670, new_n15679);
xor_4  g13331(new_n15679, new_n7029, new_n15680);
not_10 g13332(new_n7033, new_n15681);
xor_4  g13333(new_n15676, new_n15673, new_n15682);
nor_5  g13334(new_n15682, new_n15681, new_n15683);
xnor_4 g13335(new_n15682, new_n7033, new_n15684);
nor_5  g13336(new_n11952, new_n7037, new_n15685);
nor_5  g13337(new_n11974, new_n11953, new_n15686);
nor_5  g13338(new_n15686, new_n15685, new_n15687);
and_5  g13339(new_n15687, new_n15684, new_n15688);
nor_5  g13340(new_n15688, new_n15683, new_n15689);
xor_4  g13341(new_n15689, new_n15680, new_n15690);
xor_4  g13342(n21997, n5400, new_n15691);
not_10 g13343(n23923, new_n15692);
nor_5  g13344(n25119, new_n15692, new_n15693);
xor_4  g13345(n25119, n23923, new_n15694);
not_10 g13346(n329, new_n15695);
nor_5  g13347(n1163, new_n15695, new_n15696);
nor_5  g13348(new_n11995, new_n11976, new_n15697);
nor_5  g13349(new_n15697, new_n15696, new_n15698);
nor_5  g13350(new_n15698, new_n15694, new_n15699);
nor_5  g13351(new_n15699, new_n15693, new_n15700);
xor_4  g13352(new_n15700, new_n15691, new_n15701);
xnor_4 g13353(new_n15701, new_n15690, new_n15702);
xor_4  g13354(new_n15698, new_n15694, new_n15703);
xor_4  g13355(new_n15687, new_n15684, new_n15704);
and_5  g13356(new_n15704, new_n15703, new_n15705);
xnor_4 g13357(new_n15704, new_n15703, new_n15706);
not_10 g13358(new_n11975, new_n15707);
nor_5  g13359(new_n11996, new_n15707, new_n15708);
nor_5  g13360(new_n12025, new_n11997, new_n15709);
or_5   g13361(new_n15709, new_n15708, new_n15710);
nor_5  g13362(new_n15710, new_n15706, new_n15711);
nor_5  g13363(new_n15711, new_n15705, new_n15712);
xor_4  g13364(new_n15712, new_n15702, n4215);
or_5   g13365(new_n12902, n2145, new_n15714);
xor_4  g13366(new_n15714, n3582, new_n15715);
xor_4  g13367(new_n15715, n3740, new_n15716_1);
and_5  g13368(new_n12903, n2858, new_n15717);
or_5   g13369(new_n12903, n2858, new_n15718);
and_5  g13370(new_n12927, new_n15718, new_n15719);
nor_5  g13371(new_n15719, new_n15717, new_n15720);
xnor_4 g13372(new_n15720, new_n15716_1, new_n15721);
or_5   g13373(new_n8747, n27089, new_n15722);
xor_4  g13374(new_n15722, n21839, new_n15723);
xor_4  g13375(new_n15723, n22626, new_n15724);
nor_5  g13376(new_n8748, n14440, new_n15725);
xnor_4 g13377(new_n8748, n14440, new_n15726);
nor_5  g13378(new_n8750, n1654, new_n15727);
nor_5  g13379(new_n14308, new_n14305, new_n15728);
nor_5  g13380(new_n15728, new_n15727, new_n15729);
nor_5  g13381(new_n15729, new_n15726, new_n15730);
nor_5  g13382(new_n15730, new_n15725, new_n15731);
xnor_4 g13383(new_n15731, new_n15724, new_n15732);
xor_4  g13384(new_n15732, new_n15721, new_n15733);
xor_4  g13385(new_n15729, new_n15726, new_n15734);
nor_5  g13386(new_n15734, new_n12928, new_n15735);
and_5  g13387(new_n14309, new_n12930, new_n15736);
xnor_4 g13388(new_n14309, new_n12930, new_n15737);
and_5  g13389(new_n12932, new_n9607, new_n15738);
xnor_4 g13390(new_n12932, new_n9607, new_n15739);
or_5   g13391(new_n12936, new_n9609, new_n15740);
xnor_4 g13392(new_n12936, new_n9609, new_n15741);
and_5  g13393(new_n12939, new_n9615, new_n15742);
xnor_4 g13394(new_n12939, new_n9615, new_n15743_1);
and_5  g13395(new_n8582, new_n8570, new_n15744);
nor_5  g13396(new_n8598, new_n8583, new_n15745);
nor_5  g13397(new_n15745, new_n15744, new_n15746);
nor_5  g13398(new_n15746, new_n15743_1, new_n15747);
nor_5  g13399(new_n15747, new_n15742, new_n15748);
not_10 g13400(new_n15748, new_n15749_1);
or_5   g13401(new_n15749_1, new_n15741, new_n15750);
and_5  g13402(new_n15750, new_n15740, new_n15751);
nor_5  g13403(new_n15751, new_n15739, new_n15752);
nor_5  g13404(new_n15752, new_n15738, new_n15753);
nor_5  g13405(new_n15753, new_n15737, new_n15754);
or_5   g13406(new_n15754, new_n15736, new_n15755);
xnor_4 g13407(new_n15734, new_n12928, new_n15756);
nor_5  g13408(new_n15756, new_n15755, new_n15757);
nor_5  g13409(new_n15757, new_n15735, new_n15758);
xnor_4 g13410(new_n15758, new_n15733, new_n15759);
not_10 g13411(n23166, new_n15760);
or_5   g13412(new_n13604, n10611, new_n15761_1);
or_5   g13413(new_n15761_1, n3164, new_n15762_1);
or_5   g13414(new_n15762_1, n11356, new_n15763);
or_5   g13415(new_n15763, n14345, new_n15764);
or_5   g13416(new_n15764, n6381, new_n15765);
or_5   g13417(new_n15765, n10577, new_n15766_1);
xnor_4 g13418(new_n15766_1, new_n15760, new_n15767);
xnor_4 g13419(new_n15767, n9554, new_n15768);
xnor_4 g13420(new_n15765, new_n8268, new_n15769);
nor_5  g13421(new_n15769, n26408, new_n15770);
xnor_4 g13422(new_n15769, n26408, new_n15771);
xnor_4 g13423(new_n15764, new_n8271, new_n15772);
nor_5  g13424(new_n15772, n18227, new_n15773);
xnor_4 g13425(new_n15772, n18227, new_n15774);
xnor_4 g13426(new_n15763, new_n8274, new_n15775);
nor_5  g13427(new_n15775, n7377, new_n15776);
xnor_4 g13428(new_n15775, n7377, new_n15777);
xnor_4 g13429(new_n15762_1, new_n8277, new_n15778);
nor_5  g13430(new_n15778, n11630, new_n15779);
xnor_4 g13431(new_n15761_1, new_n8280, new_n15780_1);
or_5   g13432(new_n15780_1, n13453, new_n15781);
xnor_4 g13433(new_n15780_1, n13453, new_n15782);
and_5  g13434(new_n13605, n7421, new_n15783);
nor_5  g13435(new_n13617, new_n13606, new_n15784);
nor_5  g13436(new_n15784, new_n15783, new_n15785);
not_10 g13437(new_n15785, new_n15786);
or_5   g13438(new_n15786, new_n15782, new_n15787);
and_5  g13439(new_n15787, new_n15781, new_n15788);
xnor_4 g13440(new_n15778, n11630, new_n15789);
nor_5  g13441(new_n15789, new_n15788, new_n15790);
nor_5  g13442(new_n15790, new_n15779, new_n15791);
nor_5  g13443(new_n15791, new_n15777, new_n15792);
nor_5  g13444(new_n15792, new_n15776, new_n15793_1);
nor_5  g13445(new_n15793_1, new_n15774, new_n15794);
nor_5  g13446(new_n15794, new_n15773, new_n15795);
nor_5  g13447(new_n15795, new_n15771, new_n15796);
or_5   g13448(new_n15796, new_n15770, new_n15797);
xnor_4 g13449(new_n15797, new_n15768, new_n15798);
xnor_4 g13450(new_n15798, new_n15759, new_n15799);
xnor_4 g13451(new_n15795, new_n15771, new_n15800);
xor_4  g13452(new_n15756, new_n15755, new_n15801);
nor_5  g13453(new_n15801, new_n15800, new_n15802);
xnor_4 g13454(new_n15801, new_n15800, new_n15803);
xnor_4 g13455(new_n15793_1, new_n15774, new_n15804);
xnor_4 g13456(new_n15753, new_n15737, new_n15805);
nor_5  g13457(new_n15805, new_n15804, new_n15806);
xnor_4 g13458(new_n15805, new_n15804, new_n15807);
xnor_4 g13459(new_n15791, new_n15777, new_n15808);
xnor_4 g13460(new_n15751, new_n15739, new_n15809);
nor_5  g13461(new_n15809, new_n15808, new_n15810);
xnor_4 g13462(new_n15809, new_n15808, new_n15811);
xor_4  g13463(new_n15748, new_n15741, new_n15812_1);
xnor_4 g13464(new_n15789, new_n15788, new_n15813);
nor_5  g13465(new_n15813, new_n15812_1, new_n15814);
xnor_4 g13466(new_n15813, new_n15812_1, new_n15815_1);
xnor_4 g13467(new_n15785, new_n15782, new_n15816_1);
xor_4  g13468(new_n15746, new_n15743_1, new_n15817);
not_10 g13469(new_n15817, new_n15818);
and_5  g13470(new_n15818, new_n15816_1, new_n15819);
xor_4  g13471(new_n15817, new_n15816_1, new_n15820);
nor_5  g13472(new_n13618, new_n8599, new_n15821);
xor_4  g13473(new_n13618, new_n8599, new_n15822);
nor_5  g13474(new_n13620, new_n8614_1, new_n15823);
xnor_4 g13475(new_n13620, new_n8614_1, new_n15824);
nor_5  g13476(new_n13624, new_n8625, new_n15825);
or_5   g13477(new_n13626_1, new_n8620_1, new_n15826);
xnor_4 g13478(new_n13624, new_n8625, new_n15827);
nor_5  g13479(new_n15827, new_n15826, new_n15828);
nor_5  g13480(new_n15828, new_n15825, new_n15829);
nor_5  g13481(new_n15829, new_n15824, new_n15830);
nor_5  g13482(new_n15830, new_n15823, new_n15831_1);
and_5  g13483(new_n15831_1, new_n15822, new_n15832);
nor_5  g13484(new_n15832, new_n15821, new_n15833);
nor_5  g13485(new_n15833, new_n15820, new_n15834);
nor_5  g13486(new_n15834, new_n15819, new_n15835);
nor_5  g13487(new_n15835, new_n15815_1, new_n15836);
nor_5  g13488(new_n15836, new_n15814, new_n15837);
nor_5  g13489(new_n15837, new_n15811, new_n15838);
nor_5  g13490(new_n15838, new_n15810, new_n15839);
nor_5  g13491(new_n15839, new_n15807, new_n15840);
nor_5  g13492(new_n15840, new_n15806, new_n15841);
nor_5  g13493(new_n15841, new_n15803, new_n15842);
or_5   g13494(new_n15842, new_n15802, new_n15843);
xor_4  g13495(new_n15843, new_n15799, n4221);
xor_4  g13496(new_n9526, n18227, new_n15845);
and_5  g13497(new_n9528, n7377, new_n15846_1);
xnor_4 g13498(new_n9528, n7377, new_n15847);
and_5  g13499(new_n9531, n11630, new_n15848);
and_5  g13500(new_n9534, n13453, new_n15849);
nor_5  g13501(new_n11701, new_n11698, new_n15850);
nor_5  g13502(new_n15850, new_n15849, new_n15851);
xnor_4 g13503(new_n9531, n11630, new_n15852);
nor_5  g13504(new_n15852, new_n15851, new_n15853);
nor_5  g13505(new_n15853, new_n15848, new_n15854);
nor_5  g13506(new_n15854, new_n15847, new_n15855);
nor_5  g13507(new_n15855, new_n15846_1, new_n15856);
xor_4  g13508(new_n15856, new_n15845, new_n15857);
xnor_4 g13509(new_n15857, new_n14691, new_n15858);
xor_4  g13510(new_n15854, new_n15847, new_n15859_1);
and_5  g13511(new_n15859_1, new_n14695, new_n15860);
xor_4  g13512(new_n15859_1, new_n7736, new_n15861);
xor_4  g13513(new_n15852, new_n15851, new_n15862);
and_5  g13514(new_n15862, new_n7761, new_n15863);
xnor_4 g13515(new_n15862, new_n7761, new_n15864);
nor_5  g13516(new_n11702, new_n7766, new_n15865);
xnor_4 g13517(new_n11702, new_n7766, new_n15866);
nor_5  g13518(new_n7770, new_n6011, new_n15867);
xnor_4 g13519(new_n7770, new_n6011, new_n15868);
not_10 g13520(new_n6038, new_n15869_1);
nor_5  g13521(new_n7774, new_n15869_1, new_n15870);
xor_4  g13522(new_n7774, new_n6038, new_n15871);
nor_5  g13523(new_n7778, new_n6042, new_n15872);
nor_5  g13524(new_n7781, new_n6046_1, new_n15873);
xnor_4 g13525(new_n7777, new_n6042, new_n15874);
and_5  g13526(new_n15874, new_n15873, new_n15875);
nor_5  g13527(new_n15875, new_n15872, new_n15876);
nor_5  g13528(new_n15876, new_n15871, new_n15877);
nor_5  g13529(new_n15877, new_n15870, new_n15878);
nor_5  g13530(new_n15878, new_n15868, new_n15879);
nor_5  g13531(new_n15879, new_n15867, new_n15880);
nor_5  g13532(new_n15880, new_n15866, new_n15881);
nor_5  g13533(new_n15881, new_n15865, new_n15882);
nor_5  g13534(new_n15882, new_n15864, new_n15883);
nor_5  g13535(new_n15883, new_n15863, new_n15884_1);
nor_5  g13536(new_n15884_1, new_n15861, new_n15885_1);
nor_5  g13537(new_n15885_1, new_n15860, new_n15886);
xnor_4 g13538(new_n15886, new_n15858, n4224);
xor_4  g13539(new_n9652, new_n9651, n4231);
xnor_4 g13540(new_n12779, n9934, new_n15889_1);
nor_5  g13541(new_n12782, n18496, new_n15890);
nor_5  g13542(new_n15268, new_n15261, new_n15891);
nor_5  g13543(new_n15891, new_n15890, new_n15892);
xnor_4 g13544(new_n15892, new_n15889_1, new_n15893);
xnor_4 g13545(new_n15893, n2979, new_n15894);
nor_5  g13546(new_n15269, new_n5385, new_n15895);
nor_5  g13547(new_n15278, new_n15270, new_n15896);
nor_5  g13548(new_n15896, new_n15895, new_n15897);
xor_4  g13549(new_n15897, new_n15894, new_n15898);
xor_4  g13550(new_n15898, new_n10720, new_n15899);
not_10 g13551(new_n10723, new_n15900);
nor_5  g13552(new_n15279, new_n15900, new_n15901);
nor_5  g13553(new_n15289_1, new_n15280, new_n15902);
nor_5  g13554(new_n15902, new_n15901, new_n15903);
xnor_4 g13555(new_n15903, new_n15899, n4266);
xnor_4 g13556(new_n6298, new_n6276_1, n4340);
xnor_4 g13557(new_n14889, new_n12147, new_n15906);
xnor_4 g13558(new_n15906, new_n11791, new_n15907);
nor_5  g13559(new_n14890, new_n11796, new_n15908);
nor_5  g13560(new_n14891_1, new_n14887, new_n15909);
nor_5  g13561(new_n15909, new_n15908, new_n15910);
xor_4  g13562(new_n15910, new_n15907, new_n15911);
xnor_4 g13563(new_n15911, new_n4620, new_n15912);
nor_5  g13564(new_n14892, new_n14886, new_n15913);
nor_5  g13565(new_n15913, new_n14885, new_n15914);
xor_4  g13566(new_n15914, new_n15912, n4374);
xnor_4 g13567(new_n10087, new_n10042, n4401);
xor_4  g13568(new_n11746, new_n11745, n4424);
not_10 g13569(new_n9721, new_n15918_1);
and_5  g13570(new_n15918_1, n1881, new_n15919);
xnor_4 g13571(new_n9721, n1881, new_n15920);
nor_5  g13572(new_n9715, n5834, new_n15921);
xor_4  g13573(new_n9714, n5834, new_n15922_1);
and_5  g13574(new_n9708, n13851, new_n15923);
xor_4  g13575(new_n9707, n13851, new_n15924);
and_5  g13576(new_n9701, n24937, new_n15925);
nor_5  g13577(new_n14794, new_n14787, new_n15926);
nor_5  g13578(new_n15926, new_n15925, new_n15927);
nor_5  g13579(new_n15927, new_n15924, new_n15928);
or_5   g13580(new_n15928, new_n15923, new_n15929);
nor_5  g13581(new_n15929, new_n15922_1, new_n15930);
nor_5  g13582(new_n15930, new_n15921, new_n15931);
and_5  g13583(new_n15931, new_n15920, new_n15932);
nor_5  g13584(new_n15932, new_n15919, new_n15933);
nor_5  g13585(n8827, n4306, new_n15934);
nor_5  g13586(new_n9720, new_n9717, new_n15935);
nor_5  g13587(new_n15935, new_n15934, new_n15936_1);
not_10 g13588(new_n15936_1, new_n15937);
xnor_4 g13589(new_n15937, new_n15933, new_n15938);
xnor_4 g13590(new_n15938, new_n9034, new_n15939);
xor_4  g13591(new_n15931, new_n15920, new_n15940);
and_5  g13592(new_n15940, new_n9038, new_n15941);
xnor_4 g13593(new_n15940, new_n9038, new_n15942);
xnor_4 g13594(new_n15929, new_n15922_1, new_n15943);
and_5  g13595(new_n15943, new_n9042_1, new_n15944);
xor_4  g13596(new_n15927, new_n15924, new_n15945);
nor_5  g13597(new_n15945, new_n9046_1, new_n15946);
xnor_4 g13598(new_n15945, new_n9046_1, new_n15947_1);
nor_5  g13599(new_n14795, new_n9050, new_n15948);
nor_5  g13600(new_n14804, new_n14796, new_n15949);
nor_5  g13601(new_n15949, new_n15948, new_n15950);
nor_5  g13602(new_n15950, new_n15947_1, new_n15951);
nor_5  g13603(new_n15951, new_n15946, new_n15952);
xor_4  g13604(new_n15929, new_n15922_1, new_n15953);
xnor_4 g13605(new_n15953, new_n9042_1, new_n15954);
and_5  g13606(new_n15954, new_n15952, new_n15955);
nor_5  g13607(new_n15955, new_n15944, new_n15956_1);
nor_5  g13608(new_n15956_1, new_n15942, new_n15957);
nor_5  g13609(new_n15957, new_n15941, new_n15958_1);
xnor_4 g13610(new_n15958_1, new_n15939, n4432);
xnor_4 g13611(new_n13348, new_n13347, n4441);
or_5   g13612(n27120, n23065, new_n15961);
nor_5  g13613(new_n15961, n24786, new_n15962);
nand_5 g13614(new_n15962, new_n7875, new_n15963);
or_5   g13615(new_n15963, n19472, new_n15964);
or_5   g13616(new_n15964, n19042, new_n15965);
nor_5  g13617(new_n15965, n1293, new_n15966);
xnor_4 g13618(new_n15966, n13775, new_n15967_1);
xnor_4 g13619(new_n15967_1, new_n15330, new_n15968);
xnor_4 g13620(new_n15965, new_n7866, new_n15969);
nor_5  g13621(new_n15969, new_n15332_1, new_n15970);
xnor_4 g13622(new_n15969, new_n15332_1, new_n15971);
xnor_4 g13623(new_n15964, new_n7869, new_n15972);
nor_5  g13624(new_n15972, new_n15336, new_n15973);
xnor_4 g13625(new_n15963, new_n7872, new_n15974);
nor_5  g13626(new_n15974, new_n7818, new_n15975);
xnor_4 g13627(new_n15974, new_n7818, new_n15976);
xnor_4 g13628(new_n15962, n25370, new_n15977);
and_5  g13629(new_n15977, new_n7820, new_n15978);
xnor_4 g13630(new_n15977, new_n7820, new_n15979_1);
xor_4  g13631(new_n15961, n24786, new_n15980);
nor_5  g13632(new_n15980, new_n7822, new_n15981);
xnor_4 g13633(new_n15980, new_n7822, new_n15982);
xor_4  g13634(n27120, n23065, new_n15983);
nor_5  g13635(new_n15983, new_n7827, new_n15984);
nor_5  g13636(new_n15984, new_n7829, new_n15985);
nor_5  g13637(new_n15985, new_n15982, new_n15986_1);
or_5   g13638(new_n15986_1, new_n15981, new_n15987);
nor_5  g13639(new_n15987, new_n15979_1, new_n15988);
or_5   g13640(new_n15988, new_n15978, new_n15989);
nor_5  g13641(new_n15989, new_n15976, new_n15990);
nor_5  g13642(new_n15990, new_n15975, new_n15991);
xnor_4 g13643(new_n15972, new_n15336, new_n15992);
nor_5  g13644(new_n15992, new_n15991, new_n15993);
nor_5  g13645(new_n15993, new_n15973, new_n15994);
nor_5  g13646(new_n15994, new_n15971, new_n15995);
or_5   g13647(new_n15995, new_n15970, new_n15996);
xor_4  g13648(new_n15996, new_n15968, new_n15997);
nor_5  g13649(new_n10883, n26318, new_n15998);
xnor_4 g13650(new_n15998, n3710, new_n15999);
xnor_4 g13651(new_n15999, new_n4929, new_n16000);
not_10 g13652(new_n4933, new_n16001);
nor_5  g13653(new_n10884, new_n16001, new_n16002);
nor_5  g13654(new_n10916, new_n10885, new_n16003);
or_5   g13655(new_n16003, new_n16002, new_n16004);
xor_4  g13656(new_n16004, new_n16000, new_n16005);
xnor_4 g13657(new_n16005, new_n15997, new_n16006);
xor_4  g13658(new_n10916, new_n10885, new_n16007);
xor_4  g13659(new_n15994, new_n15971, new_n16008);
and_5  g13660(new_n16008, new_n16007, new_n16009);
xnor_4 g13661(new_n16008, new_n16007, new_n16010);
xor_4  g13662(new_n15992, new_n15991, new_n16011);
and_5  g13663(new_n16011, new_n10949, new_n16012);
xor_4  g13664(new_n16011, new_n10949, new_n16013_1);
xor_4  g13665(new_n15989, new_n15976, new_n16014);
nor_5  g13666(new_n16014, new_n10952, new_n16015);
xnor_4 g13667(new_n10909, new_n10908, new_n16016);
xor_4  g13668(new_n15987, new_n15979_1, new_n16017);
nor_5  g13669(new_n16017, new_n16016, new_n16018);
xnor_4 g13670(new_n16017, new_n10956, new_n16019);
xor_4  g13671(new_n15985, new_n15982, new_n16020);
nor_5  g13672(new_n16020, new_n10960, new_n16021);
nand_5 g13673(new_n16020, new_n10960, new_n16022);
xnor_4 g13674(new_n10900, new_n4946, new_n16023);
xnor_4 g13675(new_n15983, new_n7830_1, new_n16024);
and_5  g13676(new_n16024, new_n16023, new_n16025);
or_5   g13677(new_n10970, new_n7846, new_n16026);
xnor_4 g13678(new_n16024, new_n10967, new_n16027);
and_5  g13679(new_n16027, new_n16026, new_n16028);
nor_5  g13680(new_n16028, new_n16025, new_n16029_1);
and_5  g13681(new_n16029_1, new_n16022, new_n16030);
nor_5  g13682(new_n16030, new_n16021, new_n16031);
and_5  g13683(new_n16031, new_n16019, new_n16032);
or_5   g13684(new_n16032, new_n16018, new_n16033);
xnor_4 g13685(new_n16014, new_n10952, new_n16034);
nor_5  g13686(new_n16034, new_n16033, new_n16035);
nor_5  g13687(new_n16035, new_n16015, new_n16036);
and_5  g13688(new_n16036, new_n16013_1, new_n16037);
nor_5  g13689(new_n16037, new_n16012, new_n16038);
nor_5  g13690(new_n16038, new_n16010, new_n16039);
nor_5  g13691(new_n16039, new_n16009, new_n16040);
xnor_4 g13692(new_n16040, new_n16006, n4451);
xnor_4 g13693(new_n11878, new_n11857, new_n16042);
xor_4  g13694(n25494, n6659, new_n16043);
nor_5  g13695(new_n14484, n10117, new_n16044);
xor_4  g13696(n23250, n10117, new_n16045);
nor_5  g13697(n13460, new_n14412_1, new_n16046);
xor_4  g13698(n13460, n11455, new_n16047);
nor_5  g13699(n6104, new_n14415, new_n16048);
xor_4  g13700(n6104, n3945, new_n16049);
nor_5  g13701(new_n14418, n4119, new_n16050);
nor_5  g13702(new_n4786, new_n4767, new_n16051);
nor_5  g13703(new_n16051, new_n16050, new_n16052);
nor_5  g13704(new_n16052, new_n16049, new_n16053);
nor_5  g13705(new_n16053, new_n16048, new_n16054);
nor_5  g13706(new_n16054, new_n16047, new_n16055);
nor_5  g13707(new_n16055, new_n16046, new_n16056);
nor_5  g13708(new_n16056, new_n16045, new_n16057);
nor_5  g13709(new_n16057, new_n16044, new_n16058);
xor_4  g13710(new_n16058, new_n16043, new_n16059);
xnor_4 g13711(new_n16059, new_n16042, new_n16060_1);
xnor_4 g13712(new_n11876, new_n11861, new_n16061);
xor_4  g13713(new_n16056, new_n16045, new_n16062_1);
nor_5  g13714(new_n16062_1, new_n16061, new_n16063);
xnor_4 g13715(new_n16062_1, new_n16061, new_n16064);
xnor_4 g13716(new_n11874, new_n11865, new_n16065);
xor_4  g13717(new_n16054, new_n16047, new_n16066);
nor_5  g13718(new_n16066, new_n16065, new_n16067);
xnor_4 g13719(new_n16066, new_n11899, new_n16068_1);
xor_4  g13720(new_n16052, new_n16049, new_n16069);
and_5  g13721(new_n16069, new_n11903, new_n16070);
xnor_4 g13722(new_n16069, new_n11903, new_n16071);
and_5  g13723(new_n4787, new_n4766_1, new_n16072);
nor_5  g13724(new_n4817, new_n4788, new_n16073);
nor_5  g13725(new_n16073, new_n16072, new_n16074);
nor_5  g13726(new_n16074, new_n16071, new_n16075);
nor_5  g13727(new_n16075, new_n16070, new_n16076);
and_5  g13728(new_n16076, new_n16068_1, new_n16077);
nor_5  g13729(new_n16077, new_n16067, new_n16078);
nor_5  g13730(new_n16078, new_n16064, new_n16079);
or_5   g13731(new_n16079, new_n16063, new_n16080_1);
xor_4  g13732(new_n16080_1, new_n16060_1, n4476);
and_5  g13733(new_n3757, new_n12570, new_n16082);
nand_5 g13734(new_n16082, new_n12567, new_n16083);
or_5   g13735(new_n16083, n18452, new_n16084);
or_5   g13736(new_n16084, n13137, new_n16085);
nor_5  g13737(new_n16085, n1831, new_n16086);
xor_4  g13738(new_n16086, new_n5689, new_n16087);
xnor_4 g13739(new_n16085, new_n12558, new_n16088);
nor_5  g13740(new_n16088, new_n5694, new_n16089);
xnor_4 g13741(new_n16084, new_n12561, new_n16090);
nor_5  g13742(new_n16090, new_n5696_1, new_n16091);
xnor_4 g13743(new_n16090, new_n5696_1, new_n16092);
xnor_4 g13744(new_n16083, new_n12564, new_n16093);
nor_5  g13745(new_n16093, new_n5700_1, new_n16094);
xnor_4 g13746(new_n16093, new_n5700_1, new_n16095);
xnor_4 g13747(new_n16082, n21317, new_n16096);
and_5  g13748(new_n16096, new_n5705, new_n16097);
xnor_4 g13749(new_n16096, new_n5705, new_n16098_1);
and_5  g13750(new_n3786, new_n3758_1, new_n16099);
nor_5  g13751(new_n3813, new_n3787, new_n16100);
nor_5  g13752(new_n16100, new_n16099, new_n16101);
nor_5  g13753(new_n16101, new_n16098_1, new_n16102);
or_5   g13754(new_n16102, new_n16097, new_n16103);
nor_5  g13755(new_n16103, new_n16095, new_n16104);
nor_5  g13756(new_n16104, new_n16094, new_n16105);
nor_5  g13757(new_n16105, new_n16092, new_n16106);
nor_5  g13758(new_n16106, new_n16091, new_n16107);
xnor_4 g13759(new_n16088, new_n5694, new_n16108);
nor_5  g13760(new_n16108, new_n16107, new_n16109);
nor_5  g13761(new_n16109, new_n16089, new_n16110_1);
xnor_4 g13762(new_n16110_1, new_n16087, new_n16111);
xnor_4 g13763(new_n16111, new_n10516, new_n16112);
xor_4  g13764(new_n16108, new_n16107, new_n16113);
and_5  g13765(new_n16113, new_n10520, new_n16114);
xnor_4 g13766(new_n16113, new_n10520, new_n16115);
xor_4  g13767(new_n16105, new_n16092, new_n16116);
and_5  g13768(new_n16116, new_n10523, new_n16117);
xnor_4 g13769(new_n16116, new_n10523, new_n16118);
xor_4  g13770(new_n16103, new_n16095, new_n16119);
and_5  g13771(new_n16119, new_n10528, new_n16120);
xnor_4 g13772(new_n16119, new_n10528, new_n16121);
xor_4  g13773(new_n16101, new_n16098_1, new_n16122);
nor_5  g13774(new_n16122, new_n10533, new_n16123);
xnor_4 g13775(new_n16122, new_n10533, new_n16124);
nor_5  g13776(new_n3814, new_n3751, new_n16125);
nor_5  g13777(new_n3840, new_n3815, new_n16126);
nor_5  g13778(new_n16126, new_n16125, new_n16127);
nor_5  g13779(new_n16127, new_n16124, new_n16128);
nor_5  g13780(new_n16128, new_n16123, new_n16129);
nor_5  g13781(new_n16129, new_n16121, new_n16130);
nor_5  g13782(new_n16130, new_n16120, new_n16131);
nor_5  g13783(new_n16131, new_n16118, new_n16132);
nor_5  g13784(new_n16132, new_n16117, new_n16133);
nor_5  g13785(new_n16133, new_n16115, new_n16134);
nor_5  g13786(new_n16134, new_n16114, new_n16135);
xnor_4 g13787(new_n16135, new_n16112, n4478);
xnor_4 g13788(new_n11282, new_n11252, n4529);
xnor_4 g13789(new_n5618, new_n5579_1, n4552);
xnor_4 g13790(new_n5614, new_n5587, n4595);
xnor_4 g13791(new_n12884, new_n12850, n4624);
not_10 g13792(new_n7021, new_n16141);
or_5   g13793(new_n15668, n2659, new_n16142_1);
xor_4  g13794(new_n16142_1, n2858, new_n16143);
nor_5  g13795(new_n16143, n14899, new_n16144);
xnor_4 g13796(new_n16143, n14899, new_n16145);
nor_5  g13797(new_n15669, n18444, new_n16146);
nor_5  g13798(new_n15678, new_n15670, new_n16147);
nor_5  g13799(new_n16147, new_n16146, new_n16148);
nor_5  g13800(new_n16148, new_n16145, new_n16149);
or_5   g13801(new_n16149, new_n16144, new_n16150);
or_5   g13802(new_n16142_1, n2858, new_n16151);
xor_4  g13803(new_n16151, n3740, new_n16152);
xnor_4 g13804(new_n16152, n3506, new_n16153);
xnor_4 g13805(new_n16153, new_n16150, new_n16154);
nor_5  g13806(new_n16154, new_n16141, new_n16155);
xor_4  g13807(new_n16154, new_n7021, new_n16156);
not_10 g13808(new_n7025, new_n16157);
xor_4  g13809(new_n16148, new_n16145, new_n16158_1);
nor_5  g13810(new_n16158_1, new_n16157, new_n16159);
xor_4  g13811(new_n16158_1, new_n7025, new_n16160);
not_10 g13812(new_n7029, new_n16161);
nor_5  g13813(new_n15679, new_n16161, new_n16162);
nor_5  g13814(new_n15689, new_n15680, new_n16163);
nor_5  g13815(new_n16163, new_n16162, new_n16164);
nor_5  g13816(new_n16164, new_n16160, new_n16165);
nor_5  g13817(new_n16165, new_n16159, new_n16166);
nor_5  g13818(new_n16166, new_n16156, new_n16167_1);
or_5   g13819(new_n16167_1, new_n16155, new_n16168);
nor_5  g13820(new_n16151, n3740, new_n16169);
and_5  g13821(new_n16152, n3506, new_n16170);
nor_5  g13822(new_n16152, n3506, new_n16171);
nor_5  g13823(new_n16171, new_n16150, new_n16172);
or_5   g13824(new_n16172, new_n16170, new_n16173);
or_5   g13825(new_n16173, new_n16169, new_n16174);
xnor_4 g13826(new_n16174, new_n16168, new_n16175);
xnor_4 g13827(new_n16175, new_n6970, new_n16176);
xnor_4 g13828(new_n16176, new_n12311, new_n16177);
xor_4  g13829(new_n16166, new_n16156, new_n16178);
nor_5  g13830(new_n16178, new_n7141, new_n16179);
xor_4  g13831(new_n16164, new_n16160, new_n16180);
nor_5  g13832(new_n16180, new_n7146, new_n16181);
xnor_4 g13833(new_n16180, new_n7146, new_n16182);
nor_5  g13834(new_n15690, new_n7151, new_n16183);
xnor_4 g13835(new_n15690, new_n7151, new_n16184);
nor_5  g13836(new_n15704, new_n7155, new_n16185_1);
xor_4  g13837(new_n15704, new_n7155, new_n16186);
nor_5  g13838(new_n11975, new_n7159, new_n16187);
and_5  g13839(new_n11999, new_n7163, new_n16188);
nor_5  g13840(new_n15542, new_n15529, new_n16189);
or_5   g13841(new_n16189, new_n16188, new_n16190);
xnor_4 g13842(new_n11975, new_n7159, new_n16191);
nor_5  g13843(new_n16191, new_n16190, new_n16192);
nor_5  g13844(new_n16192, new_n16187, new_n16193);
and_5  g13845(new_n16193, new_n16186, new_n16194);
nor_5  g13846(new_n16194, new_n16185_1, new_n16195);
nor_5  g13847(new_n16195, new_n16184, new_n16196_1);
nor_5  g13848(new_n16196_1, new_n16183, new_n16197);
nor_5  g13849(new_n16197, new_n16182, new_n16198);
nor_5  g13850(new_n16198, new_n16181, new_n16199);
xnor_4 g13851(new_n16178, new_n7141, new_n16200);
nor_5  g13852(new_n16200, new_n16199, new_n16201);
or_5   g13853(new_n16201, new_n16179, new_n16202);
xor_4  g13854(new_n16202, new_n16177, n4646);
xnor_4 g13855(new_n12892_1, new_n12834, n4674);
xor_4  g13856(n7057, n3480, new_n16205);
nor_5  g13857(new_n6945, n8381, new_n16206_1);
nor_5  g13858(n16722, new_n8602, new_n16207);
nor_5  g13859(n20235, new_n6948, new_n16208);
or_5   g13860(new_n4660, n11486, new_n16209);
nor_5  g13861(new_n6951, n12495, new_n16210);
and_5  g13862(new_n16210, new_n16209, new_n16211);
nor_5  g13863(new_n16211, new_n16208, new_n16212);
nor_5  g13864(new_n16212, new_n16207, new_n16213);
nor_5  g13865(new_n16213, new_n16206_1, new_n16214);
xor_4  g13866(new_n16214, new_n16205, new_n16215_1);
xnor_4 g13867(new_n16215_1, new_n2934, new_n16216);
xnor_4 g13868(n16722, n8381, new_n16217_1);
xnor_4 g13869(new_n16217_1, new_n16212, new_n16218_1);
and_5  g13870(new_n16218_1, new_n2939, new_n16219_1);
xnor_4 g13871(new_n16218_1, new_n2939, new_n16220);
xnor_4 g13872(n13781, n12495, new_n16221);
or_5   g13873(new_n16221, new_n2945, new_n16222);
and_5  g13874(new_n16222, new_n2950, new_n16223_1);
xor_4  g13875(new_n16222, new_n2950, new_n16224);
xor_4  g13876(n20235, n11486, new_n16225);
xnor_4 g13877(new_n16225, new_n16210, new_n16226);
and_5  g13878(new_n16226, new_n16224, new_n16227);
nor_5  g13879(new_n16227, new_n16223_1, new_n16228);
nor_5  g13880(new_n16228, new_n16220, new_n16229);
or_5   g13881(new_n16229, new_n16219_1, new_n16230_1);
xor_4  g13882(new_n16230_1, new_n16216, n4693);
xnor_4 g13883(new_n9654, new_n9645, n4731);
and_5  g13884(new_n5526, n8526, new_n16233);
nor_5  g13885(new_n5569, new_n5527, new_n16234);
nor_5  g13886(new_n16234, new_n16233, new_n16235);
nor_5  g13887(n21784, n3582, new_n16236);
nor_5  g13888(new_n5525, new_n5492, new_n16237);
or_5   g13889(new_n16237, new_n16236, new_n16238);
nor_5  g13890(new_n16238, new_n16235, new_n16239);
xor_4  g13891(new_n16239, new_n13931, new_n16240);
xor_4  g13892(new_n16238, new_n16235, new_n16241);
nor_5  g13893(new_n16241, new_n13934, new_n16242);
xnor_4 g13894(new_n16241, new_n13934, new_n16243_1);
not_10 g13895(new_n5570, new_n16244);
and_5  g13896(new_n11636, new_n16244, new_n16245);
nor_5  g13897(new_n11674_1, new_n11637, new_n16246);
nor_5  g13898(new_n16246, new_n16245, new_n16247_1);
nor_5  g13899(new_n16247_1, new_n16243_1, new_n16248);
nor_5  g13900(new_n16248, new_n16242, new_n16249);
xnor_4 g13901(new_n16249, new_n16240, n4745);
xor_4  g13902(new_n5718, n6773, new_n16251);
xor_4  g13903(new_n16251, new_n8814, n4747);
xnor_4 g13904(new_n5288, new_n5287, n4766);
xnor_4 g13905(new_n12395, new_n12378, n4770);
xor_4  g13906(new_n14915, new_n14131, n4777);
xor_4  g13907(n17959, n6861, new_n16256);
and_5  g13908(n19357, new_n5039, new_n16257);
xor_4  g13909(n19357, n7566, new_n16258);
and_5  g13910(new_n5042, n2328, new_n16259);
xor_4  g13911(n7731, n2328, new_n16260);
nor_5  g13912(n15053, new_n5045, new_n16261);
nor_5  g13913(new_n14424, n12341, new_n16262);
nor_5  g13914(n25471, new_n5048, new_n16263);
or_5   g13915(new_n4682, n20986, new_n16264);
and_5  g13916(new_n4671, n12384, new_n16265);
and_5  g13917(new_n16265, new_n16264, new_n16266);
nor_5  g13918(new_n16266, new_n16263, new_n16267);
nor_5  g13919(new_n16267, new_n16262, new_n16268);
or_5   g13920(new_n16268, new_n16261, new_n16269);
nor_5  g13921(new_n16269, new_n16260, new_n16270);
nor_5  g13922(new_n16270, new_n16259, new_n16271);
nor_5  g13923(new_n16271, new_n16258, new_n16272);
nor_5  g13924(new_n16272, new_n16257, new_n16273);
xor_4  g13925(new_n16273, new_n16256, new_n16274);
not_10 g13926(n11580, new_n16275_1);
nor_5  g13927(n20077, n6794, new_n16276);
not_10 g13928(new_n16276, new_n16277);
nor_5  g13929(new_n16277, n15636, new_n16278);
and_5  g13930(new_n16278, new_n5089, new_n16279_1);
and_5  g13931(new_n16279_1, new_n5086, new_n16280);
xnor_4 g13932(new_n16280, n22660, new_n16281);
xnor_4 g13933(new_n16281, new_n16275_1, new_n16282);
not_10 g13934(n15884, new_n16283);
xnor_4 g13935(new_n16279_1, n1777, new_n16284);
nor_5  g13936(new_n16284, new_n16283, new_n16285);
xnor_4 g13937(new_n16284, new_n16283, new_n16286);
xnor_4 g13938(new_n16278, new_n5089, new_n16287);
and_5  g13939(new_n16287, n6356, new_n16288);
xnor_4 g13940(new_n16287, n6356, new_n16289);
not_10 g13941(n27104, new_n16290);
xnor_4 g13942(new_n16276, n15636, new_n16291);
nor_5  g13943(new_n16291, new_n16290, new_n16292);
xor_4  g13944(new_n16291, n27104, new_n16293);
xnor_4 g13945(n20077, n6794, new_n16294);
and_5  g13946(new_n16294, n27188, new_n16295);
or_5   g13947(n6794, new_n8174, new_n16296);
xnor_4 g13948(new_n16294, n27188, new_n16297);
nor_5  g13949(new_n16297, new_n16296, new_n16298);
nor_5  g13950(new_n16298, new_n16295, new_n16299);
nor_5  g13951(new_n16299, new_n16293, new_n16300);
nor_5  g13952(new_n16300, new_n16292, new_n16301);
nor_5  g13953(new_n16301, new_n16289, new_n16302);
nor_5  g13954(new_n16302, new_n16288, new_n16303);
nor_5  g13955(new_n16303, new_n16286, new_n16304);
nor_5  g13956(new_n16304, new_n16285, new_n16305);
xor_4  g13957(new_n16305, new_n16282, new_n16306);
xnor_4 g13958(new_n16306, new_n14395, new_n16307);
xor_4  g13959(new_n16303, new_n16286, new_n16308);
nor_5  g13960(new_n16308, new_n13833, new_n16309);
xor_4  g13961(new_n16301, new_n16289, new_n16310);
and_5  g13962(new_n16310, new_n13836, new_n16311);
xor_4  g13963(new_n16310, new_n13836, new_n16312);
xor_4  g13964(new_n16299, new_n16293, new_n16313);
nor_5  g13965(new_n16313, new_n4658, new_n16314);
xnor_4 g13966(new_n16313, new_n4658, new_n16315);
xor_4  g13967(new_n16297, new_n16296, new_n16316);
nor_5  g13968(new_n16316, new_n4665_1, new_n16317);
xnor_4 g13969(n6794, n6611, new_n16318);
or_5   g13970(new_n16318, new_n4661, new_n16319);
xnor_4 g13971(new_n16316, new_n4665_1, new_n16320);
nor_5  g13972(new_n16320, new_n16319, new_n16321);
nor_5  g13973(new_n16321, new_n16317, new_n16322_1);
nor_5  g13974(new_n16322_1, new_n16315, new_n16323);
nor_5  g13975(new_n16323, new_n16314, new_n16324);
and_5  g13976(new_n16324, new_n16312, new_n16325);
or_5   g13977(new_n16325, new_n16311, new_n16326);
xnor_4 g13978(new_n16308, new_n13833, new_n16327_1);
nor_5  g13979(new_n16327_1, new_n16326, new_n16328);
nor_5  g13980(new_n16328, new_n16309, new_n16329);
xor_4  g13981(new_n16329, new_n16307, new_n16330);
xnor_4 g13982(new_n16330, new_n16274, new_n16331);
xor_4  g13983(new_n16271, new_n16258, new_n16332);
xor_4  g13984(new_n16327_1, new_n16326, new_n16333);
nor_5  g13985(new_n16333, new_n16332, new_n16334);
xnor_4 g13986(new_n16333, new_n16332, new_n16335);
xnor_4 g13987(new_n16324, new_n16312, new_n16336);
xor_4  g13988(new_n16269, new_n16260, new_n16337);
nor_5  g13989(new_n16337, new_n16336, new_n16338);
xnor_4 g13990(new_n16337, new_n16336, new_n16339);
xor_4  g13991(new_n16322_1, new_n16315, new_n16340);
not_10 g13992(new_n16340, new_n16341);
xnor_4 g13993(n15053, n12341, new_n16342);
xnor_4 g13994(new_n16342, new_n16267, new_n16343);
and_5  g13995(new_n16343, new_n16341, new_n16344);
xor_4  g13996(new_n16343, new_n16340, new_n16345);
xnor_4 g13997(new_n16318, new_n4661, new_n16346);
xnor_4 g13998(n16502, n12384, new_n16347);
or_5   g13999(new_n16347, new_n16346, new_n16348);
xor_4  g14000(n25471, n20986, new_n16349);
xnor_4 g14001(new_n16349, new_n16265, new_n16350_1);
and_5  g14002(new_n16350_1, new_n16348, new_n16351);
xnor_4 g14003(new_n16320, new_n16319, new_n16352);
xor_4  g14004(new_n16350_1, new_n16348, new_n16353);
and_5  g14005(new_n16353, new_n16352, new_n16354);
nor_5  g14006(new_n16354, new_n16351, new_n16355);
nor_5  g14007(new_n16355, new_n16345, new_n16356);
nor_5  g14008(new_n16356, new_n16344, new_n16357);
nor_5  g14009(new_n16357, new_n16339, new_n16358);
nor_5  g14010(new_n16358, new_n16338, new_n16359);
nor_5  g14011(new_n16359, new_n16335, new_n16360);
or_5   g14012(new_n16360, new_n16334, new_n16361);
xor_4  g14013(new_n16361, new_n16331, n4785);
xnor_4 g14014(new_n12687, new_n12655, n4804);
xnor_4 g14015(new_n14140, new_n14123, n4810);
nor_5  g14016(new_n15760, n18105, new_n16365);
nor_5  g14017(new_n8309_1, new_n8267_1, new_n16366);
nor_5  g14018(new_n16366, new_n16365, new_n16367_1);
nor_5  g14019(new_n9722, new_n7239, new_n16368);
nor_5  g14020(new_n9767_1, new_n9723, new_n16369);
nor_5  g14021(new_n16369, new_n16368, new_n16370);
or_5   g14022(new_n15918_1, new_n9716, new_n16371);
and_5  g14023(new_n15936_1, new_n16371, new_n16372);
not_10 g14024(new_n15934, new_n16373);
nor_5  g14025(new_n16371, new_n16373, new_n16374);
nor_5  g14026(new_n16374, new_n16372, new_n16375);
xnor_4 g14027(new_n16375, new_n7298_1, new_n16376_1);
xnor_4 g14028(new_n16376_1, new_n16370, new_n16377);
and_5  g14029(new_n16377, new_n16367_1, new_n16378);
xnor_4 g14030(new_n16377, new_n16367_1, new_n16379_1);
and_5  g14031(new_n9768, new_n9663, new_n16380);
nor_5  g14032(new_n9812, new_n9769, new_n16381);
nor_5  g14033(new_n16381, new_n16380, new_n16382);
nor_5  g14034(new_n16382, new_n16379_1, new_n16383);
or_5   g14035(new_n16383, new_n16378, new_n16384);
or_5   g14036(new_n16375, new_n7297, new_n16385);
and_5  g14037(new_n16385, new_n16370, new_n16386);
and_5  g14038(new_n16375, new_n7297, new_n16387);
or_5   g14039(new_n16387, new_n16374, new_n16388);
nor_5  g14040(new_n16388, new_n16386, new_n16389);
or_5   g14041(new_n16389, new_n16384, n4814);
xnor_4 g14042(new_n14717, new_n14716, n4850);
xnor_4 g14043(new_n15514, new_n15480, n4891);
xnor_4 g14044(new_n15660, new_n15641, n4925);
xnor_4 g14045(new_n14723, new_n14705, n4947);
xor_4  g14046(new_n8541, new_n8539, n4952);
xor_4  g14047(n25068, n6790, new_n16396_1);
nor_5  g14048(n22879, new_n7258, new_n16397);
xor_4  g14049(n22879, n2331, new_n16398_1);
nor_5  g14050(new_n7262, n2117, new_n16399);
xor_4  g14051(n22631, n2117, new_n16400);
and_5  g14052(new_n7266, n5882, new_n16401);
nor_5  g14053(new_n7266, n5882, new_n16402);
and_5  g14054(new_n7270, n11775, new_n16403);
not_10 g14055(n27134, new_n16404);
nor_5  g14056(new_n16404, n4588, new_n16405);
or_5   g14057(new_n7270, n11775, new_n16406_1);
and_5  g14058(new_n16406_1, new_n16405, new_n16407_1);
nor_5  g14059(new_n16407_1, new_n16403, new_n16408);
nor_5  g14060(new_n16408, new_n16402, new_n16409);
or_5   g14061(new_n16409, new_n16401, new_n16410);
nor_5  g14062(new_n16410, new_n16400, new_n16411);
nor_5  g14063(new_n16411, new_n16399, new_n16412);
nor_5  g14064(new_n16412, new_n16398_1, new_n16413);
nor_5  g14065(new_n16413, new_n16397, new_n16414);
xor_4  g14066(new_n16414, new_n16396_1, new_n16415);
xnor_4 g14067(new_n16415, new_n13788, new_n16416);
xor_4  g14068(new_n16412, new_n16398_1, new_n16417);
nor_5  g14069(new_n16417, new_n13792, new_n16418);
xnor_4 g14070(new_n16417, new_n13792, new_n16419_1);
xor_4  g14071(new_n16410, new_n16400, new_n16420);
nor_5  g14072(new_n16420, new_n13796, new_n16421);
xnor_4 g14073(new_n16420, new_n13796, new_n16422);
xnor_4 g14074(n16743, n5882, new_n16423);
xnor_4 g14075(new_n16423, new_n16408, new_n16424_1);
nor_5  g14076(new_n16424_1, new_n13800, new_n16425);
xnor_4 g14077(new_n16424_1, new_n13800, new_n16426);
xor_4  g14078(n15258, n11775, new_n16427);
xnor_4 g14079(new_n16427, new_n16405, new_n16428_1);
nor_5  g14080(new_n16428_1, new_n13804, new_n16429);
or_5   g14081(new_n13600, new_n13599, new_n16430);
xnor_4 g14082(new_n16428_1, new_n13804, new_n16431);
nor_5  g14083(new_n16431, new_n16430, new_n16432);
nor_5  g14084(new_n16432, new_n16429, new_n16433_1);
nor_5  g14085(new_n16433_1, new_n16426, new_n16434);
or_5   g14086(new_n16434, new_n16425, new_n16435);
nor_5  g14087(new_n16435, new_n16422, new_n16436);
nor_5  g14088(new_n16436, new_n16421, new_n16437);
nor_5  g14089(new_n16437, new_n16419_1, new_n16438);
or_5   g14090(new_n16438, new_n16418, new_n16439_1);
xor_4  g14091(new_n16439_1, new_n16416, new_n16440_1);
xnor_4 g14092(new_n16440_1, new_n13728, new_n16441);
xnor_4 g14093(new_n16437, new_n16419_1, new_n16442);
nor_5  g14094(new_n16442, new_n13731, new_n16443);
xnor_4 g14095(new_n16442, new_n13731, new_n16444);
xor_4  g14096(new_n16435, new_n16422, new_n16445_1);
and_5  g14097(new_n16445_1, new_n12258, new_n16446);
xnor_4 g14098(new_n16445_1, new_n12258, new_n16447);
xor_4  g14099(new_n16433_1, new_n16426, new_n16448);
nor_5  g14100(new_n16448, new_n12262, new_n16449);
xnor_4 g14101(new_n16448, new_n12262, new_n16450);
nor_5  g14102(new_n13601, new_n9006, new_n16451);
nor_5  g14103(new_n16451, new_n12272, new_n16452);
xnor_4 g14104(new_n16451, new_n12272, new_n16453);
xor_4  g14105(new_n16431, new_n16430, new_n16454);
nor_5  g14106(new_n16454, new_n16453, new_n16455);
nor_5  g14107(new_n16455, new_n16452, new_n16456);
nor_5  g14108(new_n16456, new_n16450, new_n16457);
nor_5  g14109(new_n16457, new_n16449, new_n16458);
nor_5  g14110(new_n16458, new_n16447, new_n16459);
nor_5  g14111(new_n16459, new_n16446, new_n16460_1);
nor_5  g14112(new_n16460_1, new_n16444, new_n16461);
nor_5  g14113(new_n16461, new_n16443, new_n16462);
xnor_4 g14114(new_n16462, new_n16441, n4966);
xnor_4 g14115(new_n15954, new_n15952, n4972);
or_5   g14116(new_n6834, n23895, new_n16465);
xnor_4 g14117(new_n6834, n23895, new_n16466);
and_5  g14118(new_n6839, n17351, new_n16467);
xnor_4 g14119(new_n6839, n17351, new_n16468);
nor_5  g14120(new_n6845, new_n5030, new_n16469);
nor_5  g14121(new_n15358, new_n15347, new_n16470);
nor_5  g14122(new_n16470, new_n16469, new_n16471);
nor_5  g14123(new_n16471, new_n16468, new_n16472);
nor_5  g14124(new_n16472, new_n16467, new_n16473);
not_10 g14125(new_n16473, new_n16474);
or_5   g14126(new_n16474, new_n16466, new_n16475);
nand_5 g14127(new_n16475, new_n16465, new_n16476_1);
or_5   g14128(new_n16476_1, new_n6830, new_n16477);
or_5   g14129(new_n15316, n2289, new_n16478);
or_5   g14130(new_n16478, n23697, new_n16479);
xnor_4 g14131(new_n16479, new_n6744, new_n16480);
xor_4  g14132(new_n16480, n7593, new_n16481_1);
xnor_4 g14133(new_n16478, new_n6747, new_n16482_1);
and_5  g14134(new_n16482_1, n337, new_n16483);
nor_5  g14135(new_n16482_1, n337, new_n16484);
and_5  g14136(new_n15317, n3228, new_n16485);
or_5   g14137(new_n15317, n3228, new_n16486);
and_5  g14138(new_n15329, new_n16486, new_n16487);
nor_5  g14139(new_n16487, new_n16485, new_n16488);
nor_5  g14140(new_n16488, new_n16484, new_n16489);
nor_5  g14141(new_n16489, new_n16483, new_n16490);
xnor_4 g14142(new_n16490, new_n16481_1, new_n16491);
nor_5  g14143(new_n16491, n25972, new_n16492);
xnor_4 g14144(new_n16491, n25972, new_n16493_1);
xor_4  g14145(new_n16482_1, n337, new_n16494);
xnor_4 g14146(new_n16494, new_n16488, new_n16495);
nor_5  g14147(new_n16495, n21915, new_n16496);
nor_5  g14148(new_n15330, n13775, new_n16497);
nor_5  g14149(new_n15345_1, new_n15331, new_n16498);
nor_5  g14150(new_n16498, new_n16497, new_n16499);
xnor_4 g14151(new_n16495, n21915, new_n16500);
nor_5  g14152(new_n16500, new_n16499, new_n16501);
nor_5  g14153(new_n16501, new_n16496, new_n16502_1);
nor_5  g14154(new_n16502_1, new_n16493_1, new_n16503);
or_5   g14155(new_n16503, new_n16492, new_n16504);
nor_5  g14156(new_n16479, n2978, new_n16505);
and_5  g14157(new_n16480, n7593, new_n16506_1);
nor_5  g14158(new_n16480, n7593, new_n16507_1);
nor_5  g14159(new_n16490, new_n16507_1, new_n16508);
or_5   g14160(new_n16508, new_n16506_1, new_n16509);
nor_5  g14161(new_n16509, new_n16505, new_n16510);
not_10 g14162(new_n16510, new_n16511);
nor_5  g14163(new_n16511, new_n16504, new_n16512);
xor_4  g14164(new_n16476_1, new_n6830, new_n16513);
xnor_4 g14165(new_n16510, new_n16504, new_n16514);
nor_5  g14166(new_n16514, new_n16513, new_n16515);
xor_4  g14167(new_n16514, new_n16513, new_n16516_1);
xnor_4 g14168(new_n16473, new_n16466, new_n16517_1);
xor_4  g14169(new_n16502_1, new_n16493_1, new_n16518);
nor_5  g14170(new_n16518, new_n16517_1, new_n16519);
xnor_4 g14171(new_n16518, new_n16517_1, new_n16520);
xor_4  g14172(new_n16471, new_n16468, new_n16521_1);
not_10 g14173(new_n16521_1, new_n16522);
xor_4  g14174(new_n16500, new_n16499, new_n16523);
nor_5  g14175(new_n16523, new_n16522, new_n16524_1);
nor_5  g14176(new_n15359, new_n15346, new_n16525);
nor_5  g14177(new_n15375, new_n15360, new_n16526);
or_5   g14178(new_n16526, new_n16525, new_n16527_1);
xnor_4 g14179(new_n16523, new_n16522, new_n16528);
nor_5  g14180(new_n16528, new_n16527_1, new_n16529);
nor_5  g14181(new_n16529, new_n16524_1, new_n16530);
nor_5  g14182(new_n16530, new_n16520, new_n16531);
nor_5  g14183(new_n16531, new_n16519, new_n16532);
and_5  g14184(new_n16532, new_n16516_1, new_n16533);
nor_5  g14185(new_n16533, new_n16515, new_n16534);
xnor_4 g14186(new_n16534, new_n16512, new_n16535);
xnor_4 g14187(new_n16535, new_n16477, n5011);
not_10 g14188(n11220, new_n16537);
nor_5  g14189(new_n16537, n2944, new_n16538);
xor_4  g14190(n11220, n2944, new_n16539);
not_10 g14191(n22379, new_n16540);
nor_5  g14192(new_n16540, n767, new_n16541);
nor_5  g14193(new_n2806, new_n2767, new_n16542);
nor_5  g14194(new_n16542, new_n16541, new_n16543);
nor_5  g14195(new_n16543, new_n16539, new_n16544_1);
nor_5  g14196(new_n16544_1, new_n16538, new_n16545);
and_5  g14197(n16544, n2160, new_n16546);
or_5   g14198(n16544, n2160, new_n16547);
nor_5  g14199(n10763, n6814, new_n16548);
nor_5  g14200(new_n2837, new_n2808, new_n16549);
nor_5  g14201(new_n16549, new_n16548, new_n16550);
and_5  g14202(new_n16550, new_n16547, new_n16551);
nor_5  g14203(new_n16551, new_n16546, new_n16552);
nor_5  g14204(new_n16552, new_n13661, new_n16553);
xnor_4 g14205(new_n16552, new_n13661, new_n16554_1);
xnor_4 g14206(n16544, n2160, new_n16555);
xnor_4 g14207(new_n16555, new_n16550, new_n16556);
and_5  g14208(new_n16556, new_n13639, new_n16557);
xnor_4 g14209(new_n16556, new_n13639, new_n16558);
and_5  g14210(new_n2869, new_n2838, new_n16559);
nor_5  g14211(new_n2915, new_n2870, new_n16560);
nor_5  g14212(new_n16560, new_n16559, new_n16561);
nor_5  g14213(new_n16561, new_n16558, new_n16562);
nor_5  g14214(new_n16562, new_n16557, new_n16563);
nor_5  g14215(new_n16563, new_n16554_1, new_n16564);
nor_5  g14216(new_n16564, new_n16553, new_n16565);
not_10 g14217(new_n16565, new_n16566);
and_5  g14218(new_n16566, new_n16545, new_n16567);
xor_4  g14219(new_n16563, new_n16554_1, new_n16568);
nor_5  g14220(new_n16568, new_n16545, new_n16569);
and_5  g14221(new_n16568, new_n16545, new_n16570);
xor_4  g14222(new_n16543, new_n16539, new_n16571);
xor_4  g14223(new_n16561, new_n16558, new_n16572);
nor_5  g14224(new_n16572, new_n16571, new_n16573);
xnor_4 g14225(new_n16572, new_n16571, new_n16574);
nor_5  g14226(new_n2916, new_n2807, new_n16575);
nor_5  g14227(new_n2965, new_n2917, new_n16576);
nor_5  g14228(new_n16576, new_n16575, new_n16577);
nor_5  g14229(new_n16577, new_n16574, new_n16578);
nor_5  g14230(new_n16578, new_n16573, new_n16579);
nor_5  g14231(new_n16579, new_n16570, new_n16580);
nor_5  g14232(new_n16580, new_n16569, new_n16581);
nor_5  g14233(new_n16581, new_n16567, new_n16582);
nor_5  g14234(new_n16566, new_n16545, new_n16583_1);
nor_5  g14235(new_n16583_1, new_n16580, new_n16584_1);
nor_5  g14236(new_n16584_1, new_n16582, n5020);
or_5   g14237(n13781, n11486, new_n16586);
or_5   g14238(new_n16586, n16722, new_n16587);
nor_5  g14239(new_n16587, n3480, new_n16588);
xnor_4 g14240(new_n16588, n3018, new_n16589_1);
xnor_4 g14241(new_n16589_1, new_n2884, new_n16590);
xor_4  g14242(new_n16587, n3480, new_n16591);
nor_5  g14243(new_n16591, new_n2888, new_n16592);
xnor_4 g14244(new_n16591, new_n2888, new_n16593);
xor_4  g14245(new_n16586, n16722, new_n16594);
nor_5  g14246(new_n16594, new_n2892, new_n16595);
xnor_4 g14247(new_n16594, new_n2892, new_n16596_1);
xor_4  g14248(n13781, n11486, new_n16597);
nor_5  g14249(new_n16597, new_n2896, new_n16598);
or_5   g14250(new_n2899, n13781, new_n16599);
xnor_4 g14251(new_n16597, new_n2896, new_n16600);
nor_5  g14252(new_n16600, new_n16599, new_n16601);
nor_5  g14253(new_n16601, new_n16598, new_n16602);
nor_5  g14254(new_n16602, new_n16596_1, new_n16603);
nor_5  g14255(new_n16603, new_n16595, new_n16604);
nor_5  g14256(new_n16604, new_n16593, new_n16605);
or_5   g14257(new_n16605, new_n16592, new_n16606);
xor_4  g14258(new_n16606, new_n16590, new_n16607);
xor_4  g14259(new_n16607, new_n6273, new_n16608_1);
xor_4  g14260(new_n16604, new_n16593, new_n16609);
and_5  g14261(new_n16609, new_n6277, new_n16610);
xnor_4 g14262(new_n16609, new_n6277, new_n16611);
xor_4  g14263(new_n16602, new_n16596_1, new_n16612);
and_5  g14264(new_n16612, new_n14614, new_n16613);
xor_4  g14265(new_n16600, new_n16599, new_n16614);
and_5  g14266(new_n16614, new_n6286, new_n16615);
xor_4  g14267(new_n2899, n13781, new_n16616);
or_5   g14268(new_n16616, new_n6289, new_n16617_1);
xor_4  g14269(new_n16614, new_n6286, new_n16618);
and_5  g14270(new_n16618, new_n16617_1, new_n16619);
nor_5  g14271(new_n16619, new_n16615, new_n16620);
xor_4  g14272(new_n16612, new_n6282, new_n16621);
nor_5  g14273(new_n16621, new_n16620, new_n16622);
nor_5  g14274(new_n16622, new_n16613, new_n16623);
nor_5  g14275(new_n16623, new_n16611, new_n16624);
nor_5  g14276(new_n16624, new_n16610, new_n16625);
xnor_4 g14277(new_n16625, new_n16608_1, n5024);
xnor_4 g14278(new_n3508, new_n3479, n5046);
xor_4  g14279(new_n5377, new_n3570_1, n5062);
xnor_4 g14280(new_n11335, new_n11308, n5064);
xor_4  g14281(n12495, n11479, new_n16630_1);
xnor_4 g14282(new_n16630_1, new_n2380, new_n16631);
xnor_4 g14283(n9251, n7428, new_n16632);
or_5   g14284(new_n16632, new_n16631, new_n16633);
or_5   g14285(new_n2366, n7428, new_n16634);
xor_4  g14286(n20138, n10372, new_n16635);
xor_4  g14287(new_n16635, new_n16634, new_n16636);
xnor_4 g14288(new_n16636, new_n16633, new_n16637);
nor_5  g14289(new_n16630_1, new_n2461, new_n16638);
and_5  g14290(n12495, n11479, new_n16639);
xnor_4 g14291(n20235, n8259, new_n16640_1);
xor_4  g14292(new_n16640_1, new_n16639, new_n16641);
xnor_4 g14293(new_n16641, new_n2383, new_n16642);
xor_4  g14294(new_n16642, new_n16638, new_n16643);
xnor_4 g14295(new_n16643, new_n16637, n5082);
xor_4  g14296(new_n12387, new_n12386, n5120);
xnor_4 g14297(new_n13477_1, new_n13468, n5158);
xnor_4 g14298(new_n14721, new_n14708, n5168);
xnor_4 g14299(new_n15721, n6659, new_n16648);
nand_5 g14300(new_n12928, new_n14484, new_n16649);
xor_4  g14301(new_n12928, n23250, new_n16650);
nand_5 g14302(new_n12930, new_n14412_1, new_n16651);
xor_4  g14303(new_n12930, n11455, new_n16652);
nand_5 g14304(new_n12932, new_n14415, new_n16653);
xor_4  g14305(new_n12932, n3945, new_n16654);
and_5  g14306(new_n12936, n5255, new_n16655);
xnor_4 g14307(new_n12936, n5255, new_n16656_1);
and_5  g14308(new_n12939, n21649, new_n16657);
nor_5  g14309(new_n13859, new_n13845, new_n16658);
nor_5  g14310(new_n16658, new_n16657, new_n16659);
nor_5  g14311(new_n16659, new_n16656_1, new_n16660);
nor_5  g14312(new_n16660, new_n16655, new_n16661);
not_10 g14313(new_n16661, new_n16662);
or_5   g14314(new_n16662, new_n16654, new_n16663);
and_5  g14315(new_n16663, new_n16653, new_n16664);
or_5   g14316(new_n16664, new_n16652, new_n16665);
and_5  g14317(new_n16665, new_n16651, new_n16666);
or_5   g14318(new_n16666, new_n16650, new_n16667);
and_5  g14319(new_n16667, new_n16649, new_n16668);
xor_4  g14320(new_n16668, new_n16648, new_n16669);
xnor_4 g14321(new_n16669, new_n14410, new_n16670);
xor_4  g14322(new_n16666, new_n16650, new_n16671);
and_5  g14323(new_n16671, new_n14492, new_n16672);
xnor_4 g14324(new_n16671, new_n14492, new_n16673);
xor_4  g14325(new_n16664, new_n16652, new_n16674_1);
and_5  g14326(new_n16674_1, new_n14496, new_n16675);
xnor_4 g14327(new_n16674_1, new_n14496, new_n16676);
xnor_4 g14328(new_n16661, new_n16654, new_n16677);
and_5  g14329(new_n16677, new_n14500, new_n16678);
xnor_4 g14330(new_n16677, new_n14500, new_n16679);
xor_4  g14331(new_n16659, new_n16656_1, new_n16680);
nor_5  g14332(new_n16680, new_n14506, new_n16681);
xnor_4 g14333(new_n16680, new_n14506, new_n16682_1);
not_10 g14334(new_n13844, new_n16683);
nor_5  g14335(new_n13860, new_n16683, new_n16684_1);
nor_5  g14336(new_n13879, new_n13861, new_n16685);
nor_5  g14337(new_n16685, new_n16684_1, new_n16686);
nor_5  g14338(new_n16686, new_n16682_1, new_n16687);
nor_5  g14339(new_n16687, new_n16681, new_n16688_1);
nor_5  g14340(new_n16688_1, new_n16679, new_n16689);
nor_5  g14341(new_n16689, new_n16678, new_n16690);
nor_5  g14342(new_n16690, new_n16676, new_n16691);
nor_5  g14343(new_n16691, new_n16675, new_n16692);
nor_5  g14344(new_n16692, new_n16673, new_n16693);
nor_5  g14345(new_n16693, new_n16672, new_n16694);
xnor_4 g14346(new_n16694, new_n16670, n5184);
not_10 g14347(new_n4106, new_n16696);
nand_5 g14348(new_n4199, new_n16696, new_n16697);
nor_5  g14349(new_n4266_1, new_n16697, new_n16698);
nor_5  g14350(new_n4199, new_n16696, new_n16699);
and_5  g14351(new_n4266_1, new_n16699, new_n16700);
or_5   g14352(new_n16700, new_n16698, n5228);
not_10 g14353(n1314, new_n16702);
nor_5  g14354(n25494, new_n16702, new_n16703);
nor_5  g14355(new_n10193, new_n10174, new_n16704);
nor_5  g14356(new_n16704, new_n16703, new_n16705);
xnor_4 g14357(new_n16705, new_n6519, new_n16706);
not_10 g14358(new_n6446, new_n16707);
nor_5  g14359(new_n10194, new_n16707, new_n16708);
xnor_4 g14360(new_n10194, new_n16707, new_n16709);
nor_5  g14361(new_n10212, new_n11304, new_n16710);
nor_5  g14362(new_n11337, new_n11305, new_n16711);
nor_5  g14363(new_n16711, new_n16710, new_n16712);
nor_5  g14364(new_n16712, new_n16709, new_n16713);
nor_5  g14365(new_n16713, new_n16708, new_n16714);
xnor_4 g14366(new_n16714, new_n16706, n5256);
xor_4  g14367(new_n6051, new_n6041, n5265);
xnor_4 g14368(new_n15516, new_n15476, n5273);
xnor_4 g14369(new_n6636, new_n6601, new_n16718);
xor_4  g14370(n20946, n2289, new_n16719);
nor_5  g14371(new_n3056, n1112, new_n16720);
xor_4  g14372(n7751, n1112, new_n16721);
nor_5  g14373(new_n3057, n20179, new_n16722_1);
nor_5  g14374(new_n15196, new_n15181, new_n16723);
nor_5  g14375(new_n16723, new_n16722_1, new_n16724);
nor_5  g14376(new_n16724, new_n16721, new_n16725);
nor_5  g14377(new_n16725, new_n16720, new_n16726);
xor_4  g14378(new_n16726, new_n16719, new_n16727);
xnor_4 g14379(new_n16727, new_n16718, new_n16728);
xnor_4 g14380(new_n6634_1, new_n6604, new_n16729);
xor_4  g14381(new_n16724, new_n16721, new_n16730);
nor_5  g14382(new_n16730, new_n16729, new_n16731);
xnor_4 g14383(new_n16730, new_n16729, new_n16732);
nor_5  g14384(new_n15197, new_n15180_1, new_n16733_1);
nor_5  g14385(new_n15218, new_n15198, new_n16734);
nor_5  g14386(new_n16734, new_n16733_1, new_n16735);
nor_5  g14387(new_n16735, new_n16732, new_n16736);
nor_5  g14388(new_n16736, new_n16731, new_n16737);
xnor_4 g14389(new_n16737, new_n16728, n5274);
or_5   g14390(n25316, n20385, new_n16739);
or_5   g14391(new_n16739, n919, new_n16740);
or_5   g14392(new_n16740, n3918, new_n16741);
xor_4  g14393(new_n16741, n6513, new_n16742);
xnor_4 g14394(new_n16742, new_n8013, new_n16743_1);
xor_4  g14395(new_n16740, n3918, new_n16744);
nor_5  g14396(new_n16744, new_n8015, new_n16745);
xor_4  g14397(new_n16739, n919, new_n16746);
nor_5  g14398(new_n16746, new_n10071, new_n16747);
xor_4  g14399(new_n16746, new_n8021, new_n16748);
xor_4  g14400(n25316, n20385, new_n16749);
and_5  g14401(new_n16749, new_n10063, new_n16750);
nor_5  g14402(new_n8028, new_n11112, new_n16751);
xnor_4 g14403(new_n16749, new_n8026, new_n16752);
and_5  g14404(new_n16752, new_n16751, new_n16753);
or_5   g14405(new_n16753, new_n16750, new_n16754);
nor_5  g14406(new_n16754, new_n16748, new_n16755);
nor_5  g14407(new_n16755, new_n16747, new_n16756);
xnor_4 g14408(new_n16744, new_n8015, new_n16757);
nor_5  g14409(new_n16757, new_n16756, new_n16758);
nor_5  g14410(new_n16758, new_n16745, new_n16759);
xnor_4 g14411(new_n16759, new_n16743_1, new_n16760);
xnor_4 g14412(new_n14971, new_n7872, new_n16761);
nor_5  g14413(new_n14974, new_n7875, new_n16762);
xnor_4 g14414(new_n14974, new_n7875, new_n16763);
and_5  g14415(new_n3858, n24786, new_n16764);
xnor_4 g14416(new_n3858, n24786, new_n16765);
and_5  g14417(new_n3862, n27120, new_n16766);
nor_5  g14418(new_n3866, n23065, new_n16767);
xnor_4 g14419(new_n3862, n27120, new_n16768);
nor_5  g14420(new_n16768, new_n16767, new_n16769);
nor_5  g14421(new_n16769, new_n16766, new_n16770);
nor_5  g14422(new_n16770, new_n16765, new_n16771);
nor_5  g14423(new_n16771, new_n16764, new_n16772);
nor_5  g14424(new_n16772, new_n16763, new_n16773);
nor_5  g14425(new_n16773, new_n16762, new_n16774);
xor_4  g14426(new_n16774, new_n16761, new_n16775);
xnor_4 g14427(new_n16775, new_n16760, new_n16776);
xnor_4 g14428(new_n16772, new_n16763, new_n16777);
xor_4  g14429(new_n16757, new_n16756, new_n16778);
and_5  g14430(new_n16778, new_n16777, new_n16779);
xnor_4 g14431(new_n16778, new_n16777, new_n16780);
xnor_4 g14432(new_n16770, new_n16765, new_n16781);
xor_4  g14433(new_n16754, new_n16748, new_n16782);
and_5  g14434(new_n16782, new_n16781, new_n16783);
xnor_4 g14435(new_n16782, new_n16781, new_n16784);
xor_4  g14436(new_n16752, new_n16751, new_n16785);
xor_4  g14437(new_n16768, new_n16767, new_n16786);
nor_5  g14438(new_n16786, new_n16785, new_n16787);
xnor_4 g14439(new_n3866, n23065, new_n16788);
nand_5 g14440(new_n16788, new_n8104, new_n16789);
xor_4  g14441(new_n16786, new_n16785, new_n16790);
and_5  g14442(new_n16790, new_n16789, new_n16791);
nor_5  g14443(new_n16791, new_n16787, new_n16792);
nor_5  g14444(new_n16792, new_n16784, new_n16793);
nor_5  g14445(new_n16793, new_n16783, new_n16794);
nor_5  g14446(new_n16794, new_n16780, new_n16795);
nor_5  g14447(new_n16795, new_n16779, new_n16796);
xnor_4 g14448(new_n16796, new_n16776, n5300);
and_5  g14449(new_n6514_1, new_n6511, new_n16798_1);
and_5  g14450(new_n6518, new_n6515, new_n16799);
nor_5  g14451(new_n16799, new_n16798_1, new_n16800);
nor_5  g14452(new_n16800, new_n16705, new_n16801);
xnor_4 g14453(new_n16800, new_n16705, new_n16802);
nor_5  g14454(new_n16705, new_n6519, new_n16803);
nor_5  g14455(new_n16714, new_n16706, new_n16804);
or_5   g14456(new_n16804, new_n16803, new_n16805);
nor_5  g14457(new_n16805, new_n16802, new_n16806);
nor_5  g14458(new_n16806, new_n16801, n5325);
xnor_4 g14459(n25120, n17458, new_n16808);
nor_5  g14460(n8363, n1222, new_n16809);
xnor_4 g14461(n8363, n1222, new_n16810);
nor_5  g14462(n25240, n14680, new_n16811);
xnor_4 g14463(n25240, n14680, new_n16812_1);
nor_5  g14464(n17250, n10125, new_n16813);
xnor_4 g14465(n17250, n10125, new_n16814);
and_5  g14466(n23160, n8067, new_n16815);
or_5   g14467(n23160, n8067, new_n16816);
nor_5  g14468(n20923, n16524, new_n16817);
nor_5  g14469(new_n11706, new_n11703, new_n16818_1);
nor_5  g14470(new_n16818_1, new_n16817, new_n16819);
and_5  g14471(new_n16819, new_n16816, new_n16820);
or_5   g14472(new_n16820, new_n16815, new_n16821);
nor_5  g14473(new_n16821, new_n16814, new_n16822);
nor_5  g14474(new_n16822, new_n16813, new_n16823);
nor_5  g14475(new_n16823, new_n16812_1, new_n16824_1);
nor_5  g14476(new_n16824_1, new_n16811, new_n16825);
nor_5  g14477(new_n16825, new_n16810, new_n16826);
nor_5  g14478(new_n16826, new_n16809, new_n16827);
xnor_4 g14479(new_n16827, new_n16808, new_n16828);
nor_5  g14480(new_n16828, n23272, new_n16829);
xnor_4 g14481(new_n16828, n23272, new_n16830);
xnor_4 g14482(new_n16825, new_n16810, new_n16831);
nor_5  g14483(new_n16831, n11481, new_n16832);
xnor_4 g14484(new_n16831, n11481, new_n16833);
xnor_4 g14485(new_n16823, new_n16812_1, new_n16834_1);
nor_5  g14486(new_n16834_1, n16439, new_n16835);
xnor_4 g14487(new_n16834_1, n16439, new_n16836);
xnor_4 g14488(new_n16821, new_n16814, new_n16837_1);
nor_5  g14489(new_n16837_1, n15241, new_n16838);
xnor_4 g14490(new_n16837_1, n15241, new_n16839);
xnor_4 g14491(n23160, n8067, new_n16840);
xnor_4 g14492(new_n16840, new_n16819, new_n16841_1);
nor_5  g14493(new_n16841_1, n7678, new_n16842);
xnor_4 g14494(new_n16841_1, n7678, new_n16843);
nor_5  g14495(new_n11707, n3785, new_n16844);
nor_5  g14496(new_n11711, new_n11708, new_n16845);
nor_5  g14497(new_n16845, new_n16844, new_n16846);
nor_5  g14498(new_n16846, new_n16843, new_n16847);
nor_5  g14499(new_n16847, new_n16842, new_n16848);
nor_5  g14500(new_n16848, new_n16839, new_n16849);
nor_5  g14501(new_n16849, new_n16838, new_n16850);
nor_5  g14502(new_n16850, new_n16836, new_n16851);
nor_5  g14503(new_n16851, new_n16835, new_n16852);
nor_5  g14504(new_n16852, new_n16833, new_n16853);
nor_5  g14505(new_n16853, new_n16832, new_n16854);
nor_5  g14506(new_n16854, new_n16830, new_n16855);
nor_5  g14507(new_n16855, new_n16829, new_n16856);
nor_5  g14508(n25120, n17458, new_n16857);
nor_5  g14509(new_n16827, new_n16808, new_n16858);
nor_5  g14510(new_n16858, new_n16857, new_n16859);
nand_5 g14511(new_n16859, new_n16856, new_n16860);
xnor_4 g14512(n12702, n12507, new_n16861);
nor_5  g14513(n26797, n15077, new_n16862);
xnor_4 g14514(n26797, n15077, new_n16863);
nor_5  g14515(n23913, n3710, new_n16864);
xnor_4 g14516(n23913, n3710, new_n16865);
nor_5  g14517(n26318, n22554, new_n16866);
xnor_4 g14518(n26318, n22554, new_n16867);
nor_5  g14519(n26054, n20429, new_n16868);
xnor_4 g14520(n26054, n20429, new_n16869);
nor_5  g14521(n19081, n3909, new_n16870);
xnor_4 g14522(n19081, n3909, new_n16871);
nor_5  g14523(n23974, n8309, new_n16872);
xnor_4 g14524(n23974, n8309, new_n16873);
and_5  g14525(n19144, n2146, new_n16874);
or_5   g14526(n19144, n2146, new_n16875);
nor_5  g14527(n22173, n12593, new_n16876);
nor_5  g14528(new_n15174, new_n15173, new_n16877);
nor_5  g14529(new_n16877, new_n16876, new_n16878);
and_5  g14530(new_n16878, new_n16875, new_n16879);
or_5   g14531(new_n16879, new_n16874, new_n16880);
nor_5  g14532(new_n16880, new_n16873, new_n16881);
nor_5  g14533(new_n16881, new_n16872, new_n16882);
nor_5  g14534(new_n16882, new_n16871, new_n16883);
nor_5  g14535(new_n16883, new_n16870, new_n16884);
nor_5  g14536(new_n16884, new_n16869, new_n16885_1);
nor_5  g14537(new_n16885_1, new_n16868, new_n16886);
nor_5  g14538(new_n16886, new_n16867, new_n16887);
nor_5  g14539(new_n16887, new_n16866, new_n16888);
nor_5  g14540(new_n16888, new_n16865, new_n16889);
nor_5  g14541(new_n16889, new_n16864, new_n16890);
nor_5  g14542(new_n16890, new_n16863, new_n16891);
nor_5  g14543(new_n16891, new_n16862, new_n16892);
xnor_4 g14544(new_n16892, new_n16861, new_n16893);
nor_5  g14545(new_n16893, n12650, new_n16894);
xnor_4 g14546(new_n16893, n12650, new_n16895);
xnor_4 g14547(new_n16890, new_n16863, new_n16896);
nor_5  g14548(new_n16896, n10201, new_n16897);
xnor_4 g14549(new_n16896, n10201, new_n16898);
xnor_4 g14550(new_n16888, new_n16865, new_n16899);
nor_5  g14551(new_n16899, n10593, new_n16900);
xnor_4 g14552(new_n16899, n10593, new_n16901);
xnor_4 g14553(new_n16886, new_n16867, new_n16902);
nor_5  g14554(new_n16902, n18290, new_n16903);
xnor_4 g14555(new_n16884, new_n16869, new_n16904);
nor_5  g14556(new_n16904, n11580, new_n16905_1);
xnor_4 g14557(new_n16904, n11580, new_n16906);
xnor_4 g14558(new_n16882, new_n16871, new_n16907);
nor_5  g14559(new_n16907, n15884, new_n16908);
xnor_4 g14560(new_n16907, n15884, new_n16909);
xnor_4 g14561(new_n16880, new_n16873, new_n16910);
or_5   g14562(new_n16910, n6356, new_n16911_1);
xnor_4 g14563(n19144, n2146, new_n16912);
xnor_4 g14564(new_n16912, new_n16878, new_n16913);
and_5  g14565(new_n16913, n27104, new_n16914);
xnor_4 g14566(new_n16913, n27104, new_n16915);
nor_5  g14567(new_n15175, n27188, new_n16916);
nor_5  g14568(new_n15176_1, new_n15172, new_n16917);
or_5   g14569(new_n16917, new_n16916, new_n16918);
nor_5  g14570(new_n16918, new_n16915, new_n16919);
nor_5  g14571(new_n16919, new_n16914, new_n16920);
not_10 g14572(new_n16920, new_n16921);
xnor_4 g14573(new_n16910, n6356, new_n16922);
or_5   g14574(new_n16922, new_n16921, new_n16923);
and_5  g14575(new_n16923, new_n16911_1, new_n16924);
nor_5  g14576(new_n16924, new_n16909, new_n16925);
nor_5  g14577(new_n16925, new_n16908, new_n16926);
nor_5  g14578(new_n16926, new_n16906, new_n16927);
nor_5  g14579(new_n16927, new_n16905_1, new_n16928);
xnor_4 g14580(new_n16902, n18290, new_n16929);
nor_5  g14581(new_n16929, new_n16928, new_n16930);
nor_5  g14582(new_n16930, new_n16903, new_n16931);
nor_5  g14583(new_n16931, new_n16901, new_n16932);
nor_5  g14584(new_n16932, new_n16900, new_n16933);
nor_5  g14585(new_n16933, new_n16898, new_n16934);
nor_5  g14586(new_n16934, new_n16897, new_n16935);
nor_5  g14587(new_n16935, new_n16895, new_n16936);
or_5   g14588(new_n16936, new_n16894, new_n16937);
nor_5  g14589(n12702, n12507, new_n16938);
nor_5  g14590(new_n16892, new_n16861, new_n16939);
or_5   g14591(new_n16939, new_n16938, new_n16940);
nor_5  g14592(new_n16940, new_n16937, new_n16941);
xnor_4 g14593(new_n16941, new_n16860, new_n16942);
xor_4  g14594(new_n16859, new_n16856, new_n16943);
not_10 g14595(new_n16943, new_n16944);
xor_4  g14596(new_n16940, new_n16937, new_n16945);
nor_5  g14597(new_n16945, new_n16944, new_n16946);
xnor_4 g14598(new_n16945, new_n16944, new_n16947);
xnor_4 g14599(new_n16854, new_n16830, new_n16948);
xor_4  g14600(new_n16935, new_n16895, new_n16949);
and_5  g14601(new_n16949, new_n16948, new_n16950);
xnor_4 g14602(new_n16949, new_n16948, new_n16951_1);
xor_4  g14603(new_n16852, new_n16833, new_n16952);
not_10 g14604(new_n16952, new_n16953);
xor_4  g14605(new_n16933, new_n16898, new_n16954_1);
and_5  g14606(new_n16954_1, new_n16953, new_n16955);
xnor_4 g14607(new_n16954_1, new_n16953, new_n16956);
xnor_4 g14608(new_n16850, new_n16836, new_n16957);
xor_4  g14609(new_n16931, new_n16901, new_n16958);
and_5  g14610(new_n16958, new_n16957, new_n16959);
xnor_4 g14611(new_n16958, new_n16957, new_n16960);
xnor_4 g14612(new_n16848, new_n16839, new_n16961);
xor_4  g14613(new_n16929, new_n16928, new_n16962);
and_5  g14614(new_n16962, new_n16961, new_n16963);
xnor_4 g14615(new_n16962, new_n16961, new_n16964);
xnor_4 g14616(new_n16926, new_n16906, new_n16965);
xor_4  g14617(new_n16846, new_n16843, new_n16966);
nor_5  g14618(new_n16966, new_n16965, new_n16967);
xnor_4 g14619(new_n16966, new_n16965, new_n16968_1);
xor_4  g14620(new_n16924, new_n16909, new_n16969);
and_5  g14621(new_n16969, new_n11712_1, new_n16970);
xnor_4 g14622(new_n16969, new_n11712_1, new_n16971_1);
xnor_4 g14623(new_n16922, new_n16920, new_n16972);
and_5  g14624(new_n16972, new_n11714, new_n16973);
xor_4  g14625(new_n16918, new_n16915, new_n16974);
nor_5  g14626(new_n16974, new_n6039, new_n16975);
xor_4  g14627(new_n16974, new_n6039, new_n16976);
nor_5  g14628(new_n15177, new_n15171, new_n16977);
nor_5  g14629(new_n15178, new_n6043, new_n16978);
nor_5  g14630(new_n16978, new_n16977, new_n16979);
and_5  g14631(new_n16979, new_n16976, new_n16980);
nor_5  g14632(new_n16980, new_n16975, new_n16981);
xnor_4 g14633(new_n16972, new_n11714, new_n16982);
nor_5  g14634(new_n16982, new_n16981, new_n16983);
nor_5  g14635(new_n16983, new_n16973, new_n16984);
nor_5  g14636(new_n16984, new_n16971_1, new_n16985);
nor_5  g14637(new_n16985, new_n16970, new_n16986);
nor_5  g14638(new_n16986, new_n16968_1, new_n16987);
nor_5  g14639(new_n16987, new_n16967, new_n16988_1);
nor_5  g14640(new_n16988_1, new_n16964, new_n16989_1);
nor_5  g14641(new_n16989_1, new_n16963, new_n16990);
nor_5  g14642(new_n16990, new_n16960, new_n16991);
nor_5  g14643(new_n16991, new_n16959, new_n16992);
nor_5  g14644(new_n16992, new_n16956, new_n16993);
nor_5  g14645(new_n16993, new_n16955, new_n16994_1);
nor_5  g14646(new_n16994_1, new_n16951_1, new_n16995);
nor_5  g14647(new_n16995, new_n16950, new_n16996);
nor_5  g14648(new_n16996, new_n16947, new_n16997);
nor_5  g14649(new_n16997, new_n16946, new_n16998);
xnor_4 g14650(new_n16998, new_n16942, n5351);
nor_5  g14651(new_n14879, new_n14873, n5353);
nor_5  g14652(new_n10657, n2160, new_n17001);
nor_5  g14653(new_n10700, new_n10658, new_n17002);
nor_5  g14654(new_n17002, new_n17001, new_n17003);
nor_5  g14655(n9934, n2272, new_n17004);
nor_5  g14656(new_n10656, new_n10623, new_n17005);
or_5   g14657(new_n17005, new_n17004, new_n17006_1);
and_5  g14658(new_n17006_1, new_n17003, new_n17007);
nor_5  g14659(new_n10704, n21784, new_n17008);
or_5   g14660(new_n17008, new_n6588, new_n17009);
nor_5  g14661(new_n10705, new_n6591, new_n17010);
nor_5  g14662(new_n10719, new_n10706, new_n17011);
nor_5  g14663(new_n17011, new_n17010, new_n17012);
nor_5  g14664(new_n17012, new_n17009, new_n17013);
xnor_4 g14665(new_n17013, new_n17007, new_n17014);
xor_4  g14666(new_n17006_1, new_n17003, new_n17015);
xnor_4 g14667(new_n17008, new_n6588, new_n17016);
xnor_4 g14668(new_n17016, new_n17012, new_n17017);
and_5  g14669(new_n17017, new_n17015, new_n17018);
xnor_4 g14670(new_n17017, new_n17015, new_n17019);
and_5  g14671(new_n10720, new_n10701_1, new_n17020);
nor_5  g14672(new_n10765, new_n10721, new_n17021);
nor_5  g14673(new_n17021, new_n17020, new_n17022);
nor_5  g14674(new_n17022, new_n17019, new_n17023);
nor_5  g14675(new_n17023, new_n17018, new_n17024);
xnor_4 g14676(new_n17024, new_n17014, n5399);
and_5  g14677(new_n15893, n2979, new_n17026);
nor_5  g14678(new_n15897, new_n15894, new_n17027);
nor_5  g14679(new_n17027, new_n17026, new_n17028);
and_5  g14680(new_n12779, n9934, new_n17029);
or_5   g14681(new_n12779, n9934, new_n17030);
and_5  g14682(new_n15892, new_n17030, new_n17031);
or_5   g14683(new_n17031, new_n12821_1, new_n17032);
or_5   g14684(new_n17032, new_n17029, new_n17033);
nor_5  g14685(new_n17033, new_n17028, new_n17034);
xnor_4 g14686(new_n17034, new_n17013, new_n17035_1);
not_10 g14687(new_n17017, new_n17036);
xor_4  g14688(new_n17033, new_n17028, new_n17037_1);
nor_5  g14689(new_n17037_1, new_n17036, new_n17038);
not_10 g14690(new_n10720, new_n17039);
nor_5  g14691(new_n15898, new_n17039, new_n17040);
nor_5  g14692(new_n15903, new_n15899, new_n17041);
nor_5  g14693(new_n17041, new_n17040, new_n17042);
xor_4  g14694(new_n17037_1, new_n17017, new_n17043);
nor_5  g14695(new_n17043, new_n17042, new_n17044);
nor_5  g14696(new_n17044, new_n17038, new_n17045);
xnor_4 g14697(new_n17045, new_n17035_1, n5403);
xnor_4 g14698(new_n14144, new_n14115, n5430);
and_5  g14699(new_n13184, new_n13179, new_n17048);
nand_5 g14700(new_n13175, new_n9432, new_n17049);
nor_5  g14701(new_n13175, new_n9432, new_n17050);
or_5   g14702(new_n13185, new_n17050, new_n17051);
nand_5 g14703(new_n17051, new_n17049, new_n17052);
or_5   g14704(new_n17052, new_n9308_1, new_n17053);
nor_5  g14705(new_n17053, new_n17048, n5439);
xnor_4 g14706(new_n11068, new_n11050, n5472);
xnor_4 g14707(new_n7628, new_n7591, n5485);
xnor_4 g14708(new_n16532, new_n16516_1, n5524);
nand_5 g14709(new_n14889, new_n5462, new_n17058);
or_5   g14710(new_n17058, new_n5459, new_n17059);
or_5   g14711(new_n17059, new_n12140, new_n17060);
or_5   g14712(new_n17060, new_n12136, new_n17061);
or_5   g14713(new_n17061, new_n12132, new_n17062);
or_5   g14714(new_n17062, new_n12128, new_n17063);
or_5   g14715(new_n17063, new_n5434, new_n17064);
xnor_4 g14716(new_n17064, new_n5430_1, new_n17065);
nor_5  g14717(new_n17065, new_n12426, new_n17066);
xnor_4 g14718(new_n17065, new_n12426, new_n17067);
xor_4  g14719(new_n17063, new_n5434, new_n17068_1);
nor_5  g14720(new_n17068_1, new_n12429, new_n17069_1);
xnor_4 g14721(new_n17068_1, new_n12429, new_n17070_1);
xnor_4 g14722(new_n17062, new_n5439_1, new_n17071);
nor_5  g14723(new_n17071, new_n12432, new_n17072);
xnor_4 g14724(new_n17071, new_n12432, new_n17073);
xnor_4 g14725(new_n17061, new_n5444, new_n17074);
nor_5  g14726(new_n17074, new_n12435, new_n17075_1);
xnor_4 g14727(new_n17074, new_n12435, new_n17076);
xnor_4 g14728(new_n17060, new_n5448, new_n17077_1);
nor_5  g14729(new_n17077_1, new_n12438, new_n17078);
xnor_4 g14730(new_n17077_1, new_n12438, new_n17079);
xnor_4 g14731(new_n17059, new_n5453, new_n17080);
nor_5  g14732(new_n17080, new_n12441, new_n17081);
xnor_4 g14733(new_n17080, new_n12441, new_n17082);
xnor_4 g14734(new_n17058, new_n5457, new_n17083);
nor_5  g14735(new_n15906, new_n11791, new_n17084_1);
nor_5  g14736(new_n15910, new_n15907, new_n17085);
nor_5  g14737(new_n17085, new_n17084_1, new_n17086);
nor_5  g14738(new_n17086, new_n17083, new_n17087);
xnor_4 g14739(new_n17086, new_n17083, new_n17088);
nor_5  g14740(new_n17088, new_n11789, new_n17089);
nor_5  g14741(new_n17089, new_n17087, new_n17090_1);
nor_5  g14742(new_n17090_1, new_n17082, new_n17091);
nor_5  g14743(new_n17091, new_n17081, new_n17092);
nor_5  g14744(new_n17092, new_n17079, new_n17093);
nor_5  g14745(new_n17093, new_n17078, new_n17094);
nor_5  g14746(new_n17094, new_n17076, new_n17095_1);
nor_5  g14747(new_n17095_1, new_n17075_1, new_n17096);
nor_5  g14748(new_n17096, new_n17073, new_n17097);
nor_5  g14749(new_n17097, new_n17072, new_n17098);
nor_5  g14750(new_n17098, new_n17070_1, new_n17099);
nor_5  g14751(new_n17099, new_n17069_1, new_n17100);
nor_5  g14752(new_n17100, new_n17067, new_n17101);
nor_5  g14753(new_n17101, new_n17066, new_n17102);
or_5   g14754(new_n17064, new_n12121_1, new_n17103);
and_5  g14755(new_n17103, new_n12117, new_n17104_1);
not_10 g14756(new_n12115, new_n17105);
nor_5  g14757(new_n17103, new_n17105, new_n17106_1);
nor_5  g14758(new_n17106_1, new_n17104_1, new_n17107);
xnor_4 g14759(new_n17107, new_n12464, new_n17108);
xnor_4 g14760(new_n17108, new_n17102, new_n17109);
nor_5  g14761(new_n17109, new_n4440, new_n17110);
xnor_4 g14762(new_n17109, new_n4440, new_n17111);
xor_4  g14763(new_n17100, new_n17067, new_n17112);
and_5  g14764(new_n17112, new_n4586, new_n17113);
xnor_4 g14765(new_n17112, new_n4586, new_n17114);
xor_4  g14766(new_n17098, new_n17070_1, new_n17115);
and_5  g14767(new_n17115, new_n4590_1, new_n17116);
xnor_4 g14768(new_n17115, new_n4590_1, new_n17117);
xor_4  g14769(new_n17096, new_n17073, new_n17118);
and_5  g14770(new_n17118, new_n4595_1, new_n17119_1);
xnor_4 g14771(new_n17118, new_n4595_1, new_n17120);
xor_4  g14772(new_n17094, new_n17076, new_n17121);
and_5  g14773(new_n17121, new_n4600, new_n17122);
xnor_4 g14774(new_n17121, new_n4600, new_n17123);
xor_4  g14775(new_n17092, new_n17079, new_n17124);
and_5  g14776(new_n17124, new_n4605, new_n17125);
xnor_4 g14777(new_n17124, new_n4605, new_n17126);
xor_4  g14778(new_n17090_1, new_n17082, new_n17127);
and_5  g14779(new_n17127, new_n4610, new_n17128);
xnor_4 g14780(new_n17127, new_n4610, new_n17129);
xnor_4 g14781(new_n17088, new_n11789, new_n17130_1);
nor_5  g14782(new_n17130_1, new_n4615, new_n17131);
xor_4  g14783(new_n17130_1, new_n4615, new_n17132);
nor_5  g14784(new_n15911, new_n4620, new_n17133);
nor_5  g14785(new_n15914, new_n15912, new_n17134);
nor_5  g14786(new_n17134, new_n17133, new_n17135);
and_5  g14787(new_n17135, new_n17132, new_n17136);
nor_5  g14788(new_n17136, new_n17131, new_n17137);
nor_5  g14789(new_n17137, new_n17129, new_n17138_1);
nor_5  g14790(new_n17138_1, new_n17128, new_n17139);
nor_5  g14791(new_n17139, new_n17126, new_n17140);
nor_5  g14792(new_n17140, new_n17125, new_n17141);
nor_5  g14793(new_n17141, new_n17123, new_n17142);
nor_5  g14794(new_n17142, new_n17122, new_n17143);
nor_5  g14795(new_n17143, new_n17120, new_n17144);
nor_5  g14796(new_n17144, new_n17119_1, new_n17145);
nor_5  g14797(new_n17145, new_n17117, new_n17146);
nor_5  g14798(new_n17146, new_n17116, new_n17147);
nor_5  g14799(new_n17147, new_n17114, new_n17148);
nor_5  g14800(new_n17148, new_n17113, new_n17149);
nor_5  g14801(new_n17149, new_n17111, new_n17150);
nor_5  g14802(new_n17150, new_n17110, new_n17151);
nor_5  g14803(new_n17107, new_n12464, new_n17152);
and_5  g14804(new_n17107, new_n12464, new_n17153);
nor_5  g14805(new_n17153, new_n17102, new_n17154);
nor_5  g14806(new_n17154, new_n17152, new_n17155);
or_5   g14807(new_n17155, new_n17106_1, new_n17156);
xnor_4 g14808(new_n17156, new_n17151, n5564);
xnor_4 g14809(new_n6294, new_n6284, n5593);
xnor_4 g14810(new_n15945, new_n12843_1, new_n17159);
not_10 g14811(new_n14795, new_n17160);
nor_5  g14812(new_n17160, new_n12848, new_n17161);
xor_4  g14813(new_n14795, new_n12848, new_n17162);
not_10 g14814(new_n14797, new_n17163_1);
nor_5  g14815(new_n17163_1, new_n12852, new_n17164);
xor_4  g14816(new_n14797, new_n12852, new_n17165);
not_10 g14817(new_n12856, new_n17166);
and_5  g14818(new_n13895, new_n17166, new_n17167);
xnor_4 g14819(new_n13895, new_n17166, new_n17168_1);
xnor_4 g14820(new_n12756_1, new_n12747, new_n17169);
and_5  g14821(new_n13897, new_n17169, new_n17170);
and_5  g14822(new_n15555_1, new_n15545, new_n17171);
nor_5  g14823(new_n17171, new_n17170, new_n17172);
nor_5  g14824(new_n17172, new_n17168_1, new_n17173);
nor_5  g14825(new_n17173, new_n17167, new_n17174);
nor_5  g14826(new_n17174, new_n17165, new_n17175);
nor_5  g14827(new_n17175, new_n17164, new_n17176);
nor_5  g14828(new_n17176, new_n17162, new_n17177);
nor_5  g14829(new_n17177, new_n17161, new_n17178);
xnor_4 g14830(new_n17178, new_n17159, n5603);
xor_4  g14831(n17911, n14440, new_n17180);
not_10 g14832(n21997, new_n17181);
nor_5  g14833(new_n17181, n1654, new_n17182);
xor_4  g14834(n21997, n1654, new_n17183);
not_10 g14835(n25119, new_n17184);
nor_5  g14836(new_n17184, n13783, new_n17185);
xor_4  g14837(n25119, n13783, new_n17186);
not_10 g14838(n1163, new_n17187);
nor_5  g14839(n26660, new_n17187, new_n17188);
xor_4  g14840(n26660, n1163, new_n17189);
not_10 g14841(n18537, new_n17190);
nor_5  g14842(new_n17190, n3018, new_n17191);
or_5   g14843(n18537, new_n6939, new_n17192);
not_10 g14844(n3480, new_n17193);
nor_5  g14845(n7057, new_n17193, new_n17194);
nor_5  g14846(new_n16214, new_n16205, new_n17195);
nor_5  g14847(new_n17195, new_n17194, new_n17196);
and_5  g14848(new_n17196, new_n17192, new_n17197);
nor_5  g14849(new_n17197, new_n17191, new_n17198);
nor_5  g14850(new_n17198, new_n17189, new_n17199);
nor_5  g14851(new_n17199, new_n17188, new_n17200);
nor_5  g14852(new_n17200, new_n17186, new_n17201);
nor_5  g14853(new_n17201, new_n17185, new_n17202_1);
nor_5  g14854(new_n17202_1, new_n17183, new_n17203);
nor_5  g14855(new_n17203, new_n17182, new_n17204);
xor_4  g14856(new_n17204, new_n17180, new_n17205);
xnor_4 g14857(new_n17205, new_n2916, new_n17206);
xor_4  g14858(new_n17202_1, new_n17183, new_n17207);
nor_5  g14859(new_n17207, new_n2919, new_n17208);
xnor_4 g14860(new_n17207, new_n2919, new_n17209);
not_10 g14861(new_n2923, new_n17210);
xor_4  g14862(new_n17200, new_n17186, new_n17211);
nor_5  g14863(new_n17211, new_n17210, new_n17212);
xnor_4 g14864(new_n17211, new_n17210, new_n17213);
not_10 g14865(new_n2927, new_n17214);
xor_4  g14866(new_n17198, new_n17189, new_n17215);
nor_5  g14867(new_n17215, new_n17214, new_n17216);
xnor_4 g14868(new_n17215, new_n2927, new_n17217);
not_10 g14869(new_n2931, new_n17218);
xor_4  g14870(n18537, n3018, new_n17219_1);
xnor_4 g14871(new_n17219_1, new_n17196, new_n17220);
and_5  g14872(new_n17220, new_n17218, new_n17221);
nor_5  g14873(new_n16215_1, new_n2934, new_n17222);
nor_5  g14874(new_n16230_1, new_n16216, new_n17223);
nor_5  g14875(new_n17223, new_n17222, new_n17224);
xnor_4 g14876(new_n17220, new_n17218, new_n17225);
nor_5  g14877(new_n17225, new_n17224, new_n17226);
nor_5  g14878(new_n17226, new_n17221, new_n17227);
and_5  g14879(new_n17227, new_n17217, new_n17228);
nor_5  g14880(new_n17228, new_n17216, new_n17229);
nor_5  g14881(new_n17229, new_n17213, new_n17230);
nor_5  g14882(new_n17230, new_n17212, new_n17231);
nor_5  g14883(new_n17231, new_n17209, new_n17232_1);
or_5   g14884(new_n17232_1, new_n17208, new_n17233);
xor_4  g14885(new_n17233, new_n17206, n5609);
xnor_4 g14886(new_n12066, new_n12049, n5634);
xor_4  g14887(new_n6642, new_n6589, new_n17236_1);
nor_5  g14888(new_n3073, n2978, new_n17237);
xor_4  g14889(n3425, n2978, new_n17238);
nor_5  g14890(n23697, new_n3054, new_n17239);
xor_4  g14891(n23697, n9967, new_n17240);
nor_5  g14892(new_n3055, n2289, new_n17241);
nor_5  g14893(new_n16726, new_n16719, new_n17242);
nor_5  g14894(new_n17242, new_n17241, new_n17243_1);
nor_5  g14895(new_n17243_1, new_n17240, new_n17244);
nor_5  g14896(new_n17244, new_n17239, new_n17245);
nor_5  g14897(new_n17245, new_n17238, new_n17246);
nor_5  g14898(new_n17246, new_n17237, new_n17247);
nor_5  g14899(new_n17247, new_n17236_1, new_n17248);
not_10 g14900(new_n17247, new_n17249);
or_5   g14901(new_n17249, new_n6643, new_n17250_1);
xor_4  g14902(new_n17245, new_n17238, new_n17251_1);
nor_5  g14903(new_n17251_1, new_n6685, new_n17252);
xnor_4 g14904(new_n17251_1, new_n6685, new_n17253);
xnor_4 g14905(new_n6638, new_n6597, new_n17254);
xor_4  g14906(new_n17243_1, new_n17240, new_n17255);
nor_5  g14907(new_n17255, new_n17254, new_n17256);
xnor_4 g14908(new_n17255, new_n17254, new_n17257);
nor_5  g14909(new_n16727, new_n16718, new_n17258);
nor_5  g14910(new_n16737, new_n16728, new_n17259);
nor_5  g14911(new_n17259, new_n17258, new_n17260);
nor_5  g14912(new_n17260, new_n17257, new_n17261);
nor_5  g14913(new_n17261, new_n17256, new_n17262);
nor_5  g14914(new_n17262, new_n17253, new_n17263_1);
or_5   g14915(new_n17263_1, new_n17252, new_n17264);
and_5  g14916(new_n17264, new_n17250_1, new_n17265);
nor_5  g14917(new_n17265, new_n17248, new_n17266);
and_5  g14918(new_n6588, new_n6573, new_n17267);
or_5   g14919(new_n6641, new_n6592, new_n17268);
nor_5  g14920(new_n17268, new_n6589, new_n17269);
nor_5  g14921(new_n17269, new_n17267, new_n17270);
xnor_4 g14922(new_n17270, new_n17249, new_n17271);
xnor_4 g14923(new_n17271, new_n17266, n5643);
xor_4  g14924(n18035, n5834, new_n17273);
not_10 g14925(n5077, new_n17274);
nor_5  g14926(n13851, new_n17274, new_n17275);
nor_5  g14927(new_n13972, new_n13953, new_n17276);
nor_5  g14928(new_n17276, new_n17275, new_n17277);
xor_4  g14929(new_n17277, new_n17273, new_n17278);
xnor_4 g14930(new_n17278, new_n13538, new_n17279);
nor_5  g14931(new_n13973, new_n13562, new_n17280);
xnor_4 g14932(new_n13973, new_n13562, new_n17281);
xnor_4 g14933(new_n13533, new_n13519, new_n17282);
nor_5  g14934(new_n13975, new_n17282, new_n17283);
xnor_4 g14935(new_n13975, new_n17282, new_n17284);
xor_4  g14936(new_n13570, new_n13522, new_n17285_1);
nor_5  g14937(new_n13978, new_n17285_1, new_n17286);
xnor_4 g14938(new_n13978, new_n17285_1, new_n17287);
nor_5  g14939(new_n13981, new_n13573, new_n17288);
nor_5  g14940(new_n12525, new_n12290, new_n17289);
xnor_4 g14941(new_n12525, new_n12290, new_n17290);
nor_5  g14942(new_n12538, new_n12294, new_n17291);
xnor_4 g14943(new_n12538, new_n12294, new_n17292);
nor_5  g14944(new_n12545_1, new_n12296, new_n17293);
nor_5  g14945(new_n17293, new_n12301, new_n17294);
xnor_4 g14946(new_n17293, new_n12300, new_n17295);
and_5  g14947(new_n17295, new_n12550, new_n17296);
nor_5  g14948(new_n17296, new_n17294, new_n17297);
nor_5  g14949(new_n17297, new_n17292, new_n17298);
nor_5  g14950(new_n17298, new_n17291, new_n17299);
nor_5  g14951(new_n17299, new_n17290, new_n17300);
or_5   g14952(new_n17300, new_n17289, new_n17301);
xor_4  g14953(new_n13981, new_n13573, new_n17302_1);
and_5  g14954(new_n17302_1, new_n17301, new_n17303);
nor_5  g14955(new_n17303, new_n17288, new_n17304);
nor_5  g14956(new_n17304, new_n17287, new_n17305);
nor_5  g14957(new_n17305, new_n17286, new_n17306);
nor_5  g14958(new_n17306, new_n17284, new_n17307);
nor_5  g14959(new_n17307, new_n17283, new_n17308);
nor_5  g14960(new_n17308, new_n17281, new_n17309);
or_5   g14961(new_n17309, new_n17280, new_n17310);
xor_4  g14962(new_n17310, new_n17279, n5680);
xnor_4 g14963(new_n13269, new_n13268, n5687);
xnor_4 g14964(new_n14264, new_n14257, n5700);
xor_4  g14965(new_n9487, new_n9440, n5732);
xnor_4 g14966(n23775, n8381, new_n17315);
nor_5  g14967(n20235, n8259, new_n17316);
nor_5  g14968(new_n16640_1, new_n16639, new_n17317);
nor_5  g14969(new_n17317, new_n17316, new_n17318);
xor_4  g14970(new_n17318, new_n17315, new_n17319);
xnor_4 g14971(new_n17319, new_n2455, new_n17320_1);
nor_5  g14972(new_n16641, new_n2383, new_n17321);
nor_5  g14973(new_n16642, new_n16638, new_n17322);
or_5   g14974(new_n17322, new_n17321, new_n17323);
xor_4  g14975(new_n17323, new_n17320_1, new_n17324);
xor_4  g14976(n8869, n6385, new_n17325);
nor_5  g14977(new_n2362, n10372, new_n17326);
nor_5  g14978(new_n16635, new_n16634, new_n17327);
nor_5  g14979(new_n17327, new_n17326, new_n17328);
xor_4  g14980(new_n17328, new_n17325, new_n17329);
xor_4  g14981(new_n17329, new_n17324, new_n17330);
nor_5  g14982(new_n16636, new_n16633, new_n17331);
not_10 g14983(new_n16643, new_n17332);
nor_5  g14984(new_n17332, new_n16637, new_n17333);
nor_5  g14985(new_n17333, new_n17331, new_n17334);
xnor_4 g14986(new_n17334, new_n17330, n5742);
xnor_4 g14987(new_n12307, new_n12306, n5765);
xnor_4 g14988(new_n11284, new_n11248, n5776);
xnor_4 g14989(new_n2759, new_n2725, n5782);
xnor_4 g14990(n18901, n1163, new_n17339);
nor_5  g14991(n18537, n4376, new_n17340);
xnor_4 g14992(n18537, n4376, new_n17341);
nor_5  g14993(n14570, n7057, new_n17342);
xnor_4 g14994(n14570, n7057, new_n17343);
nor_5  g14995(n23775, n8381, new_n17344_1);
nor_5  g14996(new_n17318, new_n17315, new_n17345);
nor_5  g14997(new_n17345, new_n17344_1, new_n17346);
nor_5  g14998(new_n17346, new_n17343, new_n17347);
nor_5  g14999(new_n17347, new_n17342, new_n17348);
nor_5  g15000(new_n17348, new_n17341, new_n17349);
nor_5  g15001(new_n17349, new_n17340, new_n17350);
xor_4  g15002(new_n17350, new_n17339, new_n17351_1);
xnor_4 g15003(new_n17351_1, new_n2409_1, new_n17352);
xor_4  g15004(new_n17348, new_n17341, new_n17353);
and_5  g15005(new_n17353, new_n2403, new_n17354);
xnor_4 g15006(new_n17346, new_n17343, new_n17355);
and_5  g15007(new_n17319, new_n2455, new_n17356);
nor_5  g15008(new_n17323, new_n17320_1, new_n17357);
nor_5  g15009(new_n17357, new_n17356, new_n17358);
nor_5  g15010(new_n17358, new_n17355, new_n17359_1);
xor_4  g15011(new_n17358, new_n17355, new_n17360);
and_5  g15012(new_n17360, new_n2396, new_n17361);
nor_5  g15013(new_n17361, new_n17359_1, new_n17362);
xor_4  g15014(new_n17353, new_n2402, new_n17363);
nor_5  g15015(new_n17363, new_n17362, new_n17364);
or_5   g15016(new_n17364, new_n17354, new_n17365);
xor_4  g15017(new_n17365, new_n17352, new_n17366);
xor_4  g15018(n23068, n7099, new_n17367);
nor_5  g15019(n19514, new_n13292, new_n17368);
xor_4  g15020(n19514, n12811, new_n17369);
nor_5  g15021(n10053, new_n13295, new_n17370);
xor_4  g15022(n10053, n1118, new_n17371);
nor_5  g15023(n25974, new_n3594, new_n17372);
nor_5  g15024(new_n13299, n8399, new_n17373);
nor_5  g15025(new_n3598, n1630, new_n17374);
or_5   g15026(n9507, new_n13302, new_n17375);
nor_5  g15027(new_n3602, n1451, new_n17376);
and_5  g15028(new_n17376, new_n17375, new_n17377);
nor_5  g15029(new_n17377, new_n17374, new_n17378);
nor_5  g15030(new_n17378, new_n17373, new_n17379);
or_5   g15031(new_n17379, new_n17372, new_n17380);
nor_5  g15032(new_n17380, new_n17371, new_n17381);
nor_5  g15033(new_n17381, new_n17370, new_n17382);
nor_5  g15034(new_n17382, new_n17369, new_n17383);
nor_5  g15035(new_n17383, new_n17368, new_n17384);
xor_4  g15036(new_n17384, new_n17367, new_n17385);
xor_4  g15037(new_n17385, new_n17366, new_n17386);
xnor_4 g15038(new_n17382, new_n17369, new_n17387_1);
xor_4  g15039(new_n17363, new_n17362, new_n17388);
nor_5  g15040(new_n17388, new_n17387_1, new_n17389);
xnor_4 g15041(new_n17360, new_n2395, new_n17390);
not_10 g15042(new_n17390, new_n17391_1);
xor_4  g15043(new_n17380, new_n17371, new_n17392_1);
nor_5  g15044(new_n17392_1, new_n17391_1, new_n17393);
xor_4  g15045(new_n17392_1, new_n17390, new_n17394);
xnor_4 g15046(n25974, n8399, new_n17395);
xnor_4 g15047(new_n17395, new_n17378, new_n17396);
and_5  g15048(new_n17396, new_n17324, new_n17397);
xnor_4 g15049(new_n17396, new_n17324, new_n17398);
xnor_4 g15050(n26979, n1451, new_n17399);
or_5   g15051(new_n17399, new_n16631, new_n17400);
xor_4  g15052(n9507, n1630, new_n17401);
xnor_4 g15053(new_n17401, new_n17376, new_n17402);
and_5  g15054(new_n17402, new_n17400, new_n17403);
xor_4  g15055(new_n17402, new_n17400, new_n17404);
and_5  g15056(new_n17404, new_n17332, new_n17405);
nor_5  g15057(new_n17405, new_n17403, new_n17406);
nor_5  g15058(new_n17406, new_n17398, new_n17407);
nor_5  g15059(new_n17407, new_n17397, new_n17408);
nor_5  g15060(new_n17408, new_n17394, new_n17409);
or_5   g15061(new_n17409, new_n17393, new_n17410);
xnor_4 g15062(new_n17388, new_n17387_1, new_n17411);
nor_5  g15063(new_n17411, new_n17410, new_n17412);
nor_5  g15064(new_n17412, new_n17389, new_n17413);
xnor_4 g15065(new_n17413, new_n17386, n5833);
xnor_4 g15066(new_n11280, new_n11256, n5840);
xor_4  g15067(new_n17225, new_n17224, n5841);
xnor_4 g15068(new_n11688, new_n11687, n5850);
xnor_4 g15069(new_n17299, new_n17290, n5903);
xnor_4 g15070(new_n14968, new_n7869, new_n17419);
nor_5  g15071(new_n14971, new_n7872, new_n17420);
nor_5  g15072(new_n16774, new_n16761, new_n17421_1);
nor_5  g15073(new_n17421_1, new_n17420, new_n17422);
xnor_4 g15074(new_n17422, new_n17419, new_n17423);
or_5   g15075(new_n16741, n6513, new_n17424);
xor_4  g15076(new_n17424, n26752, new_n17425);
xnor_4 g15077(new_n17425, new_n10054, new_n17426);
nor_5  g15078(new_n16742, new_n8013, new_n17427);
nor_5  g15079(new_n16759, new_n16743_1, new_n17428);
nor_5  g15080(new_n17428, new_n17427, new_n17429);
xor_4  g15081(new_n17429, new_n17426, new_n17430);
xnor_4 g15082(new_n17430, new_n17423, new_n17431);
nor_5  g15083(new_n16775, new_n16760, new_n17432_1);
nor_5  g15084(new_n16796, new_n16776, new_n17433);
nor_5  g15085(new_n17433, new_n17432_1, new_n17434);
xnor_4 g15086(new_n17434, new_n17431, n5904);
not_10 g15087(new_n9214, new_n17436_1);
xor_4  g15088(n27089, n6814, new_n17437);
nor_5  g15089(new_n8153, n11841, new_n17438);
xor_4  g15090(n19701, n11841, new_n17439);
nor_5  g15091(new_n8156, n10710, new_n17440_1);
xor_4  g15092(n23529, n10710, new_n17441);
nor_5  g15093(new_n8159_1, n20929, new_n17442);
xor_4  g15094(n24620, n20929, new_n17443);
nor_5  g15095(n8006, new_n8162, new_n17444);
xor_4  g15096(n8006, n5211, new_n17445);
nor_5  g15097(n25074, new_n8165, new_n17446);
xor_4  g15098(n25074, n12956, new_n17447);
nor_5  g15099(n18295, new_n4027, new_n17448);
nor_5  g15100(new_n8168, n16396, new_n17449);
nor_5  g15101(new_n4030, n6502, new_n17450_1);
or_5   g15102(n9399, new_n8172, new_n17451);
nor_5  g15103(n15780, new_n4033, new_n17452);
and_5  g15104(new_n17452, new_n17451, new_n17453);
nor_5  g15105(new_n17453, new_n17450_1, new_n17454);
nor_5  g15106(new_n17454, new_n17449, new_n17455);
or_5   g15107(new_n17455, new_n17448, new_n17456);
nor_5  g15108(new_n17456, new_n17447, new_n17457);
nor_5  g15109(new_n17457, new_n17446, new_n17458_1);
nor_5  g15110(new_n17458_1, new_n17445, new_n17459);
nor_5  g15111(new_n17459, new_n17444, new_n17460);
nor_5  g15112(new_n17460, new_n17443, new_n17461_1);
nor_5  g15113(new_n17461_1, new_n17442, new_n17462);
nor_5  g15114(new_n17462, new_n17441, new_n17463);
nor_5  g15115(new_n17463, new_n17440_1, new_n17464);
nor_5  g15116(new_n17464, new_n17439, new_n17465);
nor_5  g15117(new_n17465, new_n17438, new_n17466_1);
xor_4  g15118(new_n17466_1, new_n17437, new_n17467);
xnor_4 g15119(new_n17467, new_n17436_1, new_n17468);
not_10 g15120(new_n9218, new_n17469);
xor_4  g15121(new_n17464, new_n17439, new_n17470);
nor_5  g15122(new_n17470, new_n17469, new_n17471);
xnor_4 g15123(new_n17470, new_n17469, new_n17472);
not_10 g15124(new_n9222, new_n17473);
xor_4  g15125(new_n17462, new_n17441, new_n17474);
nor_5  g15126(new_n17474, new_n17473, new_n17475);
xnor_4 g15127(new_n17474, new_n17473, new_n17476);
not_10 g15128(new_n9226, new_n17477);
xor_4  g15129(new_n17460, new_n17443, new_n17478);
nor_5  g15130(new_n17478, new_n17477, new_n17479);
xor_4  g15131(new_n17458_1, new_n17445, new_n17480);
nor_5  g15132(new_n17480, new_n9229, new_n17481);
xnor_4 g15133(new_n17480, new_n9229, new_n17482);
xor_4  g15134(new_n17456, new_n17447, new_n17483);
nor_5  g15135(new_n17483, new_n9232, new_n17484);
xnor_4 g15136(n18295, n16396, new_n17485);
xnor_4 g15137(new_n17485, new_n17454, new_n17486);
and_5  g15138(new_n17486, new_n9235, new_n17487);
xnor_4 g15139(new_n17486, new_n9239, new_n17488);
xnor_4 g15140(n15780, n2088, new_n17489);
or_5   g15141(new_n17489, new_n9241, new_n17490);
xor_4  g15142(n9399, n6502, new_n17491);
xnor_4 g15143(new_n17491, new_n17452, new_n17492);
nor_5  g15144(new_n17492, new_n17490, new_n17493_1);
xnor_4 g15145(new_n17492, new_n17490, new_n17494);
nor_5  g15146(new_n17494, new_n9247, new_n17495);
nor_5  g15147(new_n17495, new_n17493_1, new_n17496);
and_5  g15148(new_n17496, new_n17488, new_n17497);
nor_5  g15149(new_n17497, new_n17487, new_n17498);
xnor_4 g15150(new_n17483, new_n9232, new_n17499);
nor_5  g15151(new_n17499, new_n17498, new_n17500_1);
nor_5  g15152(new_n17500_1, new_n17484, new_n17501);
nor_5  g15153(new_n17501, new_n17482, new_n17502);
nor_5  g15154(new_n17502, new_n17481, new_n17503);
xnor_4 g15155(new_n17478, new_n17477, new_n17504);
nor_5  g15156(new_n17504, new_n17503, new_n17505);
nor_5  g15157(new_n17505, new_n17479, new_n17506);
nor_5  g15158(new_n17506, new_n17476, new_n17507);
nor_5  g15159(new_n17507, new_n17475, new_n17508);
nor_5  g15160(new_n17508, new_n17472, new_n17509);
nor_5  g15161(new_n17509, new_n17471, new_n17510);
xnor_4 g15162(new_n17510, new_n17468, n5911);
xor_4  g15163(new_n10745, new_n3683, n5936);
xnor_4 g15164(new_n9086, new_n9052, n5943);
xnor_4 g15165(new_n12882, new_n12854, n5964);
nor_5  g15166(new_n4687, n11184, new_n17515);
nor_5  g15167(new_n4674_1, n23146, new_n17516);
nor_5  g15168(new_n4696, n17968, new_n17517);
not_10 g15169(new_n17517, new_n17518);
nor_5  g15170(new_n17518, new_n4678, new_n17519);
nor_5  g15171(new_n17519, new_n17516, new_n17520);
nor_5  g15172(new_n17520, new_n4688, new_n17521);
or_5   g15173(new_n17521, new_n17515, new_n17522);
nor_5  g15174(new_n17522, new_n14457_1, new_n17523);
nor_5  g15175(new_n17521, new_n17515, new_n17524_1);
nor_5  g15176(new_n17524_1, new_n14465, new_n17525);
nor_5  g15177(new_n17525, new_n14464_1, new_n17526);
nor_5  g15178(new_n17526, new_n17523, new_n17527);
nor_5  g15179(new_n17527, new_n14452, new_n17528);
or_5   g15180(new_n17526, new_n17523, new_n17529_1);
nor_5  g15181(new_n17529_1, new_n14455, new_n17530);
nor_5  g15182(new_n17530, new_n14454, new_n17531);
nor_5  g15183(new_n17531, new_n17528, new_n17532);
nor_5  g15184(new_n17532, new_n14447, new_n17533);
or_5   g15185(new_n17531, new_n17528, new_n17534);
nor_5  g15186(new_n17534, new_n14450, new_n17535);
nor_5  g15187(new_n17535, new_n14449, new_n17536);
nor_5  g15188(new_n17536, new_n17533, new_n17537);
nor_5  g15189(new_n17537, new_n14445, new_n17538);
or_5   g15190(new_n17536, new_n17533, new_n17539);
nor_5  g15191(new_n17539, new_n14474, new_n17540);
nor_5  g15192(new_n17540, new_n14473, new_n17541);
nor_5  g15193(new_n17541, new_n17538, new_n17542);
nor_5  g15194(new_n17542, new_n14443, new_n17543);
or_5   g15195(new_n17541, new_n17538, new_n17544);
nor_5  g15196(new_n17544, new_n14478, new_n17545);
nor_5  g15197(new_n17545, new_n14477, new_n17546);
nor_5  g15198(new_n17546, new_n17543, new_n17547);
xnor_4 g15199(new_n17547, new_n14442, new_n17548);
xnor_4 g15200(new_n17548, new_n3078, new_n17549);
xnor_4 g15201(new_n17542, new_n14478, new_n17550);
and_5  g15202(new_n17550, new_n3083, new_n17551);
xnor_4 g15203(new_n17550, new_n3083, new_n17552);
not_10 g15204(new_n3088, new_n17553);
xor_4  g15205(new_n17537, new_n14474, new_n17554);
nor_5  g15206(new_n17554, new_n17553, new_n17555);
xnor_4 g15207(new_n17554, new_n17553, new_n17556);
not_10 g15208(new_n3093, new_n17557_1);
xnor_4 g15209(new_n17532, new_n14451, new_n17558);
nor_5  g15210(new_n17558, new_n17557_1, new_n17559);
xnor_4 g15211(new_n17558, new_n17557_1, new_n17560);
xnor_4 g15212(new_n17527, new_n14455, new_n17561);
and_5  g15213(new_n17561, new_n3097, new_n17562);
xnor_4 g15214(new_n17561, new_n3097, new_n17563);
xor_4  g15215(new_n17524_1, new_n14465, new_n17564);
and_5  g15216(new_n17564, new_n3102, new_n17565);
xnor_4 g15217(new_n17564, new_n3102, new_n17566);
xor_4  g15218(new_n17520, new_n4688, new_n17567);
and_5  g15219(new_n17567, new_n3107, new_n17568);
xnor_4 g15220(new_n17567, new_n3107, new_n17569);
xnor_4 g15221(new_n17517, new_n4678, new_n17570);
and_5  g15222(new_n17570, new_n3116, new_n17571);
or_5   g15223(new_n4697, new_n3112, new_n17572);
xnor_4 g15224(new_n17570, new_n3117, new_n17573);
and_5  g15225(new_n17573, new_n17572, new_n17574);
nor_5  g15226(new_n17574, new_n17571, new_n17575);
nor_5  g15227(new_n17575, new_n17569, new_n17576);
nor_5  g15228(new_n17576, new_n17568, new_n17577);
nor_5  g15229(new_n17577, new_n17566, new_n17578);
nor_5  g15230(new_n17578, new_n17565, new_n17579);
nor_5  g15231(new_n17579, new_n17563, new_n17580);
nor_5  g15232(new_n17580, new_n17562, new_n17581);
nor_5  g15233(new_n17581, new_n17560, new_n17582);
nor_5  g15234(new_n17582, new_n17559, new_n17583_1);
nor_5  g15235(new_n17583_1, new_n17556, new_n17584);
nor_5  g15236(new_n17584, new_n17555, new_n17585);
nor_5  g15237(new_n17585, new_n17552, new_n17586);
nor_5  g15238(new_n17586, new_n17551, new_n17587);
xnor_4 g15239(new_n17587, new_n17549, n5980);
xnor_4 g15240(new_n10147, new_n10124, n6012);
and_5  g15241(new_n9166_1, new_n8147, new_n17590);
xor_4  g15242(new_n9166_1, n16544, new_n17591);
nor_5  g15243(new_n9168, n6814, new_n17592_1);
xnor_4 g15244(new_n9168, n6814, new_n17593);
nor_5  g15245(new_n9171, n19701, new_n17594);
xnor_4 g15246(new_n9171, n19701, new_n17595);
nor_5  g15247(new_n8437, n23529, new_n17596);
nor_5  g15248(new_n8465, new_n8438, new_n17597);
nor_5  g15249(new_n17597, new_n17596, new_n17598);
nor_5  g15250(new_n17598, new_n17595, new_n17599);
nor_5  g15251(new_n17599, new_n17594, new_n17600);
nor_5  g15252(new_n17600, new_n17593, new_n17601);
nor_5  g15253(new_n17601, new_n17592_1, new_n17602);
nor_5  g15254(new_n17602, new_n17591, new_n17603);
nor_5  g15255(new_n17603, new_n17590, new_n17604);
nand_5 g15256(new_n17604, new_n9160, new_n17605);
nor_5  g15257(new_n12732, n3582, new_n17606);
xnor_4 g15258(new_n12732, n3582, new_n17607);
nor_5  g15259(new_n12735, n2145, new_n17608);
xnor_4 g15260(new_n12735, n2145, new_n17609);
nor_5  g15261(new_n12737, n5031, new_n17610);
xor_4  g15262(new_n12737, n5031, new_n17611);
and_5  g15263(new_n8489_1, n11044, new_n17612);
nor_5  g15264(new_n8517, new_n8490, new_n17613);
nor_5  g15265(new_n17613, new_n17612, new_n17614);
and_5  g15266(new_n17614, new_n17611, new_n17615);
nor_5  g15267(new_n17615, new_n17610, new_n17616);
nor_5  g15268(new_n17616, new_n17609, new_n17617);
nor_5  g15269(new_n17617, new_n17608, new_n17618);
nor_5  g15270(new_n17618, new_n17607, new_n17619);
nor_5  g15271(new_n17619, new_n17606, new_n17620);
and_5  g15272(new_n17620, new_n12774, new_n17621);
xnor_4 g15273(new_n17621, new_n17605, new_n17622);
xnor_4 g15274(new_n17604, new_n9160, new_n17623);
xor_4  g15275(new_n17620, new_n12774, new_n17624);
and_5  g15276(new_n17624, new_n17623, new_n17625);
xnor_4 g15277(new_n17624, new_n17623, new_n17626);
xnor_4 g15278(new_n17602, new_n17591, new_n17627);
xor_4  g15279(new_n17618, new_n17607, new_n17628);
nor_5  g15280(new_n17628, new_n17627, new_n17629);
xnor_4 g15281(new_n17628, new_n17627, new_n17630);
xnor_4 g15282(new_n17600, new_n17593, new_n17631);
xor_4  g15283(new_n17616, new_n17609, new_n17632);
nor_5  g15284(new_n17632, new_n17631, new_n17633);
xnor_4 g15285(new_n17632, new_n17631, new_n17634);
xnor_4 g15286(new_n17598, new_n17595, new_n17635);
xor_4  g15287(new_n17614, new_n17611, new_n17636);
nor_5  g15288(new_n17636, new_n17635, new_n17637);
xnor_4 g15289(new_n17636, new_n17635, new_n17638_1);
and_5  g15290(new_n8518, new_n8466, new_n17639);
nor_5  g15291(new_n8553, new_n8519_1, new_n17640);
nor_5  g15292(new_n17640, new_n17639, new_n17641);
nor_5  g15293(new_n17641, new_n17638_1, new_n17642);
nor_5  g15294(new_n17642, new_n17637, new_n17643);
nor_5  g15295(new_n17643, new_n17634, new_n17644);
nor_5  g15296(new_n17644, new_n17633, new_n17645);
nor_5  g15297(new_n17645, new_n17630, new_n17646);
nor_5  g15298(new_n17646, new_n17629, new_n17647);
nor_5  g15299(new_n17647, new_n17626, new_n17648);
nor_5  g15300(new_n17648, new_n17625, new_n17649);
xnor_4 g15301(new_n17649, new_n17622, n6022);
xnor_4 g15302(new_n17304, new_n17287, n6031);
xnor_4 g15303(new_n7292, new_n7241, new_n17652);
nor_5  g15304(new_n15041, n1222, new_n17653);
xnor_4 g15305(new_n17653, n17458, new_n17654);
xor_4  g15306(new_n17654, n12507, new_n17655);
or_5   g15307(new_n15042, n15077, new_n17656);
or_5   g15308(new_n15080, new_n15043, new_n17657);
and_5  g15309(new_n17657, new_n17656, new_n17658);
xnor_4 g15310(new_n17658, new_n17655, new_n17659);
xnor_4 g15311(new_n17659, new_n5231, new_n17660);
and_5  g15312(new_n15081, new_n7302, new_n17661);
nor_5  g15313(new_n15123, new_n15082_1, new_n17662);
or_5   g15314(new_n17662, new_n17661, new_n17663);
xor_4  g15315(new_n17663, new_n17660, new_n17664_1);
xnor_4 g15316(new_n17664_1, new_n17652, new_n17665);
and_5  g15317(new_n15124, new_n7405, new_n17666);
nor_5  g15318(new_n15167_1, new_n15125, new_n17667);
nor_5  g15319(new_n17667, new_n17666, new_n17668);
xnor_4 g15320(new_n17668, new_n17665, n6044);
nor_5  g15321(new_n8310, new_n8266, new_n17670);
nor_5  g15322(new_n8364, new_n8311, new_n17671);
or_5   g15323(new_n17671, new_n17670, new_n17672);
nor_5  g15324(new_n8265, n4306, new_n17673);
xor_4  g15325(new_n16367_1, new_n17673, new_n17674);
xnor_4 g15326(new_n17674, new_n17672, new_n17675);
nor_5  g15327(new_n17675, new_n4201, new_n17676);
xnor_4 g15328(new_n17675, new_n4201, new_n17677);
not_10 g15329(new_n4207, new_n17678);
nor_5  g15330(new_n8365, new_n17678, new_n17679);
nor_5  g15331(new_n8410, new_n8366, new_n17680);
nor_5  g15332(new_n17680, new_n17679, new_n17681);
nor_5  g15333(new_n17681, new_n17677, new_n17682);
nor_5  g15334(new_n17682, new_n17676, new_n17683);
or_5   g15335(new_n16367_1, new_n17673, new_n17684);
nor_5  g15336(new_n17684, new_n17672, new_n17685);
nand_5 g15337(new_n17685, new_n16696, new_n17686);
nor_5  g15338(new_n17686, new_n17683, new_n17687_1);
nor_5  g15339(new_n17685, new_n16696, new_n17688);
and_5  g15340(new_n17688, new_n17683, new_n17689);
or_5   g15341(new_n17689, new_n17687_1, n6046);
xor_4  g15342(n17077, n7437, new_n17691);
nor_5  g15343(n26510, new_n15227, new_n17692);
xor_4  g15344(n26510, n20700, new_n17693);
nor_5  g15345(n23068, new_n15229, new_n17694);
nor_5  g15346(new_n17384, new_n17367, new_n17695);
nor_5  g15347(new_n17695, new_n17694, new_n17696);
nor_5  g15348(new_n17696, new_n17693, new_n17697);
nor_5  g15349(new_n17697, new_n17692, new_n17698);
xor_4  g15350(new_n17698, new_n17691, new_n17699);
xnor_4 g15351(n21997, n18483, new_n17700);
and_5  g15352(n25119, n21934, new_n17701);
or_5   g15353(n25119, n21934, new_n17702);
nor_5  g15354(n18901, n1163, new_n17703);
nor_5  g15355(new_n17350, new_n17339, new_n17704);
nor_5  g15356(new_n17704, new_n17703, new_n17705);
and_5  g15357(new_n17705, new_n17702, new_n17706);
or_5   g15358(new_n17706, new_n17701, new_n17707);
xor_4  g15359(new_n17707, new_n17700, new_n17708);
xnor_4 g15360(new_n17708, new_n6797, new_n17709);
xnor_4 g15361(n25119, n21934, new_n17710);
xnor_4 g15362(new_n17710, new_n17705, new_n17711);
or_5   g15363(new_n17711, new_n2415, new_n17712);
nor_5  g15364(new_n17351_1, new_n2409_1, new_n17713);
nor_5  g15365(new_n17365, new_n17352, new_n17714);
nor_5  g15366(new_n17714, new_n17713, new_n17715);
not_10 g15367(new_n17715, new_n17716);
xnor_4 g15368(new_n17711, new_n2415, new_n17717);
or_5   g15369(new_n17717, new_n17716, new_n17718);
nand_5 g15370(new_n17718, new_n17712, new_n17719);
xor_4  g15371(new_n17719, new_n17709, new_n17720);
xor_4  g15372(new_n17720, new_n17699, new_n17721_1);
xnor_4 g15373(new_n17696, new_n17693, new_n17722);
xnor_4 g15374(new_n17717, new_n17715, new_n17723);
nor_5  g15375(new_n17723, new_n17722, new_n17724);
nor_5  g15376(new_n17385, new_n17366, new_n17725);
and_5  g15377(new_n17413, new_n17386, new_n17726);
or_5   g15378(new_n17726, new_n17725, new_n17727);
xnor_4 g15379(new_n17723, new_n17722, new_n17728);
nor_5  g15380(new_n17728, new_n17727, new_n17729);
nor_5  g15381(new_n17729, new_n17724, new_n17730);
xnor_4 g15382(new_n17730, new_n17721_1, n6084);
xor_4  g15383(new_n17494, new_n9247, n6160);
xnor_4 g15384(new_n17499, new_n17498, n6171);
not_10 g15385(n10275, new_n17734);
nor_5  g15386(n22359, new_n17734, new_n17735_1);
not_10 g15387(new_n8971_1, new_n17736);
nor_5  g15388(new_n13722_1, new_n17736, new_n17737);
nor_5  g15389(new_n17737, new_n17735_1, new_n17738_1);
xnor_4 g15390(new_n17738_1, new_n8974, new_n17739);
xor_4  g15391(n26264, n21905, new_n17740);
nor_5  g15392(n22918, new_n7246, new_n17741);
xor_4  g15393(n22918, n7841, new_n17742);
nor_5  g15394(n25923, new_n7250, new_n17743);
xor_4  g15395(n25923, n16812, new_n17744);
nor_5  g15396(new_n7254, n6790, new_n17745);
nor_5  g15397(new_n16414, new_n16396_1, new_n17746_1);
nor_5  g15398(new_n17746_1, new_n17745, new_n17747);
nor_5  g15399(new_n17747, new_n17744, new_n17748);
nor_5  g15400(new_n17748, new_n17743, new_n17749_1);
nor_5  g15401(new_n17749_1, new_n17742, new_n17750);
nor_5  g15402(new_n17750, new_n17741, new_n17751);
xor_4  g15403(new_n17751, new_n17740, new_n17752);
xnor_4 g15404(new_n17752, new_n14017, new_n17753);
xor_4  g15405(new_n17749_1, new_n17742, new_n17754);
nor_5  g15406(new_n17754, new_n13783_1, new_n17755);
xor_4  g15407(new_n17754, new_n13783_1, new_n17756);
xor_4  g15408(new_n17747, new_n17744, new_n17757);
and_5  g15409(new_n17757, new_n13785, new_n17758);
xnor_4 g15410(new_n17757, new_n13785, new_n17759);
and_5  g15411(new_n16415, new_n13788, new_n17760);
nor_5  g15412(new_n16439_1, new_n16416, new_n17761);
nor_5  g15413(new_n17761, new_n17760, new_n17762);
nor_5  g15414(new_n17762, new_n17759, new_n17763);
nor_5  g15415(new_n17763, new_n17758, new_n17764);
and_5  g15416(new_n17764, new_n17756, new_n17765);
or_5   g15417(new_n17765, new_n17755, new_n17766);
xor_4  g15418(new_n17766, new_n17753, new_n17767);
xnor_4 g15419(new_n17767, new_n17739, new_n17768);
xnor_4 g15420(new_n17764, new_n17756, new_n17769);
nor_5  g15421(new_n17769, new_n13723, new_n17770);
xnor_4 g15422(new_n17769, new_n13723, new_n17771);
xor_4  g15423(new_n17762, new_n17759, new_n17772);
nor_5  g15424(new_n17772, new_n13725, new_n17773);
xnor_4 g15425(new_n17772, new_n13725, new_n17774);
nor_5  g15426(new_n16440_1, new_n13728, new_n17775);
nor_5  g15427(new_n16462, new_n16441, new_n17776);
nor_5  g15428(new_n17776, new_n17775, new_n17777);
nor_5  g15429(new_n17777, new_n17774, new_n17778);
nor_5  g15430(new_n17778, new_n17773, new_n17779);
nor_5  g15431(new_n17779, new_n17771, new_n17780);
nor_5  g15432(new_n17780, new_n17770, new_n17781);
xnor_4 g15433(new_n17781, new_n17768, n6183);
xnor_4 g15434(new_n8136, new_n8115, new_n17783);
xor_4  g15435(n14702, n14345, new_n17784_1);
nor_5  g15436(new_n8277, n2999, new_n17785);
xor_4  g15437(n11356, n2999, new_n17786);
nor_5  g15438(new_n8280, n2547, new_n17787);
xor_4  g15439(n3164, n2547, new_n17788);
and_5  g15440(new_n8283, n2680, new_n17789);
nor_5  g15441(new_n12702_1, new_n12693, new_n17790);
or_5   g15442(new_n17790, new_n17789, new_n17791);
nor_5  g15443(new_n17791, new_n17788, new_n17792);
nor_5  g15444(new_n17792, new_n17787, new_n17793);
nor_5  g15445(new_n17793, new_n17786, new_n17794);
nor_5  g15446(new_n17794, new_n17785, new_n17795);
xor_4  g15447(new_n17795, new_n17784_1, new_n17796);
xnor_4 g15448(new_n17796, new_n17783, new_n17797);
xnor_4 g15449(new_n8134, new_n8117, new_n17798);
xor_4  g15450(new_n17793, new_n17786, new_n17799);
nor_5  g15451(new_n17799, new_n17798, new_n17800);
xnor_4 g15452(new_n17799, new_n17798, new_n17801);
xnor_4 g15453(new_n8132, new_n8119, new_n17802);
xor_4  g15454(new_n17791, new_n17788, new_n17803);
nor_5  g15455(new_n17803, new_n17802, new_n17804);
xnor_4 g15456(new_n17803, new_n17802, new_n17805);
and_5  g15457(new_n12703, new_n8219, new_n17806);
nor_5  g15458(new_n12718, new_n12704, new_n17807);
nor_5  g15459(new_n17807, new_n17806, new_n17808);
nor_5  g15460(new_n17808, new_n17805, new_n17809);
nor_5  g15461(new_n17809, new_n17804, new_n17810);
nor_5  g15462(new_n17810, new_n17801, new_n17811);
or_5   g15463(new_n17811, new_n17800, new_n17812);
xor_4  g15464(new_n17812, new_n17797, n6189);
xor_4  g15465(n20036, n15167, new_n17814);
nor_5  g15466(new_n11109, n11192, new_n17815);
or_5   g15467(n21095, new_n3851, new_n17816);
and_5  g15468(new_n3854, n8656, new_n17817);
and_5  g15469(new_n17817, new_n17816, new_n17818);
nor_5  g15470(new_n17818, new_n17815, new_n17819);
xor_4  g15471(new_n17819, new_n17814, new_n17820_1);
xor_4  g15472(new_n17820_1, new_n16448, new_n17821);
xnor_4 g15473(n9380, n8656, new_n17822);
or_5   g15474(new_n17822, new_n13601, new_n17823);
xor_4  g15475(n21095, n11192, new_n17824);
xnor_4 g15476(new_n17824, new_n17817, new_n17825);
and_5  g15477(new_n17825, new_n17823, new_n17826);
not_10 g15478(new_n16454, new_n17827);
xor_4  g15479(new_n17825, new_n17823, new_n17828);
and_5  g15480(new_n17828, new_n17827, new_n17829);
nor_5  g15481(new_n17829, new_n17826, new_n17830);
xnor_4 g15482(new_n17830, new_n17821, n6223);
xnor_4 g15483(new_n12716, new_n12708, n6233);
xnor_4 g15484(new_n17022, new_n17019, n6245);
xnor_4 g15485(new_n9250, new_n9240, n6248);
xor_4  g15486(n21839, n16544, new_n17835);
nor_5  g15487(n27089, new_n8150, new_n17836);
nor_5  g15488(new_n17466_1, new_n17437, new_n17837);
nor_5  g15489(new_n17837, new_n17836, new_n17838);
xor_4  g15490(new_n17838, new_n17835, new_n17839);
xnor_4 g15491(new_n17839, new_n9210, new_n17840);
nor_5  g15492(new_n17467, new_n17436_1, new_n17841);
nor_5  g15493(new_n17510, new_n17468, new_n17842);
nor_5  g15494(new_n17842, new_n17841, new_n17843);
xnor_4 g15495(new_n17843, new_n17840, n6256);
xnor_4 g15496(new_n13479, new_n13464, n6271);
not_10 g15497(n14826, new_n17846);
nor_5  g15498(new_n17846, n13549, new_n17847);
not_10 g15499(new_n8977, new_n17848);
not_10 g15500(n23493, new_n17849);
nor_5  g15501(new_n17849, n8405, new_n17850);
not_10 g15502(new_n8974, new_n17851);
nor_5  g15503(new_n17738_1, new_n17851, new_n17852);
nor_5  g15504(new_n17852, new_n17850, new_n17853);
nor_5  g15505(new_n17853, new_n17848, new_n17854);
nor_5  g15506(new_n17854, new_n17847, new_n17855_1);
not_10 g15507(n2944, new_n17856);
nor_5  g15508(n13951, new_n17856, new_n17857);
xor_4  g15509(n13951, n2944, new_n17858);
not_10 g15510(n767, new_n17859);
nor_5  g15511(n22793, new_n17859, new_n17860);
nor_5  g15512(new_n13511, new_n13487_1, new_n17861);
nor_5  g15513(new_n17861, new_n17860, new_n17862);
nor_5  g15514(new_n17862, new_n17858, new_n17863);
nor_5  g15515(new_n17863, new_n17857, new_n17864);
and_5  g15516(new_n17864, new_n17855_1, new_n17865);
xor_4  g15517(new_n17862, new_n17858, new_n17866);
xnor_4 g15518(new_n17853, new_n8977, new_n17867);
nor_5  g15519(new_n17867, new_n17866, new_n17868);
xnor_4 g15520(new_n17867, new_n17866, new_n17869);
and_5  g15521(new_n17739, new_n13512, new_n17870);
xnor_4 g15522(new_n17739, new_n13512, new_n17871);
nor_5  g15523(new_n13723, new_n13514, new_n17872);
nor_5  g15524(new_n13742, new_n13724, new_n17873);
or_5   g15525(new_n17873, new_n17872, new_n17874);
nor_5  g15526(new_n17874, new_n17871, new_n17875);
or_5   g15527(new_n17875, new_n17870, new_n17876);
nor_5  g15528(new_n17876, new_n17869, new_n17877_1);
nor_5  g15529(new_n17877_1, new_n17868, new_n17878);
xnor_4 g15530(new_n17864, new_n17855_1, new_n17879);
nor_5  g15531(new_n17879, new_n17878, new_n17880);
nor_5  g15532(new_n17880, new_n17865, new_n17881);
nor_5  g15533(new_n13413, n1881, new_n17882);
xor_4  g15534(n8827, n1881, new_n17883);
not_10 g15535(n18035, new_n17884);
nor_5  g15536(new_n17884, n5834, new_n17885);
nor_5  g15537(new_n17277, new_n17273, new_n17886);
nor_5  g15538(new_n17886, new_n17885, new_n17887);
nor_5  g15539(new_n17887, new_n17883, new_n17888);
or_5   g15540(new_n17888, new_n17882, new_n17889_1);
xnor_4 g15541(new_n17889_1, new_n17881, new_n17890);
xor_4  g15542(new_n17879, new_n17878, new_n17891);
and_5  g15543(new_n17891, new_n17889_1, new_n17892);
nor_5  g15544(new_n17888, new_n17882, new_n17893);
xnor_4 g15545(new_n17891, new_n17893, new_n17894);
xnor_4 g15546(new_n17887, new_n17883, new_n17895);
xor_4  g15547(new_n17876, new_n17869, new_n17896);
nor_5  g15548(new_n17896, new_n17895, new_n17897);
xor_4  g15549(new_n17874, new_n17871, new_n17898);
nor_5  g15550(new_n17898, new_n17278, new_n17899);
xor_4  g15551(new_n17898, new_n17278, new_n17900);
and_5  g15552(new_n13973, new_n13743, new_n17901);
nor_5  g15553(new_n13992, new_n13974, new_n17902);
nor_5  g15554(new_n17902, new_n17901, new_n17903);
and_5  g15555(new_n17903, new_n17900, new_n17904);
or_5   g15556(new_n17904, new_n17899, new_n17905);
xnor_4 g15557(new_n17896, new_n17895, new_n17906);
nor_5  g15558(new_n17906, new_n17905, new_n17907);
nor_5  g15559(new_n17907, new_n17897, new_n17908);
and_5  g15560(new_n17908, new_n17894, new_n17909);
or_5   g15561(new_n17909, new_n17892, new_n17910);
xor_4  g15562(new_n17910, new_n17890, n6276);
xnor_4 g15563(new_n16982, new_n16981, n6308);
xnor_4 g15564(new_n15257, new_n15244, n6311);
xnor_4 g15565(new_n15023, new_n15009, n6323);
and_5  g15566(new_n5430_1, new_n5395, new_n17915);
nor_5  g15567(new_n5490, new_n5431, new_n17916);
nor_5  g15568(new_n17916, new_n17915, new_n17917);
nand_5 g15569(new_n12118, new_n12461_1, new_n17918);
nor_5  g15570(new_n17918, new_n17917, new_n17919);
nor_5  g15571(new_n12118, new_n12461_1, new_n17920);
and_5  g15572(new_n17920, new_n17917, new_n17921);
nor_5  g15573(new_n17921, new_n17919, new_n17922);
nor_5  g15574(new_n17922, new_n16239, new_n17923);
xnor_4 g15575(new_n17922, new_n16239, new_n17924);
xnor_4 g15576(new_n12118, new_n12461_1, new_n17925);
xnor_4 g15577(new_n17925, new_n17917, new_n17926);
nor_5  g15578(new_n17926, new_n16241, new_n17927_1);
xnor_4 g15579(new_n17926, new_n16241, new_n17928);
nor_5  g15580(new_n5570, new_n5491, new_n17929);
nor_5  g15581(new_n5622, new_n5571, new_n17930);
nor_5  g15582(new_n17930, new_n17929, new_n17931_1);
nor_5  g15583(new_n17931_1, new_n17928, new_n17932);
nor_5  g15584(new_n17932, new_n17927_1, new_n17933);
nor_5  g15585(new_n17933, new_n17924, new_n17934);
nor_5  g15586(new_n17934, new_n17923, new_n17935);
nor_5  g15587(new_n17935, new_n17919, n6330);
xnor_4 g15588(new_n7793, new_n7764, n6339);
xnor_4 g15589(new_n12685, new_n12659, n6354);
or_5   g15590(new_n3069, n7335, new_n17939);
nor_5  g15591(new_n3076_1, n5696, new_n17940);
xnor_4 g15592(new_n3076_1, n5696, new_n17941);
nor_5  g15593(new_n3081, n13367, new_n17942);
xnor_4 g15594(new_n3081, n13367, new_n17943);
nor_5  g15595(new_n3086, n932, new_n17944);
xnor_4 g15596(new_n3086, n932, new_n17945);
nor_5  g15597(new_n3091, n6691, new_n17946);
xnor_4 g15598(new_n3091, n6691, new_n17947);
nor_5  g15599(new_n3096, n3260, new_n17948_1);
xnor_4 g15600(new_n3096, n3260, new_n17949);
nor_5  g15601(new_n3101, n20489, new_n17950);
nor_5  g15602(new_n3106, n2355, new_n17951);
xnor_4 g15603(new_n3106, n2355, new_n17952);
nor_5  g15604(new_n3118, n11121, new_n17953);
nand_5 g15605(n16217, n12315, new_n17954_1);
xor_4  g15606(new_n3118, n11121, new_n17955);
and_5  g15607(new_n17955, new_n17954_1, new_n17956_1);
nor_5  g15608(new_n17956_1, new_n17953, new_n17957);
nor_5  g15609(new_n17957, new_n17952, new_n17958);
nor_5  g15610(new_n17958, new_n17951, new_n17959_1);
xnor_4 g15611(new_n3101, n20489, new_n17960);
nor_5  g15612(new_n17960, new_n17959_1, new_n17961);
nor_5  g15613(new_n17961, new_n17950, new_n17962);
nor_5  g15614(new_n17962, new_n17949, new_n17963_1);
nor_5  g15615(new_n17963_1, new_n17948_1, new_n17964);
nor_5  g15616(new_n17964, new_n17947, new_n17965);
nor_5  g15617(new_n17965, new_n17946, new_n17966);
nor_5  g15618(new_n17966, new_n17945, new_n17967);
nor_5  g15619(new_n17967, new_n17944, new_n17968_1);
nor_5  g15620(new_n17968_1, new_n17943, new_n17969);
nor_5  g15621(new_n17969, new_n17942, new_n17970);
nor_5  g15622(new_n17970, new_n17941, new_n17971);
nor_5  g15623(new_n17971, new_n17940, new_n17972);
and_5  g15624(new_n17972, new_n17939, new_n17973);
and_5  g15625(new_n3069, n7335, new_n17974);
or_5   g15626(new_n17974, new_n3074, new_n17975);
nor_5  g15627(new_n17975, new_n17973, new_n17976_1);
and_5  g15628(new_n17976_1, new_n15421, new_n17977);
nor_5  g15629(new_n17976_1, new_n15461, new_n17978);
xnor_4 g15630(new_n17976_1, new_n15461, new_n17979);
xor_4  g15631(new_n3069, n7335, new_n17980);
xnor_4 g15632(new_n17980, new_n17972, new_n17981);
and_5  g15633(new_n17981, new_n15464, new_n17982);
xnor_4 g15634(new_n17981, new_n15464, new_n17983);
xor_4  g15635(new_n17970, new_n17941, new_n17984);
and_5  g15636(new_n17984, new_n15470_1, new_n17985);
xnor_4 g15637(new_n17984, new_n15470_1, new_n17986);
xor_4  g15638(new_n17968_1, new_n17943, new_n17987);
and_5  g15639(new_n17987, new_n15474, new_n17988);
xnor_4 g15640(new_n17987, new_n15474, new_n17989);
xor_4  g15641(new_n17966, new_n17945, new_n17990);
and_5  g15642(new_n17990, new_n15478, new_n17991);
xnor_4 g15643(new_n17990, new_n15478, new_n17992);
xor_4  g15644(new_n17964, new_n17947, new_n17993);
and_5  g15645(new_n17993, new_n15482, new_n17994);
xnor_4 g15646(new_n17993, new_n15482, new_n17995);
xor_4  g15647(new_n17962, new_n17949, new_n17996);
and_5  g15648(new_n17996, new_n15486, new_n17997);
xnor_4 g15649(new_n17996, new_n15486, new_n17998_1);
xnor_4 g15650(new_n17960, new_n17959_1, new_n17999);
nor_5  g15651(new_n17999, new_n15489, new_n18000);
xor_4  g15652(new_n17999, new_n15489, new_n18001);
xor_4  g15653(new_n17957, new_n17952, new_n18002);
nor_5  g15654(new_n18002, new_n15494, new_n18003);
xnor_4 g15655(new_n18002, new_n15494, new_n18004);
nor_5  g15656(new_n17955, new_n15498, new_n18005);
xor_4  g15657(new_n17955, new_n17954_1, new_n18006);
or_5   g15658(new_n18006, new_n15497, new_n18007);
xnor_4 g15659(n16217, n12315, new_n18008);
or_5   g15660(new_n18008, new_n15503, new_n18009);
and_5  g15661(new_n18009, new_n18007, new_n18010);
or_5   g15662(new_n18010, new_n18005, new_n18011);
nor_5  g15663(new_n18011, new_n18004, new_n18012);
nor_5  g15664(new_n18012, new_n18003, new_n18013);
and_5  g15665(new_n18013, new_n18001, new_n18014);
nor_5  g15666(new_n18014, new_n18000, new_n18015);
nor_5  g15667(new_n18015, new_n17998_1, new_n18016);
nor_5  g15668(new_n18016, new_n17997, new_n18017);
nor_5  g15669(new_n18017, new_n17995, new_n18018);
nor_5  g15670(new_n18018, new_n17994, new_n18019);
nor_5  g15671(new_n18019, new_n17992, new_n18020);
nor_5  g15672(new_n18020, new_n17991, new_n18021);
nor_5  g15673(new_n18021, new_n17989, new_n18022);
nor_5  g15674(new_n18022, new_n17988, new_n18023);
nor_5  g15675(new_n18023, new_n17986, new_n18024);
nor_5  g15676(new_n18024, new_n17985, new_n18025_1);
nor_5  g15677(new_n18025_1, new_n17983, new_n18026);
nor_5  g15678(new_n18026, new_n17982, new_n18027);
nor_5  g15679(new_n18027, new_n17979, new_n18028);
nor_5  g15680(new_n18028, new_n17978, new_n18029);
nor_5  g15681(new_n18029, new_n17977, new_n18030);
nor_5  g15682(new_n17976_1, new_n15421, new_n18031);
nor_5  g15683(new_n18031, new_n18028, new_n18032);
nor_5  g15684(new_n18032, new_n18030, n6375);
xnor_4 g15685(new_n17139, new_n17126, n6383);
xnor_4 g15686(new_n13041, new_n13007, n6407);
xnor_4 g15687(new_n7785, new_n7784, n6431);
xnor_4 g15688(new_n14865, new_n14862, n6437);
xnor_4 g15689(new_n3886, new_n3885, n6457);
xnor_4 g15690(new_n11074, new_n11041, n6465);
and_5  g15691(new_n15715, n3740, new_n18040);
nor_5  g15692(new_n15714, n3582, new_n18041);
nor_5  g15693(new_n15715, n3740, new_n18042);
nor_5  g15694(new_n15720, new_n18042, new_n18043_1);
or_5   g15695(new_n18043_1, new_n18041, new_n18044);
or_5   g15696(new_n18044, new_n18040, new_n18045_1);
xnor_4 g15697(new_n18045_1, new_n7578, new_n18046);
not_10 g15698(new_n15721, new_n18047);
nor_5  g15699(new_n18047, new_n3304, new_n18048);
xnor_4 g15700(new_n15721, new_n3304, new_n18049);
not_10 g15701(new_n12928, new_n18050);
nor_5  g15702(new_n18050, new_n3306_1, new_n18051);
and_5  g15703(new_n12964, new_n12929, new_n18052);
nor_5  g15704(new_n18052, new_n18051, new_n18053);
and_5  g15705(new_n18053, new_n18049, new_n18054);
nor_5  g15706(new_n18054, new_n18048, new_n18055);
xor_4  g15707(new_n18055, new_n18046, new_n18056);
nor_5  g15708(new_n3406, n2743, new_n18057);
and_5  g15709(new_n3409, n7026, new_n18058);
nor_5  g15710(new_n3409, n7026, new_n18059_1);
nor_5  g15711(new_n12996, new_n18059_1, new_n18060);
nor_5  g15712(new_n18060, new_n18058, new_n18061_1);
nor_5  g15713(new_n18061_1, new_n18057, new_n18062);
and_5  g15714(new_n3405, new_n4441_1, new_n18063);
and_5  g15715(new_n3406, n2743, new_n18064);
or_5   g15716(new_n18064, new_n18063, new_n18065);
nor_5  g15717(new_n18065, new_n18062, new_n18066);
xnor_4 g15718(new_n18066, new_n18056, new_n18067);
xor_4  g15719(new_n18053, new_n18049, new_n18068);
xnor_4 g15720(new_n3406, new_n12179_1, new_n18069);
xnor_4 g15721(new_n18069, new_n18061_1, new_n18070);
nor_5  g15722(new_n18070, new_n18068, new_n18071_1);
xnor_4 g15723(new_n18070, new_n18068, new_n18072);
and_5  g15724(new_n12997, new_n12965, new_n18073);
and_5  g15725(new_n13045, new_n12998, new_n18074);
nor_5  g15726(new_n18074, new_n18073, new_n18075);
nor_5  g15727(new_n18075, new_n18072, new_n18076);
nor_5  g15728(new_n18076, new_n18071_1, new_n18077);
xnor_4 g15729(new_n18077, new_n18067, n6470);
xnor_4 g15730(new_n10402, new_n10380, n6476);
xnor_4 g15731(new_n16688_1, new_n16679, n6506);
xor_4  g15732(new_n8480_1, new_n8475, new_n18081);
nor_5  g15733(new_n8504, new_n8502, new_n18082);
nand_5 g15734(new_n18082, new_n18081, new_n18083);
or_5   g15735(new_n18083, new_n8497, new_n18084);
or_5   g15736(new_n18084, new_n8494, new_n18085);
or_5   g15737(new_n18085, new_n8491, new_n18086);
or_5   g15738(new_n18086, new_n8489_1, new_n18087);
or_5   g15739(new_n18087, new_n12737, new_n18088);
xor_4  g15740(new_n18088, new_n12735, new_n18089);
xnor_4 g15741(new_n18089, new_n9168, new_n18090);
xor_4  g15742(new_n18087, new_n12737, new_n18091);
nor_5  g15743(new_n18091, new_n9171, new_n18092);
xnor_4 g15744(new_n18091, new_n9171, new_n18093);
xor_4  g15745(new_n18086, new_n8489_1, new_n18094);
nor_5  g15746(new_n18094, new_n8437, new_n18095);
xnor_4 g15747(new_n18094, new_n8437, new_n18096);
xor_4  g15748(new_n18085, new_n8491, new_n18097);
nor_5  g15749(new_n18097, new_n8439_1, new_n18098);
xnor_4 g15750(new_n18097, new_n8439_1, new_n18099);
not_10 g15751(new_n8442, new_n18100);
xor_4  g15752(new_n18084, new_n8494, new_n18101);
nor_5  g15753(new_n18101, new_n18100, new_n18102);
xor_4  g15754(new_n18101, new_n8442, new_n18103);
xor_4  g15755(new_n18083, new_n8497, new_n18104);
nor_5  g15756(new_n18104, new_n8445, new_n18105_1);
xnor_4 g15757(new_n18082, new_n8500, new_n18106);
nor_5  g15758(new_n18106, new_n8448, new_n18107);
xnor_4 g15759(new_n18106, new_n8448, new_n18108);
and_5  g15760(new_n8504, new_n8452, new_n18109);
nor_5  g15761(new_n18109, new_n8450, new_n18110);
not_10 g15762(new_n8504, new_n18111);
nor_5  g15763(new_n18111, new_n8478, new_n18112);
nor_5  g15764(new_n18112, new_n18082, new_n18113);
xor_4  g15765(n27188, n4326, new_n18114);
and_5  g15766(new_n18109, new_n18114, new_n18115);
or_5   g15767(new_n18115, new_n18110, new_n18116);
nor_5  g15768(new_n18116, new_n18113, new_n18117);
nor_5  g15769(new_n18117, new_n18110, new_n18118);
nor_5  g15770(new_n18118, new_n18108, new_n18119);
nor_5  g15771(new_n18119, new_n18107, new_n18120);
xnor_4 g15772(new_n18104, new_n8445, new_n18121);
nor_5  g15773(new_n18121, new_n18120, new_n18122);
nor_5  g15774(new_n18122, new_n18105_1, new_n18123);
nor_5  g15775(new_n18123, new_n18103, new_n18124);
nor_5  g15776(new_n18124, new_n18102, new_n18125);
nor_5  g15777(new_n18125, new_n18099, new_n18126);
nor_5  g15778(new_n18126, new_n18098, new_n18127);
nor_5  g15779(new_n18127, new_n18096, new_n18128);
nor_5  g15780(new_n18128, new_n18095, new_n18129);
nor_5  g15781(new_n18129, new_n18093, new_n18130);
nor_5  g15782(new_n18130, new_n18092, new_n18131);
xor_4  g15783(new_n18131, new_n18090, new_n18132);
xnor_4 g15784(new_n18132, new_n15081, new_n18133);
xor_4  g15785(new_n18129, new_n18093, new_n18134);
and_5  g15786(new_n18134, new_n15083, new_n18135);
xnor_4 g15787(new_n18134, new_n15083, new_n18136);
not_10 g15788(new_n15087, new_n18137);
xor_4  g15789(new_n18127, new_n18096, new_n18138);
and_5  g15790(new_n18138, new_n18137, new_n18139);
xnor_4 g15791(new_n18138, new_n18137, new_n18140);
xor_4  g15792(new_n18125, new_n18099, new_n18141);
and_5  g15793(new_n18141, new_n15090, new_n18142);
xor_4  g15794(new_n18141, new_n15090, new_n18143_1);
xor_4  g15795(new_n18123, new_n18103, new_n18144);
nor_5  g15796(new_n18144, new_n15093, new_n18145_1);
xor_4  g15797(new_n18121, new_n18120, new_n18146);
nor_5  g15798(new_n18146, new_n15096, new_n18147);
xnor_4 g15799(new_n18146, new_n15096, new_n18148);
xor_4  g15800(new_n18118, new_n18108, new_n18149);
nor_5  g15801(new_n18149, new_n15099, new_n18150);
xnor_4 g15802(new_n18149, new_n15099, new_n18151_1);
xor_4  g15803(new_n18116, new_n18113, new_n18152_1);
nor_5  g15804(new_n18152_1, new_n15105, new_n18153);
xor_4  g15805(new_n8504, new_n8452, new_n18154);
nand_5 g15806(new_n18154, new_n15107, new_n18155);
xnor_4 g15807(new_n18152_1, new_n15105, new_n18156);
nor_5  g15808(new_n18156, new_n18155, new_n18157_1);
nor_5  g15809(new_n18157_1, new_n18153, new_n18158);
nor_5  g15810(new_n18158, new_n18151_1, new_n18159);
nor_5  g15811(new_n18159, new_n18150, new_n18160);
nor_5  g15812(new_n18160, new_n18148, new_n18161);
nor_5  g15813(new_n18161, new_n18147, new_n18162);
xnor_4 g15814(new_n18144, new_n15093, new_n18163);
nor_5  g15815(new_n18163, new_n18162, new_n18164);
nor_5  g15816(new_n18164, new_n18145_1, new_n18165);
and_5  g15817(new_n18165, new_n18143_1, new_n18166);
nor_5  g15818(new_n18166, new_n18142, new_n18167);
nor_5  g15819(new_n18167, new_n18140, new_n18168);
nor_5  g15820(new_n18168, new_n18139, new_n18169);
nor_5  g15821(new_n18169, new_n18136, new_n18170);
or_5   g15822(new_n18170, new_n18135, new_n18171_1);
xor_4  g15823(new_n18171_1, new_n18133, n6514);
nor_5  g15824(new_n10371, new_n10293, new_n18173);
nor_5  g15825(new_n10406, new_n10372_1, new_n18174);
nor_5  g15826(new_n18174, new_n18173, new_n18175);
xor_4  g15827(new_n10333, new_n13634, new_n18176);
and_5  g15828(new_n18176, new_n10370, new_n18177);
nor_5  g15829(new_n10333, new_n10326_1, new_n18178);
or_5   g15830(new_n10370, new_n18178, new_n18179);
nor_5  g15831(new_n18179, new_n18176, new_n18180);
or_5   g15832(new_n18180, new_n18177, new_n18181);
xnor_4 g15833(new_n18181, new_n18175, n6542);
xnor_4 g15834(new_n13877, new_n13865, n6558);
xnor_4 g15835(new_n16226, new_n16224, n6560);
xnor_4 g15836(new_n5711, n10405, new_n18185);
and_5  g15837(new_n11200, n11302, new_n18186);
xor_4  g15838(new_n5713, n11302, new_n18187);
not_10 g15839(n17090, new_n18188);
and_5  g15840(new_n5716, new_n18188, new_n18189);
nand_5 g15841(new_n5718, n6773, new_n18190);
xnor_4 g15842(new_n5716, n17090, new_n18191);
and_5  g15843(new_n18191, new_n18190, new_n18192);
or_5   g15844(new_n18192, new_n18189, new_n18193_1);
nor_5  g15845(new_n18193_1, new_n18187, new_n18194);
nor_5  g15846(new_n18194, new_n18186, new_n18195);
xor_4  g15847(new_n18195, new_n18185, new_n18196);
xnor_4 g15848(new_n18196, new_n8803_1, new_n18197);
not_10 g15849(new_n8807, new_n18198);
xor_4  g15850(new_n18193_1, new_n18187, new_n18199);
nor_5  g15851(new_n18199, new_n18198, new_n18200);
xor_4  g15852(new_n18199, new_n8807, new_n18201);
xor_4  g15853(new_n18191, new_n18190, new_n18202);
and_5  g15854(new_n18202, new_n8812, new_n18203);
nor_5  g15855(new_n16251, new_n8815, new_n18204);
xnor_4 g15856(new_n18202, new_n8811, new_n18205);
and_5  g15857(new_n18205, new_n18204, new_n18206);
nor_5  g15858(new_n18206, new_n18203, new_n18207);
nor_5  g15859(new_n18207, new_n18201, new_n18208);
nor_5  g15860(new_n18208, new_n18200, new_n18209);
xnor_4 g15861(new_n18209, new_n18197, n6567);
or_5   g15862(new_n12324_1, n8324, new_n18211);
or_5   g15863(new_n18211, n1279, new_n18212);
or_5   g15864(new_n18212, n9445, new_n18213);
nor_5  g15865(new_n18213, n19454, new_n18214);
xnor_4 g15866(new_n18214, n1536, new_n18215);
xnor_4 g15867(new_n18215, new_n4148, new_n18216);
xor_4  g15868(new_n18213, n19454, new_n18217);
nor_5  g15869(new_n18217, new_n4153_1, new_n18218);
xnor_4 g15870(new_n18217, new_n4153_1, new_n18219);
xor_4  g15871(new_n18212, n9445, new_n18220);
nor_5  g15872(new_n18220, new_n4157, new_n18221);
xnor_4 g15873(new_n18220, new_n4157, new_n18222);
xor_4  g15874(new_n18211, n1279, new_n18223);
nor_5  g15875(new_n18223, new_n4161, new_n18224);
xnor_4 g15876(new_n18223, new_n4161, new_n18225);
nor_5  g15877(new_n12325_1, new_n3725_1, new_n18226);
nor_5  g15878(new_n12347, new_n12326, new_n18227_1);
nor_5  g15879(new_n18227_1, new_n18226, new_n18228);
nor_5  g15880(new_n18228, new_n18225, new_n18229);
nor_5  g15881(new_n18229, new_n18224, new_n18230);
nor_5  g15882(new_n18230, new_n18222, new_n18231);
nor_5  g15883(new_n18231, new_n18221, new_n18232_1);
nor_5  g15884(new_n18232_1, new_n18219, new_n18233);
nor_5  g15885(new_n18233, new_n18218, new_n18234);
xor_4  g15886(new_n18234, new_n18216, new_n18235);
xnor_4 g15887(new_n7345, n23272, new_n18236);
nor_5  g15888(new_n7348, n11481, new_n18237);
xnor_4 g15889(new_n7348, n11481, new_n18238_1);
nor_5  g15890(new_n7351, n16439, new_n18239);
xnor_4 g15891(new_n7351, n16439, new_n18240);
or_5   g15892(new_n7354, n15241, new_n18241_1);
and_5  g15893(new_n7357, n7678, new_n18242);
nor_5  g15894(new_n12367, new_n12350, new_n18243);
nor_5  g15895(new_n18243, new_n18242, new_n18244);
not_10 g15896(new_n18244, new_n18245);
xnor_4 g15897(new_n7354, n15241, new_n18246);
or_5   g15898(new_n18246, new_n18245, new_n18247);
and_5  g15899(new_n18247, new_n18241_1, new_n18248);
nor_5  g15900(new_n18248, new_n18240, new_n18249);
nor_5  g15901(new_n18249, new_n18239, new_n18250);
nor_5  g15902(new_n18250, new_n18238_1, new_n18251);
or_5   g15903(new_n18251, new_n18237, new_n18252);
xor_4  g15904(new_n18252, new_n18236, new_n18253);
xnor_4 g15905(new_n18253, new_n18235, new_n18254_1);
xor_4  g15906(new_n18232_1, new_n18219, new_n18255);
xor_4  g15907(new_n18250, new_n18238_1, new_n18256);
and_5  g15908(new_n18256, new_n18255, new_n18257);
xnor_4 g15909(new_n18256, new_n18255, new_n18258);
xor_4  g15910(new_n18230, new_n18222, new_n18259);
xor_4  g15911(new_n18248, new_n18240, new_n18260);
and_5  g15912(new_n18260, new_n18259, new_n18261);
xnor_4 g15913(new_n18260, new_n18259, new_n18262);
xor_4  g15914(new_n18228, new_n18225, new_n18263);
xnor_4 g15915(new_n18246, new_n18244, new_n18264);
and_5  g15916(new_n18264, new_n18263, new_n18265);
xnor_4 g15917(new_n18264, new_n18263, new_n18266);
nor_5  g15918(new_n12368, new_n12349_1, new_n18267);
nor_5  g15919(new_n12399, new_n12369, new_n18268);
nor_5  g15920(new_n18268, new_n18267, new_n18269);
nor_5  g15921(new_n18269, new_n18266, new_n18270);
nor_5  g15922(new_n18270, new_n18265, new_n18271);
nor_5  g15923(new_n18271, new_n18262, new_n18272);
nor_5  g15924(new_n18272, new_n18261, new_n18273);
nor_5  g15925(new_n18273, new_n18258, new_n18274_1);
nor_5  g15926(new_n18274_1, new_n18257, new_n18275);
xnor_4 g15927(new_n18275, new_n18254_1, n6576);
xor_4  g15928(new_n18006, new_n15497, new_n18277);
xnor_4 g15929(new_n18277, new_n18009, n6587);
xnor_4 g15930(new_n16994_1, new_n16951_1, n6612);
nor_5  g15931(new_n15767, new_n9721, new_n18280);
xnor_4 g15932(new_n15767, new_n9721, new_n18281);
nor_5  g15933(new_n15769, new_n9714, new_n18282);
xnor_4 g15934(new_n15769, new_n9714, new_n18283);
nor_5  g15935(new_n15772, new_n9707, new_n18284);
xnor_4 g15936(new_n15772, new_n9707, new_n18285);
nor_5  g15937(new_n15775, new_n9700, new_n18286);
xnor_4 g15938(new_n15775, new_n9700, new_n18287);
nor_5  g15939(new_n15778, new_n9693, new_n18288_1);
xnor_4 g15940(new_n15778, new_n9693, new_n18289);
or_5   g15941(new_n15780_1, new_n9686, new_n18290_1);
xnor_4 g15942(new_n15780_1, new_n9686, new_n18291);
or_5   g15943(new_n13605, new_n9679, new_n18292);
xnor_4 g15944(new_n13605, new_n9679, new_n18293);
and_5  g15945(new_n13607, new_n9673, new_n18294);
nor_5  g15946(new_n9745, n18, new_n18295_1);
and_5  g15947(new_n18295_1, new_n8290, new_n18296);
not_10 g15948(new_n13610, new_n18297);
nor_5  g15949(new_n18295_1, new_n18297, new_n18298);
nor_5  g15950(new_n18298, new_n18296, new_n18299);
and_5  g15951(new_n18299, new_n9667, new_n18300);
or_5   g15952(new_n18300, new_n18296, new_n18301_1);
xnor_4 g15953(new_n13607, new_n9673, new_n18302);
nor_5  g15954(new_n18302, new_n18301_1, new_n18303);
nor_5  g15955(new_n18303, new_n18294, new_n18304_1);
not_10 g15956(new_n18304_1, new_n18305);
or_5   g15957(new_n18305, new_n18293, new_n18306);
and_5  g15958(new_n18306, new_n18292, new_n18307);
or_5   g15959(new_n18307, new_n18291, new_n18308);
and_5  g15960(new_n18308, new_n18290_1, new_n18309);
nor_5  g15961(new_n18309, new_n18289, new_n18310_1);
nor_5  g15962(new_n18310_1, new_n18288_1, new_n18311_1);
nor_5  g15963(new_n18311_1, new_n18287, new_n18312);
nor_5  g15964(new_n18312, new_n18286, new_n18313);
nor_5  g15965(new_n18313, new_n18285, new_n18314);
nor_5  g15966(new_n18314, new_n18284, new_n18315);
nor_5  g15967(new_n18315, new_n18283, new_n18316);
nor_5  g15968(new_n18316, new_n18282, new_n18317);
nor_5  g15969(new_n18317, new_n18281, new_n18318);
nor_5  g15970(new_n18318, new_n18280, new_n18319);
nor_5  g15971(new_n15766_1, n23166, new_n18320);
and_5  g15972(new_n15937, new_n18320, new_n18321);
and_5  g15973(new_n18321, new_n18319, new_n18322);
or_5   g15974(new_n15937, new_n18320, new_n18323_1);
nor_5  g15975(new_n18323_1, new_n18319, new_n18324);
nor_5  g15976(new_n18324, new_n18322, new_n18325);
xnor_4 g15977(new_n15936_1, new_n18320, new_n18326);
xnor_4 g15978(new_n18326, new_n18319, new_n18327);
nor_5  g15979(new_n18327, new_n17624, new_n18328);
xnor_4 g15980(new_n18327, new_n17624, new_n18329);
xor_4  g15981(new_n18317, new_n18281, new_n18330);
and_5  g15982(new_n18330, new_n17628, new_n18331);
xnor_4 g15983(new_n18330, new_n17628, new_n18332_1);
xor_4  g15984(new_n18315, new_n18283, new_n18333);
and_5  g15985(new_n18333, new_n17632, new_n18334);
xnor_4 g15986(new_n18333, new_n17632, new_n18335);
xor_4  g15987(new_n18313, new_n18285, new_n18336);
and_5  g15988(new_n18336, new_n17636, new_n18337);
xnor_4 g15989(new_n18336, new_n17636, new_n18338);
not_10 g15990(new_n8518, new_n18339);
xor_4  g15991(new_n18311_1, new_n18287, new_n18340);
and_5  g15992(new_n18340, new_n18339, new_n18341);
xnor_4 g15993(new_n18340, new_n18339, new_n18342);
not_10 g15994(new_n8521, new_n18343_1);
xor_4  g15995(new_n18309, new_n18289, new_n18344);
and_5  g15996(new_n18344, new_n18343_1, new_n18345_1);
xnor_4 g15997(new_n18344, new_n18343_1, new_n18346);
not_10 g15998(new_n8525, new_n18347);
xor_4  g15999(new_n18307, new_n18291, new_n18348);
and_5  g16000(new_n18348, new_n18347, new_n18349);
xnor_4 g16001(new_n18348, new_n18347, new_n18350_1);
not_10 g16002(new_n8529, new_n18351);
xnor_4 g16003(new_n18304_1, new_n18293, new_n18352);
and_5  g16004(new_n18352, new_n18351, new_n18353);
xnor_4 g16005(new_n18352, new_n18351, new_n18354);
xor_4  g16006(new_n18302, new_n18301_1, new_n18355);
nor_5  g16007(new_n18355, new_n8533, new_n18356);
xnor_4 g16008(new_n18355, new_n8533, new_n18357);
xor_4  g16009(new_n18299, new_n9667, new_n18358);
and_5  g16010(new_n18358, new_n8536, new_n18359);
xnor_4 g16011(new_n9664, n18, new_n18360);
or_5   g16012(new_n18360, new_n8540, new_n18361);
not_10 g16013(new_n8536, new_n18362_1);
xnor_4 g16014(new_n18358, new_n18362_1, new_n18363);
and_5  g16015(new_n18363, new_n18361, new_n18364);
nor_5  g16016(new_n18364, new_n18359, new_n18365);
nor_5  g16017(new_n18365, new_n18357, new_n18366);
nor_5  g16018(new_n18366, new_n18356, new_n18367);
nor_5  g16019(new_n18367, new_n18354, new_n18368);
nor_5  g16020(new_n18368, new_n18353, new_n18369);
nor_5  g16021(new_n18369, new_n18350_1, new_n18370);
nor_5  g16022(new_n18370, new_n18349, new_n18371);
nor_5  g16023(new_n18371, new_n18346, new_n18372);
nor_5  g16024(new_n18372, new_n18345_1, new_n18373);
nor_5  g16025(new_n18373, new_n18342, new_n18374);
nor_5  g16026(new_n18374, new_n18341, new_n18375);
nor_5  g16027(new_n18375, new_n18338, new_n18376);
nor_5  g16028(new_n18376, new_n18337, new_n18377_1);
nor_5  g16029(new_n18377_1, new_n18335, new_n18378);
nor_5  g16030(new_n18378, new_n18334, new_n18379);
nor_5  g16031(new_n18379, new_n18332_1, new_n18380);
nor_5  g16032(new_n18380, new_n18331, new_n18381);
nor_5  g16033(new_n18381, new_n18329, new_n18382);
nor_5  g16034(new_n18382, new_n18328, new_n18383);
xnor_4 g16035(new_n18383, new_n17621, new_n18384);
xnor_4 g16036(new_n18384, new_n18325, n6628);
xnor_4 g16037(new_n2753, new_n2737, n6630);
xnor_4 g16038(n25331, n17911, new_n18387);
nor_5  g16039(n21997, n18483, new_n18388);
nor_5  g16040(new_n17707, new_n17700, new_n18389);
nor_5  g16041(new_n18389, new_n18388, new_n18390);
xor_4  g16042(new_n18390, new_n18387, new_n18391);
xnor_4 g16043(new_n18391, new_n6803, new_n18392);
nor_5  g16044(new_n17708, new_n6797, new_n18393);
nor_5  g16045(new_n17719, new_n17709, new_n18394);
nor_5  g16046(new_n18394, new_n18393, new_n18395);
xor_4  g16047(new_n18395, new_n18392, new_n18396);
xor_4  g16048(n14130, n468, new_n18397);
not_10 g16049(n5400, new_n18398);
nor_5  g16050(n16482, new_n18398, new_n18399);
xor_4  g16051(n16482, n5400, new_n18400);
nor_5  g16052(new_n15692, n9942, new_n18401);
nor_5  g16053(n25643, new_n15695, new_n18402);
xor_4  g16054(n25643, n329, new_n18403);
nor_5  g16055(new_n11977, n9557, new_n18404);
xor_4  g16056(n24170, n9557, new_n18405_1);
nor_5  g16057(new_n6942, n2409, new_n18406);
xor_4  g16058(n3136, n2409, new_n18407);
nor_5  g16059(n8869, new_n2359, new_n18408);
nor_5  g16060(new_n17328, new_n17325, new_n18409_1);
nor_5  g16061(new_n18409_1, new_n18408, new_n18410);
nor_5  g16062(new_n18410, new_n18407, new_n18411);
or_5   g16063(new_n18411, new_n18406, new_n18412);
nor_5  g16064(new_n18412, new_n18405_1, new_n18413);
nor_5  g16065(new_n18413, new_n18404, new_n18414_1);
nor_5  g16066(new_n18414_1, new_n18403, new_n18415);
nor_5  g16067(new_n18415, new_n18402, new_n18416);
xor_4  g16068(n23923, n9942, new_n18417);
nor_5  g16069(new_n18417, new_n18416, new_n18418_1);
nor_5  g16070(new_n18418_1, new_n18401, new_n18419);
nor_5  g16071(new_n18419, new_n18400, new_n18420);
nor_5  g16072(new_n18420, new_n18399, new_n18421);
xor_4  g16073(new_n18421, new_n18397, new_n18422);
xnor_4 g16074(new_n18422, new_n18396, new_n18423);
xor_4  g16075(new_n18419, new_n18400, new_n18424);
nor_5  g16076(new_n18424, new_n17720, new_n18425);
xor_4  g16077(new_n18424, new_n17720, new_n18426);
not_10 g16078(new_n17723, new_n18427);
xor_4  g16079(new_n18417, new_n18416, new_n18428);
and_5  g16080(new_n18428, new_n18427, new_n18429);
xor_4  g16081(new_n18414_1, new_n18403, new_n18430);
nor_5  g16082(new_n18430, new_n17366, new_n18431);
xnor_4 g16083(new_n18430, new_n17366, new_n18432);
not_10 g16084(new_n17388, new_n18433);
xor_4  g16085(new_n18412, new_n18405_1, new_n18434);
nor_5  g16086(new_n18434, new_n18433, new_n18435);
xor_4  g16087(new_n18434, new_n17388, new_n18436);
xor_4  g16088(new_n18410, new_n18407, new_n18437_1);
and_5  g16089(new_n18437_1, new_n17390, new_n18438);
xnor_4 g16090(new_n18437_1, new_n17390, new_n18439_1);
and_5  g16091(new_n17329, new_n17324, new_n18440);
and_5  g16092(new_n17334, new_n17330, new_n18441);
nor_5  g16093(new_n18441, new_n18440, new_n18442);
nor_5  g16094(new_n18442, new_n18439_1, new_n18443);
nor_5  g16095(new_n18443, new_n18438, new_n18444_1);
nor_5  g16096(new_n18444_1, new_n18436, new_n18445_1);
nor_5  g16097(new_n18445_1, new_n18435, new_n18446);
nor_5  g16098(new_n18446, new_n18432, new_n18447);
or_5   g16099(new_n18447, new_n18431, new_n18448);
xor_4  g16100(new_n18428, new_n17723, new_n18449);
nor_5  g16101(new_n18449, new_n18448, new_n18450);
nor_5  g16102(new_n18450, new_n18429, new_n18451);
and_5  g16103(new_n18451, new_n18426, new_n18452_1);
or_5   g16104(new_n18452_1, new_n18425, new_n18453);
xor_4  g16105(new_n18453, new_n18423, n6634);
xnor_4 g16106(new_n5975, new_n5963, n6652);
xnor_4 g16107(new_n11328, new_n11314, n6655);
xnor_4 g16108(new_n10862, new_n10843, n6669);
xnor_4 g16109(new_n8547, new_n8531, n6671);
xnor_4 g16110(new_n12221, new_n12203, n6673);
nor_5  g16111(new_n18181, new_n18175, new_n18460);
or_5   g16112(new_n10333, new_n13634, new_n18461);
nor_5  g16113(new_n18179, new_n18461, new_n18462);
or_5   g16114(new_n18462, new_n18460, n6674);
xnor_4 g16115(new_n15021, new_n15013, n6684);
xor_4  g16116(new_n11081, new_n11034, n6706);
xnor_4 g16117(n12702, n8614, new_n18466);
nor_5  g16118(n26797, n15182, new_n18467_1);
xnor_4 g16119(n26797, n15182, new_n18468);
nor_5  g16120(n27037, n23913, new_n18469);
xnor_4 g16121(n27037, n23913, new_n18470);
nor_5  g16122(n22554, n8964, new_n18471);
xnor_4 g16123(n22554, n8964, new_n18472);
nor_5  g16124(n20429, n20151, new_n18473);
xnor_4 g16125(n20429, n20151, new_n18474);
nor_5  g16126(n7693, n3909, new_n18475);
xnor_4 g16127(n7693, n3909, new_n18476);
nor_5  g16128(n23974, n10405, new_n18477);
xnor_4 g16129(n23974, n10405, new_n18478);
and_5  g16130(n11302, n2146, new_n18479);
or_5   g16131(n11302, n2146, new_n18480);
nor_5  g16132(n22173, n17090, new_n18481);
nor_5  g16133(new_n14174_1, new_n14173, new_n18482_1);
nor_5  g16134(new_n18482_1, new_n18481, new_n18483_1);
and_5  g16135(new_n18483_1, new_n18480, new_n18484);
or_5   g16136(new_n18484, new_n18479, new_n18485);
nor_5  g16137(new_n18485, new_n18478, new_n18486);
nor_5  g16138(new_n18486, new_n18477, new_n18487);
nor_5  g16139(new_n18487, new_n18476, new_n18488);
nor_5  g16140(new_n18488, new_n18475, new_n18489);
nor_5  g16141(new_n18489, new_n18474, new_n18490);
nor_5  g16142(new_n18490, new_n18473, new_n18491);
nor_5  g16143(new_n18491, new_n18472, new_n18492);
nor_5  g16144(new_n18492, new_n18471, new_n18493);
nor_5  g16145(new_n18493, new_n18470, new_n18494);
nor_5  g16146(new_n18494, new_n18469, new_n18495);
nor_5  g16147(new_n18495, new_n18468, new_n18496_1);
nor_5  g16148(new_n18496_1, new_n18467_1, new_n18497);
xor_4  g16149(new_n18497, new_n18466, new_n18498);
and_5  g16150(new_n18498, n1831, new_n18499);
xnor_4 g16151(new_n18498, n1831, new_n18500);
xor_4  g16152(new_n18495, new_n18468, new_n18501);
and_5  g16153(new_n18501, n13137, new_n18502);
xnor_4 g16154(new_n18501, n13137, new_n18503);
xor_4  g16155(new_n18493, new_n18470, new_n18504);
and_5  g16156(new_n18504, n18452, new_n18505);
xnor_4 g16157(new_n18504, n18452, new_n18506);
xor_4  g16158(new_n18491, new_n18472, new_n18507);
and_5  g16159(new_n18507, n21317, new_n18508);
xnor_4 g16160(new_n18507, n21317, new_n18509_1);
xor_4  g16161(new_n18489, new_n18474, new_n18510);
and_5  g16162(new_n18510, n12398, new_n18511);
xnor_4 g16163(new_n18510, n12398, new_n18512);
xor_4  g16164(new_n18487, new_n18476, new_n18513_1);
and_5  g16165(new_n18513_1, n19789, new_n18514);
xnor_4 g16166(new_n18513_1, n19789, new_n18515_1);
xor_4  g16167(new_n18485, new_n18478, new_n18516);
and_5  g16168(new_n18516, n20169, new_n18517);
xnor_4 g16169(new_n18516, n20169, new_n18518);
xor_4  g16170(n11302, n2146, new_n18519);
xnor_4 g16171(new_n18519, new_n18483_1, new_n18520);
and_5  g16172(new_n18520, n8285, new_n18521);
xnor_4 g16173(new_n18520, n8285, new_n18522);
nor_5  g16174(new_n14175, new_n14172, new_n18523);
nor_5  g16175(new_n18523, new_n14171, new_n18524);
nor_5  g16176(new_n18524, new_n18522, new_n18525);
nor_5  g16177(new_n18525, new_n18521, new_n18526);
nor_5  g16178(new_n18526, new_n18518, new_n18527);
nor_5  g16179(new_n18527, new_n18517, new_n18528);
nor_5  g16180(new_n18528, new_n18515_1, new_n18529);
nor_5  g16181(new_n18529, new_n18514, new_n18530);
nor_5  g16182(new_n18530, new_n18512, new_n18531);
nor_5  g16183(new_n18531, new_n18511, new_n18532);
nor_5  g16184(new_n18532, new_n18509_1, new_n18533);
nor_5  g16185(new_n18533, new_n18508, new_n18534);
nor_5  g16186(new_n18534, new_n18506, new_n18535);
nor_5  g16187(new_n18535, new_n18505, new_n18536);
nor_5  g16188(new_n18536, new_n18503, new_n18537_1);
nor_5  g16189(new_n18537_1, new_n18502, new_n18538);
nor_5  g16190(new_n18538, new_n18500, new_n18539);
nor_5  g16191(new_n18539, new_n18499, new_n18540);
nor_5  g16192(n12702, n8614, new_n18541);
nor_5  g16193(new_n18497, new_n18466, new_n18542);
nor_5  g16194(new_n18542, new_n18541, new_n18543);
xor_4  g16195(new_n18543, new_n18540, new_n18544);
and_5  g16196(new_n18215, new_n10495, new_n18545);
and_5  g16197(new_n18234, new_n18216, new_n18546);
nor_5  g16198(new_n18546, new_n18545, new_n18547);
not_10 g16199(n1536, new_n18548);
and_5  g16200(new_n18214, new_n18548, new_n18549);
xor_4  g16201(new_n18549, new_n4135, new_n18550);
xnor_4 g16202(new_n18550, new_n18547, new_n18551);
xnor_4 g16203(new_n18551, new_n18544, new_n18552);
not_10 g16204(new_n18235, new_n18553);
xor_4  g16205(new_n18538, new_n18500, new_n18554);
and_5  g16206(new_n18554, new_n18553, new_n18555);
xor_4  g16207(new_n18554, new_n18235, new_n18556);
xor_4  g16208(new_n18536, new_n18503, new_n18557);
and_5  g16209(new_n18557, new_n18255, new_n18558_1);
xnor_4 g16210(new_n18557, new_n18255, new_n18559);
xor_4  g16211(new_n18534, new_n18506, new_n18560);
and_5  g16212(new_n18560, new_n18259, new_n18561);
xnor_4 g16213(new_n18560, new_n18259, new_n18562);
xor_4  g16214(new_n18532, new_n18509_1, new_n18563);
and_5  g16215(new_n18563, new_n18263, new_n18564);
xnor_4 g16216(new_n18563, new_n18263, new_n18565);
xor_4  g16217(new_n18530, new_n18512, new_n18566);
and_5  g16218(new_n18566, new_n12348, new_n18567);
xnor_4 g16219(new_n18566, new_n12348, new_n18568);
xor_4  g16220(new_n18528, new_n18515_1, new_n18569);
and_5  g16221(new_n18569, new_n12371, new_n18570);
xnor_4 g16222(new_n18569, new_n12371, new_n18571);
xor_4  g16223(new_n18526, new_n18518, new_n18572_1);
and_5  g16224(new_n18572_1, new_n12374, new_n18573);
xor_4  g16225(new_n18572_1, new_n12374, new_n18574_1);
xnor_4 g16226(new_n12340, new_n12334, new_n18575);
xor_4  g16227(new_n18524, new_n18522, new_n18576_1);
nor_5  g16228(new_n18576_1, new_n18575, new_n18577);
and_5  g16229(new_n14176, new_n12383_1, new_n18578_1);
and_5  g16230(new_n14177, new_n14167, new_n18579);
or_5   g16231(new_n18579, new_n18578_1, new_n18580);
xnor_4 g16232(new_n18576_1, new_n18575, new_n18581);
nor_5  g16233(new_n18581, new_n18580, new_n18582_1);
nor_5  g16234(new_n18582_1, new_n18577, new_n18583_1);
and_5  g16235(new_n18583_1, new_n18574_1, new_n18584_1);
nor_5  g16236(new_n18584_1, new_n18573, new_n18585);
nor_5  g16237(new_n18585, new_n18571, new_n18586);
nor_5  g16238(new_n18586, new_n18570, new_n18587);
nor_5  g16239(new_n18587, new_n18568, new_n18588);
nor_5  g16240(new_n18588, new_n18567, new_n18589);
nor_5  g16241(new_n18589, new_n18565, new_n18590);
nor_5  g16242(new_n18590, new_n18564, new_n18591);
nor_5  g16243(new_n18591, new_n18562, new_n18592);
nor_5  g16244(new_n18592, new_n18561, new_n18593);
nor_5  g16245(new_n18593, new_n18559, new_n18594);
nor_5  g16246(new_n18594, new_n18558_1, new_n18595);
nor_5  g16247(new_n18595, new_n18556, new_n18596);
nor_5  g16248(new_n18596, new_n18555, new_n18597);
xnor_4 g16249(new_n18597, new_n18552, n6707);
xor_4  g16250(new_n11810, new_n11592, n6736);
xor_4  g16251(n23895, n5101, new_n18600);
and_5  g16252(new_n5027, n16507, new_n18601);
xor_4  g16253(n17351, n16507, new_n18602);
and_5  g16254(n22470, new_n5030, new_n18603);
xor_4  g16255(n22470, n11736, new_n18604);
and_5  g16256(new_n5033, n19116, new_n18605);
and_5  g16257(new_n5036, n6861, new_n18606);
nor_5  g16258(new_n16273, new_n16256, new_n18607);
nor_5  g16259(new_n18607, new_n18606, new_n18608);
xor_4  g16260(n23200, n19116, new_n18609);
nor_5  g16261(new_n18609, new_n18608, new_n18610_1);
nor_5  g16262(new_n18610_1, new_n18605, new_n18611);
nor_5  g16263(new_n18611, new_n18604, new_n18612);
nor_5  g16264(new_n18612, new_n18603, new_n18613);
nor_5  g16265(new_n18613, new_n18602, new_n18614);
nor_5  g16266(new_n18614, new_n18601, new_n18615);
xor_4  g16267(new_n18615, new_n18600, new_n18616);
not_10 g16268(n12650, new_n18617);
and_5  g16269(new_n16280, new_n5083, new_n18618);
and_5  g16270(new_n18618, new_n5080, new_n18619);
and_5  g16271(new_n18619, new_n5077_1, new_n18620);
and_5  g16272(new_n18620, new_n5074, new_n18621);
xnor_4 g16273(new_n18621, n13494, new_n18622);
xnor_4 g16274(new_n18622, new_n18617, new_n18623);
not_10 g16275(n10201, new_n18624);
xnor_4 g16276(new_n18620, n25345, new_n18625);
nor_5  g16277(new_n18625, new_n18624, new_n18626);
xnor_4 g16278(new_n18625, new_n18624, new_n18627);
xnor_4 g16279(new_n18619, new_n5077_1, new_n18628);
and_5  g16280(new_n18628, n10593, new_n18629);
xnor_4 g16281(new_n18628, n10593, new_n18630);
not_10 g16282(n18290, new_n18631);
xnor_4 g16283(new_n18618, n13490, new_n18632);
nor_5  g16284(new_n18632, new_n18631, new_n18633);
xnor_4 g16285(new_n18632, new_n18631, new_n18634);
nor_5  g16286(new_n16281, new_n16275_1, new_n18635_1);
nor_5  g16287(new_n16305, new_n16282, new_n18636);
nor_5  g16288(new_n18636, new_n18635_1, new_n18637);
nor_5  g16289(new_n18637, new_n18634, new_n18638);
nor_5  g16290(new_n18638, new_n18633, new_n18639);
nor_5  g16291(new_n18639, new_n18630, new_n18640);
nor_5  g16292(new_n18640, new_n18629, new_n18641);
nor_5  g16293(new_n18641, new_n18627, new_n18642);
nor_5  g16294(new_n18642, new_n18626, new_n18643);
xor_4  g16295(new_n18643, new_n18623, new_n18644);
xnor_4 g16296(new_n18644, new_n14384, new_n18645);
xor_4  g16297(new_n18641, new_n18627, new_n18646);
nor_5  g16298(new_n18646, new_n14386, new_n18647);
xor_4  g16299(new_n18639, new_n18630, new_n18648);
nand_5 g16300(new_n18648, new_n14389, new_n18649_1);
xnor_4 g16301(new_n18648, new_n14389, new_n18650);
xor_4  g16302(new_n18637, new_n18634, new_n18651);
nor_5  g16303(new_n18651, new_n14392, new_n18652);
xnor_4 g16304(new_n18651, new_n14392, new_n18653_1);
nor_5  g16305(new_n16306, new_n14395, new_n18654);
nor_5  g16306(new_n16329, new_n16307, new_n18655);
nor_5  g16307(new_n18655, new_n18654, new_n18656);
nor_5  g16308(new_n18656, new_n18653_1, new_n18657);
nor_5  g16309(new_n18657, new_n18652, new_n18658);
not_10 g16310(new_n18658, new_n18659);
or_5   g16311(new_n18659, new_n18650, new_n18660);
nand_5 g16312(new_n18660, new_n18649_1, new_n18661);
xnor_4 g16313(new_n18646, new_n14386, new_n18662);
nor_5  g16314(new_n18662, new_n18661, new_n18663);
nor_5  g16315(new_n18663, new_n18647, new_n18664);
xor_4  g16316(new_n18664, new_n18645, new_n18665);
xnor_4 g16317(new_n18665, new_n18616, new_n18666);
xor_4  g16318(new_n18613, new_n18602, new_n18667);
xor_4  g16319(new_n18662, new_n18661, new_n18668);
nor_5  g16320(new_n18668, new_n18667, new_n18669);
xnor_4 g16321(new_n18668, new_n18667, new_n18670);
xor_4  g16322(new_n18611, new_n18604, new_n18671);
xnor_4 g16323(new_n18658, new_n18650, new_n18672);
not_10 g16324(new_n18672, new_n18673);
nor_5  g16325(new_n18673, new_n18671, new_n18674);
xnor_4 g16326(new_n18672, new_n18671, new_n18675);
xnor_4 g16327(new_n18609, new_n18608, new_n18676);
xor_4  g16328(new_n18656, new_n18653_1, new_n18677);
not_10 g16329(new_n18677, new_n18678);
nor_5  g16330(new_n18678, new_n18676, new_n18679_1);
xor_4  g16331(new_n18677, new_n18676, new_n18680);
and_5  g16332(new_n16330, new_n16274, new_n18681);
nor_5  g16333(new_n16361, new_n16331, new_n18682);
nor_5  g16334(new_n18682, new_n18681, new_n18683);
nor_5  g16335(new_n18683, new_n18680, new_n18684);
nor_5  g16336(new_n18684, new_n18679_1, new_n18685);
and_5  g16337(new_n18685, new_n18675, new_n18686);
nor_5  g16338(new_n18686, new_n18674, new_n18687);
nor_5  g16339(new_n18687, new_n18670, new_n18688);
or_5   g16340(new_n18688, new_n18669, new_n18689);
xor_4  g16341(new_n18689, new_n18666, n6791);
xnor_4 g16342(new_n3502_1, new_n3493, n6802);
xnor_4 g16343(new_n14725, new_n14701_1, n6826);
xnor_4 g16344(new_n9082, new_n9060, n6835);
and_5  g16345(new_n16556, n11220, new_n18694);
xnor_4 g16346(new_n16556, n11220, new_n18695);
and_5  g16347(new_n2838, n22379, new_n18696);
xnor_4 g16348(new_n2838, n22379, new_n18697);
and_5  g16349(new_n2871, n1662, new_n18698);
xnor_4 g16350(new_n2871, n1662, new_n18699);
and_5  g16351(new_n2875, n12875, new_n18700);
xnor_4 g16352(new_n2875, n12875, new_n18701);
and_5  g16353(new_n2879, n2035, new_n18702);
nor_5  g16354(new_n2883, n5213, new_n18703);
xnor_4 g16355(new_n2883, n5213, new_n18704);
nor_5  g16356(new_n2887_1, n4665, new_n18705);
xor_4  g16357(new_n2887_1, n4665, new_n18706);
and_5  g16358(new_n2891, n19005, new_n18707);
xnor_4 g16359(new_n2891, n19005, new_n18708_1);
and_5  g16360(new_n2898, n5438, new_n18709);
nor_5  g16361(new_n18709, n4326, new_n18710);
xnor_4 g16362(new_n18709, n4326, new_n18711);
nor_5  g16363(new_n18711, new_n2895, new_n18712);
or_5   g16364(new_n18712, new_n18710, new_n18713);
nor_5  g16365(new_n18713, new_n18708_1, new_n18714);
nor_5  g16366(new_n18714, new_n18707, new_n18715);
and_5  g16367(new_n18715, new_n18706, new_n18716);
nor_5  g16368(new_n18716, new_n18705, new_n18717);
nor_5  g16369(new_n18717, new_n18704, new_n18718);
or_5   g16370(new_n18718, new_n18703, new_n18719);
xnor_4 g16371(new_n2879, n2035, new_n18720);
nor_5  g16372(new_n18720, new_n18719, new_n18721_1);
nor_5  g16373(new_n18721_1, new_n18702, new_n18722);
nor_5  g16374(new_n18722, new_n18701, new_n18723);
nor_5  g16375(new_n18723, new_n18700, new_n18724);
nor_5  g16376(new_n18724, new_n18699, new_n18725_1);
nor_5  g16377(new_n18725_1, new_n18698, new_n18726);
nor_5  g16378(new_n18726, new_n18697, new_n18727);
nor_5  g16379(new_n18727, new_n18696, new_n18728);
nor_5  g16380(new_n18728, new_n18695, new_n18729);
nor_5  g16381(new_n18729, new_n18694, new_n18730);
nor_5  g16382(new_n18730, new_n16552, new_n18731);
xor_4  g16383(new_n18731, new_n16239, new_n18732);
not_10 g16384(new_n16241, new_n18733);
xor_4  g16385(new_n18730, new_n16552, new_n18734);
nor_5  g16386(new_n18734, new_n18733, new_n18735);
xor_4  g16387(new_n18734, new_n16241, new_n18736);
xor_4  g16388(new_n18728, new_n18695, new_n18737_1);
nor_5  g16389(new_n18737_1, new_n16244, new_n18738);
xor_4  g16390(new_n18737_1, new_n5570, new_n18739);
xor_4  g16391(new_n18726, new_n18697, new_n18740);
nor_5  g16392(new_n18740, new_n11638, new_n18741);
xor_4  g16393(new_n18740, new_n5572, new_n18742);
not_10 g16394(new_n5577, new_n18743);
xor_4  g16395(new_n18724, new_n18699, new_n18744);
nor_5  g16396(new_n18744, new_n18743, new_n18745_1);
xor_4  g16397(new_n18744, new_n5577, new_n18746);
xor_4  g16398(new_n18722, new_n18701, new_n18747);
nor_5  g16399(new_n18747, new_n11644, new_n18748);
xor_4  g16400(new_n18747, new_n5581, new_n18749);
not_10 g16401(new_n5585, new_n18750);
xor_4  g16402(new_n18720, new_n18719, new_n18751_1);
nor_5  g16403(new_n18751_1, new_n18750, new_n18752);
xor_4  g16404(new_n18751_1, new_n5585, new_n18753);
xor_4  g16405(new_n18717, new_n18704, new_n18754);
and_5  g16406(new_n18754, new_n5589, new_n18755);
xnor_4 g16407(new_n18754, new_n5589, new_n18756);
xor_4  g16408(new_n18715, new_n18706, new_n18757);
and_5  g16409(new_n18757, new_n5593_1, new_n18758);
xnor_4 g16410(new_n18757, new_n5593_1, new_n18759);
xor_4  g16411(new_n18713, new_n18708_1, new_n18760);
nor_5  g16412(new_n18760, new_n5599, new_n18761);
xor_4  g16413(new_n18760, new_n5597, new_n18762);
xor_4  g16414(new_n18711, new_n2895, new_n18763);
and_5  g16415(new_n18763, new_n11655, new_n18764);
and_5  g16416(new_n5331, new_n5330_1, new_n18765);
xnor_4 g16417(new_n18763, new_n5601, new_n18766);
and_5  g16418(new_n18766, new_n18765, new_n18767);
nor_5  g16419(new_n18767, new_n18764, new_n18768);
nor_5  g16420(new_n18768, new_n18762, new_n18769);
nor_5  g16421(new_n18769, new_n18761, new_n18770);
nor_5  g16422(new_n18770, new_n18759, new_n18771);
nor_5  g16423(new_n18771, new_n18758, new_n18772);
nor_5  g16424(new_n18772, new_n18756, new_n18773);
nor_5  g16425(new_n18773, new_n18755, new_n18774);
nor_5  g16426(new_n18774, new_n18753, new_n18775);
nor_5  g16427(new_n18775, new_n18752, new_n18776);
nor_5  g16428(new_n18776, new_n18749, new_n18777);
nor_5  g16429(new_n18777, new_n18748, new_n18778);
nor_5  g16430(new_n18778, new_n18746, new_n18779);
nor_5  g16431(new_n18779, new_n18745_1, new_n18780_1);
nor_5  g16432(new_n18780_1, new_n18742, new_n18781);
nor_5  g16433(new_n18781, new_n18741, new_n18782_1);
nor_5  g16434(new_n18782_1, new_n18739, new_n18783);
nor_5  g16435(new_n18783, new_n18738, new_n18784);
nor_5  g16436(new_n18784, new_n18736, new_n18785);
nor_5  g16437(new_n18785, new_n18735, new_n18786);
xnor_4 g16438(new_n18786, new_n18732, n6853);
xor_4  g16439(new_n10022, new_n9989, new_n18788);
xnor_4 g16440(new_n13466, new_n18788, new_n18789);
nor_5  g16441(new_n13470, new_n10052, new_n18790);
xnor_4 g16442(new_n13470, new_n10052, new_n18791);
nor_5  g16443(new_n10056, new_n11679, new_n18792);
nor_5  g16444(new_n11694, new_n11680, new_n18793);
or_5   g16445(new_n18793, new_n18792, new_n18794);
nor_5  g16446(new_n18794, new_n18791, new_n18795);
nor_5  g16447(new_n18795, new_n18790, new_n18796);
xor_4  g16448(new_n18796, new_n18789, n6862);
not_10 g16449(n22253, new_n18798);
nor_5  g16450(new_n18798, n8305, new_n18799);
nor_5  g16451(new_n14342_1, new_n14323_1, new_n18800);
nor_5  g16452(new_n18800, new_n18799, new_n18801);
not_10 g16453(n25296, new_n18802_1);
nor_5  g16454(new_n18802_1, n23717, new_n18803);
nor_5  g16455(new_n10209, new_n10195, new_n18804);
nor_5  g16456(new_n18804, new_n18803, new_n18805);
nor_5  g16457(new_n18805, new_n16705, new_n18806);
and_5  g16458(new_n10210, new_n10194, new_n18807);
nor_5  g16459(new_n10232, new_n10211, new_n18808);
nor_5  g16460(new_n18808, new_n18807, new_n18809);
xnor_4 g16461(new_n18805, new_n16705, new_n18810);
nor_5  g16462(new_n18810, new_n18809, new_n18811);
nor_5  g16463(new_n18811, new_n18806, new_n18812);
and_5  g16464(new_n18812, new_n18801, new_n18813);
and_5  g16465(new_n14343, new_n14322, new_n18814);
nor_5  g16466(new_n14362, new_n14344, new_n18815);
nor_5  g16467(new_n18815, new_n18814, new_n18816);
nor_5  g16468(new_n18816, new_n18812, new_n18817);
or_5   g16469(new_n18817, new_n18813, new_n18818);
xor_4  g16470(new_n18810, new_n18809, new_n18819);
nor_5  g16471(new_n18819, new_n18801, new_n18820);
or_5   g16472(new_n18815, new_n18814, new_n18821);
xnor_4 g16473(new_n18810, new_n18809, new_n18822);
nor_5  g16474(new_n18822, new_n18821, new_n18823);
or_5   g16475(new_n18823, new_n18820, new_n18824);
nor_5  g16476(new_n18824, new_n18818, n6863);
xnor_4 g16477(new_n5620, new_n5575, n6867);
xnor_4 g16478(new_n16193, new_n16186, n6965);
xnor_4 g16479(new_n6734, new_n6699, n6967);
xor_4  g16480(new_n13043_1, new_n13003, n6975);
xor_4  g16481(new_n18156, new_n18155, n6983);
xnor_4 g16482(new_n13448, new_n10038, new_n18831_1);
nor_5  g16483(new_n13453_1, new_n10040, new_n18832);
xnor_4 g16484(new_n13453_1, new_n10040, new_n18833);
nor_5  g16485(new_n13456_1, new_n10043, new_n18834);
xor_4  g16486(new_n13456_1, new_n10043, new_n18835);
and_5  g16487(new_n13461, new_n10046, new_n18836);
nor_5  g16488(new_n13466, new_n18788, new_n18837);
nor_5  g16489(new_n18796, new_n18789, new_n18838);
nor_5  g16490(new_n18838, new_n18837, new_n18839);
xnor_4 g16491(new_n13461, new_n10046, new_n18840);
nor_5  g16492(new_n18840, new_n18839, new_n18841);
nor_5  g16493(new_n18841, new_n18836, new_n18842);
and_5  g16494(new_n18842, new_n18835, new_n18843_1);
nor_5  g16495(new_n18843_1, new_n18834, new_n18844);
nor_5  g16496(new_n18844, new_n18833, new_n18845);
nor_5  g16497(new_n18845, new_n18832, new_n18846);
xnor_4 g16498(new_n18846, new_n18831_1, n6985);
xnor_4 g16499(new_n13283, new_n13244, n6998);
xor_4  g16500(new_n10005, new_n8080, n7032);
xnor_4 g16501(new_n18021, new_n17989, n7038);
xnor_4 g16502(new_n16027, new_n16026, n7079);
xnor_4 g16503(new_n6723, new_n6722, n7190);
xnor_4 g16504(new_n14294_1, new_n14290, n7229);
xnor_4 g16505(new_n7787, new_n7776, n7230);
xnor_4 g16506(new_n17302_1, new_n17301, n7233);
xnor_4 g16507(new_n11913, new_n11905_1, n7236);
xor_4  g16508(new_n14621, new_n6288, n7253);
and_5  g16509(new_n17653, new_n6526, new_n18858_1);
or_5   g16510(new_n17654, n12507, new_n18859_1);
and_5  g16511(new_n17654, n12507, new_n18860);
or_5   g16512(new_n17658, new_n18860, new_n18861);
and_5  g16513(new_n18861, new_n18859_1, new_n18862);
or_5   g16514(new_n18862, new_n18858_1, new_n18863);
not_10 g16515(new_n9166_1, new_n18864_1);
or_5   g16516(new_n18088, new_n12735, new_n18865_1);
xor_4  g16517(new_n18865_1, new_n12732, new_n18866);
nor_5  g16518(new_n18866, new_n18864_1, new_n18867);
xor_4  g16519(new_n18866, new_n9166_1, new_n18868);
nor_5  g16520(new_n18089, new_n9168, new_n18869);
nor_5  g16521(new_n18131, new_n18090, new_n18870);
nor_5  g16522(new_n18870, new_n18869, new_n18871);
nor_5  g16523(new_n18871, new_n18868, new_n18872);
or_5   g16524(new_n18872, new_n18867, new_n18873);
or_5   g16525(new_n18865_1, new_n12732, new_n18874);
and_5  g16526(new_n18874, new_n12774, new_n18875);
nor_5  g16527(new_n18874, new_n12772, new_n18876);
nor_5  g16528(new_n18876, new_n18875, new_n18877);
xnor_4 g16529(new_n18877, new_n9160, new_n18878);
xnor_4 g16530(new_n18878, new_n18873, new_n18879);
and_5  g16531(new_n18879, new_n18863, new_n18880_1);
nor_5  g16532(new_n18862, new_n18858_1, new_n18881);
xnor_4 g16533(new_n18879, new_n18881, new_n18882);
xor_4  g16534(new_n18871, new_n18868, new_n18883);
nor_5  g16535(new_n18883, new_n17659, new_n18884);
nor_5  g16536(new_n18132, new_n15081, new_n18885);
nor_5  g16537(new_n18171_1, new_n18133, new_n18886_1);
nor_5  g16538(new_n18886_1, new_n18885, new_n18887_1);
xnor_4 g16539(new_n18883, new_n17659, new_n18888);
nor_5  g16540(new_n18888, new_n18887_1, new_n18889);
nor_5  g16541(new_n18889, new_n18884, new_n18890);
and_5  g16542(new_n18890, new_n18882, new_n18891);
nor_5  g16543(new_n18891, new_n18880_1, new_n18892);
and_5  g16544(new_n18877, new_n9160, new_n18893);
nor_5  g16545(new_n18877, new_n9160, new_n18894);
nor_5  g16546(new_n18894, new_n18873, new_n18895);
or_5   g16547(new_n18895, new_n18876, new_n18896);
or_5   g16548(new_n18896, new_n18893, new_n18897);
xnor_4 g16549(new_n18897, new_n18892, n7256);
nor_5  g16550(new_n7204, n2416, new_n18899);
xor_4  g16551(n22764, n2416, new_n18900);
nor_5  g16552(new_n7242, n21905, new_n18901_1);
nor_5  g16553(new_n17751, new_n17740, new_n18902);
nor_5  g16554(new_n18902, new_n18901_1, new_n18903);
nor_5  g16555(new_n18903, new_n18900, new_n18904);
nor_5  g16556(new_n18904, new_n18899, new_n18905);
xor_4  g16557(new_n18903, new_n18900, new_n18906);
and_5  g16558(new_n18906, new_n14013, new_n18907_1);
xnor_4 g16559(new_n18906, new_n14013, new_n18908);
and_5  g16560(new_n17752, new_n14017, new_n18909);
nor_5  g16561(new_n17766, new_n17753, new_n18910);
nor_5  g16562(new_n18910, new_n18909, new_n18911);
nor_5  g16563(new_n18911, new_n18908, new_n18912);
nor_5  g16564(new_n18912, new_n18907_1, new_n18913);
xor_4  g16565(new_n18913, new_n18905, new_n18914);
xnor_4 g16566(new_n18914, new_n14010, new_n18915);
xnor_4 g16567(new_n18915, new_n17855_1, new_n18916);
xor_4  g16568(new_n18911, new_n18908, new_n18917);
nor_5  g16569(new_n18917, new_n17867, new_n18918);
xnor_4 g16570(new_n18917, new_n17867, new_n18919_1);
nor_5  g16571(new_n17767, new_n17739, new_n18920);
nor_5  g16572(new_n17781, new_n17768, new_n18921);
nor_5  g16573(new_n18921, new_n18920, new_n18922);
nor_5  g16574(new_n18922, new_n18919_1, new_n18923);
nor_5  g16575(new_n18923, new_n18918, new_n18924);
xnor_4 g16576(new_n18924, new_n18916, n7268);
not_10 g16577(new_n9822, new_n18926_1);
or_5   g16578(new_n18926_1, n752, new_n18927);
or_5   g16579(new_n18927, n2175, new_n18928);
or_5   g16580(new_n18928, n13026, new_n18929);
nor_5  g16581(new_n18929, n23912, new_n18930);
nor_5  g16582(new_n18928, n13026, new_n18931);
xor_4  g16583(new_n18931, n23912, new_n18932);
and_5  g16584(new_n18932, n10514, new_n18933);
xnor_4 g16585(new_n18932, n10514, new_n18934);
nor_5  g16586(new_n18927, n2175, new_n18935);
xor_4  g16587(new_n18935, n13026, new_n18936);
and_5  g16588(new_n18936, n18649, new_n18937);
xnor_4 g16589(new_n18936, n18649, new_n18938);
nor_5  g16590(new_n18926_1, n752, new_n18939);
xor_4  g16591(new_n18939, n2175, new_n18940_1);
and_5  g16592(new_n18940_1, n6218, new_n18941);
xnor_4 g16593(new_n18940_1, n6218, new_n18942);
not_10 g16594(new_n9823, new_n18943);
and_5  g16595(new_n18943, n20470, new_n18944);
xor_4  g16596(new_n9823, n20470, new_n18945_1);
not_10 g16597(n21222, new_n18946);
nor_5  g16598(new_n9826, new_n18946, new_n18947);
xnor_4 g16599(new_n9826, new_n18946, new_n18948);
and_5  g16600(new_n9829, n9832, new_n18949);
xnor_4 g16601(new_n9829, n9832, new_n18950);
and_5  g16602(new_n9834, n1558, new_n18951);
xor_4  g16603(new_n9833_1, n1558, new_n18952);
xnor_4 g16604(new_n9817, n5131, new_n18953);
and_5  g16605(new_n18953, n21749, new_n18954);
xnor_4 g16606(new_n18953, n21749, new_n18955);
and_5  g16607(new_n9840, n7769, new_n18956);
not_10 g16608(n21138, new_n18957);
nor_5  g16609(new_n18957, n15506, new_n18958);
xor_4  g16610(new_n9840, n7769, new_n18959);
and_5  g16611(new_n18959, new_n18958, new_n18960);
nor_5  g16612(new_n18960, new_n18956, new_n18961);
nor_5  g16613(new_n18961, new_n18955, new_n18962_1);
nor_5  g16614(new_n18962_1, new_n18954, new_n18963);
nor_5  g16615(new_n18963, new_n18952, new_n18964);
nor_5  g16616(new_n18964, new_n18951, new_n18965);
nor_5  g16617(new_n18965, new_n18950, new_n18966);
nor_5  g16618(new_n18966, new_n18949, new_n18967);
nor_5  g16619(new_n18967, new_n18948, new_n18968);
nor_5  g16620(new_n18968, new_n18947, new_n18969);
nor_5  g16621(new_n18969, new_n18945_1, new_n18970_1);
nor_5  g16622(new_n18970_1, new_n18944, new_n18971);
nor_5  g16623(new_n18971, new_n18942, new_n18972);
nor_5  g16624(new_n18972, new_n18941, new_n18973);
nor_5  g16625(new_n18973, new_n18938, new_n18974);
nor_5  g16626(new_n18974, new_n18937, new_n18975);
nor_5  g16627(new_n18975, new_n18934, new_n18976);
nor_5  g16628(new_n18976, new_n18933, new_n18977_1);
nand_5 g16629(new_n18977_1, new_n18930, new_n18978);
xor_4  g16630(new_n18975, new_n18934, new_n18979);
nor_5  g16631(new_n18979, n9872, new_n18980);
xnor_4 g16632(new_n18979, n9872, new_n18981);
xor_4  g16633(new_n18973, new_n18938, new_n18982_1);
nor_5  g16634(new_n18982_1, n5842, new_n18983);
xnor_4 g16635(new_n18982_1, n5842, new_n18984);
xor_4  g16636(new_n18971, new_n18942, new_n18985);
nor_5  g16637(new_n18985, n6379, new_n18986);
xnor_4 g16638(new_n18985, n6379, new_n18987);
xor_4  g16639(new_n18969, new_n18945_1, new_n18988);
nor_5  g16640(new_n18988, n2102, new_n18989);
xnor_4 g16641(new_n18988, n2102, new_n18990);
xor_4  g16642(new_n18967, new_n18948, new_n18991);
nor_5  g16643(new_n18991, n17954, new_n18992);
xor_4  g16644(new_n18965, new_n18950, new_n18993);
nor_5  g16645(new_n18993, n8256, new_n18994);
xnor_4 g16646(new_n18993, n8256, new_n18995);
xor_4  g16647(new_n18963, new_n18952, new_n18996);
nor_5  g16648(new_n18996, n24150, new_n18997);
xnor_4 g16649(new_n18996, n24150, new_n18998);
xor_4  g16650(new_n18961, new_n18955, new_n18999_1);
nor_5  g16651(new_n18999_1, n19584, new_n19000);
xnor_4 g16652(new_n18999_1, n19584, new_n19001);
xor_4  g16653(new_n18959, new_n18958, new_n19002);
and_5  g16654(new_n19002, n5060, new_n19003);
nor_5  g16655(new_n19002, n5060, new_n19004);
xnor_4 g16656(n21138, n15506, new_n19005_1);
nand_5 g16657(new_n19005_1, n15332, new_n19006);
nor_5  g16658(new_n19006, new_n19004, new_n19007);
or_5   g16659(new_n19007, new_n19003, new_n19008);
nor_5  g16660(new_n19008, new_n19001, new_n19009);
nor_5  g16661(new_n19009, new_n19000, new_n19010);
nor_5  g16662(new_n19010, new_n18998, new_n19011);
nor_5  g16663(new_n19011, new_n18997, new_n19012);
nor_5  g16664(new_n19012, new_n18995, new_n19013);
nor_5  g16665(new_n19013, new_n18994, new_n19014);
xnor_4 g16666(new_n18991, n17954, new_n19015);
nor_5  g16667(new_n19015, new_n19014, new_n19016);
nor_5  g16668(new_n19016, new_n18992, new_n19017);
nor_5  g16669(new_n19017, new_n18990, new_n19018);
nor_5  g16670(new_n19018, new_n18989, new_n19019);
nor_5  g16671(new_n19019, new_n18987, new_n19020);
nor_5  g16672(new_n19020, new_n18986, new_n19021);
nor_5  g16673(new_n19021, new_n18984, new_n19022);
nor_5  g16674(new_n19022, new_n18983, new_n19023);
nor_5  g16675(new_n19023, new_n18981, new_n19024);
nor_5  g16676(new_n19024, new_n18980, new_n19025);
nor_5  g16677(new_n19025, new_n18978, new_n19026);
nor_5  g16678(new_n18977_1, new_n18930, new_n19027);
and_5  g16679(new_n19027, new_n19025, new_n19028);
nor_5  g16680(new_n19028, new_n19026, new_n19029);
xnor_4 g16681(new_n19029, new_n13232, new_n19030);
xnor_4 g16682(new_n18977_1, new_n18930, new_n19031);
xnor_4 g16683(new_n19031, new_n19025, new_n19032);
nor_5  g16684(new_n19032, new_n13235, new_n19033_1);
xnor_4 g16685(new_n19032, new_n13235, new_n19034);
xor_4  g16686(new_n19023, new_n18981, new_n19035);
nor_5  g16687(new_n19035, new_n14291, new_n19036);
xnor_4 g16688(new_n19035, new_n14291, new_n19037);
xor_4  g16689(new_n19021, new_n18984, new_n19038);
nor_5  g16690(new_n19038, new_n2712, new_n19039);
xor_4  g16691(new_n2608, new_n2574, new_n19040);
xor_4  g16692(new_n19019, new_n18987, new_n19041);
nor_5  g16693(new_n19041, new_n19040, new_n19042_1);
xnor_4 g16694(new_n19041, new_n19040, new_n19043);
xor_4  g16695(new_n19017, new_n18990, new_n19044_1);
nor_5  g16696(new_n19044_1, new_n2724, new_n19045);
xnor_4 g16697(new_n19044_1, new_n2724, new_n19046);
xnor_4 g16698(new_n2603, new_n2579, new_n19047);
xor_4  g16699(new_n19015, new_n19014, new_n19048);
nor_5  g16700(new_n19048, new_n19047, new_n19049);
xnor_4 g16701(new_n19048, new_n19047, new_n19050);
xor_4  g16702(new_n19012, new_n18995, new_n19051);
nor_5  g16703(new_n19051, new_n13254, new_n19052);
xnor_4 g16704(new_n19051, new_n13254, new_n19053);
xor_4  g16705(new_n19010, new_n18998, new_n19054);
nor_5  g16706(new_n19054, new_n2735, new_n19055);
xnor_4 g16707(new_n19054, new_n2735, new_n19056);
xor_4  g16708(new_n19008, new_n19001, new_n19057);
nor_5  g16709(new_n19057, new_n2739, new_n19058);
xnor_4 g16710(new_n19057, new_n2739, new_n19059);
xor_4  g16711(new_n19002, n5060, new_n19060);
xnor_4 g16712(new_n19060, new_n19006, new_n19061);
and_5  g16713(new_n19061, new_n2743_1, new_n19062);
xor_4  g16714(new_n19005_1, n15332, new_n19063);
or_5   g16715(new_n19063, new_n2746, new_n19064);
xnor_4 g16716(new_n19061, new_n2744, new_n19065);
and_5  g16717(new_n19065, new_n19064, new_n19066);
nor_5  g16718(new_n19066, new_n19062, new_n19067);
nor_5  g16719(new_n19067, new_n19059, new_n19068);
nor_5  g16720(new_n19068, new_n19058, new_n19069);
nor_5  g16721(new_n19069, new_n19056, new_n19070);
nor_5  g16722(new_n19070, new_n19055, new_n19071);
nor_5  g16723(new_n19071, new_n19053, new_n19072);
nor_5  g16724(new_n19072, new_n19052, new_n19073);
nor_5  g16725(new_n19073, new_n19050, new_n19074);
nor_5  g16726(new_n19074, new_n19049, new_n19075);
nor_5  g16727(new_n19075, new_n19046, new_n19076);
nor_5  g16728(new_n19076, new_n19045, new_n19077);
nor_5  g16729(new_n19077, new_n19043, new_n19078);
nor_5  g16730(new_n19078, new_n19042_1, new_n19079);
xnor_4 g16731(new_n19038, new_n2712, new_n19080);
nor_5  g16732(new_n19080, new_n19079, new_n19081_1);
nor_5  g16733(new_n19081_1, new_n19039, new_n19082);
nor_5  g16734(new_n19082, new_n19037, new_n19083);
nor_5  g16735(new_n19083, new_n19036, new_n19084);
nor_5  g16736(new_n19084, new_n19034, new_n19085);
nor_5  g16737(new_n19085, new_n19033_1, new_n19086);
xnor_4 g16738(new_n19086, new_n19030, n7277);
xor_4  g16739(new_n12062, new_n12055, n7280);
xnor_4 g16740(new_n5294, new_n5271, n7298);
xnor_4 g16741(new_n17643, new_n17634, n7308);
xnor_4 g16742(new_n17864, new_n6573, new_n19091);
and_5  g16743(new_n17866, new_n6590_1, new_n19092);
xnor_4 g16744(new_n17866, new_n6590_1, new_n19093);
and_5  g16745(new_n13512, new_n6594, new_n19094);
nor_5  g16746(new_n13537, new_n13513, new_n19095);
nor_5  g16747(new_n19095, new_n19094, new_n19096);
nor_5  g16748(new_n19096, new_n19093, new_n19097);
nor_5  g16749(new_n19097, new_n19092, new_n19098);
xnor_4 g16750(new_n19098, new_n19091, new_n19099);
xnor_4 g16751(new_n19099, new_n17889_1, new_n19100);
xor_4  g16752(new_n17887, new_n17883, new_n19101);
xor_4  g16753(new_n19096, new_n19093, new_n19102);
nor_5  g16754(new_n19102, new_n19101, new_n19103);
and_5  g16755(new_n17278, new_n13538, new_n19104);
nor_5  g16756(new_n17310, new_n17279, new_n19105);
nor_5  g16757(new_n19105, new_n19104, new_n19106);
xnor_4 g16758(new_n19102, new_n17895, new_n19107_1);
and_5  g16759(new_n19107_1, new_n19106, new_n19108);
nor_5  g16760(new_n19108, new_n19103, new_n19109);
xnor_4 g16761(new_n19109, new_n19100, n7313);
xnor_4 g16762(new_n3506_1, new_n3483, n7346);
xor_4  g16763(new_n18805, new_n12646, new_n19112);
nor_5  g16764(new_n18805, new_n12649, new_n19113);
xnor_4 g16765(new_n18805, new_n12649, new_n19114);
not_10 g16766(new_n10210, new_n19115);
and_5  g16767(new_n12653, new_n19115, new_n19116_1);
xnor_4 g16768(new_n12653, new_n19115, new_n19117);
not_10 g16769(new_n10213, new_n19118);
and_5  g16770(new_n12657_1, new_n19118, new_n19119);
xnor_4 g16771(new_n12657_1, new_n19118, new_n19120);
nor_5  g16772(new_n12661, new_n10217, new_n19121);
nor_5  g16773(new_n5951, new_n5845, new_n19122);
nor_5  g16774(new_n5981, new_n5952, new_n19123);
nor_5  g16775(new_n19123, new_n19122, new_n19124);
xor_4  g16776(new_n12661, new_n10217, new_n19125_1);
and_5  g16777(new_n19125_1, new_n19124, new_n19126);
nor_5  g16778(new_n19126, new_n19121, new_n19127);
nor_5  g16779(new_n19127, new_n19120, new_n19128);
nor_5  g16780(new_n19128, new_n19119, new_n19129);
nor_5  g16781(new_n19129, new_n19117, new_n19130);
nor_5  g16782(new_n19130, new_n19116_1, new_n19131);
nor_5  g16783(new_n19131, new_n19114, new_n19132);
or_5   g16784(new_n19132, new_n19113, new_n19133);
xor_4  g16785(new_n19133, new_n19112, n7349);
xnor_4 g16786(new_n19082, new_n19037, n7363);
nor_5  g16787(n21839, new_n8147, new_n19136);
nor_5  g16788(new_n17838, new_n17835, new_n19137);
nor_5  g16789(new_n19137, new_n19136, new_n19138);
xnor_4 g16790(new_n19138, new_n9207, new_n19139);
nor_5  g16791(new_n17839, new_n9210, new_n19140);
nor_5  g16792(new_n17843, new_n17840, new_n19141_1);
nor_5  g16793(new_n19141_1, new_n19140, new_n19142);
xnor_4 g16794(new_n19142, new_n19139, n7390);
xnor_4 g16795(new_n8240, new_n8239, n7403);
xnor_4 g16796(new_n8408_1, new_n8370, n7408);
xnor_4 g16797(new_n18165, new_n18143_1, n7432);
not_10 g16798(new_n16239, new_n19147);
and_5  g16799(new_n19147, new_n13931, new_n19148);
nor_5  g16800(new_n16249, new_n16240, new_n19149);
or_5   g16801(new_n19149, new_n19148, n7475);
xnor_4 g16802(new_n4809, new_n4808, n7477);
xnor_4 g16803(new_n8092, new_n8069, n7507);
xnor_4 g16804(new_n15586, new_n10325, new_n19153);
and_5  g16805(new_n10773, n23895, new_n19154);
xnor_4 g16806(new_n10773, n23895, new_n19155);
and_5  g16807(new_n6222, n17351, new_n19156);
nor_5  g16808(new_n6258, new_n6223_1, new_n19157);
nor_5  g16809(new_n19157, new_n19156, new_n19158);
nor_5  g16810(new_n19158, new_n19155, new_n19159);
nor_5  g16811(new_n19159, new_n19154, new_n19160);
xnor_4 g16812(new_n19160, new_n10819, new_n19161);
xnor_4 g16813(new_n19161, new_n19153, new_n19162);
xnor_4 g16814(new_n15584, new_n15581, new_n19163_1);
xor_4  g16815(new_n19158, new_n19155, new_n19164_1);
nor_5  g16816(new_n19164_1, new_n19163_1, new_n19165);
xnor_4 g16817(new_n19164_1, new_n19163_1, new_n19166);
nor_5  g16818(new_n6259, new_n6197, new_n19167);
nor_5  g16819(new_n6306, new_n6260, new_n19168);
nor_5  g16820(new_n19168, new_n19167, new_n19169);
nor_5  g16821(new_n19169, new_n19166, new_n19170);
nor_5  g16822(new_n19170, new_n19165, new_n19171);
xnor_4 g16823(new_n19171, new_n19162, n7514);
xnor_4 g16824(new_n9804, new_n9781, n7558);
xnor_4 g16825(new_n10856, new_n10855, n7572);
xnor_4 g16826(new_n5710, n7693, new_n19175);
and_5  g16827(new_n5711, n10405, new_n19176_1);
nor_5  g16828(new_n18195, new_n18185, new_n19177);
nor_5  g16829(new_n19177, new_n19176_1, new_n19178);
xor_4  g16830(new_n19178, new_n19175, new_n19179);
xnor_4 g16831(new_n19179, new_n8798, new_n19180);
nor_5  g16832(new_n18196, new_n8803_1, new_n19181);
nor_5  g16833(new_n18209, new_n18197, new_n19182);
nor_5  g16834(new_n19182, new_n19181, new_n19183);
xnor_4 g16835(new_n19183, new_n19180, n7575);
xnor_4 g16836(new_n18936, new_n8742, new_n19185);
xnor_4 g16837(new_n8739, new_n8713, new_n19186);
nor_5  g16838(new_n18940_1, new_n19186, new_n19187);
xnor_4 g16839(new_n18940_1, new_n19186, new_n19188);
nor_5  g16840(new_n18943, new_n8789, new_n19189);
nor_5  g16841(new_n9854, new_n9824, new_n19190);
nor_5  g16842(new_n19190, new_n19189, new_n19191);
nor_5  g16843(new_n19191, new_n19188, new_n19192);
nor_5  g16844(new_n19192, new_n19187, new_n19193);
xor_4  g16845(new_n19193, new_n19185, new_n19194);
xnor_4 g16846(new_n19194, new_n10378, new_n19195);
xor_4  g16847(new_n19191, new_n19188, new_n19196_1);
and_5  g16848(new_n19196_1, new_n10383, new_n19197);
xnor_4 g16849(new_n19196_1, new_n10383, new_n19198);
nor_5  g16850(new_n9864, new_n9855, new_n19199);
nor_5  g16851(new_n9895, new_n9865, new_n19200);
or_5   g16852(new_n19200, new_n19199, new_n19201);
nor_5  g16853(new_n19201, new_n19198, new_n19202_1);
nor_5  g16854(new_n19202_1, new_n19197, new_n19203);
xor_4  g16855(new_n19203, new_n19195, n7585);
xnor_4 g16856(new_n18665, new_n7020, new_n19205);
nor_5  g16857(new_n18668, new_n7024, new_n19206);
xnor_4 g16858(new_n18668, new_n7024, new_n19207);
xnor_4 g16859(new_n7012, new_n6979, new_n19208);
and_5  g16860(new_n18672, new_n19208, new_n19209);
xnor_4 g16861(new_n18672, new_n19208, new_n19210);
nor_5  g16862(new_n18677, new_n7032_1, new_n19211);
xnor_4 g16863(new_n18677, new_n7032_1, new_n19212);
nor_5  g16864(new_n16330, new_n7036, new_n19213);
xnor_4 g16865(new_n16330, new_n7036, new_n19214);
nor_5  g16866(new_n16333, new_n7040, new_n19215);
xnor_4 g16867(new_n16333, new_n7040, new_n19216);
nor_5  g16868(new_n16336, new_n7044, new_n19217);
xnor_4 g16869(new_n16336, new_n7044, new_n19218);
and_5  g16870(new_n16341, new_n7049, new_n19219);
xor_4  g16871(new_n16340, new_n7049, new_n19220_1);
or_5   g16872(new_n16346, new_n7059, new_n19221_1);
and_5  g16873(new_n19221_1, new_n7055, new_n19222);
xor_4  g16874(new_n19221_1, new_n7055, new_n19223_1);
and_5  g16875(new_n19223_1, new_n16352, new_n19224_1);
nor_5  g16876(new_n19224_1, new_n19222, new_n19225);
nor_5  g16877(new_n19225, new_n19220_1, new_n19226);
nor_5  g16878(new_n19226, new_n19219, new_n19227);
nor_5  g16879(new_n19227, new_n19218, new_n19228_1);
nor_5  g16880(new_n19228_1, new_n19217, new_n19229);
nor_5  g16881(new_n19229, new_n19216, new_n19230);
nor_5  g16882(new_n19230, new_n19215, new_n19231);
nor_5  g16883(new_n19231, new_n19214, new_n19232);
nor_5  g16884(new_n19232, new_n19213, new_n19233_1);
nor_5  g16885(new_n19233_1, new_n19212, new_n19234_1);
nor_5  g16886(new_n19234_1, new_n19211, new_n19235);
nor_5  g16887(new_n19235, new_n19210, new_n19236);
nor_5  g16888(new_n19236, new_n19209, new_n19237);
nor_5  g16889(new_n19237, new_n19207, new_n19238);
nor_5  g16890(new_n19238, new_n19206, new_n19239);
xnor_4 g16891(new_n19239, new_n19205, n7588);
or_5   g16892(new_n6059, n21832, new_n19241);
or_5   g16893(new_n19241, n21753, new_n19242);
or_5   g16894(new_n19242, n10739, new_n19243);
nor_5  g16895(new_n19243, n13074, new_n19244_1);
xnor_4 g16896(new_n19244_1, n23463, new_n19245);
xnor_4 g16897(new_n19245, n23250, new_n19246);
xnor_4 g16898(new_n19243, new_n10095, new_n19247);
nor_5  g16899(new_n19247, n11455, new_n19248);
xnor_4 g16900(new_n19247, n11455, new_n19249);
xnor_4 g16901(new_n19242, new_n10098, new_n19250);
nor_5  g16902(new_n19250, n3945, new_n19251);
xnor_4 g16903(new_n19250, n3945, new_n19252);
xnor_4 g16904(new_n19241, new_n2350, new_n19253);
nor_5  g16905(new_n19253, n5255, new_n19254);
xnor_4 g16906(new_n19253, n5255, new_n19255);
nor_5  g16907(new_n6060, n21649, new_n19256);
xnor_4 g16908(new_n6060, n21649, new_n19257);
nor_5  g16909(new_n6077, n18274, new_n19258);
nor_5  g16910(new_n6093, n3828, new_n19259);
xnor_4 g16911(new_n6093, n3828, new_n19260);
nor_5  g16912(new_n6088, n23842, new_n19261);
nand_5 g16913(n21654, n2387, new_n19262);
xor_4  g16914(new_n6088, n23842, new_n19263);
and_5  g16915(new_n19263, new_n19262, new_n19264);
nor_5  g16916(new_n19264, new_n19261, new_n19265);
nor_5  g16917(new_n19265, new_n19260, new_n19266);
nor_5  g16918(new_n19266, new_n19259, new_n19267);
xnor_4 g16919(new_n6077, n18274, new_n19268);
nor_5  g16920(new_n19268, new_n19267, new_n19269);
nor_5  g16921(new_n19269, new_n19258, new_n19270_1);
nor_5  g16922(new_n19270_1, new_n19257, new_n19271);
nor_5  g16923(new_n19271, new_n19256, new_n19272);
nor_5  g16924(new_n19272, new_n19255, new_n19273);
nor_5  g16925(new_n19273, new_n19254, new_n19274);
nor_5  g16926(new_n19274, new_n19252, new_n19275);
nor_5  g16927(new_n19275, new_n19251, new_n19276);
nor_5  g16928(new_n19276, new_n19249, new_n19277);
nor_5  g16929(new_n19277, new_n19248, new_n19278);
xor_4  g16930(new_n19278, new_n19246, new_n19279);
xnor_4 g16931(new_n19279, new_n12965, new_n19280);
xnor_4 g16932(new_n19276, new_n19249, new_n19281);
nor_5  g16933(new_n19281, new_n12999, new_n19282_1);
xor_4  g16934(new_n19281, new_n12999, new_n19283);
xor_4  g16935(new_n19274, new_n19252, new_n19284);
nor_5  g16936(new_n19284, new_n13005_1, new_n19285);
xnor_4 g16937(new_n19284, new_n13005_1, new_n19286);
xor_4  g16938(new_n19272, new_n19255, new_n19287);
nor_5  g16939(new_n19287, new_n13009, new_n19288);
xor_4  g16940(new_n19270_1, new_n19257, new_n19289);
nor_5  g16941(new_n19289, new_n13013, new_n19290);
xor_4  g16942(new_n19268, new_n19267, new_n19291);
nor_5  g16943(new_n19291, new_n13016, new_n19292);
xnor_4 g16944(new_n19291, new_n13016, new_n19293);
not_10 g16945(new_n13020, new_n19294);
xor_4  g16946(new_n19265, new_n19260, new_n19295);
nor_5  g16947(new_n19295, new_n19294, new_n19296);
xor_4  g16948(new_n19295, new_n13020, new_n19297);
nor_5  g16949(new_n19263, new_n13023, new_n19298);
xor_4  g16950(new_n19263, new_n19262, new_n19299);
or_5   g16951(new_n19299, new_n13025, new_n19300);
xnor_4 g16952(n21654, n2387, new_n19301);
or_5   g16953(new_n19301, new_n13029, new_n19302);
and_5  g16954(new_n19302, new_n19300, new_n19303);
or_5   g16955(new_n19303, new_n19298, new_n19304);
nor_5  g16956(new_n19304, new_n19297, new_n19305);
nor_5  g16957(new_n19305, new_n19296, new_n19306);
nor_5  g16958(new_n19306, new_n19293, new_n19307);
nor_5  g16959(new_n19307, new_n19292, new_n19308);
xnor_4 g16960(new_n19289, new_n13013, new_n19309);
nor_5  g16961(new_n19309, new_n19308, new_n19310);
nor_5  g16962(new_n19310, new_n19290, new_n19311);
xnor_4 g16963(new_n19287, new_n13009, new_n19312);
nor_5  g16964(new_n19312, new_n19311, new_n19313);
nor_5  g16965(new_n19313, new_n19288, new_n19314_1);
nor_5  g16966(new_n19314_1, new_n19286, new_n19315_1);
nor_5  g16967(new_n19315_1, new_n19285, new_n19316);
and_5  g16968(new_n19316, new_n19283, new_n19317);
or_5   g16969(new_n19317, new_n19282_1, new_n19318);
xor_4  g16970(new_n19318, new_n19280, n7598);
xnor_4 g16971(new_n16247_1, new_n16243_1, n7607);
xnor_4 g16972(new_n4638, new_n4614, n7610);
xnor_4 g16973(new_n3225, new_n3214, n7616);
xnor_4 g16974(n10514, n6105, new_n19323_1);
nor_5  g16975(n18649, n3795, new_n19324);
xnor_4 g16976(n18649, n3795, new_n19325);
nor_5  g16977(n25464, n6218, new_n19326);
xnor_4 g16978(n25464, n6218, new_n19327_1);
nor_5  g16979(n20470, n4590, new_n19328);
xnor_4 g16980(n20470, n4590, new_n19329);
nor_5  g16981(n26752, n21222, new_n19330);
xnor_4 g16982(n26752, n21222, new_n19331);
nor_5  g16983(n9832, n6513, new_n19332);
xnor_4 g16984(n9832, n6513, new_n19333_1);
and_5  g16985(n3918, n1558, new_n19334);
or_5   g16986(n3918, n1558, new_n19335);
nor_5  g16987(n21749, n919, new_n19336);
nor_5  g16988(new_n14901, new_n14896, new_n19337);
nor_5  g16989(new_n19337, new_n19336, new_n19338);
and_5  g16990(new_n19338, new_n19335, new_n19339);
or_5   g16991(new_n19339, new_n19334, new_n19340);
nor_5  g16992(new_n19340, new_n19333_1, new_n19341);
nor_5  g16993(new_n19341, new_n19332, new_n19342);
nor_5  g16994(new_n19342, new_n19331, new_n19343);
nor_5  g16995(new_n19343, new_n19330, new_n19344);
nor_5  g16996(new_n19344, new_n19329, new_n19345);
nor_5  g16997(new_n19345, new_n19328, new_n19346);
nor_5  g16998(new_n19346, new_n19327_1, new_n19347);
nor_5  g16999(new_n19347, new_n19326, new_n19348_1);
nor_5  g17000(new_n19348_1, new_n19325, new_n19349);
nor_5  g17001(new_n19349, new_n19324, new_n19350);
xor_4  g17002(new_n19350, new_n19323_1, new_n19351);
and_5  g17003(new_n19351, n9872, new_n19352);
xnor_4 g17004(new_n19351, n9872, new_n19353);
xor_4  g17005(new_n19348_1, new_n19325, new_n19354_1);
and_5  g17006(new_n19354_1, n5842, new_n19355);
xnor_4 g17007(new_n19354_1, n5842, new_n19356);
xor_4  g17008(new_n19346, new_n19327_1, new_n19357_1);
and_5  g17009(new_n19357_1, n6379, new_n19358);
xnor_4 g17010(new_n19357_1, n6379, new_n19359);
xor_4  g17011(new_n19344, new_n19329, new_n19360);
and_5  g17012(new_n19360, n2102, new_n19361_1);
xnor_4 g17013(new_n19360, n2102, new_n19362);
xor_4  g17014(new_n19342, new_n19331, new_n19363);
and_5  g17015(new_n19363, n17954, new_n19364);
xnor_4 g17016(new_n19363, n17954, new_n19365);
xor_4  g17017(new_n19340, new_n19333_1, new_n19366);
and_5  g17018(new_n19366, n8256, new_n19367_1);
xnor_4 g17019(new_n19366, n8256, new_n19368);
xor_4  g17020(n3918, n1558, new_n19369);
xnor_4 g17021(new_n19369, new_n19338, new_n19370);
and_5  g17022(new_n19370, n24150, new_n19371);
xnor_4 g17023(new_n19370, n24150, new_n19372);
and_5  g17024(new_n14902, n19584, new_n19373);
and_5  g17025(new_n14910, new_n14903, new_n19374);
nor_5  g17026(new_n19374, new_n19373, new_n19375);
nor_5  g17027(new_n19375, new_n19372, new_n19376);
nor_5  g17028(new_n19376, new_n19371, new_n19377);
nor_5  g17029(new_n19377, new_n19368, new_n19378);
nor_5  g17030(new_n19378, new_n19367_1, new_n19379);
nor_5  g17031(new_n19379, new_n19365, new_n19380);
nor_5  g17032(new_n19380, new_n19364, new_n19381);
nor_5  g17033(new_n19381, new_n19362, new_n19382);
nor_5  g17034(new_n19382, new_n19361_1, new_n19383);
nor_5  g17035(new_n19383, new_n19359, new_n19384);
nor_5  g17036(new_n19384, new_n19358, new_n19385_1);
nor_5  g17037(new_n19385_1, new_n19356, new_n19386);
nor_5  g17038(new_n19386, new_n19355, new_n19387);
nor_5  g17039(new_n19387, new_n19353, new_n19388);
nor_5  g17040(new_n19388, new_n19352, new_n19389_1);
nor_5  g17041(n10514, n6105, new_n19390);
nor_5  g17042(new_n19350, new_n19323_1, new_n19391);
nor_5  g17043(new_n19391, new_n19390, new_n19392);
nor_5  g17044(new_n19392, new_n19389_1, new_n19393);
xnor_4 g17045(new_n19393, new_n14158, new_n19394);
xnor_4 g17046(new_n19392, new_n19389_1, new_n19395);
nor_5  g17047(new_n19395, new_n14055, new_n19396);
xnor_4 g17048(new_n19395, new_n14055, new_n19397);
xor_4  g17049(new_n14096, new_n14051, new_n19398);
xor_4  g17050(new_n19387, new_n19353, new_n19399);
and_5  g17051(new_n19399, new_n19398, new_n19400);
xnor_4 g17052(new_n19399, new_n19398, new_n19401_1);
xnor_4 g17053(new_n14049, new_n14019, new_n19402);
xor_4  g17054(new_n19385_1, new_n19356, new_n19403);
and_5  g17055(new_n19403, new_n19402, new_n19404);
xnor_4 g17056(new_n19403, new_n19402, new_n19405);
not_10 g17057(new_n14105, new_n19406);
xor_4  g17058(new_n19383, new_n19359, new_n19407);
and_5  g17059(new_n19407, new_n19406, new_n19408);
xor_4  g17060(new_n19407, new_n14105, new_n19409);
not_10 g17061(new_n14109, new_n19410);
xor_4  g17062(new_n19381, new_n19362, new_n19411);
and_5  g17063(new_n19411, new_n19410, new_n19412);
xor_4  g17064(new_n19411, new_n14109, new_n19413);
not_10 g17065(new_n14113, new_n19414_1);
xor_4  g17066(new_n19379, new_n19365, new_n19415);
and_5  g17067(new_n19415, new_n19414_1, new_n19416);
xor_4  g17068(new_n19415, new_n14113, new_n19417);
not_10 g17069(new_n14117, new_n19418);
xor_4  g17070(new_n19377, new_n19368, new_n19419);
and_5  g17071(new_n19419, new_n19418, new_n19420);
xor_4  g17072(new_n19419, new_n14117, new_n19421);
xor_4  g17073(new_n19375, new_n19372, new_n19422);
and_5  g17074(new_n19422, new_n14121_1, new_n19423);
xnor_4 g17075(new_n19422, new_n14121_1, new_n19424_1);
and_5  g17076(new_n14911, new_n14137, new_n19425);
nor_5  g17077(new_n14919, new_n14912, new_n19426);
nor_5  g17078(new_n19426, new_n19425, new_n19427);
nor_5  g17079(new_n19427, new_n19424_1, new_n19428);
nor_5  g17080(new_n19428, new_n19423, new_n19429);
nor_5  g17081(new_n19429, new_n19421, new_n19430);
nor_5  g17082(new_n19430, new_n19420, new_n19431);
nor_5  g17083(new_n19431, new_n19417, new_n19432);
nor_5  g17084(new_n19432, new_n19416, new_n19433);
nor_5  g17085(new_n19433, new_n19413, new_n19434);
nor_5  g17086(new_n19434, new_n19412, new_n19435);
nor_5  g17087(new_n19435, new_n19409, new_n19436);
nor_5  g17088(new_n19436, new_n19408, new_n19437);
nor_5  g17089(new_n19437, new_n19405, new_n19438);
nor_5  g17090(new_n19438, new_n19404, new_n19439);
nor_5  g17091(new_n19439, new_n19401_1, new_n19440);
nor_5  g17092(new_n19440, new_n19400, new_n19441);
nor_5  g17093(new_n19441, new_n19397, new_n19442);
or_5   g17094(new_n19442, new_n19396, new_n19443);
xnor_4 g17095(new_n19443, new_n19394, n7630);
nor_5  g17096(new_n17034, new_n17013, new_n19445);
nor_5  g17097(new_n17045, new_n17035_1, new_n19446);
nor_5  g17098(new_n19446, new_n19445, n7643);
xnor_4 g17099(new_n10978, new_n10955, n7647);
xnor_4 g17100(new_n9084, new_n9056, n7679);
xnor_4 g17101(new_n18371, new_n18346, n7686);
xnor_4 g17102(new_n16565, new_n16545, new_n19451);
xnor_4 g17103(new_n19451, new_n16581, n7698);
xnor_4 g17104(new_n17645, new_n17630, n7708);
xor_4  g17105(new_n16556, n3324, new_n19454_1);
and_5  g17106(new_n2838, n17911, new_n19455);
xnor_4 g17107(new_n2838, n17911, new_n19456);
nor_5  g17108(new_n2871, n21997, new_n19457);
xnor_4 g17109(new_n2871, n21997, new_n19458_1);
nor_5  g17110(new_n2875, n25119, new_n19459);
and_5  g17111(new_n7758, new_n7737, new_n19460);
nor_5  g17112(new_n19460, new_n19459, new_n19461);
nor_5  g17113(new_n19461, new_n19458_1, new_n19462);
or_5   g17114(new_n19462, new_n19457, new_n19463);
nor_5  g17115(new_n19463, new_n19456, new_n19464);
nor_5  g17116(new_n19464, new_n19455, new_n19465);
xor_4  g17117(new_n19465, new_n19454_1, new_n19466);
xor_4  g17118(new_n5526, n3740, new_n19467_1);
nor_5  g17119(new_n5528, n2858, new_n19468);
and_5  g17120(new_n14688, new_n14681, new_n19469);
nor_5  g17121(new_n19469, new_n19468, new_n19470);
xor_4  g17122(new_n19470, new_n19467_1, new_n19471);
xnor_4 g17123(new_n19471, new_n19466, new_n19472_1);
xor_4  g17124(new_n19463, new_n19456, new_n19473);
nor_5  g17125(new_n19473, new_n14689, new_n19474);
xnor_4 g17126(new_n19473, new_n14689, new_n19475);
xor_4  g17127(new_n19461, new_n19458_1, new_n19476);
and_5  g17128(new_n19476, new_n14691, new_n19477_1);
xnor_4 g17129(new_n19476, new_n14691, new_n19478);
and_5  g17130(new_n7759_1, new_n7736, new_n19479);
nor_5  g17131(new_n7795, new_n7760, new_n19480);
nor_5  g17132(new_n19480, new_n19479, new_n19481);
nor_5  g17133(new_n19481, new_n19478, new_n19482);
nor_5  g17134(new_n19482, new_n19477_1, new_n19483);
nor_5  g17135(new_n19483, new_n19475, new_n19484);
nor_5  g17136(new_n19484, new_n19474, new_n19485);
xnor_4 g17137(new_n19485, new_n19472_1, n7780);
and_5  g17138(new_n2567, n18880, new_n19487);
xnor_4 g17139(new_n2567, n18880, new_n19488);
and_5  g17140(new_n2569, n25475, new_n19489);
nor_5  g17141(new_n8741, new_n8711, new_n19490);
nor_5  g17142(new_n19490, new_n19489, new_n19491);
nor_5  g17143(new_n19491, new_n19488, new_n19492);
nor_5  g17144(new_n19492, new_n19487, new_n19493);
xor_4  g17145(new_n19493, new_n13231, new_n19494_1);
and_5  g17146(new_n15723, new_n2657, new_n19495);
xnor_4 g17147(new_n15723, new_n2657, new_n19496_1);
and_5  g17148(new_n8748, new_n2660, new_n19497);
nor_5  g17149(new_n8782_1, new_n8749, new_n19498);
nor_5  g17150(new_n19498, new_n19497, new_n19499);
nor_5  g17151(new_n19499, new_n19496_1, new_n19500);
nor_5  g17152(new_n19500, new_n19495, new_n19501);
nor_5  g17153(new_n15722, n21839, new_n19502);
xor_4  g17154(new_n19502, new_n9163, new_n19503);
xnor_4 g17155(new_n19503, new_n19501, new_n19504);
xnor_4 g17156(new_n19504, new_n19494_1, new_n19505);
xor_4  g17157(new_n19491, new_n19488, new_n19506);
xor_4  g17158(new_n19499, new_n19496_1, new_n19507);
nor_5  g17159(new_n19507, new_n19506, new_n19508);
xnor_4 g17160(new_n19507, new_n19506, new_n19509);
xor_4  g17161(new_n8741, new_n8711, new_n19510);
nor_5  g17162(new_n8783, new_n19510, new_n19511);
and_5  g17163(new_n8832, new_n8784, new_n19512);
nor_5  g17164(new_n19512, new_n19511, new_n19513);
nor_5  g17165(new_n19513, new_n19509, new_n19514_1);
nor_5  g17166(new_n19514_1, new_n19508, new_n19515_1);
xnor_4 g17167(new_n19515_1, new_n19505, n7794);
xnor_4 g17168(new_n15876, new_n15871, n7811);
xor_4  g17169(new_n15829, new_n15824, n7830);
xnor_4 g17170(new_n19235, new_n19210, n7834);
xnor_4 g17171(new_n9889, new_n9876, n7884);
xnor_4 g17172(new_n2951, new_n2950, n7937);
xnor_4 g17173(new_n2963, new_n2921, n7943);
xor_4  g17174(new_n8826, new_n8797, n7950);
not_10 g17175(new_n14010, new_n19524);
xnor_4 g17176(new_n17891, new_n19524, new_n19525);
and_5  g17177(new_n17896, new_n14012, new_n19526);
nor_5  g17178(new_n17898, new_n14017, new_n19527);
xnor_4 g17179(new_n17898, new_n14017, new_n19528);
nor_5  g17180(new_n13783_1, new_n13743, new_n19529);
nor_5  g17181(new_n13822, new_n13784, new_n19530);
nor_5  g17182(new_n19530, new_n19529, new_n19531_1);
nor_5  g17183(new_n19531_1, new_n19528, new_n19532);
or_5   g17184(new_n19532, new_n19527, new_n19533);
xnor_4 g17185(new_n17896, new_n14013, new_n19534);
and_5  g17186(new_n19534, new_n19533, new_n19535);
or_5   g17187(new_n19535, new_n19526, new_n19536);
xor_4  g17188(new_n19536, new_n19525, n7959);
xnor_4 g17189(new_n15880, new_n15866, n7968);
xnor_4 g17190(new_n16790, new_n16789, n7992);
xnor_4 g17191(new_n11625, n9554, new_n19540);
nand_5 g17192(new_n11628, n26408, new_n19541);
xnor_4 g17193(new_n11628, n26408, new_n19542);
nor_5  g17194(new_n9526, n18227, new_n19543);
and_5  g17195(new_n15856, new_n15845, new_n19544);
nor_5  g17196(new_n19544, new_n19543, new_n19545);
not_10 g17197(new_n19545, new_n19546);
or_5   g17198(new_n19546, new_n19542, new_n19547);
and_5  g17199(new_n19547, new_n19541, new_n19548);
xnor_4 g17200(new_n19548, new_n19540, new_n19549);
xnor_4 g17201(new_n19549, new_n16948, new_n19550);
xnor_4 g17202(new_n19545, new_n19542, new_n19551);
and_5  g17203(new_n19551, new_n16952, new_n19552);
xnor_4 g17204(new_n19551, new_n16952, new_n19553);
nor_5  g17205(new_n16957, new_n15857, new_n19554);
xnor_4 g17206(new_n16957, new_n15857, new_n19555);
not_10 g17207(new_n15859_1, new_n19556);
nor_5  g17208(new_n16961, new_n19556, new_n19557);
xor_4  g17209(new_n16961, new_n15859_1, new_n19558);
and_5  g17210(new_n16966, new_n15862, new_n19559);
xnor_4 g17211(new_n16966, new_n15862, new_n19560);
nor_5  g17212(new_n11712_1, new_n11702, new_n19561);
nor_5  g17213(new_n11717, new_n11713, new_n19562);
nor_5  g17214(new_n19562, new_n19561, new_n19563);
nor_5  g17215(new_n19563, new_n19560, new_n19564);
nor_5  g17216(new_n19564, new_n19559, new_n19565);
nor_5  g17217(new_n19565, new_n19558, new_n19566);
nor_5  g17218(new_n19566, new_n19557, new_n19567);
nor_5  g17219(new_n19567, new_n19555, new_n19568);
nor_5  g17220(new_n19568, new_n19554, new_n19569);
nor_5  g17221(new_n19569, new_n19553, new_n19570_1);
nor_5  g17222(new_n19570_1, new_n19552, new_n19571);
xnor_4 g17223(new_n19571, new_n19550, n7999);
xnor_4 g17224(new_n16458, new_n16447, n8027);
nor_5  g17225(new_n19493, new_n13231, new_n19574);
and_5  g17226(new_n5692, n8614, new_n19575_1);
xnor_4 g17227(new_n5692, n8614, new_n19576);
and_5  g17228(new_n5697, n15182, new_n19577);
nor_5  g17229(new_n5701, n27037, new_n19578);
xnor_4 g17230(new_n5701, n27037, new_n19579);
or_5   g17231(new_n5704_1, n8964, new_n19580);
xnor_4 g17232(new_n5704_1, n8964, new_n19581);
and_5  g17233(new_n5707, n20151, new_n19582);
and_5  g17234(new_n5710, n7693, new_n19583);
nor_5  g17235(new_n19178, new_n19175, new_n19584_1);
nor_5  g17236(new_n19584_1, new_n19583, new_n19585);
xnor_4 g17237(new_n5707, n20151, new_n19586);
nor_5  g17238(new_n19586, new_n19585, new_n19587);
nor_5  g17239(new_n19587, new_n19582, new_n19588);
not_10 g17240(new_n19588, new_n19589);
or_5   g17241(new_n19589, new_n19581, new_n19590);
and_5  g17242(new_n19590, new_n19580, new_n19591);
nor_5  g17243(new_n19591, new_n19579, new_n19592);
or_5   g17244(new_n19592, new_n19578, new_n19593);
xnor_4 g17245(new_n5697, n15182, new_n19594);
nor_5  g17246(new_n19594, new_n19593, new_n19595);
nor_5  g17247(new_n19595, new_n19577, new_n19596);
nor_5  g17248(new_n19596, new_n19576, new_n19597);
nor_5  g17249(new_n19597, new_n19575_1, new_n19598);
or_5   g17250(new_n19598, new_n11295, new_n19599);
and_5  g17251(new_n19599, new_n19574, new_n19600);
nor_5  g17252(new_n19599, new_n19574, new_n19601);
xnor_4 g17253(new_n19493, new_n13231, new_n19602_1);
xnor_4 g17254(new_n19598, new_n5660, new_n19603);
nor_5  g17255(new_n19603, new_n19602_1, new_n19604);
xnor_4 g17256(new_n19603, new_n19602_1, new_n19605);
xnor_4 g17257(new_n19491, new_n19488, new_n19606);
xor_4  g17258(new_n19596, new_n19576, new_n19607);
nor_5  g17259(new_n19607, new_n19606, new_n19608_1);
xnor_4 g17260(new_n19607, new_n19606, new_n19609);
xor_4  g17261(new_n19594, new_n19593, new_n19610);
nor_5  g17262(new_n19610, new_n8742, new_n19611);
xnor_4 g17263(new_n19610, new_n8742, new_n19612);
xor_4  g17264(new_n19591, new_n19579, new_n19613);
and_5  g17265(new_n19613, new_n8785, new_n19614);
xnor_4 g17266(new_n19613, new_n8785, new_n19615);
xnor_4 g17267(new_n19588, new_n19581, new_n19616);
and_5  g17268(new_n19616, new_n8792, new_n19617_1);
xnor_4 g17269(new_n19616, new_n8792, new_n19618_1);
xor_4  g17270(new_n19586, new_n19585, new_n19619);
nor_5  g17271(new_n19619, new_n8794, new_n19620);
xnor_4 g17272(new_n19619, new_n8794, new_n19621);
nor_5  g17273(new_n19179, new_n8798, new_n19622);
nor_5  g17274(new_n19183, new_n19180, new_n19623_1);
nor_5  g17275(new_n19623_1, new_n19622, new_n19624);
nor_5  g17276(new_n19624, new_n19621, new_n19625);
nor_5  g17277(new_n19625, new_n19620, new_n19626);
nor_5  g17278(new_n19626, new_n19618_1, new_n19627);
nor_5  g17279(new_n19627, new_n19617_1, new_n19628);
nor_5  g17280(new_n19628, new_n19615, new_n19629);
nor_5  g17281(new_n19629, new_n19614, new_n19630);
nor_5  g17282(new_n19630, new_n19612, new_n19631);
nor_5  g17283(new_n19631, new_n19611, new_n19632);
nor_5  g17284(new_n19632, new_n19609, new_n19633);
nor_5  g17285(new_n19633, new_n19608_1, new_n19634);
nor_5  g17286(new_n19634, new_n19605, new_n19635);
nor_5  g17287(new_n19635, new_n19604, new_n19636);
nor_5  g17288(new_n19636, new_n19601, new_n19637);
or_5   g17289(new_n19637, new_n19600, n8031);
and_5  g17290(new_n15723, n22626, new_n19639);
or_5   g17291(new_n15723, n22626, new_n19640);
and_5  g17292(new_n15731, new_n19640, new_n19641_1);
or_5   g17293(new_n19641_1, new_n19502, new_n19642);
nor_5  g17294(new_n19642, new_n19639, new_n19643);
not_10 g17295(new_n19643, new_n19644);
nor_5  g17296(new_n19644, new_n18045_1, new_n19645);
xor_4  g17297(new_n19643, new_n18045_1, new_n19646);
and_5  g17298(new_n15732, new_n18047, new_n19647);
or_5   g17299(new_n15757, new_n15735, new_n19648_1);
nor_5  g17300(new_n19648_1, new_n15733, new_n19649);
nor_5  g17301(new_n19649, new_n19647, new_n19650);
nor_5  g17302(new_n19650, new_n19646, new_n19651);
or_5   g17303(new_n19651, new_n19645, new_n19652_1);
nor_5  g17304(new_n15767, n9554, new_n19653);
nor_5  g17305(new_n15797, new_n19653, new_n19654);
and_5  g17306(new_n15767, n9554, new_n19655);
or_5   g17307(new_n19655, new_n18320, new_n19656);
nor_5  g17308(new_n19656, new_n19654, new_n19657);
nor_5  g17309(new_n19657, new_n19652_1, new_n19658);
nor_5  g17310(new_n19651, new_n19645, new_n19659);
or_5   g17311(new_n19656, new_n19654, new_n19660);
xnor_4 g17312(new_n19660, new_n19659, new_n19661);
xor_4  g17313(new_n19650, new_n19646, new_n19662);
nor_5  g17314(new_n19662, new_n19660, new_n19663);
xnor_4 g17315(new_n19650, new_n19646, new_n19664_1);
xnor_4 g17316(new_n19664_1, new_n19657, new_n19665);
nor_5  g17317(new_n15798, new_n15759, new_n19666);
nor_5  g17318(new_n15843, new_n15799, new_n19667);
nor_5  g17319(new_n19667, new_n19666, new_n19668);
nor_5  g17320(new_n19668, new_n19665, new_n19669);
nor_5  g17321(new_n19669, new_n19663, new_n19670);
nor_5  g17322(new_n19670, new_n19661, new_n19671);
nor_5  g17323(new_n19671, new_n19658, n8042);
nor_5  g17324(new_n9031, new_n8943_1, new_n19673);
nor_5  g17325(new_n9096, new_n9032_1, new_n19674);
or_5   g17326(new_n19674, new_n19673, n8095);
nor_5  g17327(new_n15760, n4306, new_n19676);
xor_4  g17328(n23166, n4306, new_n19677);
nor_5  g17329(new_n8268, n3279, new_n19678);
xor_4  g17330(n10577, n3279, new_n19679);
nor_5  g17331(n13914, new_n8271, new_n19680_1);
xor_4  g17332(n13914, n6381, new_n19681);
nor_5  g17333(n14702, new_n8274, new_n19682);
nor_5  g17334(new_n17795, new_n17784_1, new_n19683);
nor_5  g17335(new_n19683, new_n19682, new_n19684);
nor_5  g17336(new_n19684, new_n19681, new_n19685);
nor_5  g17337(new_n19685, new_n19680_1, new_n19686);
nor_5  g17338(new_n19686, new_n19679, new_n19687);
nor_5  g17339(new_n19687, new_n19678, new_n19688);
nor_5  g17340(new_n19688, new_n19677, new_n19689);
nor_5  g17341(new_n19689, new_n19676, new_n19690);
xnor_4 g17342(new_n19690, new_n8146, new_n19691);
xor_4  g17343(new_n19688, new_n19677, new_n19692);
nor_5  g17344(new_n19692, new_n8196, new_n19693);
xnor_4 g17345(new_n19692, new_n8196, new_n19694);
xnor_4 g17346(new_n8140, new_n8111, new_n19695);
xor_4  g17347(new_n19686, new_n19679, new_n19696);
nor_5  g17348(new_n19696, new_n19695, new_n19697);
xnor_4 g17349(new_n19696, new_n19695, new_n19698);
xnor_4 g17350(new_n8138, new_n8113, new_n19699);
xor_4  g17351(new_n19684, new_n19681, new_n19700);
nor_5  g17352(new_n19700, new_n19699, new_n19701_1);
xor_4  g17353(new_n19700, new_n19699, new_n19702);
and_5  g17354(new_n17796, new_n17783, new_n19703);
nor_5  g17355(new_n17812, new_n17797, new_n19704);
nor_5  g17356(new_n19704, new_n19703, new_n19705);
and_5  g17357(new_n19705, new_n19702, new_n19706);
nor_5  g17358(new_n19706, new_n19701_1, new_n19707);
nor_5  g17359(new_n19707, new_n19698, new_n19708);
nor_5  g17360(new_n19708, new_n19697, new_n19709);
nor_5  g17361(new_n19709, new_n19694, new_n19710);
nor_5  g17362(new_n19710, new_n19693, new_n19711);
xnor_4 g17363(new_n19711, new_n19691, n8103);
xnor_4 g17364(new_n17176, new_n17162, n8109);
and_5  g17365(new_n17621, new_n17605, new_n19714);
nor_5  g17366(new_n17649, new_n17622, new_n19715);
or_5   g17367(new_n19715, new_n19714, n8127);
xnor_4 g17368(new_n15287, new_n15284, n8130);
nor_5  g17369(n8856, new_n10596, new_n19718);
xor_4  g17370(n8856, n4319, new_n19719);
nor_5  g17371(new_n10599, n14130, new_n19720);
xor_4  g17372(n23463, n14130, new_n19721);
nor_5  g17373(n16482, new_n10095, new_n19722);
xor_4  g17374(n16482, n13074, new_n19723);
nor_5  g17375(new_n10098, n9942, new_n19724);
nor_5  g17376(new_n2378, new_n2349, new_n19725);
nor_5  g17377(new_n19725, new_n19724, new_n19726);
nor_5  g17378(new_n19726, new_n19723, new_n19727);
nor_5  g17379(new_n19727, new_n19722, new_n19728);
nor_5  g17380(new_n19728, new_n19721, new_n19729);
nor_5  g17381(new_n19729, new_n19720, new_n19730);
nor_5  g17382(new_n19730, new_n19719, new_n19731);
nor_5  g17383(new_n19731, new_n19718, new_n19732);
xnor_4 g17384(new_n19732, new_n6859, new_n19733);
nor_5  g17385(new_n19732, new_n6862_1, new_n19734);
xnor_4 g17386(new_n19732, new_n6862_1, new_n19735);
not_10 g17387(new_n6866, new_n19736_1);
xor_4  g17388(new_n19730, new_n19719, new_n19737);
nor_5  g17389(new_n19737, new_n19736_1, new_n19738);
xor_4  g17390(new_n19737, new_n6866, new_n19739);
xnor_4 g17391(new_n19728, new_n19721, new_n19740);
and_5  g17392(new_n19740, new_n6870, new_n19741);
xor_4  g17393(new_n19740, new_n6870, new_n19742);
xnor_4 g17394(new_n19726, new_n19723, new_n19743);
nor_5  g17395(new_n19743, new_n6874, new_n19744);
xnor_4 g17396(new_n19743, new_n6874, new_n19745);
nor_5  g17397(new_n2485, new_n2379, new_n19746);
nor_5  g17398(new_n2521, new_n2486, new_n19747);
nor_5  g17399(new_n19747, new_n19746, new_n19748);
nor_5  g17400(new_n19748, new_n19745, new_n19749_1);
nor_5  g17401(new_n19749_1, new_n19744, new_n19750);
and_5  g17402(new_n19750, new_n19742, new_n19751);
nor_5  g17403(new_n19751, new_n19741, new_n19752);
nor_5  g17404(new_n19752, new_n19739, new_n19753);
nor_5  g17405(new_n19753, new_n19738, new_n19754);
nor_5  g17406(new_n19754, new_n19735, new_n19755);
nor_5  g17407(new_n19755, new_n19734, new_n19756_1);
xnor_4 g17408(new_n19756_1, new_n19733, n8135);
xnor_4 g17409(new_n6902, new_n2510, n8139);
nand_5 g17410(new_n16588, new_n6939, new_n19759);
or_5   g17411(new_n19759, n26660, new_n19760);
xor_4  g17412(new_n19760, n13783, new_n19761);
xnor_4 g17413(new_n19761, new_n2876, new_n19762);
xor_4  g17414(new_n19759, n26660, new_n19763);
and_5  g17415(new_n19763, new_n2880, new_n19764);
xnor_4 g17416(new_n19763, new_n2880, new_n19765);
and_5  g17417(new_n16589_1, new_n2884, new_n19766);
nor_5  g17418(new_n16606, new_n16590, new_n19767_1);
nor_5  g17419(new_n19767_1, new_n19766, new_n19768);
nor_5  g17420(new_n19768, new_n19765, new_n19769);
nor_5  g17421(new_n19769, new_n19764, new_n19770_1);
xor_4  g17422(new_n19770_1, new_n19762, new_n19771);
xnor_4 g17423(new_n19771, new_n6266, new_n19772);
xor_4  g17424(new_n19768, new_n19765, new_n19773);
nor_5  g17425(new_n19773, new_n6270, new_n19774);
xnor_4 g17426(new_n19773, new_n6270, new_n19775);
not_10 g17427(new_n6273, new_n19776);
nor_5  g17428(new_n16607, new_n19776, new_n19777);
nor_5  g17429(new_n16625, new_n16608_1, new_n19778);
nor_5  g17430(new_n19778, new_n19777, new_n19779);
nor_5  g17431(new_n19779, new_n19775, new_n19780_1);
nor_5  g17432(new_n19780_1, new_n19774, new_n19781);
xnor_4 g17433(new_n19781, new_n19772, n8148);
xor_4  g17434(new_n16034, new_n16033, n8149);
xnor_4 g17435(new_n3689, new_n3673, n8159);
xor_4  g17436(new_n10550, new_n2531, n8179);
xnor_4 g17437(new_n13475, new_n13472, n8215);
xnor_4 g17438(new_n17174, new_n17165, n8267);
xnor_4 g17439(new_n18205, new_n18204, n8276);
not_10 g17440(n1654, new_n19789_1);
nor_5  g17441(new_n19760, n13783, new_n19790);
nand_5 g17442(new_n19790, new_n19789_1, new_n19791);
or_5   g17443(new_n19791, n14440, new_n19792_1);
xor_4  g17444(new_n19792_1, n22626, new_n19793);
nor_5  g17445(new_n19793, new_n13639, new_n19794);
xnor_4 g17446(new_n19793, new_n13639, new_n19795);
xor_4  g17447(new_n19791, n14440, new_n19796);
or_5   g17448(new_n19796, new_n2869, new_n19797);
xnor_4 g17449(new_n19796, new_n2869, new_n19798_1);
xnor_4 g17450(new_n19790, n1654, new_n19799);
and_5  g17451(new_n19799, new_n2872, new_n19800);
and_5  g17452(new_n19761, new_n2876, new_n19801);
nor_5  g17453(new_n19770_1, new_n19762, new_n19802);
nor_5  g17454(new_n19802, new_n19801, new_n19803_1);
xnor_4 g17455(new_n19799, new_n2872, new_n19804);
nor_5  g17456(new_n19804, new_n19803_1, new_n19805);
nor_5  g17457(new_n19805, new_n19800, new_n19806);
not_10 g17458(new_n19806, new_n19807);
or_5   g17459(new_n19807, new_n19798_1, new_n19808);
and_5  g17460(new_n19808, new_n19797, new_n19809);
nor_5  g17461(new_n19809, new_n19795, new_n19810);
nor_5  g17462(new_n19810, new_n19794, new_n19811);
nor_5  g17463(new_n19792_1, n22626, new_n19812);
xnor_4 g17464(new_n19812, new_n13661, new_n19813);
xnor_4 g17465(new_n19813, new_n19811, new_n19814);
nor_5  g17466(new_n19814, new_n15639, new_n19815);
xnor_4 g17467(new_n19814, new_n15639, new_n19816);
xor_4  g17468(new_n19809, new_n19795, new_n19817);
and_5  g17469(new_n19817, new_n19163_1, new_n19818);
xnor_4 g17470(new_n19817, new_n19163_1, new_n19819);
xnor_4 g17471(new_n19806, new_n19798_1, new_n19820);
and_5  g17472(new_n19820, new_n6197, new_n19821);
xor_4  g17473(new_n19804, new_n19803_1, new_n19822);
nor_5  g17474(new_n19822, new_n6262, new_n19823);
xnor_4 g17475(new_n19822, new_n6262, new_n19824);
nor_5  g17476(new_n19771, new_n6266, new_n19825);
nor_5  g17477(new_n19781, new_n19772, new_n19826);
nor_5  g17478(new_n19826, new_n19825, new_n19827);
nor_5  g17479(new_n19827, new_n19824, new_n19828);
nor_5  g17480(new_n19828, new_n19823, new_n19829);
xnor_4 g17481(new_n19820, new_n6197, new_n19830);
nor_5  g17482(new_n19830, new_n19829, new_n19831);
nor_5  g17483(new_n19831, new_n19821, new_n19832);
nor_5  g17484(new_n19832, new_n19819, new_n19833);
nor_5  g17485(new_n19833, new_n19818, new_n19834);
nor_5  g17486(new_n19834, new_n19816, new_n19835);
nor_5  g17487(new_n19835, new_n19815, new_n19836);
and_5  g17488(new_n19836, new_n15587, new_n19837);
or_5   g17489(new_n19812, new_n13662, new_n19838);
nor_5  g17490(new_n19838, new_n19811, new_n19839);
or_5   g17491(new_n19836, new_n15587, new_n19840);
and_5  g17492(new_n19812, new_n13662, new_n19841);
and_5  g17493(new_n19841, new_n19811, new_n19842);
nor_5  g17494(new_n19842, new_n19840, new_n19843);
nor_5  g17495(new_n19843, new_n19839, new_n19844);
nor_5  g17496(new_n19844, new_n19837, n8288);
xor_4  g17497(new_n10151, new_n6717, n8306);
xor_4  g17498(new_n7196, new_n7153, n8320);
xnor_4 g17499(new_n11278, new_n11260, n8321);
xnor_4 g17500(new_n14869, new_n14856, n8339);
xnor_4 g17501(new_n8248, new_n8206, n8376);
xor_4  g17502(new_n17489, new_n9241, n8408);
xor_4  g17503(new_n13029, new_n13028, n8417);
xnor_4 g17504(new_n11664, new_n11650, n8432);
not_10 g17505(new_n9160, new_n19854);
nor_5  g17506(new_n9163, new_n19854, new_n19855);
nor_5  g17507(new_n9206, new_n9164_1, new_n19856);
nor_5  g17508(new_n19856, new_n19855, new_n19857);
not_10 g17509(new_n19857, new_n19858);
and_5  g17510(new_n19858, new_n9145, new_n19859);
nor_5  g17511(new_n9207, new_n9145, new_n19860);
nor_5  g17512(new_n9268, new_n9208, new_n19861);
nor_5  g17513(new_n19861, new_n19860, new_n19862);
nor_5  g17514(new_n19862, new_n19859, new_n19863);
nor_5  g17515(new_n19858, new_n9145, new_n19864);
nor_5  g17516(new_n19864, new_n19861, new_n19865);
nor_5  g17517(new_n19865, new_n19863, n8453);
xor_4  g17518(new_n14166, new_n12387, n8480);
xnor_4 g17519(new_n15025, new_n15005, n8489);
xnor_4 g17520(new_n19752, new_n19739, n8505);
xnor_4 g17521(new_n17908, new_n17894, n8510);
xor_4  g17522(new_n10970, new_n7846, n8519);
xnor_4 g17523(new_n8818, new_n8817, n8535);
xnor_4 g17524(new_n17641, new_n17638_1, n8550);
xnor_4 g17525(new_n18768, new_n18762, n8563);
xnor_4 g17526(new_n12060, new_n12059, n8594);
xnor_4 g17527(new_n6296, new_n6280, n8608);
xor_4  g17528(new_n4243, new_n4242, n8620);
xnor_4 g17529(new_n6738, new_n6691_1, n8637);
xnor_4 g17530(new_n15654, new_n15653, n8662);
xnor_4 g17531(new_n17227, new_n17217, n8716);
xnor_4 g17532(new_n7155, new_n7154, new_n19881);
xnor_4 g17533(new_n19881, new_n7194, n8744);
nand_5 g17534(new_n11625, n9554, new_n19883);
or_5   g17535(new_n19548, new_n19540, new_n19884);
and_5  g17536(new_n19884, new_n19883, new_n19885);
xnor_4 g17537(new_n19885, new_n13930, new_n19886);
and_5  g17538(new_n5526, n3740, new_n19887);
and_5  g17539(new_n19470, new_n19467_1, new_n19888);
nor_5  g17540(new_n19888, new_n19887, new_n19889);
xor_4  g17541(new_n19889, new_n16238, new_n19890);
xnor_4 g17542(new_n19890, new_n19886, new_n19891);
nor_5  g17543(new_n19549, new_n19471, new_n19892);
xor_4  g17544(new_n19549, new_n19471, new_n19893);
nor_5  g17545(new_n19551, new_n14689, new_n19894);
xnor_4 g17546(new_n19551, new_n14689, new_n19895);
nor_5  g17547(new_n15857, new_n14691, new_n19896);
nor_5  g17548(new_n15886, new_n15858, new_n19897);
or_5   g17549(new_n19897, new_n19896, new_n19898);
nor_5  g17550(new_n19898, new_n19895, new_n19899);
nor_5  g17551(new_n19899, new_n19894, new_n19900);
and_5  g17552(new_n19900, new_n19893, new_n19901);
nor_5  g17553(new_n19901, new_n19892, new_n19902);
xnor_4 g17554(new_n19902, new_n19891, n8803);
and_5  g17555(new_n18621, new_n5071, new_n19904);
nor_5  g17556(new_n18622, new_n18617, new_n19905_1);
nor_5  g17557(new_n18643, new_n18623, new_n19906);
nor_5  g17558(new_n19906, new_n19905_1, new_n19907);
xor_4  g17559(new_n19907, new_n19904, new_n19908);
nor_5  g17560(n16544, n4319, new_n19909_1);
nor_5  g17561(new_n14383, new_n14364_1, new_n19910);
nor_5  g17562(new_n19910, new_n19909_1, new_n19911_1);
xor_4  g17563(new_n19911_1, new_n19908, new_n19912);
nor_5  g17564(new_n18644, new_n14384, new_n19913);
nor_5  g17565(new_n18664, new_n18645, new_n19914);
nor_5  g17566(new_n19914, new_n19913, new_n19915);
xnor_4 g17567(new_n19915, new_n19912, new_n19916_1);
xnor_4 g17568(new_n19916_1, new_n7018, new_n19917);
nor_5  g17569(new_n18665, new_n7020, new_n19918);
nor_5  g17570(new_n19239, new_n19205, new_n19919);
nor_5  g17571(new_n19919, new_n19918, new_n19920);
xnor_4 g17572(new_n19920, new_n19917, n8809);
nor_5  g17573(new_n19889, new_n16238, new_n19922_1);
nor_5  g17574(new_n16556, n3324, new_n19923_1);
and_5  g17575(new_n19465, new_n19454_1, new_n19924);
or_5   g17576(new_n19924, new_n19923_1, new_n19925);
nor_5  g17577(new_n19925, new_n16552, new_n19926);
xor_4  g17578(new_n19926, new_n19922_1, new_n19927);
not_10 g17579(new_n19890, new_n19928);
xor_4  g17580(new_n19925, new_n16552, new_n19929);
nor_5  g17581(new_n19929, new_n19928, new_n19930_1);
xor_4  g17582(new_n19929, new_n19890, new_n19931);
and_5  g17583(new_n19471, new_n19466, new_n19932);
nor_5  g17584(new_n19485, new_n19472_1, new_n19933);
nor_5  g17585(new_n19933, new_n19932, new_n19934);
nor_5  g17586(new_n19934, new_n19931, new_n19935);
nor_5  g17587(new_n19935, new_n19930_1, new_n19936);
xnor_4 g17588(new_n19936, new_n19927, n8821);
xnor_4 g17589(new_n14138, new_n14136_1, n8824);
xor_4  g17590(new_n16191, new_n16190, n8849);
xnor_4 g17591(new_n12499, new_n12491, n8861);
xor_4  g17592(n22442, n8856, new_n19941_1);
not_10 g17593(n468, new_n19942);
nor_5  g17594(n14130, new_n19942, new_n19943);
nor_5  g17595(new_n18421, new_n18397, new_n19944);
nor_5  g17596(new_n19944, new_n19943, new_n19945);
xnor_4 g17597(new_n19945, new_n19941_1, new_n19946);
xnor_4 g17598(n3324, n2272, new_n19947);
nor_5  g17599(n25331, n17911, new_n19948);
nor_5  g17600(new_n18390, new_n18387, new_n19949);
nor_5  g17601(new_n19949, new_n19948, new_n19950);
xor_4  g17602(new_n19950, new_n19947, new_n19951);
xnor_4 g17603(new_n19951, new_n6809, new_n19952);
nor_5  g17604(new_n18391, new_n6803, new_n19953);
nor_5  g17605(new_n18395, new_n18392, new_n19954);
nor_5  g17606(new_n19954, new_n19953, new_n19955);
xnor_4 g17607(new_n19955, new_n19952, new_n19956);
xnor_4 g17608(new_n19956, new_n19946, new_n19957);
and_5  g17609(new_n18422, new_n18396, new_n19958);
nor_5  g17610(new_n18453, new_n18423, new_n19959);
nor_5  g17611(new_n19959, new_n19958, new_n19960);
xor_4  g17612(new_n19960, new_n19957, n8862);
xor_4  g17613(new_n12393, new_n12392, n8884);
xor_4  g17614(new_n17399, new_n16631, n8909);
xnor_4 g17615(new_n10568, new_n10527, n8911);
xnor_4 g17616(new_n10090, new_n10089, n8971);
xnor_4 g17617(new_n19632, new_n19609, n8982);
xnor_4 g17618(new_n5012, new_n4996, n8993);
xor_4  g17619(new_n13037, new_n13036, n9012);
nor_5  g17620(new_n18543, new_n18540, new_n19969);
or_5   g17621(new_n18546, new_n18545, new_n19970);
or_5   g17622(new_n18549, new_n4135, new_n19971);
nor_5  g17623(new_n19971, new_n19970, new_n19972);
xnor_4 g17624(new_n19972, new_n19969, new_n19973);
and_5  g17625(new_n18551, new_n18544, new_n19974);
nor_5  g17626(new_n18597, new_n18552, new_n19975);
nor_5  g17627(new_n19975, new_n19974, new_n19976);
xnor_4 g17628(new_n19976, new_n19973, n9032);
xor_4  g17629(new_n14623, new_n14622, n9042);
xnor_4 g17630(new_n15837, new_n15811, n9046);
xnor_4 g17631(new_n7455, new_n7404, n9047);
xnor_4 g17632(new_n13872, new_n13871, n9104);
nor_5  g17633(new_n18913, new_n18905, new_n19982);
nor_5  g17634(new_n19982, new_n19524, new_n19983);
and_5  g17635(new_n18913, new_n18905, new_n19984);
nor_5  g17636(new_n19984, new_n14010, new_n19985);
nor_5  g17637(new_n19985, new_n19983, new_n19986);
xnor_4 g17638(new_n19986, new_n17855_1, new_n19987);
nor_5  g17639(new_n18915, new_n17855_1, new_n19988_1);
nor_5  g17640(new_n18924, new_n18916, new_n19989);
or_5   g17641(new_n19989, new_n19988_1, new_n19990);
xor_4  g17642(new_n19990, new_n19987, n9129);
xnor_4 g17643(new_n17585, new_n17552, n9146);
xor_4  g17644(new_n7846, new_n6082, n9164);
xor_4  g17645(new_n11594, new_n11593, n9166);
xnor_4 g17646(new_n16568, new_n16545, new_n19995);
xnor_4 g17647(new_n19995, new_n16579, n9182);
xnor_4 g17648(new_n6494, new_n6464, n9191);
xnor_4 g17649(new_n10573, new_n10519, n9217);
xor_4  g17650(new_n14779, new_n14778, n9220);
xnor_4 g17651(new_n17575, new_n17569, n9261);
xor_4  g17652(n22626, n3324, new_n20001);
not_10 g17653(n17911, new_n20002);
nor_5  g17654(new_n20002, n14440, new_n20003);
nor_5  g17655(new_n17204, new_n17180, new_n20004_1);
nor_5  g17656(new_n20004_1, new_n20003, new_n20005);
xor_4  g17657(new_n20005, new_n20001, new_n20006);
and_5  g17658(new_n20006, new_n16572, new_n20007);
xnor_4 g17659(new_n20006, new_n16572, new_n20008);
and_5  g17660(new_n17205, new_n2916, new_n20009);
nor_5  g17661(new_n17233, new_n17206, new_n20010);
nor_5  g17662(new_n20010, new_n20009, new_n20011);
nor_5  g17663(new_n20011, new_n20008, new_n20012);
nor_5  g17664(new_n20012, new_n20007, new_n20013_1);
not_10 g17665(new_n16568, new_n20014);
not_10 g17666(n3324, new_n20015);
nor_5  g17667(n22626, new_n20015, new_n20016);
nor_5  g17668(new_n20005, new_n20001, new_n20017_1);
nor_5  g17669(new_n20017_1, new_n20016, new_n20018);
xnor_4 g17670(new_n20018, new_n20014, new_n20019);
xnor_4 g17671(new_n20019, new_n20013_1, n9287);
xor_4  g17672(new_n12876, new_n12866, n9308);
xnor_4 g17673(new_n4642, new_n4604, n9344);
xnor_4 g17674(new_n3504, new_n3488, n9364);
or_5   g17675(new_n20018, new_n20014, new_n20024);
nor_5  g17676(new_n20024, new_n20013_1, new_n20025);
and_5  g17677(new_n20025, new_n16565, new_n20026);
and_5  g17678(new_n20018, new_n20014, new_n20027);
and_5  g17679(new_n20027, new_n20013_1, new_n20028);
and_5  g17680(new_n20028, new_n16566, new_n20029);
or_5   g17681(new_n20029, new_n20026, n9371);
xor_4  g17682(new_n9242, new_n9241, n9382);
xor_4  g17683(new_n19670, new_n19661, n9403);
xnor_4 g17684(new_n11600, new_n11578, n9419);
xnor_4 g17685(new_n19435, new_n19409, n9423);
xnor_4 g17686(new_n17229, new_n17213, n9430);
xor_4  g17687(n25120, n23272, new_n20036_1);
nor_5  g17688(n11481, new_n6974, new_n20037);
xor_4  g17689(n11481, n8363, new_n20038);
nor_5  g17690(n16439, new_n6977, new_n20039);
nor_5  g17691(new_n14303, new_n14300, new_n20040_1);
nor_5  g17692(new_n20040_1, new_n20039, new_n20041);
nor_5  g17693(new_n20041, new_n20038, new_n20042);
nor_5  g17694(new_n20042, new_n20037, new_n20043);
xor_4  g17695(new_n20043, new_n20036_1, new_n20044);
xor_4  g17696(new_n20044, new_n15732, new_n20045);
xor_4  g17697(new_n20041, new_n20038, new_n20046);
not_10 g17698(new_n20046, new_n20047);
nor_5  g17699(new_n20047, new_n15734, new_n20048);
xor_4  g17700(new_n20046, new_n15734, new_n20049);
not_10 g17701(new_n14304, new_n20050);
nor_5  g17702(new_n14309, new_n20050, new_n20051);
nor_5  g17703(new_n14314, new_n14310_1, new_n20052);
nor_5  g17704(new_n20052, new_n20051, new_n20053);
nor_5  g17705(new_n20053, new_n20049, new_n20054);
nor_5  g17706(new_n20054, new_n20048, new_n20055);
xnor_4 g17707(new_n20055, new_n20045, new_n20056);
xnor_4 g17708(new_n20056, new_n15798, new_n20057);
xor_4  g17709(new_n20053, new_n20049, new_n20058);
nor_5  g17710(new_n20058, new_n15800, new_n20059);
xnor_4 g17711(new_n20058, new_n15800, new_n20060);
nor_5  g17712(new_n15804, new_n14315, new_n20061_1);
xnor_4 g17713(new_n15804, new_n14315, new_n20062);
xor_4  g17714(new_n15791, new_n15777, new_n20063);
and_5  g17715(new_n20063, new_n9635_1, new_n20064);
xnor_4 g17716(new_n20063, new_n9635_1, new_n20065);
nor_5  g17717(new_n15813, new_n9637, new_n20066);
xor_4  g17718(new_n15813, new_n9637, new_n20067);
nor_5  g17719(new_n15816_1, new_n9640, new_n20068);
and_5  g17720(new_n13618, new_n9643, new_n20069_1);
nor_5  g17721(new_n13631, new_n13619, new_n20070);
nor_5  g17722(new_n20070, new_n20069_1, new_n20071);
xnor_4 g17723(new_n15816_1, new_n9640, new_n20072);
nor_5  g17724(new_n20072, new_n20071, new_n20073);
nor_5  g17725(new_n20073, new_n20068, new_n20074);
and_5  g17726(new_n20074, new_n20067, new_n20075);
nor_5  g17727(new_n20075, new_n20066, new_n20076);
nor_5  g17728(new_n20076, new_n20065, new_n20077_1);
nor_5  g17729(new_n20077_1, new_n20064, new_n20078);
nor_5  g17730(new_n20078, new_n20062, new_n20079);
nor_5  g17731(new_n20079, new_n20061_1, new_n20080);
nor_5  g17732(new_n20080, new_n20060, new_n20081);
or_5   g17733(new_n20081, new_n20059, new_n20082);
xor_4  g17734(new_n20082, new_n20057, n9435);
xnor_4 g17735(new_n14727, new_n14698, n9451);
xor_4  g17736(n12657, n10763, new_n20085);
nor_5  g17737(n17077, new_n15224, new_n20086_1);
nor_5  g17738(new_n17698, new_n17691, new_n20087);
nor_5  g17739(new_n20087, new_n20086_1, new_n20088);
xor_4  g17740(new_n20088, new_n20085, new_n20089);
xnor_4 g17741(new_n20089, new_n18396, new_n20090);
nor_5  g17742(new_n17720, new_n17699, new_n20091);
and_5  g17743(new_n17730, new_n17721_1, new_n20092);
nor_5  g17744(new_n20092, new_n20091, new_n20093);
xnor_4 g17745(new_n20093, new_n20090, n9458);
nor_5  g17746(n12507, new_n16537, new_n20095);
xor_4  g17747(n12507, n11220, new_n20096_1);
nor_5  g17748(new_n16540, n15077, new_n20097);
nor_5  g17749(new_n13558, new_n13539, new_n20098);
nor_5  g17750(new_n20098, new_n20097, new_n20099);
nor_5  g17751(new_n20099, new_n20096_1, new_n20100);
nor_5  g17752(new_n20100, new_n20095, new_n20101);
not_10 g17753(new_n20101, new_n20102);
xnor_4 g17754(new_n20102, new_n19099, new_n20103_1);
xor_4  g17755(new_n20099, new_n20096_1, new_n20104);
nor_5  g17756(new_n20104, new_n19102, new_n20105);
xnor_4 g17757(new_n20104, new_n19102, new_n20106);
nor_5  g17758(new_n13559, new_n13538, new_n20107);
nor_5  g17759(new_n13590, new_n13560, new_n20108);
nor_5  g17760(new_n20108, new_n20107, new_n20109);
nor_5  g17761(new_n20109, new_n20106, new_n20110);
nor_5  g17762(new_n20110, new_n20105, new_n20111);
xnor_4 g17763(new_n20111, new_n20103_1, n9459);
xnor_4 g17764(new_n13820, new_n13819, n9508);
xnor_4 g17765(new_n11604, new_n11570, n9552);
xnor_4 g17766(new_n4245, new_n4244, n9556);
xor_4  g17767(new_n10064, new_n8028, n9558);
xor_4  g17768(new_n19301, new_n13029, n9616);
xnor_4 g17769(new_n7791, new_n7768, n9622);
xnor_4 g17770(new_n15216, new_n15202, n9626);
xnor_4 g17771(new_n4250, new_n4233, n9633);
nor_5  g17772(new_n6971_1, n23272, new_n20121);
nor_5  g17773(new_n20043, new_n20036_1, new_n20122);
nor_5  g17774(new_n20122, new_n20121, new_n20123);
and_5  g17775(new_n20123, new_n19643, new_n20124);
xnor_4 g17776(new_n20123, new_n19643, new_n20125);
not_10 g17777(new_n20044, new_n20126_1);
nor_5  g17778(new_n20126_1, new_n15732, new_n20127);
nor_5  g17779(new_n20055, new_n20045, new_n20128);
or_5   g17780(new_n20128, new_n20127, new_n20129);
nor_5  g17781(new_n20129, new_n20125, new_n20130);
nor_5  g17782(new_n20130, new_n20124, new_n20131);
and_5  g17783(new_n20131, new_n5117, new_n20132);
xnor_4 g17784(new_n20131, new_n5117, new_n20133);
xor_4  g17785(new_n20129, new_n20125, new_n20134);
nor_5  g17786(new_n20134, new_n5117, new_n20135);
xnor_4 g17787(new_n20134, new_n5117, new_n20136);
xor_4  g17788(new_n20055, new_n20045, new_n20137);
nor_5  g17789(new_n20137, new_n5118, new_n20138_1);
and_5  g17790(new_n20058, new_n5174, new_n20139);
xnor_4 g17791(new_n20058, new_n5174, new_n20140);
and_5  g17792(new_n14315, new_n5178, new_n20141);
nor_5  g17793(new_n14319, new_n14316, new_n20142);
nor_5  g17794(new_n20142, new_n20141, new_n20143);
nor_5  g17795(new_n20143, new_n20140, new_n20144);
nor_5  g17796(new_n20144, new_n20139, new_n20145);
xnor_4 g17797(new_n20056, new_n5118, new_n20146);
and_5  g17798(new_n20146, new_n20145, new_n20147);
or_5   g17799(new_n20147, new_n20138_1, new_n20148);
nor_5  g17800(new_n20148, new_n20136, new_n20149_1);
nor_5  g17801(new_n20149_1, new_n20135, new_n20150);
nor_5  g17802(new_n20150, new_n20133, new_n20151_1);
nor_5  g17803(new_n20151_1, new_n20132, n9635);
xnor_4 g17804(new_n17931_1, new_n17928, n9648);
xor_4  g17805(new_n4626, new_n4625, n9689);
xnor_4 g17806(new_n9802, new_n9784, n9695);
xnor_4 g17807(new_n6916, new_n6872, n9699);
xnor_4 g17808(new_n15302, new_n14733, new_n20157);
and_5  g17809(new_n14744, new_n14733, new_n20158);
nor_5  g17810(new_n14785, new_n14745, new_n20159);
or_5   g17811(new_n20159, new_n20158, new_n20160);
xor_4  g17812(new_n20160, new_n20157, n9726);
xnor_4 g17813(new_n12071, new_n9073, n9753);
xnor_4 g17814(new_n3227, new_n3210, n9761);
xnor_4 g17815(new_n9088, new_n9048, n9763);
xnor_4 g17816(new_n12390, new_n12388, n9767);
xor_4  g17817(new_n12545_1, new_n12296, n9771);
xor_4  g17818(new_n19748, new_n19745, n9778);
xnor_4 g17819(new_n14520, new_n14511, n9783);
xnor_4 g17820(new_n6117, new_n6115, n9803);
not_10 g17821(new_n3177, new_n20170);
and_5  g17822(new_n19244_1, new_n10599, new_n20171);
and_5  g17823(new_n20171, new_n10596, new_n20172);
not_10 g17824(new_n16517_1, new_n20173);
xnor_4 g17825(new_n20171, n4319, new_n20174);
and_5  g17826(new_n20174, new_n20173, new_n20175);
nor_5  g17827(new_n20174, new_n20173, new_n20176);
and_5  g17828(new_n19245, new_n16521_1, new_n20177);
nor_5  g17829(new_n19245, new_n16521_1, new_n20178);
and_5  g17830(new_n19247, new_n15359, new_n20179_1);
or_5   g17831(new_n19247, new_n15359, new_n20180);
nor_5  g17832(new_n19250, new_n15362, new_n20181);
and_5  g17833(new_n19253, new_n15365, new_n20182);
xnor_4 g17834(new_n19253, new_n15365, new_n20183);
and_5  g17835(new_n6075, new_n6060, new_n20184);
nor_5  g17836(new_n6101, new_n6076, new_n20185);
nor_5  g17837(new_n20185, new_n20184, new_n20186);
nor_5  g17838(new_n20186, new_n20183, new_n20187_1);
or_5   g17839(new_n20187_1, new_n20182, new_n20188);
xnor_4 g17840(new_n19250, new_n15362, new_n20189);
nor_5  g17841(new_n20189, new_n20188, new_n20190);
nor_5  g17842(new_n20190, new_n20181, new_n20191);
and_5  g17843(new_n20191, new_n20180, new_n20192);
nor_5  g17844(new_n20192, new_n20179_1, new_n20193);
nor_5  g17845(new_n20193, new_n20178, new_n20194);
nor_5  g17846(new_n20194, new_n20177, new_n20195);
nor_5  g17847(new_n20195, new_n20176, new_n20196);
nor_5  g17848(new_n20196, new_n20175, new_n20197);
xnor_4 g17849(new_n20197, new_n16513, new_n20198);
xor_4  g17850(new_n20198, new_n20172, new_n20199);
and_5  g17851(new_n20199, new_n20170, new_n20200);
xnor_4 g17852(new_n20199, new_n20170, new_n20201);
not_10 g17853(new_n3184, new_n20202);
xnor_4 g17854(new_n20174, new_n16517_1, new_n20203);
xnor_4 g17855(new_n20203, new_n20195, new_n20204);
nor_5  g17856(new_n20204, new_n20202, new_n20205);
xnor_4 g17857(new_n20204, new_n20202, new_n20206);
not_10 g17858(new_n3188, new_n20207);
xor_4  g17859(new_n19245, new_n16521_1, new_n20208);
xnor_4 g17860(new_n20208, new_n20193, new_n20209);
nor_5  g17861(new_n20209, new_n20207, new_n20210);
xnor_4 g17862(new_n20209, new_n20207, new_n20211);
not_10 g17863(new_n3192, new_n20212);
xnor_4 g17864(new_n19247, new_n15359, new_n20213_1);
xnor_4 g17865(new_n20213_1, new_n20191, new_n20214);
nor_5  g17866(new_n20214, new_n20212, new_n20215);
xnor_4 g17867(new_n20214, new_n20212, new_n20216);
xor_4  g17868(new_n20189, new_n20188, new_n20217);
and_5  g17869(new_n20217, new_n3196, new_n20218);
xnor_4 g17870(new_n20217, new_n3196, new_n20219);
not_10 g17871(new_n3200, new_n20220);
xor_4  g17872(new_n20186, new_n20183, new_n20221);
nor_5  g17873(new_n20221, new_n20220, new_n20222);
xnor_4 g17874(new_n20221, new_n20220, new_n20223);
nor_5  g17875(new_n6102, new_n6055, new_n20224);
nor_5  g17876(new_n6124, new_n6103, new_n20225);
nor_5  g17877(new_n20225, new_n20224, new_n20226);
nor_5  g17878(new_n20226, new_n20223, new_n20227);
nor_5  g17879(new_n20227, new_n20222, new_n20228);
nor_5  g17880(new_n20228, new_n20219, new_n20229);
nor_5  g17881(new_n20229, new_n20218, new_n20230);
nor_5  g17882(new_n20230, new_n20216, new_n20231);
nor_5  g17883(new_n20231, new_n20215, new_n20232);
nor_5  g17884(new_n20232, new_n20211, new_n20233);
nor_5  g17885(new_n20233, new_n20210, new_n20234);
nor_5  g17886(new_n20234, new_n20206, new_n20235_1);
nor_5  g17887(new_n20235_1, new_n20205, new_n20236);
nor_5  g17888(new_n20236, new_n20201, new_n20237);
or_5   g17889(new_n20237, new_n20200, new_n20238);
or_5   g17890(new_n20196, new_n20175, new_n20239);
nor_5  g17891(new_n20239, new_n16513, new_n20240);
xor_4  g17892(new_n20172, new_n16477, new_n20241);
and_5  g17893(new_n20241, new_n20240, new_n20242);
nor_5  g17894(new_n20241, new_n20197, new_n20243);
or_5   g17895(new_n20243, new_n20242, new_n20244);
nor_5  g17896(new_n20244, new_n20238, new_n20245);
or_5   g17897(new_n20172, new_n16477, new_n20246);
or_5   g17898(new_n20246, new_n20239, new_n20247);
xnor_4 g17899(new_n20247, new_n20245, n9833);
and_5  g17900(new_n15966, new_n7863, new_n20249);
and_5  g17901(new_n20249, new_n7860, new_n20250_1);
and_5  g17902(new_n20250_1, new_n15560, new_n20251);
or_5   g17903(new_n20251, new_n16510, new_n20252);
xnor_4 g17904(new_n20250_1, n25972, new_n20253);
and_5  g17905(new_n20253, new_n16491, new_n20254);
xnor_4 g17906(new_n20253, new_n16491, new_n20255);
xnor_4 g17907(new_n20249, n21915, new_n20256);
and_5  g17908(new_n20256, new_n16495, new_n20257);
xnor_4 g17909(new_n20256, new_n16495, new_n20258);
and_5  g17910(new_n15967_1, new_n15330, new_n20259_1);
nor_5  g17911(new_n15996, new_n15968, new_n20260);
nor_5  g17912(new_n20260, new_n20259_1, new_n20261);
nor_5  g17913(new_n20261, new_n20258, new_n20262);
nor_5  g17914(new_n20262, new_n20257, new_n20263);
nor_5  g17915(new_n20263, new_n20255, new_n20264);
or_5   g17916(new_n20264, new_n20254, new_n20265);
or_5   g17917(new_n20265, new_n20252, new_n20266);
nand_5 g17918(new_n15998, new_n9104_1, new_n20267);
nor_5  g17919(new_n20267, n15077, new_n20268);
and_5  g17920(new_n20268, new_n9098, new_n20269);
xnor_4 g17921(new_n20269, new_n15298, new_n20270);
xnor_4 g17922(new_n20268, n12507, new_n20271);
nor_5  g17923(new_n20271, new_n11759, new_n20272);
xnor_4 g17924(new_n20267, new_n9101, new_n20273);
nor_5  g17925(new_n20273, new_n4895, new_n20274);
xnor_4 g17926(new_n20273, new_n4895, new_n20275);
and_5  g17927(new_n15999, new_n4929, new_n20276);
nor_5  g17928(new_n16004, new_n16000, new_n20277);
or_5   g17929(new_n20277, new_n20276, new_n20278);
nor_5  g17930(new_n20278, new_n20275, new_n20279_1);
nor_5  g17931(new_n20279_1, new_n20274, new_n20280);
xnor_4 g17932(new_n20271, new_n11759, new_n20281);
nor_5  g17933(new_n20281, new_n20280, new_n20282);
nor_5  g17934(new_n20282, new_n20272, new_n20283);
xnor_4 g17935(new_n20283, new_n20270, new_n20284);
xor_4  g17936(new_n20251, new_n16510, new_n20285);
xnor_4 g17937(new_n20285, new_n20265, new_n20286);
nor_5  g17938(new_n20286, new_n20284, new_n20287_1);
xnor_4 g17939(new_n20286, new_n20284, new_n20288);
xnor_4 g17940(new_n20263, new_n20255, new_n20289);
xor_4  g17941(new_n20281, new_n20280, new_n20290);
and_5  g17942(new_n20290, new_n20289, new_n20291);
xnor_4 g17943(new_n20290, new_n20289, new_n20292);
nor_5  g17944(new_n20277, new_n20276, new_n20293);
xor_4  g17945(new_n20293, new_n20275, new_n20294);
xor_4  g17946(new_n20261, new_n20258, new_n20295);
nor_5  g17947(new_n20295, new_n20294, new_n20296);
xnor_4 g17948(new_n20295, new_n20294, new_n20297);
nor_5  g17949(new_n16005, new_n15997, new_n20298);
nor_5  g17950(new_n16040, new_n16006, new_n20299);
nor_5  g17951(new_n20299, new_n20298, new_n20300);
nor_5  g17952(new_n20300, new_n20297, new_n20301_1);
nor_5  g17953(new_n20301_1, new_n20296, new_n20302);
nor_5  g17954(new_n20302, new_n20292, new_n20303);
nor_5  g17955(new_n20303, new_n20291, new_n20304);
nor_5  g17956(new_n20304, new_n20288, new_n20305);
nor_5  g17957(new_n20305, new_n20287_1, new_n20306);
nor_5  g17958(new_n20306, new_n20266, new_n20307);
xor_4  g17959(new_n20306, new_n20266, new_n20308);
or_5   g17960(new_n20269, new_n14736, new_n20309);
nor_5  g17961(new_n20283, new_n20309, new_n20310);
not_10 g17962(new_n20310, new_n20311);
nor_5  g17963(new_n20311, new_n20308, new_n20312);
or_5   g17964(new_n20312, new_n20307, n9838);
xnor_4 g17965(new_n18075, new_n18072, n9867);
nor_5  g17966(new_n17659, new_n5231, new_n20315);
nor_5  g17967(new_n17663, new_n17660, new_n20316);
nor_5  g17968(new_n20316, new_n20315, new_n20317);
nor_5  g17969(new_n20317, new_n18863, new_n20318);
xnor_4 g17970(new_n20317, new_n18881, new_n20319);
nor_5  g17971(new_n20319, new_n7397, new_n20320);
nor_5  g17972(new_n17664_1, new_n17652, new_n20321);
nor_5  g17973(new_n17668, new_n17665, new_n20322);
or_5   g17974(new_n20322, new_n20321, new_n20323);
xor_4  g17975(new_n20319, new_n7397, new_n20324);
and_5  g17976(new_n20324, new_n20323, new_n20325);
nor_5  g17977(new_n20325, new_n20320, new_n20326);
nor_5  g17978(new_n20326, new_n20318, new_n20327);
nor_5  g17979(new_n20327, new_n7299, n9890);
xor_4  g17980(new_n16530, new_n16520, n9917);
xnor_4 g17981(new_n19127, new_n19120, n9919);
xnor_4 g17982(new_n16690, new_n16676, n9938);
xnor_4 g17983(new_n16353, new_n16352, n9946);
xnor_4 g17984(n21784, n3740, new_n20333_1);
nor_5  g17985(n5521, n2858, new_n20334);
xnor_4 g17986(n5521, n2858, new_n20335);
nor_5  g17987(n11926, n2659, new_n20336);
xnor_4 g17988(n11926, n2659, new_n20337);
nor_5  g17989(n24327, n4325, new_n20338);
xnor_4 g17990(n24327, n4325, new_n20339);
and_5  g17991(n22198, n5337, new_n20340);
or_5   g17992(n22198, n5337, new_n20341);
nor_5  g17993(n20826, n626, new_n20342);
nor_5  g17994(new_n11736_1, new_n11733, new_n20343);
nor_5  g17995(new_n20343, new_n20342, new_n20344);
and_5  g17996(new_n20344, new_n20341, new_n20345);
or_5   g17997(new_n20345, new_n20340, new_n20346);
nor_5  g17998(new_n20346, new_n20339, new_n20347);
nor_5  g17999(new_n20347, new_n20338, new_n20348);
nor_5  g18000(new_n20348, new_n20337, new_n20349_1);
nor_5  g18001(new_n20349_1, new_n20336, new_n20350);
nor_5  g18002(new_n20350, new_n20335, new_n20351);
nor_5  g18003(new_n20351, new_n20334, new_n20352);
xor_4  g18004(new_n20352, new_n20333_1, new_n20353);
xnor_4 g18005(new_n20353, new_n4476_1, new_n20354);
xor_4  g18006(new_n20350, new_n20335, new_n20355_1);
and_5  g18007(new_n20355_1, new_n4480, new_n20356);
xor_4  g18008(new_n20355_1, new_n4479, new_n20357);
xor_4  g18009(new_n20348, new_n20337, new_n20358);
and_5  g18010(new_n20358, new_n4484, new_n20359_1);
xor_4  g18011(new_n20346, new_n20339, new_n20360);
and_5  g18012(new_n20360, new_n4488, new_n20361);
xor_4  g18013(new_n20360, new_n4487, new_n20362);
xnor_4 g18014(n22198, n5337, new_n20363);
xnor_4 g18015(new_n20363, new_n20344, new_n20364);
nor_5  g18016(new_n20364, new_n4491, new_n20365);
nor_5  g18017(new_n11737, new_n11732, new_n20366_1);
and_5  g18018(new_n11738, new_n4495, new_n20367);
or_5   g18019(new_n20367, new_n20366_1, new_n20368);
xnor_4 g18020(new_n20364, new_n4491, new_n20369);
nor_5  g18021(new_n20369, new_n20368, new_n20370);
nor_5  g18022(new_n20370, new_n20365, new_n20371);
nor_5  g18023(new_n20371, new_n20362, new_n20372);
nor_5  g18024(new_n20372, new_n20361, new_n20373);
xor_4  g18025(new_n20358, new_n4483, new_n20374);
nor_5  g18026(new_n20374, new_n20373, new_n20375);
nor_5  g18027(new_n20375, new_n20359_1, new_n20376);
nor_5  g18028(new_n20376, new_n20357, new_n20377);
nor_5  g18029(new_n20377, new_n20356, new_n20378);
xor_4  g18030(new_n20378, new_n20354, new_n20379);
xnor_4 g18031(new_n20379, new_n15893, new_n20380);
xor_4  g18032(new_n20376, new_n20357, new_n20381);
and_5  g18033(new_n20381, new_n15269, new_n20382);
xnor_4 g18034(new_n20381, new_n15269, new_n20383);
xor_4  g18035(new_n20374, new_n20373, new_n20384);
and_5  g18036(new_n20384, new_n15271_1, new_n20385_1);
xnor_4 g18037(new_n20384, new_n15271_1, new_n20386);
xnor_4 g18038(new_n20371, new_n20362, new_n20387);
nor_5  g18039(new_n20387, new_n3551, new_n20388_1);
xor_4  g18040(new_n20387, new_n3551, new_n20389);
xor_4  g18041(new_n20369, new_n20368, new_n20390);
nor_5  g18042(new_n20390, new_n3554, new_n20391);
and_5  g18043(new_n11739, new_n3557, new_n20392);
nor_5  g18044(new_n11748, new_n11740, new_n20393);
nor_5  g18045(new_n20393, new_n20392, new_n20394);
xnor_4 g18046(new_n20390, new_n3554, new_n20395);
nor_5  g18047(new_n20395, new_n20394, new_n20396);
nor_5  g18048(new_n20396, new_n20391, new_n20397);
and_5  g18049(new_n20397, new_n20389, new_n20398);
nor_5  g18050(new_n20398, new_n20388_1, new_n20399);
nor_5  g18051(new_n20399, new_n20386, new_n20400);
nor_5  g18052(new_n20400, new_n20385_1, new_n20401);
nor_5  g18053(new_n20401, new_n20383, new_n20402_1);
or_5   g18054(new_n20402_1, new_n20382, new_n20403_1);
xor_4  g18055(new_n20403_1, new_n20380, n9968);
nor_5  g18056(new_n18812, new_n12594, new_n20405);
xnor_4 g18057(new_n18812, new_n12594, new_n20406);
nor_5  g18058(new_n18819, new_n12594, new_n20407);
xnor_4 g18059(new_n18822, new_n12594, new_n20408);
nor_5  g18060(new_n10233, new_n10173, new_n20409_1);
nor_5  g18061(new_n10274, new_n10234, new_n20410);
nor_5  g18062(new_n20410, new_n20409_1, new_n20411_1);
and_5  g18063(new_n20411_1, new_n20408, new_n20412);
or_5   g18064(new_n20412, new_n20407, new_n20413);
nor_5  g18065(new_n20413, new_n20406, new_n20414);
nor_5  g18066(new_n20414, new_n20405, n10009);
xnor_4 g18067(new_n19513, new_n19509, n10010);
and_5  g18068(new_n13382, new_n9971, new_n20417);
and_5  g18069(new_n13411, new_n13383, new_n20418);
nor_5  g18070(new_n20418, new_n20417, new_n20419);
not_10 g18071(new_n20419, new_n20420);
nor_5  g18072(new_n20420, new_n13448, new_n20421);
xnor_4 g18073(new_n20420, new_n13448, new_n20422);
and_5  g18074(new_n13448, new_n13412, new_n20423);
nor_5  g18075(new_n13485, new_n13449, new_n20424_1);
nor_5  g18076(new_n20424_1, new_n20423, new_n20425);
nor_5  g18077(new_n20425, new_n20422, new_n20426);
nor_5  g18078(new_n20426, new_n20421, n10019);
xnor_4 g18079(new_n13287, new_n13237, n10021);
xor_4  g18080(new_n8705, new_n8697, n10055);
xnor_4 g18081(new_n9659, new_n9639, n10101);
xnor_4 g18082(new_n4258, new_n4217, n10111);
nor_5  g18083(n16544, new_n20015, new_n20432);
xor_4  g18084(n16544, n3324, new_n20433);
nor_5  g18085(new_n20002, n6814, new_n20434);
xor_4  g18086(n17911, n6814, new_n20435);
nor_5  g18087(new_n17181, n19701, new_n20436_1);
xor_4  g18088(n21997, n19701, new_n20437);
nor_5  g18089(new_n17184, n23529, new_n20438);
xor_4  g18090(n25119, n23529, new_n20439);
nor_5  g18091(n24620, new_n17187, new_n20440);
xor_4  g18092(n24620, n1163, new_n20441_1);
nor_5  g18093(new_n17190, n5211, new_n20442);
or_5   g18094(n18537, new_n8162, new_n20443);
nor_5  g18095(new_n8165, n7057, new_n20444);
nor_5  g18096(new_n8611, new_n8600, new_n20445_1);
nor_5  g18097(new_n20445_1, new_n20444, new_n20446);
and_5  g18098(new_n20446, new_n20443, new_n20447);
nor_5  g18099(new_n20447, new_n20442, new_n20448);
nor_5  g18100(new_n20448, new_n20441_1, new_n20449);
nor_5  g18101(new_n20449, new_n20440, new_n20450_1);
nor_5  g18102(new_n20450_1, new_n20439, new_n20451);
nor_5  g18103(new_n20451, new_n20438, new_n20452);
nor_5  g18104(new_n20452, new_n20437, new_n20453);
nor_5  g18105(new_n20453, new_n20436_1, new_n20454);
nor_5  g18106(new_n20454, new_n20435, new_n20455_1);
nor_5  g18107(new_n20455_1, new_n20434, new_n20456);
nor_5  g18108(new_n20456, new_n20433, new_n20457);
nor_5  g18109(new_n20457, new_n20432, new_n20458);
xnor_4 g18110(new_n20458, new_n19659, new_n20459);
and_5  g18111(new_n20458, new_n19664_1, new_n20460);
nor_5  g18112(new_n20458, new_n19664_1, new_n20461);
xor_4  g18113(new_n15758, new_n15733, new_n20462);
xor_4  g18114(new_n20456, new_n20433, new_n20463);
nor_5  g18115(new_n20463, new_n20462, new_n20464);
xnor_4 g18116(new_n20463, new_n20462, new_n20465);
xor_4  g18117(new_n20454, new_n20435, new_n20466);
nor_5  g18118(new_n20466, new_n15801, new_n20467);
xnor_4 g18119(new_n20466, new_n15801, new_n20468);
xor_4  g18120(new_n20452, new_n20437, new_n20469);
nor_5  g18121(new_n20469, new_n15805, new_n20470_1);
xnor_4 g18122(new_n20469, new_n15805, new_n20471);
xor_4  g18123(new_n20450_1, new_n20439, new_n20472);
nor_5  g18124(new_n20472, new_n15809, new_n20473);
xnor_4 g18125(new_n20472, new_n15809, new_n20474);
xor_4  g18126(new_n20448, new_n20441_1, new_n20475);
nor_5  g18127(new_n20475, new_n15812_1, new_n20476);
xor_4  g18128(n18537, n5211, new_n20477);
xnor_4 g18129(new_n20477, new_n20446, new_n20478_1);
and_5  g18130(new_n20478_1, new_n15817, new_n20479);
xnor_4 g18131(new_n20478_1, new_n15817, new_n20480);
not_10 g18132(new_n8599, new_n20481);
nor_5  g18133(new_n8612, new_n20481, new_n20482);
nor_5  g18134(new_n8630, new_n8613, new_n20483);
nor_5  g18135(new_n20483, new_n20482, new_n20484);
nor_5  g18136(new_n20484, new_n20480, new_n20485);
nor_5  g18137(new_n20485, new_n20479, new_n20486);
xor_4  g18138(new_n20475, new_n15812_1, new_n20487);
and_5  g18139(new_n20487, new_n20486, new_n20488);
nor_5  g18140(new_n20488, new_n20476, new_n20489_1);
nor_5  g18141(new_n20489_1, new_n20474, new_n20490_1);
nor_5  g18142(new_n20490_1, new_n20473, new_n20491);
nor_5  g18143(new_n20491, new_n20471, new_n20492);
nor_5  g18144(new_n20492, new_n20470_1, new_n20493);
nor_5  g18145(new_n20493, new_n20468, new_n20494);
nor_5  g18146(new_n20494, new_n20467, new_n20495_1);
nor_5  g18147(new_n20495_1, new_n20465, new_n20496);
or_5   g18148(new_n20496, new_n20464, new_n20497);
nor_5  g18149(new_n20497, new_n20461, new_n20498);
nor_5  g18150(new_n20498, new_n20460, new_n20499);
xnor_4 g18151(new_n20499, new_n20459, n10165);
xnor_4 g18152(new_n11812, new_n11811, n10236);
xnor_4 g18153(new_n13165, new_n13141_1, n10239);
xnor_4 g18154(new_n5830, new_n5793, n10244);
xnor_4 g18155(new_n16623, new_n16611, n10261);
xnor_4 g18156(new_n14360, new_n14347, n10262);
xor_4  g18157(new_n15503, new_n15502, n10287);
nor_5  g18158(new_n19885, new_n13930, new_n20507);
xor_4  g18159(new_n19922_1, new_n20507, new_n20508);
nor_5  g18160(new_n19890, new_n19886, new_n20509);
nor_5  g18161(new_n19902, new_n19891, new_n20510);
nor_5  g18162(new_n20510, new_n20509, new_n20511);
xnor_4 g18163(new_n20511, new_n20508, n10295);
xnor_4 g18164(new_n13581, new_n13577, n10321);
xnor_4 g18165(new_n13167, new_n13138, n10326);
xor_4  g18166(new_n2751, new_n2741, n10327);
xnor_4 g18167(new_n18822, new_n18801, new_n20516);
xnor_4 g18168(new_n20516, new_n18816, n10330);
xnor_4 g18169(new_n19439, new_n19401_1, n10340);
xor_4  g18170(new_n15500, new_n15497, new_n20519);
xnor_4 g18171(new_n20519, new_n15504, n10345);
or_5   g18172(new_n4533, new_n4530, new_n20521);
and_5  g18173(new_n17621, new_n20521, new_n20522);
nor_5  g18174(new_n17624, new_n4534, new_n20523);
xnor_4 g18175(new_n17624, new_n4534, new_n20524);
and_5  g18176(new_n17628, new_n4537, new_n20525);
xnor_4 g18177(new_n17628, new_n4537, new_n20526);
xor_4  g18178(new_n4526, new_n4482, new_n20527);
and_5  g18179(new_n17632, new_n20527, new_n20528);
xnor_4 g18180(new_n17632, new_n20527, new_n20529);
xor_4  g18181(new_n4524, new_n4486, new_n20530);
and_5  g18182(new_n17636, new_n20530, new_n20531);
xnor_4 g18183(new_n17636, new_n20530, new_n20532);
nor_5  g18184(new_n8518, new_n4545, new_n20533_1);
xnor_4 g18185(new_n8518, new_n4545, new_n20534);
nor_5  g18186(new_n8521, new_n4548, new_n20535);
xnor_4 g18187(new_n8521, new_n4548, new_n20536);
nor_5  g18188(new_n8525, new_n4551, new_n20537);
xnor_4 g18189(new_n8525, new_n4551, new_n20538);
nor_5  g18190(new_n8529, new_n4554, new_n20539);
xnor_4 g18191(new_n8529, new_n4554, new_n20540);
nor_5  g18192(new_n8533, new_n4556, new_n20541);
xnor_4 g18193(new_n8533, new_n4556, new_n20542);
nor_5  g18194(new_n8539, new_n4562, new_n20543);
and_5  g18195(new_n20543, new_n8536, new_n20544);
not_10 g18196(new_n4559, new_n20545);
xnor_4 g18197(new_n20543, new_n18362_1, new_n20546);
and_5  g18198(new_n20546, new_n20545, new_n20547);
nor_5  g18199(new_n20547, new_n20544, new_n20548);
nor_5  g18200(new_n20548, new_n20542, new_n20549);
nor_5  g18201(new_n20549, new_n20541, new_n20550);
nor_5  g18202(new_n20550, new_n20540, new_n20551);
nor_5  g18203(new_n20551, new_n20539, new_n20552);
nor_5  g18204(new_n20552, new_n20538, new_n20553);
nor_5  g18205(new_n20553, new_n20537, new_n20554);
nor_5  g18206(new_n20554, new_n20536, new_n20555);
nor_5  g18207(new_n20555, new_n20535, new_n20556);
nor_5  g18208(new_n20556, new_n20534, new_n20557);
nor_5  g18209(new_n20557, new_n20533_1, new_n20558);
nor_5  g18210(new_n20558, new_n20532, new_n20559);
nor_5  g18211(new_n20559, new_n20531, new_n20560);
nor_5  g18212(new_n20560, new_n20529, new_n20561);
nor_5  g18213(new_n20561, new_n20528, new_n20562);
nor_5  g18214(new_n20562, new_n20526, new_n20563);
nor_5  g18215(new_n20563, new_n20525, new_n20564);
nor_5  g18216(new_n20564, new_n20524, new_n20565);
or_5   g18217(new_n20565, new_n20523, new_n20566);
xnor_4 g18218(new_n17621, new_n20521, new_n20567);
nor_5  g18219(new_n20567, new_n20566, new_n20568);
nor_5  g18220(new_n20568, new_n20522, n10356);
xor_4  g18221(new_n18163, new_n18162, n10385);
nor_5  g18222(new_n18383, new_n17621, new_n20571);
nand_5 g18223(new_n18383, new_n17621, new_n20572);
and_5  g18224(new_n20572, new_n18324, new_n20573);
nor_5  g18225(new_n20573, new_n20571, new_n20574);
nor_5  g18226(new_n20574, new_n18322, n10387);
xnor_4 g18227(new_n18585, new_n18571, n10388);
xnor_4 g18228(new_n14148_1, new_n14107_1, n10390);
xor_4  g18229(new_n8620_1, new_n8619, n10404);
xnor_4 g18230(new_n14518, new_n14515, n10409);
xnor_4 g18231(new_n14715, new_n7781, n10420);
xnor_4 g18232(new_n16616, new_n6288, n10432);
xnor_4 g18233(new_n19606, new_n18932, new_n20582_1);
nor_5  g18234(new_n18936, new_n8742, new_n20583);
nor_5  g18235(new_n19193, new_n19185, new_n20584);
nor_5  g18236(new_n20584, new_n20583, new_n20585);
xor_4  g18237(new_n20585, new_n20582_1, new_n20586);
xnor_4 g18238(new_n20586, new_n10374, new_n20587);
and_5  g18239(new_n19194, new_n10378, new_n20588);
nor_5  g18240(new_n19203, new_n19195, new_n20589);
nor_5  g18241(new_n20589, new_n20588, new_n20590_1);
xor_4  g18242(new_n20590_1, new_n20587, n10484);
xnor_4 g18243(new_n10263, new_n10250_1, n10489);
xnor_4 g18244(new_n12213, new_n3442, n10525);
xnor_4 g18245(new_n16020, new_n10960, new_n20594);
xnor_4 g18246(new_n20594, new_n16029_1, n10540);
xnor_4 g18247(new_n14631, new_n14607, n10561);
xnor_4 g18248(new_n14152, new_n14099, n10564);
xor_4  g18249(new_n9073, new_n9072, n10588);
xnor_4 g18250(new_n9076, new_n9075, n10595);
xor_4  g18251(new_n19306, new_n19293, n10617);
xnor_4 g18252(new_n11290_1, new_n11236, n10628);
xor_4  g18253(new_n9613, new_n5269, new_n20602_1);
nor_5  g18254(new_n9618, new_n5272, new_n20603);
xnor_4 g18255(new_n9618, new_n5272, new_n20604_1);
and_5  g18256(new_n9621, new_n5276, new_n20605);
xnor_4 g18257(new_n9621, new_n5276, new_n20606);
or_5   g18258(new_n5310, new_n5281, new_n20607);
and_5  g18259(new_n20607, new_n5318, new_n20608);
xor_4  g18260(new_n20607, new_n5318, new_n20609_1);
and_5  g18261(new_n20609_1, new_n5287, new_n20610);
nor_5  g18262(new_n20610, new_n20608, new_n20611);
nor_5  g18263(new_n20611, new_n20606, new_n20612);
nor_5  g18264(new_n20612, new_n20605, new_n20613);
nor_5  g18265(new_n20613, new_n20604_1, new_n20614);
nor_5  g18266(new_n20614, new_n20603, new_n20615);
xnor_4 g18267(new_n20615, new_n20602_1, n10647);
or_5   g18268(new_n7571, new_n7570, new_n20617);
or_5   g18269(new_n7578, new_n20617, new_n20618);
and_5  g18270(new_n3406, new_n3396, new_n20619);
nor_5  g18271(new_n3461, new_n3407, new_n20620);
or_5   g18272(new_n20620, new_n18063, new_n20621);
or_5   g18273(new_n20621, new_n20619, new_n20622);
nor_5  g18274(new_n20622, new_n12182, new_n20623_1);
xnor_4 g18275(new_n20623_1, new_n20618, new_n20624);
xor_4  g18276(new_n7578, new_n7572_1, new_n20625);
xor_4  g18277(new_n20622, new_n12182, new_n20626);
nor_5  g18278(new_n20626, new_n20625, new_n20627);
nor_5  g18279(new_n3462, new_n3351, new_n20628);
nor_5  g18280(new_n3516_1, new_n3463, new_n20629_1);
or_5   g18281(new_n20629_1, new_n20628, new_n20630);
xnor_4 g18282(new_n20626, new_n20625, new_n20631);
nor_5  g18283(new_n20631, new_n20630, new_n20632);
nor_5  g18284(new_n20632, new_n20627, new_n20633);
xnor_4 g18285(new_n20633, new_n20624, n10653);
xor_4  g18286(new_n8229, new_n8228, n10692);
xor_4  g18287(new_n13336, new_n3997, n10694);
xnor_4 g18288(new_n18451, new_n18426, n10701);
xnor_4 g18289(new_n5610, new_n5595, n10756);
not_10 g18290(n6659, new_n20639);
nor_5  g18291(new_n20639, n5101, new_n20640);
nor_5  g18292(new_n14487, new_n14483, new_n20641);
nor_5  g18293(new_n20641, new_n20640, new_n20642);
not_10 g18294(new_n20642, new_n20643);
not_10 g18295(n13419, new_n20644);
and_5  g18296(new_n14488, new_n20644, new_n20645);
nor_5  g18297(new_n14488, new_n20644, new_n20646);
not_10 g18298(n4967, new_n20647);
and_5  g18299(new_n14440_1, new_n20647, new_n20648);
nor_5  g18300(new_n14440_1, new_n20647, new_n20649);
or_5   g18301(new_n17546, new_n17543, new_n20650);
nor_5  g18302(new_n20650, new_n20649, new_n20651);
nor_5  g18303(new_n20651, new_n20648, new_n20652);
nor_5  g18304(new_n20652, new_n20646, new_n20653);
nor_5  g18305(new_n20653, new_n20645, new_n20654);
and_5  g18306(new_n20654, new_n20643, new_n20655);
xnor_4 g18307(new_n20655, new_n3053, new_n20656);
xnor_4 g18308(new_n20654, new_n20642, new_n20657);
and_5  g18309(new_n20657, new_n3179, new_n20658_1);
xnor_4 g18310(new_n20657, new_n3179, new_n20659);
xnor_4 g18311(new_n20652, new_n14489, new_n20660);
nor_5  g18312(new_n20660, new_n3071, new_n20661_1);
xnor_4 g18313(new_n20660, new_n3071, new_n20662);
nor_5  g18314(new_n17548, new_n3078, new_n20663);
nor_5  g18315(new_n17587, new_n17549, new_n20664);
or_5   g18316(new_n20664, new_n20663, new_n20665);
nor_5  g18317(new_n20665, new_n20662, new_n20666);
nor_5  g18318(new_n20666, new_n20661_1, new_n20667);
nor_5  g18319(new_n20667, new_n20659, new_n20668);
nor_5  g18320(new_n20668, new_n20658_1, new_n20669);
xnor_4 g18321(new_n20669, new_n20656, n10775);
xnor_4 g18322(new_n19225, new_n19220_1, n10780);
xnor_4 g18323(n17095, n1689, new_n20672);
nor_5  g18324(n22591, n22274, new_n20673_1);
and_5  g18325(n26167, n24129, new_n20674);
xnor_4 g18326(n22591, n22274, new_n20675);
nor_5  g18327(new_n20675, new_n20674, new_n20676);
nor_5  g18328(new_n20676, new_n20673_1, new_n20677);
xor_4  g18329(new_n20677, new_n20672, new_n20678_1);
xnor_4 g18330(new_n20678_1, n21749, new_n20679);
and_5  g18331(new_n8105, n21138, new_n20680_1);
nor_5  g18332(new_n20680_1, n7769, new_n20681);
xor_4  g18333(new_n20675, new_n20674, new_n20682);
xnor_4 g18334(new_n20680_1, n7769, new_n20683);
nor_5  g18335(new_n20683, new_n20682, new_n20684);
nor_5  g18336(new_n20684, new_n20681, new_n20685_1);
xnor_4 g18337(new_n20685_1, new_n20679, new_n20686);
xnor_4 g18338(new_n20686, new_n16782, new_n20687);
xor_4  g18339(new_n20683, new_n20682, new_n20688);
and_5  g18340(new_n20688, new_n16785, new_n20689);
nand_5 g18341(new_n8106, new_n8104, new_n20690);
xnor_4 g18342(new_n20688, new_n16785, new_n20691_1);
nor_5  g18343(new_n20691_1, new_n20690, new_n20692);
nor_5  g18344(new_n20692, new_n20689, new_n20693);
xor_4  g18345(new_n20693, new_n20687, n10817);
and_5  g18346(new_n19911_1, new_n19908, new_n20695);
and_5  g18347(new_n19907, new_n19904, new_n20696_1);
nor_5  g18348(new_n19911_1, new_n19908, new_n20697);
nor_5  g18349(new_n19915, new_n20697, new_n20698);
or_5   g18350(new_n20698, new_n20696_1, new_n20699);
nor_5  g18351(new_n20699, new_n20695, new_n20700_1);
nor_5  g18352(new_n20700_1, new_n7018, new_n20701);
nor_5  g18353(new_n19916_1, new_n7018, new_n20702);
nor_5  g18354(new_n19920, new_n19917, new_n20703);
or_5   g18355(new_n20703, new_n20702, new_n20704_1);
xnor_4 g18356(new_n20700_1, new_n7018, new_n20705_1);
nor_5  g18357(new_n20705_1, new_n20704_1, new_n20706);
nor_5  g18358(new_n20706, new_n20701, n10834);
xor_4  g18359(new_n20150, new_n20133, n10851);
xnor_4 g18360(new_n19707, new_n19698, n10874);
xor_4  g18361(new_n20326, new_n20318, new_n20710);
xnor_4 g18362(new_n20710, new_n7299, n10924);
nor_5  g18363(new_n10036, new_n10033, new_n20712);
nor_5  g18364(new_n10092, new_n10037, new_n20713_1);
nor_5  g18365(new_n20713_1, new_n20712, n10943);
xnor_4 g18366(new_n10761, new_n10729, n10961);
xnor_4 g18367(new_n9568, new_n9557_1, n11005);
xnor_4 g18368(new_n19483, new_n19475, n11023);
nor_5  g18369(new_n16480, new_n6590_1, new_n20718);
xnor_4 g18370(new_n16480, new_n6590_1, new_n20719);
nor_5  g18371(new_n16482_1, new_n6594, new_n20720);
xnor_4 g18372(new_n16482_1, new_n6594, new_n20721);
and_5  g18373(new_n15317, new_n6598, new_n20722_1);
xnor_4 g18374(new_n15317, new_n6598, new_n20723_1);
and_5  g18375(new_n10920, new_n6602, new_n20724);
nor_5  g18376(new_n10945, new_n10921, new_n20725);
nor_5  g18377(new_n20725, new_n20724, new_n20726);
nor_5  g18378(new_n20726, new_n20723_1, new_n20727);
or_5   g18379(new_n20727, new_n20722_1, new_n20728);
nor_5  g18380(new_n20728, new_n20721, new_n20729);
nor_5  g18381(new_n20729, new_n20720, new_n20730);
nor_5  g18382(new_n20730, new_n20719, new_n20731);
nor_5  g18383(new_n20731, new_n20718, new_n20732);
or_5   g18384(new_n20732, new_n6573, new_n20733);
or_5   g18385(new_n20733, new_n16505, new_n20734);
xor_4  g18386(new_n20283, new_n20270, new_n20735);
xnor_4 g18387(new_n20732, new_n6573, new_n20736);
xnor_4 g18388(new_n20736, new_n16505, new_n20737);
and_5  g18389(new_n20737, new_n20735, new_n20738);
xnor_4 g18390(new_n20737, new_n20735, new_n20739);
xor_4  g18391(new_n20730, new_n20719, new_n20740);
and_5  g18392(new_n20740, new_n20290, new_n20741);
xnor_4 g18393(new_n20740, new_n20290, new_n20742);
xnor_4 g18394(new_n20293, new_n20275, new_n20743);
xor_4  g18395(new_n20728, new_n20721, new_n20744);
and_5  g18396(new_n20744, new_n20743, new_n20745);
xnor_4 g18397(new_n20744, new_n20743, new_n20746);
xor_4  g18398(new_n20726, new_n20723_1, new_n20747);
nor_5  g18399(new_n20747, new_n16005, new_n20748_1);
xnor_4 g18400(new_n20747, new_n16005, new_n20749);
nor_5  g18401(new_n10946, new_n10917, new_n20750);
nor_5  g18402(new_n10982, new_n10947, new_n20751);
nor_5  g18403(new_n20751, new_n20750, new_n20752);
nor_5  g18404(new_n20752, new_n20749, new_n20753);
nor_5  g18405(new_n20753, new_n20748_1, new_n20754);
nor_5  g18406(new_n20754, new_n20746, new_n20755);
nor_5  g18407(new_n20755, new_n20745, new_n20756);
nor_5  g18408(new_n20756, new_n20742, new_n20757);
nor_5  g18409(new_n20757, new_n20741, new_n20758);
nor_5  g18410(new_n20758, new_n20739, new_n20759);
nor_5  g18411(new_n20759, new_n20738, new_n20760);
nor_5  g18412(new_n20760, new_n20734, new_n20761_1);
xor_4  g18413(new_n20760, new_n20734, new_n20762);
nor_5  g18414(new_n20762, new_n20311, new_n20763);
or_5   g18415(new_n20763, new_n20761_1, n11025);
xnor_4 g18416(new_n14959, new_n7860, new_n20765);
nor_5  g18417(new_n14962, new_n7863, new_n20766);
xnor_4 g18418(new_n14962, new_n7863, new_n20767);
nor_5  g18419(new_n14965, new_n7866, new_n20768);
xnor_4 g18420(new_n14965, new_n7866, new_n20769);
nor_5  g18421(new_n14968, new_n7869, new_n20770);
nor_5  g18422(new_n17422, new_n17419, new_n20771);
nor_5  g18423(new_n20771, new_n20770, new_n20772);
nor_5  g18424(new_n20772, new_n20769, new_n20773);
nor_5  g18425(new_n20773, new_n20768, new_n20774_1);
nor_5  g18426(new_n20774_1, new_n20767, new_n20775);
nor_5  g18427(new_n20775, new_n20766, new_n20776);
xnor_4 g18428(new_n20776, new_n20765, new_n20777);
or_5   g18429(new_n17424, n26752, new_n20778);
or_5   g18430(new_n20778, n4590, new_n20779);
or_5   g18431(new_n20779, n25464, new_n20780);
xor_4  g18432(new_n20780, n3795, new_n20781);
xnor_4 g18433(new_n20781, new_n7992_1, new_n20782);
xor_4  g18434(new_n20779, n25464, new_n20783);
nor_5  g18435(new_n20783, new_n7997, new_n20784);
xnor_4 g18436(new_n20783, new_n7997, new_n20785);
xor_4  g18437(new_n20778, n4590, new_n20786);
nor_5  g18438(new_n20786, new_n8002, new_n20787);
xnor_4 g18439(new_n20786, new_n8002, new_n20788_1);
nor_5  g18440(new_n17425, new_n10054, new_n20789);
nor_5  g18441(new_n17429, new_n17426, new_n20790);
nor_5  g18442(new_n20790, new_n20789, new_n20791);
nor_5  g18443(new_n20791, new_n20788_1, new_n20792);
nor_5  g18444(new_n20792, new_n20787, new_n20793);
nor_5  g18445(new_n20793, new_n20785, new_n20794_1);
nor_5  g18446(new_n20794_1, new_n20784, new_n20795_1);
xor_4  g18447(new_n20795_1, new_n20782, new_n20796);
xnor_4 g18448(new_n20796, new_n20777, new_n20797);
xnor_4 g18449(new_n20774_1, new_n20767, new_n20798);
xor_4  g18450(new_n20793, new_n20785, new_n20799);
and_5  g18451(new_n20799, new_n20798, new_n20800);
xnor_4 g18452(new_n20799, new_n20798, new_n20801);
xnor_4 g18453(new_n20772, new_n20769, new_n20802);
xor_4  g18454(new_n20791, new_n20788_1, new_n20803_1);
and_5  g18455(new_n20803_1, new_n20802, new_n20804);
xnor_4 g18456(new_n20803_1, new_n20802, new_n20805);
and_5  g18457(new_n17430, new_n17423, new_n20806);
nor_5  g18458(new_n17434, new_n17431, new_n20807);
nor_5  g18459(new_n20807, new_n20806, new_n20808);
nor_5  g18460(new_n20808, new_n20805, new_n20809);
nor_5  g18461(new_n20809, new_n20804, new_n20810);
nor_5  g18462(new_n20810, new_n20801, new_n20811);
nor_5  g18463(new_n20811, new_n20800, new_n20812);
xnor_4 g18464(new_n20812, new_n20797, n11063);
xnor_4 g18465(new_n18583_1, new_n18574_1, n11078);
xnor_4 g18466(new_n19227, new_n19218, n11080);
xnor_4 g18467(new_n12501, new_n12487, n11094);
xnor_4 g18468(new_n20487, new_n20486, n11101);
xnor_4 g18469(new_n19299, new_n13023, new_n20818);
xnor_4 g18470(new_n20818, new_n19302, n11103);
xnor_4 g18471(new_n5979, new_n5955, n11120);
xor_4  g18472(new_n4632, new_n4629, n11127);
xnor_4 g18473(new_n13584, new_n13583, n11132);
xnor_4 g18474(new_n10085, new_n10045, n11134);
xnor_4 g18475(new_n3500, new_n3499, n11138);
xnor_4 g18476(new_n9473, new_n9463, n11182);
xnor_4 g18477(new_n12511, new_n12467_1, n11234);
xnor_4 g18478(new_n19886, new_n16943, new_n20827);
nor_5  g18479(new_n19549, new_n16948, new_n20828);
nor_5  g18480(new_n19571, new_n19550, new_n20829);
nor_5  g18481(new_n20829, new_n20828, new_n20830);
xnor_4 g18482(new_n20830, new_n20827, n11245);
xnor_4 g18483(new_n7855, new_n7843, n11261);
xnor_4 g18484(new_n20810, new_n20801, n11275);
or_5   g18485(new_n12235_1, new_n12177, n11290);
xnor_4 g18486(new_n8543, new_n8542, n11313);
xnor_4 g18487(new_n15297, new_n14744, new_n20836);
xnor_4 g18488(new_n20836, new_n15309, n11325);
xnor_4 g18489(new_n12551, new_n12550, n11326);
xnor_4 g18490(new_n15512, new_n15484, n11330);
xnor_4 g18491(new_n10079, new_n10055_1, n11347);
xnor_4 g18492(new_n20548, new_n20542, n11348);
xnor_4 g18493(new_n13690, new_n13682, n11352);
not_10 g18494(n22442, new_n20843);
nor_5  g18495(new_n20843, n3324, new_n20844);
xor_4  g18496(n22442, n3324, new_n20845);
nor_5  g18497(n17911, new_n19942, new_n20846);
nor_5  g18498(n21997, new_n18398, new_n20847);
nor_5  g18499(new_n15700, new_n15691, new_n20848);
nor_5  g18500(new_n20848, new_n20847, new_n20849);
xor_4  g18501(n17911, n468, new_n20850);
nor_5  g18502(new_n20850, new_n20849, new_n20851);
nor_5  g18503(new_n20851, new_n20846, new_n20852);
nor_5  g18504(new_n20852, new_n20845, new_n20853);
or_5   g18505(new_n20853, new_n20844, new_n20854);
nor_5  g18506(new_n16174, new_n16168, new_n20855);
nor_5  g18507(new_n20855, new_n6970, new_n20856);
nand_5 g18508(new_n16174, new_n16168, new_n20857);
and_5  g18509(new_n20857, new_n6970, new_n20858);
nor_5  g18510(new_n20858, new_n20856, new_n20859);
xnor_4 g18511(new_n20859, new_n20854, new_n20860);
nor_5  g18512(new_n20854, new_n16176, new_n20861);
and_5  g18513(new_n20854, new_n16176, new_n20862);
xor_4  g18514(new_n20852, new_n20845, new_n20863);
nor_5  g18515(new_n20863, new_n16178, new_n20864);
xor_4  g18516(new_n20863, new_n16178, new_n20865);
xor_4  g18517(new_n20850, new_n20849, new_n20866);
and_5  g18518(new_n20866, new_n16180, new_n20867);
xnor_4 g18519(new_n20866, new_n16180, new_n20868);
and_5  g18520(new_n15701, new_n15690, new_n20869_1);
nor_5  g18521(new_n15712, new_n15702, new_n20870);
nor_5  g18522(new_n20870, new_n20869_1, new_n20871);
nor_5  g18523(new_n20871, new_n20868, new_n20872);
nor_5  g18524(new_n20872, new_n20867, new_n20873);
and_5  g18525(new_n20873, new_n20865, new_n20874);
or_5   g18526(new_n20874, new_n20864, new_n20875);
nor_5  g18527(new_n20875, new_n20862, new_n20876);
nor_5  g18528(new_n20876, new_n20861, new_n20877);
xnor_4 g18529(new_n20877, new_n20860, n11375);
xor_4  g18530(new_n11321, new_n6484, n11379);
not_10 g18531(n10250, new_n20880);
nor_5  g18532(new_n20880, n2570, new_n20881);
nor_5  g18533(new_n14956, new_n14923, new_n20882);
nor_5  g18534(new_n20882, new_n20881, new_n20883);
xnor_4 g18535(new_n20883, new_n10819, new_n20884);
nor_5  g18536(new_n14957, new_n10773, new_n20885);
nor_5  g18537(new_n14991, new_n14958, new_n20886);
nor_5  g18538(new_n20886, new_n20885, new_n20887);
xor_4  g18539(new_n20887, new_n20884, new_n20888);
xnor_4 g18540(new_n20888, new_n5779, new_n20889);
and_5  g18541(new_n14992, new_n14922, new_n20890);
nor_5  g18542(new_n15031_1, new_n14993, new_n20891);
nor_5  g18543(new_n20891, new_n20890, new_n20892);
xnor_4 g18544(new_n20892, new_n20889, n11386);
xnor_4 g18545(new_n17577, new_n17566, n11391);
xnor_4 g18546(new_n19534, new_n19533, n11398);
xor_4  g18547(new_n11592, new_n11590, n11403);
xnor_4 g18548(new_n11062, new_n11057, n11419);
xnor_4 g18549(new_n17408, new_n17394, n11439);
xnor_4 g18550(n7569, n2570, new_n20899);
nor_5  g18551(n19033, n17037, new_n20900);
xnor_4 g18552(n19033, n17037, new_n20901);
nor_5  g18553(n5386, n655, new_n20902);
xnor_4 g18554(n5386, n655, new_n20903);
nor_5  g18555(n26191, n18145, new_n20904);
xnor_4 g18556(n26191, n18145, new_n20905);
nor_5  g18557(n26512, n10712, new_n20906);
xnor_4 g18558(n26512, n10712, new_n20907);
nor_5  g18559(n25126, n19575, new_n20908);
xnor_4 g18560(n25126, n19575, new_n20909);
and_5  g18561(n19608, n15378, new_n20910);
or_5   g18562(n19608, n15378, new_n20911);
nor_5  g18563(n17095, n1689, new_n20912);
nor_5  g18564(new_n20677, new_n20672, new_n20913);
nor_5  g18565(new_n20913, new_n20912, new_n20914);
and_5  g18566(new_n20914, new_n20911, new_n20915_1);
or_5   g18567(new_n20915_1, new_n20910, new_n20916);
nor_5  g18568(new_n20916, new_n20909, new_n20917);
nor_5  g18569(new_n20917, new_n20908, new_n20918);
nor_5  g18570(new_n20918, new_n20907, new_n20919);
nor_5  g18571(new_n20919, new_n20906, new_n20920);
nor_5  g18572(new_n20920, new_n20905, new_n20921);
nor_5  g18573(new_n20921, new_n20904, new_n20922);
nor_5  g18574(new_n20922, new_n20903, new_n20923_1);
nor_5  g18575(new_n20923_1, new_n20902, new_n20924);
nor_5  g18576(new_n20924, new_n20901, new_n20925);
nor_5  g18577(new_n20925, new_n20900, new_n20926);
xor_4  g18578(new_n20926, new_n20899, new_n20927);
nor_5  g18579(new_n20927, n10514, new_n20928);
xor_4  g18580(new_n20927, n10514, new_n20929_1);
xor_4  g18581(new_n20924, new_n20901, new_n20930);
and_5  g18582(new_n20930, n18649, new_n20931);
xnor_4 g18583(new_n20930, n18649, new_n20932);
xor_4  g18584(new_n20922, new_n20903, new_n20933);
and_5  g18585(new_n20933, n6218, new_n20934);
xnor_4 g18586(new_n20933, n6218, new_n20935_1);
xor_4  g18587(new_n20920, new_n20905, new_n20936_1);
and_5  g18588(new_n20936_1, n20470, new_n20937);
xnor_4 g18589(new_n20936_1, n20470, new_n20938);
xor_4  g18590(new_n20918, new_n20907, new_n20939);
and_5  g18591(new_n20939, n21222, new_n20940);
xnor_4 g18592(new_n20939, n21222, new_n20941);
xor_4  g18593(new_n20916, new_n20909, new_n20942);
and_5  g18594(new_n20942, n9832, new_n20943);
xnor_4 g18595(new_n20942, n9832, new_n20944);
xor_4  g18596(n19608, n15378, new_n20945);
xnor_4 g18597(new_n20945, new_n20914, new_n20946_1);
nor_5  g18598(new_n20946_1, n1558, new_n20947);
xnor_4 g18599(new_n20946_1, n1558, new_n20948);
nor_5  g18600(new_n20678_1, n21749, new_n20949);
nor_5  g18601(new_n20685_1, new_n20679, new_n20950);
nor_5  g18602(new_n20950, new_n20949, new_n20951);
nor_5  g18603(new_n20951, new_n20948, new_n20952);
or_5   g18604(new_n20952, new_n20947, new_n20953);
nor_5  g18605(new_n20953, new_n20944, new_n20954);
nor_5  g18606(new_n20954, new_n20943, new_n20955);
nor_5  g18607(new_n20955, new_n20941, new_n20956);
nor_5  g18608(new_n20956, new_n20940, new_n20957);
nor_5  g18609(new_n20957, new_n20938, new_n20958);
nor_5  g18610(new_n20958, new_n20937, new_n20959);
nor_5  g18611(new_n20959, new_n20935_1, new_n20960);
nor_5  g18612(new_n20960, new_n20934, new_n20961);
nor_5  g18613(new_n20961, new_n20932, new_n20962);
nor_5  g18614(new_n20962, new_n20931, new_n20963);
and_5  g18615(new_n20963, new_n20929_1, new_n20964);
nor_5  g18616(new_n20964, new_n20928, new_n20965);
nor_5  g18617(n7569, n2570, new_n20966);
nor_5  g18618(new_n20926, new_n20899, new_n20967);
or_5   g18619(new_n20967, new_n20966, new_n20968);
xor_4  g18620(new_n20968, new_n20965, new_n20969);
or_5   g18621(new_n20780, n3795, new_n20970);
nor_5  g18622(new_n20970, n6105, new_n20971);
xnor_4 g18623(new_n20971, new_n10036, new_n20972);
xor_4  g18624(new_n20970, n6105, new_n20973);
nor_5  g18625(new_n20973, new_n7937_1, new_n20974);
xnor_4 g18626(new_n20973, new_n7937_1, new_n20975);
nor_5  g18627(new_n20781, new_n7992_1, new_n20976);
nor_5  g18628(new_n20795_1, new_n20782, new_n20977);
nor_5  g18629(new_n20977, new_n20976, new_n20978);
nor_5  g18630(new_n20978, new_n20975, new_n20979);
nor_5  g18631(new_n20979, new_n20974, new_n20980);
xnor_4 g18632(new_n20980, new_n20972, new_n20981);
xnor_4 g18633(new_n20981, new_n20969, new_n20982);
xnor_4 g18634(new_n20963, new_n20929_1, new_n20983);
xor_4  g18635(new_n20978, new_n20975, new_n20984);
and_5  g18636(new_n20984, new_n20983, new_n20985);
xnor_4 g18637(new_n20984, new_n20983, new_n20986_1);
xor_4  g18638(new_n20961, new_n20932, new_n20987);
and_5  g18639(new_n20987, new_n20796, new_n20988);
xnor_4 g18640(new_n20987, new_n20796, new_n20989);
xor_4  g18641(new_n20959, new_n20935_1, new_n20990);
and_5  g18642(new_n20990, new_n20799, new_n20991);
xnor_4 g18643(new_n20990, new_n20799, new_n20992);
xor_4  g18644(new_n20957, new_n20938, new_n20993);
and_5  g18645(new_n20993, new_n20803_1, new_n20994);
xnor_4 g18646(new_n20993, new_n20803_1, new_n20995);
xor_4  g18647(new_n20955, new_n20941, new_n20996);
and_5  g18648(new_n20996, new_n17430, new_n20997);
xnor_4 g18649(new_n20996, new_n17430, new_n20998);
xor_4  g18650(new_n16759, new_n16743_1, new_n20999);
xor_4  g18651(new_n20953, new_n20944, new_n21000);
and_5  g18652(new_n21000, new_n20999, new_n21001);
xnor_4 g18653(new_n21000, new_n20999, new_n21002);
xnor_4 g18654(new_n16757, new_n16756, new_n21003);
xor_4  g18655(new_n20951, new_n20948, new_n21004);
nor_5  g18656(new_n21004, new_n21003, new_n21005);
nor_5  g18657(new_n20686, new_n16782, new_n21006);
nor_5  g18658(new_n20693, new_n20687, new_n21007);
nor_5  g18659(new_n21007, new_n21006, new_n21008_1);
xor_4  g18660(new_n21004, new_n21003, new_n21009);
and_5  g18661(new_n21009, new_n21008_1, new_n21010);
nor_5  g18662(new_n21010, new_n21005, new_n21011);
nor_5  g18663(new_n21011, new_n21002, new_n21012);
nor_5  g18664(new_n21012, new_n21001, new_n21013);
nor_5  g18665(new_n21013, new_n20998, new_n21014);
nor_5  g18666(new_n21014, new_n20997, new_n21015);
nor_5  g18667(new_n21015, new_n20995, new_n21016);
nor_5  g18668(new_n21016, new_n20994, new_n21017_1);
nor_5  g18669(new_n21017_1, new_n20992, new_n21018);
nor_5  g18670(new_n21018, new_n20991, new_n21019);
nor_5  g18671(new_n21019, new_n20989, new_n21020);
nor_5  g18672(new_n21020, new_n20988, new_n21021);
nor_5  g18673(new_n21021, new_n20986_1, new_n21022);
nor_5  g18674(new_n21022, new_n20985, new_n21023);
xnor_4 g18675(new_n21023, new_n20982, n11462);
xnor_4 g18676(new_n18589, new_n18565, n11470);
xnor_4 g18677(new_n13990, new_n13977, n11472);
xnor_4 g18678(new_n17247, new_n6643, new_n21027);
xnor_4 g18679(new_n21027, new_n17264, n11496);
xnor_4 g18680(new_n18375, new_n18338, n11506);
xnor_4 g18681(new_n5226_1, new_n5177, new_n21030);
xnor_4 g18682(new_n20046, new_n21030, new_n21031);
xnor_4 g18683(new_n5224, new_n5181, new_n21032);
nor_5  g18684(new_n14304, new_n21032, new_n21033);
xnor_4 g18685(new_n14304, new_n21032, new_n21034_1);
xnor_4 g18686(new_n5222, new_n5186, new_n21035);
nor_5  g18687(new_n9594, new_n21035, new_n21036);
xnor_4 g18688(new_n9594, new_n21035, new_n21037);
xnor_4 g18689(new_n5220, new_n5190, new_n21038);
nor_5  g18690(new_n9610, new_n21038, new_n21039);
xnor_4 g18691(new_n9610, new_n21038, new_n21040);
not_10 g18692(new_n5269, new_n21041);
nor_5  g18693(new_n9613, new_n21041, new_n21042);
nor_5  g18694(new_n20615, new_n20602_1, new_n21043);
nor_5  g18695(new_n21043, new_n21042, new_n21044);
nor_5  g18696(new_n21044, new_n21040, new_n21045);
nor_5  g18697(new_n21045, new_n21039, new_n21046_1);
nor_5  g18698(new_n21046_1, new_n21037, new_n21047);
nor_5  g18699(new_n21047, new_n21036, new_n21048);
nor_5  g18700(new_n21048, new_n21034_1, new_n21049);
nor_5  g18701(new_n21049, new_n21033, new_n21050);
xnor_4 g18702(new_n21050, new_n21031, n11515);
xnor_4 g18703(new_n19237, new_n19207, n11538);
xnor_4 g18704(new_n17043, new_n17042, n11548);
xnor_4 g18705(new_n17297, new_n17292, n11564);
nor_5  g18706(new_n20843, n8856, new_n21055);
nor_5  g18707(new_n19945, new_n19941_1, new_n21056);
nor_5  g18708(new_n21056, new_n21055, new_n21057);
nor_5  g18709(n3324, n2272, new_n21058);
nor_5  g18710(new_n19950, new_n19947, new_n21059);
nor_5  g18711(new_n21059, new_n21058, new_n21060);
nor_5  g18712(new_n21060, new_n6813, new_n21061);
nor_5  g18713(new_n19951, new_n6809, new_n21062_1);
nor_5  g18714(new_n19955, new_n19952, new_n21063);
or_5   g18715(new_n21063, new_n21062_1, new_n21064);
xnor_4 g18716(new_n21060, new_n6813, new_n21065);
nor_5  g18717(new_n21065, new_n21064, new_n21066);
nor_5  g18718(new_n21066, new_n21061, new_n21067);
xor_4  g18719(new_n21067, new_n21057, new_n21068);
nor_5  g18720(new_n21063, new_n21062_1, new_n21069);
xor_4  g18721(new_n21065, new_n21069, new_n21070);
nor_5  g18722(new_n21070, new_n21057, new_n21071);
xnor_4 g18723(new_n21065, new_n21069, new_n21072);
xnor_4 g18724(new_n21072, new_n21057, new_n21073);
nor_5  g18725(new_n19956, new_n19946, new_n21074);
nor_5  g18726(new_n19960, new_n19957, new_n21075);
nor_5  g18727(new_n21075, new_n21074, new_n21076);
and_5  g18728(new_n21076, new_n21073, new_n21077);
nor_5  g18729(new_n21077, new_n21071, new_n21078_1);
xnor_4 g18730(new_n21078_1, new_n21068, n11591);
nor_5  g18731(new_n7567, new_n7561, new_n21080);
and_5  g18732(new_n7579, new_n7568, new_n21081);
nor_5  g18733(new_n7579, new_n7568, new_n21082);
or_5   g18734(new_n7634, new_n21082, new_n21083);
nand_5 g18735(new_n21083, new_n20618, new_n21084);
or_5   g18736(new_n21084, new_n21081, new_n21085);
nor_5  g18737(new_n21085, new_n21080, n11607);
xnor_4 g18738(new_n16988_1, new_n16964, n11647);
xor_4  g18739(new_n20871, new_n20868, n11674);
xnor_4 g18740(new_n17881, new_n19524, new_n21089);
nor_5  g18741(new_n17891, new_n19524, new_n21090);
nor_5  g18742(new_n19536, new_n19525, new_n21091);
nor_5  g18743(new_n21091, new_n21090, new_n21092);
xor_4  g18744(new_n21092, new_n21089, n11682);
xor_4  g18745(new_n20148, new_n20136, n11710);
xnor_4 g18746(new_n12505, new_n12479, n11712);
xnor_4 g18747(new_n19832, new_n19819, n11724);
xnor_4 g18748(new_n16454, new_n16453, n11741);
xor_4  g18749(new_n16221, new_n2945, n11770);
xnor_4 g18750(new_n7621, new_n7620, n11771);
xnor_4 g18751(new_n17145, new_n17117, n11818);
xnor_4 g18752(new_n20611, new_n20606, n11837);
and_5  g18753(new_n14642, new_n3353, new_n21102);
xnor_4 g18754(new_n21102, n2743, new_n21103);
and_5  g18755(new_n21103, new_n5430_1, new_n21104);
xnor_4 g18756(new_n21103, new_n5430_1, new_n21105);
nor_5  g18757(new_n14643, new_n5434, new_n21106);
nor_5  g18758(new_n14679, new_n14644, new_n21107);
nor_5  g18759(new_n21107, new_n21106, new_n21108);
nor_5  g18760(new_n21108, new_n21105, new_n21109);
nor_5  g18761(new_n21109, new_n21104, new_n21110);
nand_5 g18762(new_n21102, new_n12179_1, new_n21111);
xnor_4 g18763(new_n21111, new_n12117, new_n21112);
xnor_4 g18764(new_n21112, new_n21110, new_n21113);
xnor_4 g18765(new_n21113, new_n19890, new_n21114);
xor_4  g18766(new_n21108, new_n21105, new_n21115);
nor_5  g18767(new_n21115, new_n19471, new_n21116);
xnor_4 g18768(new_n21115, new_n19471, new_n21117);
and_5  g18769(new_n14689, new_n14680_1, new_n21118);
nor_5  g18770(new_n14731, new_n14690, new_n21119);
nor_5  g18771(new_n21119, new_n21118, new_n21120);
nor_5  g18772(new_n21120, new_n21117, new_n21121);
nor_5  g18773(new_n21121, new_n21116, new_n21122);
xnor_4 g18774(new_n21122, new_n21114, n11842);
xnor_4 g18775(new_n14269, new_n14251, n11843);
xnor_4 g18776(new_n16794, new_n16780, n11905);
xnor_4 g18777(new_n10258, new_n10253, n11965);
xnor_4 g18778(new_n16686, new_n16682_1, n12000);
xor_4  g18779(new_n14802, new_n14799, n12003);
xnor_4 g18780(new_n15371, new_n15370, n12011);
xnor_4 g18781(new_n15833, new_n15820, n12072);
xor_4  g18782(new_n9657, new_n9656, n12131);
xor_4  g18783(new_n14781, new_n14750, n12146);
xnor_4 g18784(new_n15019_1, new_n15016, n12157);
xnor_4 g18785(new_n9264, new_n9216, n12158);
xnor_4 g18786(new_n20232, new_n20211, n12179);
xnor_4 g18787(new_n5832, new_n5789, n12192);
xnor_4 g18788(new_n20550, new_n20540, n12223);
xnor_4 g18789(new_n9262, new_n9220_1, n12225);
xnor_4 g18790(new_n20613, new_n20604_1, n12228);
xnor_4 g18791(new_n12058, new_n6523, n12235);
xnor_4 g18792(new_n8242, new_n8218, n12302);
xnor_4 g18793(new_n15163, new_n15133, n12304);
xor_4  g18794(n19196, n1742, new_n21143);
nor_5  g18795(new_n14933, n4858, new_n21144);
xor_4  g18796(n23586, n4858, new_n21145);
nor_5  g18797(new_n14936, n8244, new_n21146);
xor_4  g18798(n21226, n8244, new_n21147);
nor_5  g18799(n9493, new_n14939, new_n21148);
nor_5  g18800(n20036, new_n11106, new_n21149);
nor_5  g18801(new_n17819, new_n17814, new_n21150);
or_5   g18802(new_n21150, new_n21149, new_n21151);
xor_4  g18803(n9493, n4426, new_n21152);
nor_5  g18804(new_n21152, new_n21151, new_n21153);
nor_5  g18805(new_n21153, new_n21148, new_n21154_1);
nor_5  g18806(new_n21154_1, new_n21147, new_n21155);
nor_5  g18807(new_n21155, new_n21146, new_n21156);
nor_5  g18808(new_n21156, new_n21145, new_n21157_1);
nor_5  g18809(new_n21157_1, new_n21144, new_n21158);
xor_4  g18810(new_n21158, new_n21143, new_n21159);
xnor_4 g18811(new_n21159, new_n17772, new_n21160);
xor_4  g18812(new_n21156, new_n21145, new_n21161);
nor_5  g18813(new_n21161, new_n16440_1, new_n21162);
xnor_4 g18814(new_n21161, new_n16440_1, new_n21163);
xor_4  g18815(new_n21154_1, new_n21147, new_n21164);
nor_5  g18816(new_n21164, new_n16442, new_n21165);
xnor_4 g18817(new_n21164, new_n16442, new_n21166);
not_10 g18818(new_n16445_1, new_n21167);
xor_4  g18819(new_n21152, new_n21151, new_n21168_1);
nor_5  g18820(new_n21168_1, new_n21167, new_n21169);
xor_4  g18821(new_n21168_1, new_n16445_1, new_n21170);
not_10 g18822(new_n16448, new_n21171);
and_5  g18823(new_n17820_1, new_n21171, new_n21172);
nor_5  g18824(new_n17830, new_n17821, new_n21173_1);
nor_5  g18825(new_n21173_1, new_n21172, new_n21174);
nor_5  g18826(new_n21174, new_n21170, new_n21175);
nor_5  g18827(new_n21175, new_n21169, new_n21176_1);
nor_5  g18828(new_n21176_1, new_n21166, new_n21177);
nor_5  g18829(new_n21177, new_n21165, new_n21178);
nor_5  g18830(new_n21178, new_n21163, new_n21179);
nor_5  g18831(new_n21179, new_n21162, new_n21180);
xnor_4 g18832(new_n21180, new_n21160, n12324);
xnor_4 g18833(new_n19531_1, new_n19528, n12325);
xor_4  g18834(new_n9475, new_n9458_1, n12329);
xnor_4 g18835(new_n7853, new_n7852, n12330);
xnor_4 g18836(new_n5300_1, new_n5259, n12346);
xnor_4 g18837(new_n6908, new_n6888, n12349);
xnor_4 g18838(new_n17573, new_n17572, n12364);
not_10 g18839(new_n20123, new_n21188);
and_5  g18840(new_n21188, new_n5242, new_n21189);
xnor_4 g18841(new_n21188, new_n5242, new_n21190);
nor_5  g18842(new_n20123, new_n5245, new_n21191);
xnor_4 g18843(new_n20123, new_n5245, new_n21192);
xnor_4 g18844(new_n5228_1, new_n5173, new_n21193_1);
nor_5  g18845(new_n20044, new_n21193_1, new_n21194);
xnor_4 g18846(new_n20044, new_n21193_1, new_n21195);
nor_5  g18847(new_n20046, new_n21030, new_n21196);
nor_5  g18848(new_n21050, new_n21031, new_n21197);
nor_5  g18849(new_n21197, new_n21196, new_n21198);
nor_5  g18850(new_n21198, new_n21195, new_n21199);
nor_5  g18851(new_n21199, new_n21194, new_n21200);
nor_5  g18852(new_n21200, new_n21192, new_n21201);
or_5   g18853(new_n21201, new_n21191, new_n21202);
nor_5  g18854(new_n21202, new_n21190, new_n21203_1);
nor_5  g18855(new_n21203_1, new_n21189, n12383);
xor_4  g18856(new_n7783, new_n7781, n12397);
xor_4  g18857(new_n15506_1, new_n15496_1, n12408);
and_5  g18858(new_n17881, new_n19524, new_n21207);
nor_5  g18859(new_n21092, new_n21089, new_n21208);
nor_5  g18860(new_n21208, new_n21207, n12449);
xnor_4 g18861(new_n19316, new_n19283, n12461);
or_5   g18862(new_n19160, new_n10815, new_n21211);
and_5  g18863(new_n21211, new_n15587, new_n21212);
nor_5  g18864(new_n21211, new_n15587, new_n21213);
nor_5  g18865(new_n19161, new_n19153, new_n21214);
nor_5  g18866(new_n19171, new_n19162, new_n21215);
nor_5  g18867(new_n21215, new_n21214, new_n21216);
nor_5  g18868(new_n21216, new_n21213, new_n21217);
or_5   g18869(new_n21217, new_n21212, n12462);
xor_4  g18870(new_n20244, new_n20238, n12467);
nor_5  g18871(new_n14384, n3324, new_n21220);
nor_5  g18872(new_n14409, new_n14385, new_n21221);
or_5   g18873(new_n21221, new_n21220, new_n21222_1);
nor_5  g18874(new_n21222_1, new_n19911_1, new_n21223);
nor_5  g18875(new_n14489, new_n14482, new_n21224);
nor_5  g18876(new_n14488, n13419, new_n21225_1);
or_5   g18877(new_n21225_1, new_n21224, new_n21226_1);
nor_5  g18878(new_n21226_1, new_n20643, new_n21227);
xor_4  g18879(new_n21222_1, new_n19911_1, new_n21228);
xnor_4 g18880(new_n21226_1, new_n20642, new_n21229);
nor_5  g18881(new_n21229, new_n21228, new_n21230);
xor_4  g18882(new_n21229, new_n21228, new_n21231);
nor_5  g18883(new_n14490, new_n14410, new_n21232);
nor_5  g18884(new_n14530, new_n14491, new_n21233);
nor_5  g18885(new_n21233, new_n21232, new_n21234);
and_5  g18886(new_n21234, new_n21231, new_n21235);
nor_5  g18887(new_n21235, new_n21230, new_n21236);
xor_4  g18888(new_n21236, new_n21227, new_n21237);
xnor_4 g18889(new_n21237, new_n21223, n12469);
xnor_4 g18890(new_n9893, new_n9870, n12515);
nor_5  g18891(new_n20880, n5140, new_n21240);
xor_4  g18892(n10250, n5140, new_n21241);
nor_5  g18893(new_n14924, n6204, new_n21242);
xor_4  g18894(n7674, n6204, new_n21243);
nor_5  g18895(new_n14927, n3349, new_n21244);
xor_4  g18896(n6397, n3349, new_n21245);
nor_5  g18897(new_n14930, n1742, new_n21246);
nor_5  g18898(new_n21158, new_n21143, new_n21247);
nor_5  g18899(new_n21247, new_n21246, new_n21248);
nor_5  g18900(new_n21248, new_n21245, new_n21249);
nor_5  g18901(new_n21249, new_n21244, new_n21250);
nor_5  g18902(new_n21250, new_n21243, new_n21251);
nor_5  g18903(new_n21251, new_n21242, new_n21252);
nor_5  g18904(new_n21252, new_n21241, new_n21253);
nor_5  g18905(new_n21253, new_n21240, new_n21254_1);
not_10 g18906(new_n21254_1, new_n21255);
xnor_4 g18907(new_n21255, new_n19986, new_n21256);
and_5  g18908(new_n21254_1, new_n18915, new_n21257);
nor_5  g18909(new_n21254_1, new_n18915, new_n21258);
xor_4  g18910(new_n21252, new_n21241, new_n21259);
nor_5  g18911(new_n21259, new_n18917, new_n21260);
xnor_4 g18912(new_n21259, new_n18917, new_n21261);
xor_4  g18913(new_n21250, new_n21243, new_n21262);
nor_5  g18914(new_n21262, new_n17767, new_n21263);
xnor_4 g18915(new_n21262, new_n17767, new_n21264);
xor_4  g18916(new_n21248, new_n21245, new_n21265);
nor_5  g18917(new_n21265, new_n17769, new_n21266);
xnor_4 g18918(new_n21265, new_n17769, new_n21267);
nor_5  g18919(new_n21159, new_n17772, new_n21268);
nor_5  g18920(new_n21180, new_n21160, new_n21269);
nor_5  g18921(new_n21269, new_n21268, new_n21270);
nor_5  g18922(new_n21270, new_n21267, new_n21271);
nor_5  g18923(new_n21271, new_n21266, new_n21272);
nor_5  g18924(new_n21272, new_n21264, new_n21273);
nor_5  g18925(new_n21273, new_n21263, new_n21274);
nor_5  g18926(new_n21274, new_n21261, new_n21275);
or_5   g18927(new_n21275, new_n21260, new_n21276_1);
nor_5  g18928(new_n21276_1, new_n21258, new_n21277);
nor_5  g18929(new_n21277, new_n21257, new_n21278);
xnor_4 g18930(new_n21278, new_n21256, n12516);
xnor_4 g18931(new_n6725, new_n6715, n12540);
xnor_4 g18932(new_n10555, new_n10554, n12545);
xnor_4 g18933(new_n18587, new_n18568, n12552);
xnor_4 g18934(new_n7445, new_n7424, n12566);
xnor_4 g18935(new_n12021, new_n12005, n12569);
xnor_4 g18936(new_n5836, new_n5781, n12607);
xnor_4 g18937(new_n9094, new_n9036, n12620);
xnor_4 g18938(new_n3510, new_n3475, n12621);
xnor_4 g18939(new_n16618, new_n16617_1, n12654);
xor_4  g18940(new_n17822, new_n13601, n12665);
xnor_4 g18941(new_n15540, new_n15531, n12670);
xor_4  g18942(new_n6897, new_n2505, n12707);
xnor_4 g18943(new_n6487, new_n6477, n12725);
xnor_4 g18944(new_n14528, new_n14495, n12727);
xor_4  g18945(new_n8824_1, new_n8801, n12740);
xor_4  g18946(new_n18888, new_n18887_1, n12742);
xor_4  g18947(new_n19063, new_n2746, n12746);
xor_4  g18948(new_n8394, new_n8393, n12756);
xnor_4 g18949(new_n6500, new_n6452, n12783);
xnor_4 g18950(new_n21255, new_n18915, new_n21299);
xnor_4 g18951(new_n21299, new_n21276_1, n12801);
xnor_4 g18952(new_n16127, new_n16124, n12812);
xnor_4 g18953(new_n14729, new_n14694, n12816);
nor_5  g18954(new_n15721, n6659, new_n21303);
nor_5  g18955(new_n16668, new_n16648, new_n21304);
or_5   g18956(new_n21304, new_n21303, new_n21305);
nor_5  g18957(new_n21305, new_n18045_1, new_n21306);
xor_4  g18958(new_n21305, new_n18045_1, new_n21307);
nor_5  g18959(new_n21307, new_n21228, new_n21308);
xnor_4 g18960(new_n21307, new_n21228, new_n21309);
and_5  g18961(new_n16669, new_n14410, new_n21310);
nor_5  g18962(new_n16694, new_n16670, new_n21311);
nor_5  g18963(new_n21311, new_n21310, new_n21312);
nor_5  g18964(new_n21312, new_n21309, new_n21313);
nor_5  g18965(new_n21313, new_n21308, new_n21314);
nor_5  g18966(new_n21314, new_n21306, new_n21315);
nor_5  g18967(new_n21315, new_n21223, n12843);
xnor_4 g18968(new_n19107_1, new_n19106, n12864);
not_10 g18969(new_n4476_1, new_n21318);
nor_5  g18970(new_n20353, new_n21318, new_n21319);
and_5  g18971(new_n20378, new_n20354, new_n21320);
nor_5  g18972(new_n21320, new_n21319, new_n21321);
nor_5  g18973(n21784, n3740, new_n21322);
nor_5  g18974(new_n20352, new_n20333_1, new_n21323);
nor_5  g18975(new_n21323, new_n21322, new_n21324);
xnor_4 g18976(new_n21324, new_n4533, new_n21325);
xnor_4 g18977(new_n21325, new_n21321, new_n21326);
nor_5  g18978(new_n21326, new_n17033, new_n21327);
and_5  g18979(new_n20379, new_n15893, new_n21328);
nor_5  g18980(new_n20403_1, new_n20380, new_n21329);
nor_5  g18981(new_n21329, new_n21328, new_n21330);
xnor_4 g18982(new_n21326, new_n17033, new_n21331);
nor_5  g18983(new_n21331, new_n21330, new_n21332);
nor_5  g18984(new_n21332, new_n21327, new_n21333);
and_5  g18985(new_n21324, new_n4533, new_n21334);
nor_5  g18986(new_n21324, new_n4533, new_n21335);
nor_5  g18987(new_n21335, new_n21321, new_n21336);
nor_5  g18988(new_n21336, new_n21334, new_n21337);
and_5  g18989(new_n21337, new_n21333, n12865);
xnor_4 g18990(new_n11666, new_n11648, n12870);
xnor_4 g18991(new_n19071, new_n19053, n12873);
and_5  g18992(new_n20507, new_n16860, new_n21341);
xnor_4 g18993(new_n20507, new_n16860, new_n21342);
nor_5  g18994(new_n19886, new_n16943, new_n21343);
nor_5  g18995(new_n20830, new_n20827, new_n21344);
nor_5  g18996(new_n21344, new_n21343, new_n21345);
nor_5  g18997(new_n21345, new_n21342, new_n21346);
or_5   g18998(new_n21346, new_n21341, n12904);
xor_4  g18999(new_n9480, new_n9479, n12941);
xnor_4 g19000(new_n10141, new_n10133, n12942);
xnor_4 g19001(new_n5373, new_n3568, new_n21350);
xnor_4 g19002(new_n21350, new_n5378, n12978);
xor_4  g19003(new_n8837, new_n7178, n12980);
xor_4  g19004(new_n5967, new_n4361, n12985);
xnor_4 g19005(new_n13169, new_n13134, n12987);
not_10 g19006(n2160, new_n21355);
nor_5  g19007(n11220, new_n21355, new_n21356);
nor_5  g19008(new_n15239, new_n15220, new_n21357);
nor_5  g19009(new_n21357, new_n21356, new_n21358);
xor_4  g19010(new_n21358, new_n13412, new_n21359);
and_5  g19011(new_n15240, new_n13450, new_n21360);
nor_5  g19012(new_n15259, new_n15241_1, new_n21361);
nor_5  g19013(new_n21361, new_n21360, new_n21362);
xnor_4 g19014(new_n21362, new_n21359, n12992);
nor_5  g19015(new_n20174, n6659, new_n21364);
nor_5  g19016(new_n19245, n23250, new_n21365_1);
nor_5  g19017(new_n19278, new_n19246, new_n21366);
nor_5  g19018(new_n21366, new_n21365_1, new_n21367_1);
and_5  g19019(new_n20174, n6659, new_n21368);
nor_5  g19020(new_n21368, new_n21367_1, new_n21369);
nor_5  g19021(new_n21369, new_n21364, new_n21370);
nor_5  g19022(new_n21370, new_n20172, new_n21371);
not_10 g19023(new_n21371, new_n21372);
xnor_4 g19024(new_n21372, new_n18056, new_n21373);
not_10 g19025(new_n18068, new_n21374);
xnor_4 g19026(new_n20174, new_n20639, new_n21375);
xnor_4 g19027(new_n21375, new_n21367_1, new_n21376);
nor_5  g19028(new_n21376, new_n21374, new_n21377);
nor_5  g19029(new_n19279, new_n12965, new_n21378);
nor_5  g19030(new_n19318, new_n19280, new_n21379);
nor_5  g19031(new_n21379, new_n21378, new_n21380);
xor_4  g19032(new_n21376, new_n18068, new_n21381);
nor_5  g19033(new_n21381, new_n21380, new_n21382);
nor_5  g19034(new_n21382, new_n21377, new_n21383);
xnor_4 g19035(new_n21383, new_n21373, n13005);
xor_4  g19036(new_n18154, new_n15107, n13043);
xnor_4 g19037(new_n16200, new_n16199, n13048);
xnor_4 g19038(new_n13945, new_n13944, n13054);
xnor_4 g19039(new_n16355, new_n16345, n13082);
xnor_4 g19040(new_n6492, new_n6468, n13096);
xnor_4 g19041(new_n16357, new_n16339, n13116);
xnor_4 g19042(new_n18169, new_n18136, n13122);
xnor_4 g19043(new_n5818, new_n5817, n13141);
xor_4  g19044(new_n18011, new_n18004, n13144);
xnor_4 g19045(new_n18593, new_n18559, n13168);
xnor_4 g19046(new_n19231, new_n19214, n13198);
xnor_4 g19047(new_n13163, new_n13145, n13199);
xnor_4 g19048(new_n13273_1, new_n13261, n13204);
xnor_4 g19049(new_n9255, new_n9231, n13209);
xnor_4 g19050(new_n17810, new_n17801, n13270);
xnor_4 g19051(new_n11917, new_n11897, n13273);
xnor_4 g19052(new_n20234, new_n20206, n13285);
xnor_4 g19053(new_n19630, new_n19612, n13338);
xnor_4 g19054(new_n7190_1, new_n7167, n13407);
xor_4  g19055(new_n5001, new_n3965, new_n21404_1);
xnor_4 g19056(new_n21404_1, new_n14764, n13409);
xnor_4 g19057(new_n5016, new_n4988, n13456);
nor_5  g19058(new_n19574, new_n18930, new_n21407);
nor_5  g19059(new_n19606, new_n18932, new_n21408);
nor_5  g19060(new_n20585, new_n20582_1, new_n21409);
nor_5  g19061(new_n21409, new_n21408, new_n21410);
or_5   g19062(new_n19602_1, new_n18930, new_n21411);
and_5  g19063(new_n21411, new_n21410, new_n21412);
and_5  g19064(new_n21412, new_n21407, new_n21413);
xnor_4 g19065(new_n19602_1, new_n18930, new_n21414);
xor_4  g19066(new_n21414, new_n21410, new_n21415);
nor_5  g19067(new_n21415, new_n10293, new_n21416);
xor_4  g19068(new_n21415, new_n10293, new_n21417);
and_5  g19069(new_n20586, new_n10374, new_n21418);
nor_5  g19070(new_n20590_1, new_n20587, new_n21419);
nor_5  g19071(new_n21419, new_n21418, new_n21420);
and_5  g19072(new_n21420, new_n21417, new_n21421);
nor_5  g19073(new_n21421, new_n21416, new_n21422);
xor_4  g19074(new_n19574, new_n18930, new_n21423);
and_5  g19075(new_n21423, new_n21410, new_n21424);
nor_5  g19076(new_n21423, new_n21412, new_n21425);
nor_5  g19077(new_n21425, new_n21424, new_n21426);
nor_5  g19078(new_n21426, new_n21422, new_n21427);
or_5   g19079(new_n21427, new_n21413, n13457);
xnor_4 g19080(new_n11011_1, new_n11003, n13477);
xnor_4 g19081(new_n11333, new_n11332, n13484);
xnor_4 g19082(new_n18776, new_n18749, n13486);
xnor_4 g19083(new_n20134, new_n19660, new_n21432);
nor_5  g19084(new_n20056, new_n15798, new_n21433);
nor_5  g19085(new_n20082, new_n20057, new_n21434);
nor_5  g19086(new_n21434, new_n21433, new_n21435);
xor_4  g19087(new_n21435, new_n21432, n13487);
xnor_4 g19088(new_n4813, new_n4796, n13500);
xor_4  g19089(new_n4248, new_n4247, n13501);
xnor_4 g19090(new_n5824, new_n5805, n13506);
xnor_4 g19091(new_n5608, new_n5600, n13548);
xnor_4 g19092(new_n21015, new_n20995, n13551);
xnor_4 g19093(new_n4636, new_n4618, n13602);
xnor_4 g19094(new_n15878, new_n15868, n13626);
xnor_4 g19095(new_n7441, new_n7433, n13683);
xnor_4 g19096(new_n18377_1, new_n18335, n13710);
xnor_4 g19097(new_n18015, new_n17998_1, n13722);
xnor_4 g19098(new_n12826, new_n12775, new_n21447);
xnor_4 g19099(new_n21447, new_n12894, n13754);
xor_4  g19100(new_n2757, new_n2729, n13764);
xnor_4 g19101(new_n13026_1, new_n13023, new_n21450);
xnor_4 g19102(new_n21450, new_n13030, n13798);
xnor_4 g19103(new_n15882, new_n15864, n13835);
xnor_4 g19104(new_n14358, new_n14357, n13850);
xor_4  g19105(new_n16346, new_n7059, n13922);
xnor_4 g19106(new_n17779, new_n17771, n13923);
xnor_4 g19107(new_n10560, new_n10559, n14004);
xnor_4 g19108(new_n10763_1, new_n10725, n14036);
xnor_4 g19109(new_n19709, new_n19694, n14059);
xor_4  g19110(new_n15710, new_n15706, n14081);
xnor_4 g19111(new_n17260, new_n17257, n14095);
xor_4  g19112(new_n6112, new_n3215, n14107);
xnor_4 g19113(new_n8094, new_n8065, n14121);
xor_4  g19114(new_n10970, new_n10969, n14126);
xnor_4 g19115(new_n18019, new_n17992, n14136);
and_5  g19116(new_n21358, new_n13412, new_n21465);
nor_5  g19117(new_n21358, new_n13412, new_n21466);
nor_5  g19118(new_n21362, new_n21466, new_n21467);
nor_5  g19119(new_n21467, new_n21465, new_n21468);
xnor_4 g19120(new_n21358, new_n20419, new_n21469);
xnor_4 g19121(new_n21469, new_n21468, n14147);
xnor_4 g19122(new_n19441, new_n19397, n14174);
xnor_4 g19123(new_n15027, new_n15001, n14190);
xnor_4 g19124(new_n5014, new_n4992, n14211);
xnor_4 g19125(new_n15211, new_n15208, n14222);
xnor_4 g19126(new_n12231, new_n12187, n14267);
xnor_4 g19127(new_n5290, new_n5280, n14271);
xnor_4 g19128(new_n8545, new_n8535_1, n14277);
xnor_4 g19129(new_n7616_1, new_n7615, n14294);
xnor_4 g19130(new_n21021, new_n20986_1, n14310);
xnor_4 g19131(new_n21044, new_n21040, n14326);
xnor_4 g19132(new_n11286, new_n11244, n14342);
xnor_4 g19133(new_n16792, new_n16784, n14353);
and_5  g19134(new_n19690, new_n10582, new_n21483);
nor_5  g19135(new_n19690, new_n8146, new_n21484);
nor_5  g19136(new_n19711, new_n19691, new_n21485);
nor_5  g19137(new_n21485, new_n21484, new_n21486);
nor_5  g19138(new_n21486, new_n21483, new_n21487);
nor_5  g19139(new_n19690, new_n10582, new_n21488);
nor_5  g19140(new_n21488, new_n21485, new_n21489_1);
nor_5  g19141(new_n21489_1, new_n21487, n14364);
xor_4  g19142(new_n20143, new_n20140, n14375);
xnor_4 g19143(new_n20558, new_n20532, n14412);
nor_5  g19144(new_n10514_1, new_n4136, new_n21493);
or_5   g19145(new_n16086, new_n5689, new_n21494);
nor_5  g19146(new_n16110_1, new_n21494, new_n21495);
xnor_4 g19147(new_n21495, new_n21493, new_n21496);
nor_5  g19148(new_n16111, new_n10516, new_n21497);
nor_5  g19149(new_n16135, new_n16112, new_n21498);
nor_5  g19150(new_n21498, new_n21497, new_n21499);
xnor_4 g19151(new_n21499, new_n21496, n14414);
xor_4  g19152(new_n14132, new_n14131, n14457);
xnor_4 g19153(new_n4640, new_n4609, n14464);
xnor_4 g19154(new_n9891, new_n9873, n14471);
and_5  g19155(new_n18045_1, new_n7578, new_n21504);
nor_5  g19156(new_n18055, new_n18046, new_n21505);
nor_5  g19157(new_n21505, new_n21504, new_n21506);
xnor_4 g19158(new_n21506, new_n21372, new_n21507);
and_5  g19159(new_n21371, new_n18056, new_n21508);
nor_5  g19160(new_n21371, new_n18056, new_n21509);
nor_5  g19161(new_n21383, new_n21509, new_n21510);
nor_5  g19162(new_n21510, new_n21508, new_n21511);
xnor_4 g19163(new_n21511, new_n21507, n14475);
xnor_4 g19164(new_n11274, new_n11273_1, n14541);
not_10 g19165(new_n19922_1, new_n21514);
nor_5  g19166(new_n19926, new_n21514, new_n21515);
nor_5  g19167(new_n19936, new_n19927, new_n21516);
or_5   g19168(new_n21516, new_n21515, n14546);
xor_4  g19169(new_n10068, new_n10067, n14547);
xnor_4 g19170(new_n11598, new_n11582, n14593);
xnor_4 g19171(new_n8549, new_n8527, n14636);
xnor_4 g19172(new_n21178, new_n21163, n14701);
xnor_4 g19173(new_n11064, new_n11055, n14734);
xnor_4 g19174(new_n6498, new_n6456_1, n14746);
xnor_4 g19175(new_n8816, new_n8814, n14763);
xnor_4 g19176(new_n20754, new_n20746, n14772);
xnor_4 g19177(new_n20146, new_n20145, n14801);
xnor_4 g19178(new_n19754, new_n19735, n14819);
xnor_4 g19179(new_n13281, new_n13247, n14827);
xnor_4 g19180(new_n19169, new_n19166, n14839);
xnor_4 g19181(new_n15874, new_n15873, n14849);
nor_5  g19182(new_n19029, new_n13232, new_n21531);
nor_5  g19183(new_n19086, new_n19030, new_n21532);
nor_5  g19184(new_n21532, new_n21531, new_n21533);
nor_5  g19185(new_n21533, new_n19026, n14891);
xor_4  g19186(new_n5932, new_n4387, n14931);
nand_5 g19187(new_n21495, new_n10515, new_n21536);
nor_5  g19188(new_n21499, new_n21536, new_n21537);
nor_5  g19189(new_n21495, new_n10515, new_n21538_1);
and_5  g19190(new_n21499, new_n21538_1, new_n21539);
or_5   g19191(new_n21539, new_n21537, n14944);
xor_4  g19192(new_n16788, new_n8104, n14977);
xnor_4 g19193(new_n11606, new_n11566_1, n14989);
xnor_4 g19194(new_n9797, new_n9790, n15002);
xnor_4 g19195(new_n20609_1, new_n5287, n15004);
xnor_4 g19196(new_n8246, new_n8210, n15011);
xor_4  g19197(new_n20665, new_n20662, n15019);
and_5  g19198(new_n13931, new_n13924, new_n21547);
nor_5  g19199(new_n13951_1, new_n13932, new_n21548);
or_5   g19200(new_n21548, new_n21547, n15031);
xor_4  g19201(new_n16347, new_n16346, n15033);
xor_4  g19202(new_n10854, new_n6523, n15052);
xnor_4 g19203(new_n17933, new_n17924, n15082);
xnor_4 g19204(new_n7443, new_n7428_1, n15094);
xor_4  g19205(new_n10613, new_n10610, n15118);
xnor_4 g19206(new_n21345, new_n21342, n15128);
xnor_4 g19207(new_n17149, new_n17111, n15139);
xnor_4 g19208(new_n15302, new_n15304, new_n21557);
xnor_4 g19209(new_n21557, new_n15311, n15145);
xnor_4 g19210(new_n13483, new_n13455, n15165);
xor_4  g19211(new_n13870, new_n4695, n15176);
xor_4  g19212(new_n18581, new_n18580, n15180);
xnor_4 g19213(new_n14783, new_n14748, n15205);
xor_4  g19214(new_n5007, new_n3967, n15230);
xor_4  g19215(new_n15536, new_n15535, n15255);
xnor_4 g19216(new_n8828, new_n8793, n15275);
xnor_4 g19217(new_n12676, new_n12673, n15300);
and_5  g19218(new_n21111, new_n12117, new_n21567);
and_5  g19219(new_n21567, new_n21110, new_n21568);
or_5   g19220(new_n21111, new_n12117, new_n21569);
nor_5  g19221(new_n21569, new_n21110, new_n21570);
nor_5  g19222(new_n21570, new_n21568, new_n21571);
xor_4  g19223(new_n21571, new_n19922_1, new_n21572);
nor_5  g19224(new_n21113, new_n19890, new_n21573);
nor_5  g19225(new_n21122, new_n21114, new_n21574);
or_5   g19226(new_n21574, new_n21573, new_n21575);
xnor_4 g19227(new_n21575, new_n21572, n15307);
xnor_4 g19228(new_n18379, new_n18332_1, n15327);
xnor_4 g19229(new_n18365, new_n18357, n15345);
xnor_4 g19230(new_n11596, new_n11586, n15353);
xor_4  g19231(new_n21202, new_n21190, n15366);
xnor_4 g19232(new_n21337, new_n21333, n15382);
xnor_4 g19233(new_n8400, new_n8382, n15407);
xor_4  g19234(new_n13599, new_n12297, n15428);
and_5  g19235(new_n20968, new_n20965, new_n21584);
and_5  g19236(new_n20981, new_n20969, new_n21585);
nor_5  g19237(new_n21023, new_n20982, new_n21586);
nor_5  g19238(new_n21586, new_n21585, new_n21587);
nor_5  g19239(new_n21587, new_n21584, new_n21588);
or_5   g19240(new_n20971, new_n10036, new_n21589);
or_5   g19241(new_n20980, new_n21589, new_n21590);
nor_5  g19242(new_n21590, new_n21584, new_n21591);
nor_5  g19243(new_n21591, new_n21586, new_n21592);
nor_5  g19244(new_n21592, new_n21588, n15435);
or_5   g19245(new_n20623_1, new_n20618, new_n21594);
nor_5  g19246(new_n20633, new_n21594, new_n21595);
and_5  g19247(new_n20623_1, new_n20618, new_n21596);
and_5  g19248(new_n20633, new_n21596, new_n21597);
or_5   g19249(new_n21597, new_n21595, n15438);
xnor_4 g19250(new_n21017_1, new_n20992, n15465);
xor_4  g19251(new_n7781, new_n6045, n15467);
xnor_4 g19252(new_n7200, new_n7143, n15470);
xnor_4 g19253(new_n13285_1, new_n13240, n15477);
xnor_4 g19254(new_n21272, new_n21264, n15481);
xnor_4 g19255(new_n13688, new_n13685, n15496);
xnor_4 g19256(new_n10980, new_n10951, n15501);
xnor_4 g19257(new_n17262, new_n17253, n15555);
xnor_4 g19258(new_n19569, new_n19553, n15558);
and_5  g19259(new_n21514, new_n20507, new_n21608);
nor_5  g19260(new_n20511, new_n20508, new_n21609);
or_5   g19261(new_n21609, new_n21608, n15559);
and_5  g19262(new_n5024_1, n5101, new_n21611);
nor_5  g19263(new_n18615, new_n18600, new_n21612);
nor_5  g19264(new_n21612, new_n21611, new_n21613);
and_5  g19265(new_n21613, new_n20700_1, new_n21614);
and_5  g19266(new_n18665, new_n18616, new_n21615_1);
nor_5  g19267(new_n18689, new_n18666, new_n21616);
nor_5  g19268(new_n21616, new_n21615_1, new_n21617);
nor_5  g19269(new_n21613, new_n19916_1, new_n21618);
or_5   g19270(new_n21618, new_n21617, new_n21619);
nor_5  g19271(new_n21619, new_n20700_1, new_n21620);
nor_5  g19272(new_n21618, new_n21617, new_n21621);
not_10 g19273(new_n21613, new_n21622);
nor_5  g19274(new_n21622, new_n19916_1, new_n21623);
nor_5  g19275(new_n21623, new_n21621, new_n21624);
or_5   g19276(new_n21624, new_n21620, new_n21625);
nor_5  g19277(new_n21625, new_n21614, n15570);
xnor_4 g19278(new_n11292, new_n11232, n15573);
xnor_4 g19279(new_n10571, new_n10570, n15588);
xnor_4 g19280(new_n19750, new_n19742, n15590);
xnor_4 g19281(new_n20302, new_n20292, n15598);
xnor_4 g19282(new_n8551, new_n8523, n15614);
xnor_4 g19283(new_n20758, new_n20739, n15662);
xnor_4 g19284(new_n3231, new_n3202, n15716);
xnor_4 g19285(new_n13171, new_n13131, n15749);
xnor_4 g19286(new_n17172, new_n17168_1, n15762);
xor_4  g19287(new_n7179, new_n7178, n15793);
xnor_4 g19288(new_n20552, new_n20538, n15812);
xnor_4 g19289(new_n11288, new_n11240, n15815);
xnor_4 g19290(new_n7613, new_n7612, n15816);
xnor_4 g19291(new_n10860, new_n10847, n15831);
xnor_4 g19292(new_n8703, new_n8702, n15846);
xnor_4 g19293(new_n7670_1, new_n7669, n15859);
and_5  g19294(new_n7345, n23272, new_n21643);
nor_5  g19295(new_n18252, new_n18236, new_n21644);
nor_5  g19296(new_n21644, new_n21643, new_n21645_1);
nor_5  g19297(new_n21645_1, new_n7344, new_n21646);
xnor_4 g19298(new_n21646, new_n19972, new_n21647);
xor_4  g19299(new_n18550, new_n18547, new_n21648);
xor_4  g19300(new_n21645_1, new_n7344, new_n21649_1);
nor_5  g19301(new_n21649_1, new_n21648, new_n21650);
nor_5  g19302(new_n18253, new_n18235, new_n21651);
nor_5  g19303(new_n18275, new_n18254_1, new_n21652);
or_5   g19304(new_n21652, new_n21651, new_n21653);
xnor_4 g19305(new_n21649_1, new_n18551, new_n21654_1);
and_5  g19306(new_n21654_1, new_n21653, new_n21655);
nor_5  g19307(new_n21655, new_n21650, new_n21656);
xnor_4 g19308(new_n21656, new_n21647, n15869);
xnor_4 g19309(new_n17308, new_n17281, n15885);
or_5   g19310(new_n19393, new_n14158, new_n21659);
nor_5  g19311(new_n19443, new_n21659, new_n21660);
and_5  g19312(new_n19442, new_n19393, new_n21661);
or_5   g19313(new_n21661, new_n21660, n15889);
xnor_4 g19314(new_n17295, new_n12550, n15917);
xor_4  g19315(new_n12545_1, new_n12544, n15922);
xor_4  g19316(new_n6479, new_n6478, n15947);
and_5  g19317(new_n17864, new_n6573, new_n21666);
or_5   g19318(new_n19097, new_n19092, new_n21667);
nor_5  g19319(new_n21667, new_n19091, new_n21668);
nor_5  g19320(new_n21668, new_n21666, new_n21669);
xnor_4 g19321(new_n21669, new_n17889_1, new_n21670);
xor_4  g19322(new_n19098, new_n19091, new_n21671);
nor_5  g19323(new_n21671, new_n17893, new_n21672);
nor_5  g19324(new_n19109, new_n19100, new_n21673);
or_5   g19325(new_n21673, new_n21672, new_n21674_1);
xor_4  g19326(new_n21674_1, new_n21670, n15956);
xor_4  g19327(new_n12316, new_n12313, n15958);
nor_5  g19328(new_n15571, new_n11033, new_n21677);
and_5  g19329(new_n15571, new_n15565, new_n21678);
nor_5  g19330(new_n21678, new_n21677, new_n21679);
nor_5  g19331(new_n15566, new_n11033, new_n21680_1);
or_5   g19332(new_n15568, new_n21680_1, new_n21681);
nor_5  g19333(new_n21681, new_n21679, n15986);
xnor_4 g19334(new_n21120, new_n21117, n16013);
nor_5  g19335(new_n20101, new_n21671, new_n21684);
nor_5  g19336(new_n20102, new_n19099, new_n21685_1);
nor_5  g19337(new_n20111, new_n21685_1, new_n21686);
nor_5  g19338(new_n21686, new_n21684, new_n21687_1);
xnor_4 g19339(new_n21669, new_n20102, new_n21688);
xnor_4 g19340(new_n21688, new_n21687_1, n16060);
nor_5  g19341(new_n14957, new_n15560, new_n21690);
xnor_4 g19342(new_n14957, new_n15560, new_n21691);
nor_5  g19343(new_n14959, new_n7860, new_n21692);
nor_5  g19344(new_n20776, new_n20765, new_n21693);
nor_5  g19345(new_n21693, new_n21692, new_n21694);
nor_5  g19346(new_n21694, new_n21691, new_n21695);
nor_5  g19347(new_n21695, new_n21690, new_n21696);
nor_5  g19348(new_n21696, new_n20883, new_n21697);
xor_4  g19349(new_n20980, new_n20972, new_n21698);
xor_4  g19350(new_n21696, new_n20883, new_n21699);
nor_5  g19351(new_n21699, new_n21698, new_n21700);
xnor_4 g19352(new_n21699, new_n21698, new_n21701);
xnor_4 g19353(new_n20978, new_n20975, new_n21702);
xor_4  g19354(new_n21694, new_n21691, new_n21703);
nor_5  g19355(new_n21703, new_n21702, new_n21704);
xnor_4 g19356(new_n21703, new_n21702, new_n21705);
and_5  g19357(new_n20796, new_n20777, new_n21706);
nor_5  g19358(new_n20812, new_n20797, new_n21707);
nor_5  g19359(new_n21707, new_n21706, new_n21708);
nor_5  g19360(new_n21708, new_n21705, new_n21709);
nor_5  g19361(new_n21709, new_n21704, new_n21710);
nor_5  g19362(new_n21710, new_n21701, new_n21711);
nor_5  g19363(new_n21711, new_n21700, new_n21712);
xnor_4 g19364(new_n21712, new_n21697, new_n21713);
xnor_4 g19365(new_n21713, new_n21590, n16062);
xnor_4 g19366(new_n21200, new_n21192, n16068);
xnor_4 g19367(new_n21420, new_n21417, n16080);
and_5  g19368(new_n20888, new_n5779, new_n21717_1);
nor_5  g19369(new_n20892, new_n20889, new_n21718);
nor_5  g19370(new_n21718, new_n21717_1, new_n21719_1);
nor_5  g19371(new_n20883, new_n10819, new_n21720);
nor_5  g19372(new_n20887, new_n20884, new_n21721);
nor_5  g19373(new_n21721, new_n21720, new_n21722);
xnor_4 g19374(new_n21722, new_n21719_1, n16098);
xnor_4 g19375(new_n16076, new_n16068_1, n16110);
xnor_4 g19376(new_n13817, new_n13791, n16142);
xnor_4 g19377(new_n15157, new_n15145_1, n16185);
xnor_4 g19378(new_n11330_1, new_n11312, n16196);
xnor_4 g19379(new_n19125_1, new_n19124, n16206);
xor_4  g19380(new_n19201, new_n19198, n16215);
xnor_4 g19381(new_n17406, new_n17398, n16218);
xor_4  g19382(new_n3683, new_n3681, n16219);
xnor_4 g19383(new_n6292, new_n6291, n16230);
xor_4  g19384(new_n7667, new_n7659, n16243);
xnor_4 g19385(new_n15831_1, new_n15822, n16275);
xnor_4 g19386(new_n9258, new_n9257, n16279);
nor_5  g19387(new_n18731, new_n19147, new_n21736);
nor_5  g19388(new_n18786, new_n18732, new_n21737);
or_5   g19389(new_n21737, new_n21736, n16322);
xnor_4 g19390(new_n15839, new_n15807, n16327);
xnor_4 g19391(new_n19565, new_n19558, n16350);
xor_4  g19392(new_n6047, new_n6045, n16367);
xnor_4 g19393(new_n17504, new_n17503, n16379);
xnor_4 g19394(new_n18369, new_n18350_1, n16398);
xnor_4 g19395(new_n12304_1, new_n12303, n16406);
xnor_4 g19396(new_n20304, new_n20288, n16407);
xnor_4 g19397(new_n21710, new_n21701, n16419);
xnor_4 g19398(new_n7630_1, new_n7587, n16424);
xor_4  g19399(new_n12649, new_n12590, new_n21748);
xnor_4 g19400(new_n21748, new_n12689, n16428);
xnor_4 g19401(new_n10876, new_n10818, n16433);
xnor_4 g19402(new_n10872, new_n10826, n16440);
xnor_4 g19403(new_n16078, new_n16064, n16445);
xnor_4 g19404(new_n12890, new_n12838, n16460);
xnor_4 g19405(new_n18271, new_n18262, n16481);
nor_5  g19406(new_n13448, new_n10033, new_n21755);
nor_5  g19407(new_n13448, new_n10038, new_n21756);
nor_5  g19408(new_n18846, new_n18831_1, new_n21757);
or_5   g19409(new_n21757, new_n21756, new_n21758);
xnor_4 g19410(new_n13448, new_n10033, new_n21759);
nor_5  g19411(new_n21759, new_n21758, new_n21760);
nor_5  g19412(new_n21760, new_n21755, n16493);
xnor_4 g19413(new_n4400, new_n4377, n16506);
xnor_4 g19414(new_n11658, new_n11657, n16516);
xor_4  g19415(new_n20395, new_n20394, n16517);
xnor_4 g19416(new_n14262, new_n14261, n16527);
xnor_4 g19417(new_n9791, new_n8344, n16554);
xor_4  g19418(new_n5604, new_n5330_1, n16583);
xnor_4 g19419(new_n19857, new_n9145, new_n21768);
xnor_4 g19420(new_n21768, new_n19862, n16584);
xnor_4 g19421(new_n17581, new_n17560, n16589);
xor_4  g19422(new_n17906, new_n17905, n16596);
xnor_4 g19423(new_n20564, new_n20524, n16617);
xnor_4 g19424(new_n6912, new_n6880, n16630);
xor_4  g19425(new_n20546, new_n4559, n16640);
xor_4  g19426(new_n2505, new_n2504, n16656);
xnor_4 g19427(new_n6304, new_n6264, n16674);
xnor_4 g19428(new_n12888, new_n12842, n16682);
xnor_4 g19429(new_n20491, new_n20471, n16684);
xnor_4 g19430(new_n9566, new_n9562, n16688);
xnor_4 g19431(new_n5820, new_n5813, n16733);
xor_4  g19432(new_n7186, new_n7185, n16798);
xnor_4 g19433(new_n15255_1, new_n15254, n16834);
xnor_4 g19434(new_n2961_1, new_n2925, n16837);
xnor_4 g19435(new_n20109, new_n20106, n16841);
xnor_4 g19436(new_n4699, new_n4698, n16885);
xnor_4 g19437(new_n7457, new_n7400, n16905);
nor_5  g19438(new_n20028, new_n20025, new_n21787);
xnor_4 g19439(new_n21787, new_n16565, n16951);
xor_4  g19440(new_n14768, new_n14759, n16954);
xor_4  g19441(new_n7611, new_n3497, n16989);
xnor_4 g19442(new_n17506, new_n17476, n17006);
xnor_4 g19443(new_n12215, new_n12214, n17068);
xnor_4 g19444(new_n13808, new_n13806, n17070);
xnor_4 g19445(new_n18782_1, new_n18739, n17075);
xnor_4 g19446(new_n15508_1, new_n15492, n17084);
xnor_4 g19447(new_n4393, new_n4392, n17104);
xnor_4 g19448(new_n12023, new_n12001, n17106);
xor_4  g19449(new_n8820, new_n8809_1, n17119);
xnor_4 g19450(new_n11921, new_n11889, n17130);
xnor_4 g19451(new_n21013, new_n20998, n17138);
xnor_4 g19452(new_n20397, new_n20389, n17163);
xor_4  g19453(new_n18449, new_n18448, n17168);
xnor_4 g19454(new_n10398, new_n10389, n17202);
xor_4  g19455(new_n17728, new_n17727, n17219);
xnor_4 g19456(new_n16990, new_n16960, n17232);
xnor_4 g19457(new_n13906, new_n13902, n17236);
xor_4  g19458(new_n9485, new_n9484, n17243);
xnor_4 g19459(new_n10074, new_n10060, n17263);
and_5  g19460(new_n17889_1, new_n17881, new_n21809);
nor_5  g19461(new_n17910, new_n17890, new_n21810);
nor_5  g19462(new_n21810, new_n21809, n17285);
xnor_4 g19463(new_n10564_1, new_n10536, n17320);
xnor_4 g19464(new_n2761_1, new_n2719, n17337);
xnor_4 g19465(new_n20228, new_n20219, n17344);
xnor_4 g19466(new_n20236, new_n20201, n17359);
xnor_4 g19467(new_n12870_1, new_n12071, n17387);
xor_4  g19468(new_n4697, new_n4695, n17391);
xnor_4 g19469(new_n17501, new_n17482, n17392);
xnor_4 g19470(new_n20493, new_n20468, n17421);
xnor_4 g19471(new_n11009, new_n5970, n17432);
xnor_4 g19472(new_n19433, new_n19413, n17436);
xor_4  g19473(new_n6478, new_n4360, n17440);
xnor_4 g19474(new_n7699, new_n5330_1, n17450);
or_5   g19475(new_n17269, new_n17267, new_n21824);
nor_5  g19476(new_n21824, new_n6682, new_n21825);
nor_5  g19477(new_n6681, new_n17236_1, new_n21826);
nor_5  g19478(new_n6682, new_n6643, new_n21827);
nor_5  g19479(new_n6742, new_n21827, new_n21828);
nor_5  g19480(new_n21828, new_n21826, new_n21829);
nor_5  g19481(new_n21829, new_n21825, new_n21830);
nor_5  g19482(new_n17270, new_n6681, new_n21831);
nor_5  g19483(new_n21831, new_n21828, new_n21832_1);
nor_5  g19484(new_n21832_1, new_n21830, n17461);
xor_4  g19485(new_n21381, new_n21380, n17466);
xnor_4 g19486(new_n12229, new_n12190, n17493);
xor_4  g19487(new_n19898, new_n19895, n17500);
xnor_4 g19488(new_n20752, new_n20749, n17524);
xnor_4 g19489(new_n5298, new_n5263, n17529);
xnor_4 g19490(new_n13624, new_n5327, new_n21839_1);
xnor_4 g19491(new_n21839_1, new_n13627, n17557);
xnor_4 g19492(new_n15165_1, new_n15129, n17583);
xnor_4 g19493(new_n12880, new_n12858, n17592);
xnor_4 g19494(new_n7618, new_n7606, n17638);
xnor_4 g19495(new_n18273, new_n18258, n17687);
xnor_4 g19496(new_n12509, new_n12471, n17721);
xnor_4 g19497(new_n20080, new_n20060, n17735);
not_10 g19498(new_n19502, new_n21847);
or_5   g19499(new_n21847, new_n9163, new_n21848);
nor_5  g19500(new_n21848, new_n19501, new_n21849);
and_5  g19501(new_n21847, new_n9163, new_n21850);
and_5  g19502(new_n21850, new_n19501, new_n21851);
nor_5  g19503(new_n21851, new_n21849, new_n21852);
and_5  g19504(new_n21852, new_n19574, new_n21853);
or_5   g19505(new_n21852, new_n19574, new_n21854);
nor_5  g19506(new_n19504, new_n19494_1, new_n21855);
nor_5  g19507(new_n19515_1, new_n19505, new_n21856);
nor_5  g19508(new_n21856, new_n21855, new_n21857);
and_5  g19509(new_n21857, new_n21854, new_n21858);
or_5   g19510(new_n21858, new_n21849, new_n21859);
nor_5  g19511(new_n21859, new_n21853, n17738);
xor_4  g19512(new_n13986, new_n13983, n17746);
xnor_4 g19513(new_n21174, new_n21170, n17749);
xnor_4 g19514(new_n17141, new_n17123, n17820);
xnor_4 g19515(new_n12878, new_n12862, n17855);
and_5  g19516(new_n4533, new_n4530, new_n21865);
and_5  g19517(new_n4583, new_n21865, new_n21866);
nor_5  g19518(new_n4583, new_n20521, new_n21867);
or_5   g19519(new_n21867, new_n21866, new_n21868);
and_5  g19520(new_n4584, new_n4440, new_n21869);
nor_5  g19521(new_n4650, new_n4585, new_n21870);
nor_5  g19522(new_n21870, new_n21869, new_n21871);
nor_5  g19523(new_n21871, new_n21868, new_n21872);
nor_5  g19524(new_n21872, new_n21866, n17877);
xnor_4 g19525(new_n14155, new_n14154, n17889);
and_5  g19526(new_n21067, new_n21057, new_n21875);
nor_5  g19527(new_n21078_1, new_n21875, new_n21876);
nor_5  g19528(new_n21067, new_n21057, new_n21877);
nor_5  g19529(new_n21077, new_n21877, new_n21878);
nor_5  g19530(new_n21878, new_n21876, n17912);
xor_4  g19531(new_n20484, new_n20480, n17927);
xnor_4 g19532(new_n20556, new_n20534, n17931);
xnor_4 g19533(new_n7181, new_n7180, n17948);
xor_4  g19534(new_n14355, new_n14352, n17956);
nor_5  g19535(new_n11614, new_n11423, new_n21884);
nor_5  g19536(new_n11549, new_n11423, new_n21885);
nor_5  g19537(new_n11613, new_n21885, new_n21886);
nor_5  g19538(new_n21886, new_n21884, n17963);
nor_5  g19539(n25494, new_n20639, new_n21888);
nor_5  g19540(new_n16058, new_n16043, new_n21889);
nor_5  g19541(new_n21889, new_n21888, new_n21890);
not_10 g19542(new_n21890, new_n21891);
nor_5  g19543(new_n21891, new_n11884, new_n21892);
nor_5  g19544(new_n21890, new_n11887, new_n21893);
xor_4  g19545(new_n21890, new_n11887, new_n21894);
and_5  g19546(new_n16059, new_n16042, new_n21895);
nor_5  g19547(new_n16080_1, new_n16060_1, new_n21896);
nor_5  g19548(new_n21896, new_n21895, new_n21897);
and_5  g19549(new_n21897, new_n21894, new_n21898_1);
nor_5  g19550(new_n21898_1, new_n21893, new_n21899);
nor_5  g19551(new_n21899, new_n21892, new_n21900);
and_5  g19552(new_n21891, new_n11884, new_n21901);
nor_5  g19553(new_n21901, new_n21898_1, new_n21902);
nor_5  g19554(new_n21902, new_n21900, n17976);
xnor_4 g19555(new_n6496, new_n6460, n17998);
xnor_4 g19556(new_n13267, new_n2746, n18025);
xnor_4 g19557(new_n19080, new_n19079, n18043);
xnor_4 g19558(new_n20411_1, new_n20408, n18045);
xnor_4 g19559(new_n3687, new_n3677, n18059);
xnor_4 g19560(new_n18780_1, new_n18742, n18061);
xnor_4 g19561(new_n3239, new_n3186, n18071);
xnor_4 g19562(new_n9092, new_n9040, n18143);
xnor_4 g19563(new_n19900, new_n19893, n18152);
xnor_4 g19564(new_n6904, new_n6896, n18193);
xor_4  g19565(new_n10604, new_n10595_1, new_n21914);
xnor_4 g19566(new_n21914, new_n10617_1, n18232);
xnor_4 g19567(new_n15510, new_n15488, n18238);
xnor_4 g19568(new_n16979, new_n16976, n18241);
xnor_4 g19569(new_n19429, new_n19421, n18254);
xnor_4 g19570(new_n20078, new_n20062, n18288);
xnor_4 g19571(new_n11079, new_n11038, n18301);
xnor_4 g19572(new_n20399, new_n20386, n18304);
xnor_4 g19573(new_n12233, new_n12184, n18310);
xnor_4 g19574(new_n6049, new_n6048, n18311);
xnor_4 g19575(new_n16197, new_n16182, n18323);
xnor_4 g19576(new_n5018, new_n4984, n18332);
xor_4  g19577(new_n20567, new_n20566, n18343);
xnor_4 g19578(new_n17808, new_n17805, n18350);
xnor_4 g19579(new_n16621, new_n16620, n18362);
xnor_4 g19580(new_n4646_1, new_n4594, n18377);
xnor_4 g19581(new_n3838, new_n3819, n18405);
xnor_4 g19582(new_n15373, new_n15364, n18414);
xnor_4 g19583(new_n13343, new_n13335, n18418);
xnor_4 g19584(new_n7451, new_n7412, n18437);
xnor_4 g19585(new_n18595, new_n18556, n18439);
xnor_4 g19586(new_n10139, new_n10138, n18445);
xnor_4 g19587(new_n6302, new_n6268, n18467);
xnor_4 g19588(new_n16996, new_n16947, n18482);
xnor_4 g19589(new_n17306, new_n17284, n18509);
xnor_4 g19590(new_n12714, new_n8234, n18513);
xnor_4 g19591(new_n13815, new_n13814, n18515);
xnor_4 g19592(new_n14629, new_n14610, n18572);
and_5  g19593(new_n21712, new_n21697, new_n21942);
nor_5  g19594(new_n21942, new_n21590, new_n21943_1);
or_5   g19595(new_n21712, new_n21697, new_n21944);
and_5  g19596(new_n21944, new_n21590, new_n21945);
nor_5  g19597(new_n21945, new_n21943_1, n18574);
xnor_4 g19598(new_n19563, new_n19560, n18576);
xnor_4 g19599(new_n20873, new_n20865, n18582);
xnor_4 g19600(new_n18367, new_n18354, n18583);
xnor_4 g19601(new_n18766, new_n18765, n18610);
xor_4  g19602(new_n20425, new_n20422, n18635);
xnor_4 g19603(new_n6122, new_n6121, n18653);
xnor_4 g19604(new_n3514, new_n3467, n18679);
xnor_4 g19605(new_n18890, new_n18882, n18693);
xnor_4 g19606(new_n2959, new_n2929_1, n18708);
xnor_4 g19607(new_n21211, new_n15587, new_n21956);
xnor_4 g19608(new_n21956, new_n21216, n18721);
xnor_4 g19609(new_n17147, new_n17114, n18725);
xnor_4 g19610(new_n19233_1, new_n19212, n18751);
xnor_4 g19611(new_n15159, new_n15141, n18780);
xnor_4 g19612(new_n18025_1, new_n17983, n18782);
not_10 g19613(new_n6789, new_n21962);
nor_5  g19614(new_n6859, new_n21962, new_n21963);
nor_5  g19615(new_n6922, new_n21963, new_n21964);
and_5  g19616(new_n6859, new_n21962, new_n21965);
nor_5  g19617(new_n6921, new_n21965, new_n21966);
nor_5  g19618(new_n21966, new_n21964, n18802);
xor_4  g19619(new_n9887, new_n9886, n18830);
xor_4  g19620(new_n11690, new_n11684, n18831);
xnor_4 g19621(new_n10858, new_n10850, n18843);
xnor_4 g19622(new_n2955, new_n2938, n18858);
xnor_4 g19623(new_n9080, new_n9064, n18859);
xnor_4 g19624(new_n15841, new_n15803, n18864);
xnor_4 g19625(new_n4264, new_n4205_1, n18865);
xnor_4 g19626(new_n19830, new_n19829, n18886);
xnor_4 g19627(new_n15155, new_n15154, n18887);
xnor_4 g19628(new_n8096, new_n8061, n18919);
xnor_4 g19629(new_n11276, new_n11265, n18940);
xor_4  g19630(new_n21331, new_n21330, n18945);
xnor_4 g19631(new_n21048, new_n21034_1, n18970);
xnor_4 g19632(new_n15566, new_n11036, new_n21981_1);
xnor_4 g19633(new_n21981_1, new_n15571, n18977);
xnor_4 g19634(new_n13908, new_n13899, n18982);
xor_4  g19635(new_n19312, new_n19311, n18999);
xnor_4 g19636(new_n5304, new_n5251, n19044);
xor_4  g19637(new_n13629, new_n13622, n19125);
xnor_4 g19638(new_n5302_1, new_n5255_1, n19141);
xnor_4 g19639(new_n15940, new_n12835, new_n21988);
nor_5  g19640(new_n15953, new_n12840, new_n21989);
xnor_4 g19641(new_n15953, new_n12840, new_n21990);
and_5  g19642(new_n15945, new_n12843_1, new_n21991);
nor_5  g19643(new_n17178, new_n17159, new_n21992);
nor_5  g19644(new_n21992, new_n21991, new_n21993_1);
nor_5  g19645(new_n21993_1, new_n21990, new_n21994);
nor_5  g19646(new_n21994, new_n21989, new_n21995);
xnor_4 g19647(new_n21995, new_n21988, n19164);
xnor_4 g19648(new_n7626, new_n7625, n19174);
xnor_4 g19649(new_n19481, new_n19478, n19176);
xnor_4 g19650(new_n20401, new_n20383, n19202);
xnor_4 g19651(new_n18685, new_n18675, n19220);
xor_4  g19652(new_n7198, new_n7148, n19221);
xnor_4 g19653(new_n10261_1, new_n10260, n19223);
xor_4  g19654(new_n15827, new_n15826, n19224);
xnor_4 g19655(new_n14296, new_n14286, n19233);
xnor_4 g19656(new_n11672, new_n11641, n19244);
xnor_4 g19657(new_n8098, new_n8057, n19314);
xnor_4 g19658(new_n9800, new_n9799, n19315);
xnor_4 g19659(new_n12225_1, new_n12196, n19323);
xnor_4 g19660(new_n20226, new_n20223, n19333);
nor_5  g19661(new_n15937, new_n15933, new_n22010);
nor_5  g19662(new_n22010, new_n9031, new_n22011);
nor_5  g19663(new_n15938, new_n9034, new_n22012);
nor_5  g19664(new_n15958_1, new_n15939, new_n22013);
or_5   g19665(new_n22013, new_n22012, new_n22014);
xnor_4 g19666(new_n22010, new_n9031, new_n22015);
nor_5  g19667(new_n22015, new_n22014, new_n22016_1);
nor_5  g19668(new_n22016_1, new_n22011, n19348);
xnor_4 g19669(new_n15522, new_n15463, n19354);
xnor_4 g19670(new_n10081, new_n10051, n19367);
xnor_4 g19671(new_n17647, new_n17626, n19385);
or_5   g19672(new_n15586, new_n10325, new_n22021);
xnor_4 g19673(new_n15636_1, new_n22021, new_n22022);
xnor_4 g19674(new_n22022, new_n15662_1, n19389);
xnor_4 g19675(new_n15029, new_n14997, n19401);
xor_4  g19676(new_n20667, new_n20659, n19414);
xor_4  g19677(new_n17828, new_n16454, n19424);
xnor_4 g19678(new_n19834, new_n19816, n19450);
not_10 g19679(new_n22010, new_n22028);
nor_5  g19680(new_n22028, new_n12775, new_n22029);
xor_4  g19681(new_n22010, new_n12775, new_n22030);
nor_5  g19682(new_n15938, new_n12830, new_n22031);
xnor_4 g19683(new_n15938, new_n12830, new_n22032);
and_5  g19684(new_n15940, new_n12835, new_n22033);
nor_5  g19685(new_n21995, new_n21988, new_n22034);
nor_5  g19686(new_n22034, new_n22033, new_n22035);
nor_5  g19687(new_n22035, new_n22032, new_n22036);
nor_5  g19688(new_n22036, new_n22031, new_n22037);
nor_5  g19689(new_n22037, new_n22030, new_n22038);
or_5   g19690(new_n22038, new_n22029, n19458);
xnor_4 g19691(new_n13988, new_n13980, n19467);
xnor_4 g19692(new_n7453, new_n7408_1, n19496);
xor_4  g19693(new_n13947, new_n13939, n19523);
xnor_4 g19694(new_n4256_1, new_n4221_1, n19570);
xnor_4 g19695(new_n10974, new_n10965, n19602);
xnor_4 g19696(new_n11323, new_n11317, n19617);
xnor_4 g19697(new_n12507_1, new_n12475, n19623);
xor_4  g19698(new_n20705_1, new_n20704_1, n19641);
xnor_4 g19699(new_n20495_1, new_n20465, n19648);
xnor_4 g19700(new_n14627, new_n14613, n19664);
xnor_4 g19701(new_n18446, new_n18432, n19736);
nor_5  g19702(new_n20669, new_n20655, new_n22051);
nor_5  g19703(new_n20655, new_n3053, new_n22052);
nor_5  g19704(new_n20668, new_n22052, new_n22053);
nor_5  g19705(new_n22053, new_n22051, n19749);
xnor_4 g19706(new_n13692, new_n13679, n19756);
xnor_4 g19707(new_n10972, new_n10971, n19767);
xnor_4 g19708(new_n3180, new_n20170, new_n22057);
xnor_4 g19709(new_n22057, new_n3241, n19780);
xnor_4 g19710(new_n21234, new_n21231, n19792);
xnor_4 g19711(new_n19069, new_n19056, n19798);
xor_4  g19712(new_n15252, new_n15249, n19873);
nor_5  g19713(new_n17024, new_n17007, new_n22062);
not_10 g19714(new_n17013, new_n22063_1);
nor_5  g19715(new_n22063_1, new_n17007, new_n22064);
nor_5  g19716(new_n17023, new_n22064, new_n22065);
nor_5  g19717(new_n22065, new_n22062, n19909);
xnor_4 g19718(new_n18444_1, new_n18436, n19916);
xnor_4 g19719(new_n19073, new_n19050, n19923);
xnor_4 g19720(new_n17508, new_n17472, n19930);
xnor_4 g19721(new_n5838, new_n5747, n19968);
xnor_4 g19722(new_n18013, new_n18001, n19988);
and_5  g19723(new_n19858, new_n19138, new_n22072_1);
nor_5  g19724(new_n19138, new_n9207, new_n22073);
nor_5  g19725(new_n19142, new_n19139, new_n22074);
nor_5  g19726(new_n22074, new_n22073, new_n22075);
nor_5  g19727(new_n22075, new_n22072_1, new_n22076_1);
nor_5  g19728(new_n19858, new_n19138, new_n22077);
nor_5  g19729(new_n22077, new_n22074, new_n22078);
nor_5  g19730(new_n22078, new_n22076_1, n20004);
xnor_4 g19731(new_n19229, new_n19216, n20017);
xnor_4 g19732(new_n16992, new_n16956, n20033);
xnor_4 g19733(new_n12681, new_n12680, n20061);
xnor_4 g19734(new_n16577, new_n16574, n20069);
and_5  g19735(new_n13232, new_n13225, new_n22084);
nor_5  g19736(new_n13289, new_n13233, new_n22085);
or_5   g19737(new_n22085, new_n22084, n20086);
xnor_4 g19738(new_n17903, new_n17900, n20096);
xnor_4 g19739(new_n12217, new_n12210, n20103);
xnor_4 g19740(new_n10566, new_n10532, n20126);
xnor_4 g19741(new_n19634, new_n19605, n20149);
xnor_4 g19742(new_n10870, new_n10830, n20187);
xnor_4 g19743(new_n16038, new_n16010, n20279);
or_5   g19744(new_n20858, new_n20856, new_n22093);
nor_5  g19745(new_n22093, new_n20854, new_n22094);
or_5   g19746(new_n20862, new_n22094, new_n22095);
nor_5  g19747(new_n20875, new_n20859, new_n22096);
nor_5  g19748(new_n20874, new_n20864, new_n22097);
nor_5  g19749(new_n22097, new_n16176, new_n22098);
or_5   g19750(new_n22098, new_n22096, new_n22099);
nor_5  g19751(new_n22099, new_n22095, n20287);
xnor_4 g19752(new_n18922, new_n18919_1, n20301);
nor_5  g19753(new_n7459, new_n7396, new_n22102);
nor_5  g19754(new_n22102, new_n7299, n20330);
xnor_4 g19755(new_n10866, new_n10836, n20333);
not_10 g19756(new_n9308_1, new_n22105);
nand_5 g19757(new_n9430_1, new_n22105, new_n22106);
nor_5  g19758(new_n9491, new_n22106, new_n22107_1);
nor_5  g19759(new_n9430_1, new_n22105, new_n22108);
and_5  g19760(new_n9491, new_n22108, new_n22109);
or_5   g19761(new_n22109, new_n22107_1, n20355);
xor_4  g19762(new_n7660, new_n4803, n20366);
xnor_4 g19763(new_n17681, new_n17677, n20388);
xnor_4 g19764(new_n20554, new_n20536, n20402);
xnor_4 g19765(new_n14142, new_n14119, n20403);
xor_4  g19766(new_n2945, new_n2944_1, n20424);
xnor_4 g19767(new_n18770, new_n18759, n20436);
xor_4  g19768(new_n7439, new_n7438, n20441);
xnor_4 g19769(new_n6920, new_n6864, n20445);
xnor_4 g19770(new_n4648, new_n4589, n20450);
xnor_4 g19771(new_n15170, new_n6047, n20490);
xor_4  g19772(new_n18683, new_n18680, n20495);
nor_5  g19773(new_n14159, new_n14158, new_n22122);
and_5  g19774(new_n22122, new_n14157, new_n22123);
nand_5 g19775(new_n14159, new_n14158, new_n22124_1);
nor_5  g19776(new_n22124_1, new_n14157, new_n22125);
or_5   g19777(new_n22125, new_n22123, n20515);
nor_5  g19778(new_n21236, new_n21227, new_n22127);
nor_5  g19779(new_n22127, new_n21223, n20533);
xnor_4 g19780(new_n16456, new_n16450, n20582);
xnor_4 g19781(new_n18167, new_n18140, n20590);
xnor_4 g19782(new_n3223, new_n3220, n20602);
xnor_4 g19783(new_n15152, new_n15151, n20609);
xnor_4 g19784(new_n5973, new_n5966, n20623);
xnor_4 g19785(new_n19084, new_n19034, n20629);
xnor_4 g19786(new_n12678, new_n12669, n20661);
xnor_4 g19787(new_n7702, new_n7701, n20673);
xnor_4 g19788(new_n19077, new_n19043, n20678);
nor_5  g19789(new_n13667, new_n13634, new_n22138);
nor_5  g19790(new_n13698, new_n22138, new_n22139);
and_5  g19791(new_n13667, new_n13634, new_n22140);
or_5   g19792(new_n22140, new_n13664, new_n22141);
nor_5  g19793(new_n22141, new_n22139, n20680);
xnor_4 g19794(new_n5816, new_n3883, n20685);
xnor_4 g19795(new_n21890, new_n11884, new_n22144_1);
xnor_4 g19796(new_n22144_1, new_n21899, n20691);
xnor_4 g19797(new_n14625, new_n14617, n20696);
xnor_4 g19798(new_n21011, new_n21002, n20704);
xor_4  g19799(new_n20072, new_n20071, n20705);
xnor_4 g19800(new_n9090_1, new_n9044, n20709);
xnor_4 g19801(new_n13588, new_n13564, n20713);
xnor_4 g19802(new_n7848, new_n7847, n20722);
not_10 g19803(new_n21506, new_n22152);
and_5  g19804(new_n22152, new_n18066, new_n22153);
nor_5  g19805(new_n18066, new_n18056, new_n22154);
and_5  g19806(new_n18066, new_n18056, new_n22155);
nor_5  g19807(new_n18077, new_n22155, new_n22156);
nor_5  g19808(new_n22156, new_n22154, new_n22157_1);
nor_5  g19809(new_n22157_1, new_n22153, new_n22158);
nor_5  g19810(new_n22152, new_n18066, new_n22159);
nor_5  g19811(new_n22159, new_n22156, new_n22160);
nor_5  g19812(new_n22160, new_n22158, n20723);
xnor_4 g19813(new_n20854, new_n16176, new_n22162);
xnor_4 g19814(new_n22162, new_n22097, n20748);
xor_4  g19815(new_n5010, new_n5000, n20761);
xnor_4 g19816(new_n18778, new_n18746, n20774);
xnor_4 g19817(new_n22037, new_n22030, n20788);
nor_5  g19818(new_n21358, new_n20419, new_n22167);
nor_5  g19819(new_n22167, new_n21468, new_n22168);
and_5  g19820(new_n21358, new_n20419, new_n22169);
nor_5  g19821(new_n22169, new_n21467, new_n22170);
nor_5  g19822(new_n22170, new_n22168, n20795);
xnor_4 g19823(new_n18812, new_n18801, new_n22172);
and_5  g19824(new_n18819, new_n18801, new_n22173_1);
nor_5  g19825(new_n22173_1, new_n18821, new_n22174);
nor_5  g19826(new_n22174, new_n18820, new_n22175);
xnor_4 g19827(new_n22175, new_n22172, n20803);
xor_4  g19828(new_n21871, new_n21868, n20869);
xnor_4 g19829(new_n21176_1, new_n21166, n20879);
xnor_4 g19830(new_n5826, new_n5801, n20915);
xor_4  g19831(new_n19955, new_n19952, new_n22180);
xor_4  g19832(n19282, n2160, new_n22181);
nor_5  g19833(n12657, new_n15221, new_n22182);
nor_5  g19834(new_n20088, new_n20085, new_n22183);
nor_5  g19835(new_n22183, new_n22182, new_n22184);
xor_4  g19836(new_n22184, new_n22181, new_n22185);
nor_5  g19837(new_n22185, new_n22180, new_n22186);
nor_5  g19838(new_n20089, new_n18396, new_n22187);
nor_5  g19839(new_n20093, new_n20090, new_n22188);
nor_5  g19840(new_n22188, new_n22187, new_n22189);
xnor_4 g19841(new_n22185, new_n22180, new_n22190);
nor_5  g19842(new_n22190, new_n22189, new_n22191);
nor_5  g19843(new_n22191, new_n22186, new_n22192);
nor_5  g19844(n19282, new_n21355, new_n22193);
nor_5  g19845(new_n22184, new_n22181, new_n22194);
nor_5  g19846(new_n22194, new_n22193, new_n22195);
nand_5 g19847(new_n22195, new_n21072, new_n22196);
nor_5  g19848(new_n22196, new_n22192, new_n22197);
and_5  g19849(new_n22197, new_n21067, new_n22198_1);
or_5   g19850(new_n21066, new_n21061, new_n22199);
nor_5  g19851(new_n22195, new_n21072, new_n22200);
and_5  g19852(new_n22200, new_n22192, new_n22201_1);
and_5  g19853(new_n22201_1, new_n22199, new_n22202);
or_5   g19854(new_n22202, new_n22198_1, n20935);
xnor_4 g19855(new_n20489_1, new_n20474, n20936);
xnor_4 g19856(new_n15551, new_n15550, n21008);
xnor_4 g19857(new_n18023, new_n17986, n21017);
and_5  g19858(new_n21571, new_n19922_1, new_n22207);
nor_5  g19859(new_n21571, new_n19922_1, new_n22208);
nor_5  g19860(new_n21575, new_n22208, new_n22209);
or_5   g19861(new_n22209, new_n21570, new_n22210);
nor_5  g19862(new_n22210, new_n22207, n21034);
xor_4  g19863(new_n20631, new_n20630, n21046);
xnor_4 g19864(new_n7789, new_n7772, n21062);
xor_4  g19865(new_n21314, new_n21306, new_n22214);
xnor_4 g19866(new_n22214, new_n21223, n21093);
xnor_4 g19867(new_n8853, new_n7174, n21094);
xnor_4 g19868(new_n13481, new_n13459, n21123);
xor_4  g19869(new_n17404, new_n16643, n21154);
xnor_4 g19870(new_n14271_1, new_n14248, n21157);
xnor_4 g19871(new_n19626, new_n19618_1, n21168);
xor_4  g19872(new_n6717, new_n6716, n21173);
xnor_4 g19873(new_n4252, new_n4229, n21176);
xnor_4 g19874(new_n13159, new_n13152, n21182);
not_10 g19875(new_n20458, new_n22224);
nor_5  g19876(new_n22224, new_n19659, new_n22225);
nor_5  g19877(new_n20497, new_n19652_1, new_n22226);
or_5   g19878(new_n22226, new_n22225, new_n22227);
nor_5  g19879(new_n20496, new_n20464, new_n22228);
nor_5  g19880(new_n22228, new_n19662, new_n22229);
or_5   g19881(new_n22229, new_n20461, new_n22230);
nor_5  g19882(new_n22230, new_n22227, n21193);
xnor_4 g19883(new_n8626, new_n8625, n21203);
xor_4  g19884(new_n15150, new_n2524, n21225);
xnor_4 g19885(new_n18381, new_n18329, n21238);
xnor_4 g19886(new_n12683, new_n12663, n21254);
xnor_4 g19887(new_n18591, new_n18562, n21298);
xnor_4 g19888(new_n18360, new_n8539, n21302);
xnor_4 g19889(new_n18442, new_n18439_1, n21349);
xnor_4 g19890(new_n14772_1, new_n14770, n21365);
xnor_4 g19891(new_n13949, new_n13936, n21367);
xnor_4 g19892(new_n10759, new_n10732, n21396);
xnor_4 g19893(new_n6918, new_n6868, n21399);
xor_4  g19894(new_n3248, new_n3243, n21404);
xnor_4 g19895(new_n7704, new_n7695, n21446);
xnor_4 g19896(new_n10615, new_n10607, n21472);
xnor_4 g19897(new_n6736_1, new_n6695, n21525);
xnor_4 g19898(new_n15884_1, new_n15861, n21549);
xnor_4 g19899(new_n18269, new_n18266, n21615);
nor_5  g19900(new_n20859, new_n7137, new_n22249);
xnor_4 g19901(new_n20859, new_n7137, new_n22250);
nor_5  g19902(new_n16176, new_n12311, new_n22251);
nor_5  g19903(new_n16202, new_n16177, new_n22252);
nor_5  g19904(new_n22252, new_n22251, new_n22253_1);
nor_5  g19905(new_n22253_1, new_n22250, new_n22254);
nor_5  g19906(new_n22254, new_n22249, n21628);
and_5  g19907(new_n20131, new_n19660, new_n22256);
xnor_4 g19908(new_n20131, new_n19660, new_n22257);
nor_5  g19909(new_n20134, new_n19660, new_n22258);
nor_5  g19910(new_n21435, new_n21432, new_n22259);
nor_5  g19911(new_n22259, new_n22258, new_n22260);
nor_5  g19912(new_n22260, new_n22257, new_n22261);
nor_5  g19913(new_n22261, new_n22256, n21637);
xnor_4 g19914(new_n20074, new_n20067, n21645);
xor_4  g19915(new_n11004, new_n5967, n21665);
xnor_4 g19916(new_n13696, new_n13673, n21680);
xnor_4 g19917(new_n20562, new_n20526, n21685);
xnor_4 g19918(new_n17143, new_n17120, n21717);
xnor_4 g19919(new_n15538, new_n15533, n21719);
xnor_4 g19920(new_n17135, new_n17132, n21750);
xnor_4 g19921(new_n20324, new_n20323, n21765);
xnor_4 g19922(new_n22190, new_n22189, n21800);
xnor_4 g19923(new_n3994, new_n3990, new_n22272);
xnor_4 g19924(new_n22272, new_n3998, n21820);
xnor_4 g19925(new_n18017, new_n17995, n21874);
xnor_4 g19926(new_n12219, new_n12207, n21943);
xnor_4 g19927(new_n14776, new_n14754, n21960);
xor_4  g19928(new_n6485_1, new_n6484, n21976);
xnor_4 g19929(new_n10270, new_n10242, n21986);
xnor_4 g19930(new_n10083, new_n10048, n22016);
xnor_4 g19931(new_n17137, new_n17129, n22027);
xnor_4 g19932(new_n12019, new_n12011_1, n22050);
xnor_4 g19933(new_n3884, new_n3883, n22063);
xnor_4 g19934(new_n19624, new_n19621, n22076);
or_5   g19935(new_n12645, new_n12643, new_n22284);
nor_5  g19936(new_n18805, new_n22284, new_n22285);
nor_5  g19937(new_n19133, new_n19112, new_n22286);
nor_5  g19938(new_n22286, new_n22285, n22090);
xnor_4 g19939(new_n21046_1, new_n21037, n22107);
xnor_4 g19940(new_n16359, new_n16335, n22113);
nor_5  g19941(new_n12646, new_n12590, new_n22290_1);
nor_5  g19942(new_n12691, new_n22290_1, new_n22291);
and_5  g19943(new_n12646, new_n12590, new_n22292);
nor_5  g19944(new_n12690, new_n22292, new_n22293);
nor_5  g19945(new_n22293, new_n22291, n22124);
or_5   g19946(new_n21668, new_n21666, new_n22295);
nor_5  g19947(new_n22295, new_n17893, new_n22296);
nor_5  g19948(new_n21674_1, new_n21670, new_n22297);
nor_5  g19949(new_n22297, new_n22296, n22126);
nor_5  g19950(new_n22201_1, new_n22197, new_n22299);
xnor_4 g19951(new_n22299, new_n22199, n22130);
xor_4  g19952(new_n16528, new_n16527_1, n22144);
xnor_4 g19953(new_n21426, new_n21422, n22150);
xnor_4 g19954(new_n18207, new_n18201, n22157);
xnor_4 g19955(new_n21993_1, new_n21990, n22213);
xnor_4 g19956(new_n9471, new_n9470, n22283);
xor_4  g19957(new_n18840, new_n18839, n22311);
xnor_4 g19958(new_n8100, new_n8053, n22317);
xnor_4 g19959(new_n16131, new_n16118, n22341);
not_10 g19960(new_n6519, new_n22309_1);
nor_5  g19961(new_n22309_1, new_n6508, new_n22310);
and_5  g19962(new_n22310, new_n6504, new_n22311_1);
nand_5 g19963(new_n22309_1, new_n6508, new_n22312);
nor_5  g19964(new_n22312, new_n6504, new_n22313);
nor_5  g19965(new_n22313, new_n22311_1, new_n22314);
xnor_4 g19966(new_n22314, new_n16800, n22353);
xnor_4 g19967(new_n16129, new_n16121, n22444);
xor_4  g19968(new_n9248, new_n9247, n22467);
xor_4  g19969(new_n8080, new_n8079, n22484);
xnor_4 g19970(new_n4262, new_n4209, n22489);
xnor_4 g19971(new_n7632, new_n7583, n22494);
xnor_4 g19972(new_n9477, new_n9454, n22533);
xnor_4 g19973(new_n21009, new_n21008_1, n22584);
or_5   g19974(new_n16534, new_n16512, new_n22323);
and_5  g19975(new_n22323, new_n16477, n22589);
xnor_4 g19976(new_n22035, new_n22032, n22620);
xnor_4 g19977(new_n7700, new_n7699, n22623);
xnor_4 g19978(new_n15658, new_n15645, n22697);
xnor_4 g19979(new_n8090, new_n8073, n22714);
xnor_4 g19980(new_n10874_1, new_n10822, n22761);
xnor_4 g19981(new_n17579, new_n17563, n22779);
xnor_4 g19982(new_n21019, new_n20989, n22787);
xnor_4 g19983(new_n2519, new_n2490, n22819);
xor_4  g19984(new_n8392, new_n4243, n22858);
xor_4  g19985(new_n19690, new_n10582, new_n22334);
xnor_4 g19986(new_n22334, new_n21486, n22870);
xor_4  g19987(new_n8822, new_n8805, n22891);
xor_4  g19988(new_n18160, new_n18148, n22897);
xnor_4 g19989(new_n9266, new_n9212, n22903);
xnor_4 g19990(new_n13173, new_n13127, n22907);
xnor_4 g19991(new_n6490, new_n6489, n22910);
xnor_4 g19992(new_n11301, new_n11294, n22914);
xor_4  g19993(new_n5310, new_n5281, n22939);
xnor_4 g19994(new_n17685, new_n4106, new_n22343);
xnor_4 g19995(new_n22343, new_n17683, n22998);
xnor_4 g19996(new_n8086, new_n8085, n23006);
xnor_4 g19997(new_n11692, new_n11682_1, n23007);
xnor_4 g19998(new_n16712, new_n16709, n23009);
xnor_4 g19999(new_n15520, new_n15468, n23014);
xor_4  g20000(new_n22260, new_n22257, n23047);
xnor_4 g20001(new_n16195, new_n16184, n23058);
nor_5  g20002(new_n17156, new_n17151, n23066);
or_5   g20003(new_n17051, new_n22105, new_n22352);
and_5  g20004(new_n22352, new_n17053, new_n22353_1);
xnor_4 g20005(new_n22353_1, new_n17048, n23067);
xor_4  g20006(new_n14766, new_n14761, n23238);
xnor_4 g20007(new_n15956_1, new_n15942, n23247);
xor_4  g20008(new_n13810, new_n13802, n23248);
xnor_4 g20009(new_n16031, new_n16019, n23270);
xnor_4 g20010(new_n21076, new_n21073, n23289);
xnor_4 g20011(new_n5020_1, new_n4980, n23305);
xnor_4 g20012(new_n19427, new_n19424_1, n23341);
xor_4  g20013(new_n8539, new_n4561, n23342);
not_10 g20014(new_n19732, new_n22363);
nor_5  g20015(new_n22363, new_n6859, new_n22364);
nor_5  g20016(new_n19756_1, new_n22364, new_n22365);
and_5  g20017(new_n22363, new_n6859, new_n22366);
nor_5  g20018(new_n19755, new_n22366, new_n22367);
nor_5  g20019(new_n22367, new_n22365, n23355);
xnor_4 g20020(new_n17777, new_n17774, n23371);
xnor_4 g20021(new_n14146, new_n14111, n23401);
xnor_4 g20022(new_n12017, new_n12016, n23414);
xnor_4 g20023(new_n16036, new_n16013_1, n23429);
nor_5  g20024(new_n19976, new_n19969, new_n22373);
or_5   g20025(new_n19971, new_n19970, new_n22374);
nor_5  g20026(new_n22374, new_n19969, new_n22375);
nor_5  g20027(new_n22375, new_n19975, new_n22376);
nor_5  g20028(new_n22376, new_n22373, n23433);
xnor_4 g20029(new_n16984, new_n16971_1, n23434);
nor_5  g20030(new_n22295, new_n20102, new_n22379_1);
nor_5  g20031(new_n22379_1, new_n21687_1, new_n22380);
nor_5  g20032(new_n21669, new_n20101, new_n22381);
nor_5  g20033(new_n22381, new_n21686, new_n22382);
nor_5  g20034(new_n22382, new_n22380, n23450);
xnor_4 g20035(new_n15518, new_n15472, n23471);
xnor_4 g20036(new_n19437, new_n19405, n23480);
xor_4  g20037(new_n16389, new_n16384, n23546);
xnor_4 g20038(new_n19067, new_n19059, n23550);
xnor_4 g20039(new_n6730, new_n6707_1, n23585);
xor_4  g20040(new_n18158, new_n18151_1, n23588);
xor_4  g20041(new_n19309, new_n19308, n23619);
xnor_4 g20042(new_n2953, new_n2943, n23624);
xnor_4 g20043(new_n10751, new_n10744, n23628);
xnor_4 g20044(new_n20230, new_n20216, n23637);
xnor_4 g20045(new_n20808, new_n20805, n23663);
xnor_4 g20046(new_n10753, new_n10741, n23669);
xnor_4 g20047(new_n11919, new_n11893, n23684);
xnor_4 g20048(new_n17496, new_n17488, n23690);
xnor_4 g20049(new_n20560, new_n20529, n23714);
nor_5  g20050(new_n21722, new_n21719_1, n23719);
xnor_4 g20051(new_n19705, new_n19702, n23748);
xnor_4 g20052(new_n9882, new_n6522, n23856);
xnor_4 g20053(new_n6728, new_n6727, n23883);
xnor_4 g20054(new_n13153, new_n5341, new_n22403);
xnor_4 g20055(new_n22403, new_n13155, n23888);
xnor_4 g20056(new_n3229, new_n3206, n23899);
xor_4  g20057(new_n13626_1, new_n8620_1, n23903);
xnor_4 g20058(new_n11670, new_n11643, n23924);
xnor_4 g20059(new_n15214, new_n15213, n23935);
xnor_4 g20060(new_n11915, new_n11901, n23942);
xnor_4 g20061(new_n16228, new_n16220, n23954);
xnor_4 g20062(new_n17231, new_n17209, n23958);
xor_4  g20063(new_n20691_1, new_n20690, n23986);
xor_4  g20064(new_n15553, new_n15548, n24002);
xnor_4 g20065(new_n11814, new_n11807, n24039);
xnor_4 g20066(new_n21654_1, new_n21653, n24052);
xnor_4 g20067(new_n18772, new_n18756, n24092);
xnor_4 g20068(new_n14267_1, new_n14266, n24096);
xnor_4 g20069(new_n11072, new_n11044_1, n24097);
xnor_4 g20070(new_n10757, new_n10735, n24105);
xnor_4 g20071(new_n16692, new_n16673, n24119);
xnor_4 g20072(new_n13694, new_n13676, n24133);
xnor_4 g20073(new_n18373, new_n18342, n24141);
xnor_4 g20074(new_n19599, new_n19574, new_n22423);
xnor_4 g20075(new_n22423, new_n19636, n24145);
xnor_4 g20076(new_n20300, new_n20297, n24146);
xnor_4 g20077(new_n11608, new_n11562, n24155);
xnor_4 g20078(new_n21897, new_n21894, n24160);
xnor_4 g20079(new_n8406, new_n8373, n24167);
nor_5  g20080(new_n18897, new_n18892, n24172);
xnor_4 g20081(new_n13161, new_n13149, n24177);
xor_4  g20082(new_n21759, new_n21758, n24228);
xnor_4 g20083(new_n16133, new_n16115, n24258);
nor_5  g20084(new_n16800, new_n6508, new_n22433_1);
or_5   g20085(new_n22312, new_n6504, new_n22434);
nor_5  g20086(new_n22434, new_n16800, new_n22435);
nor_5  g20087(new_n22435, new_n22311_1, new_n22436);
nor_5  g20088(new_n22436, new_n22433_1, n24260);
xnor_4 g20089(new_n17583_1, new_n17556, n24289);
xnor_4 g20090(new_n4395, new_n4385, n24297);
xor_4  g20091(new_n10749, new_n3678, n24307);
xnor_4 g20092(new_n2513_1, new_n2503, n24342);
xnor_4 g20093(new_n14774, new_n14756, n24345);
xnor_4 g20094(new_n8628, new_n8618, n24347);
xnor_4 g20095(new_n4644, new_n4599, n24373);
xor_4  g20096(new_n16632, new_n16631, n24406);
xnor_4 g20097(new_n12553, new_n12543, n24415);
xnor_4 g20098(new_n9795, new_n9794, n24421);
xnor_4 g20099(new_n12397_1, new_n12373, n24431);
xnor_4 g20100(new_n10864, new_n10840, n24472);
or_5   g20101(new_n21083, new_n20618, new_n22450);
and_5  g20102(new_n22450, new_n21085, new_n22451);
xnor_4 g20103(new_n22451, new_n21080, n24476);
xnor_4 g20104(new_n9260, new_n9224, n24483);
xor_4  g20105(new_n12297, new_n12296, n24501);
xnor_4 g20106(new_n16735, new_n16732, n24512);
xnor_4 g20107(new_n4398, new_n4397, n24558);
xor_4  g20108(new_n2747, new_n2746, n24576);
xnor_4 g20109(new_n2749, new_n2748, n24579);
xnor_4 g20110(new_n18844, new_n18833, n24602);
xnor_4 g20111(new_n13039, new_n13011, n24604);
xnor_4 g20112(new_n21198, new_n21195, n24626);
xnor_4 g20113(new_n20310, new_n20308, n24629);
xnor_4 g20114(new_n20076, new_n20065, n24636);
xnor_4 g20115(new_n19827, new_n19824, n24715);
xnor_4 g20116(new_n18784, new_n18736, n24723);
xnor_4 g20117(new_n15459, new_n15420, new_n22466);
xnor_4 g20118(new_n22466, new_n15524, n24749);
xnor_4 g20119(new_n18774, new_n18753, n24758);
xnor_4 g20120(new_n21270, new_n21267, n24784);
xnor_4 g20121(new_n14917, new_n14916, n24807);
xor_4  g20122(new_n8848, new_n7179, n24826);
xnor_4 g20123(new_n6914, new_n6876, n24840);
xnor_4 g20124(new_n9078, new_n9068, n24841);
xnor_4 g20125(new_n4811, new_n4801, n24853);
xnor_4 g20126(new_n2957, new_n2933, n24857);
xnor_4 g20127(new_n5822_1, new_n5810, n24887);
xor_4  g20128(new_n8396, new_n8388, n24934);
xnor_4 g20129(new_n6740, new_n6687, n24998);
xnor_4 g20130(new_n10557, new_n10545, n25006);
xnor_4 g20131(new_n19129, new_n19117, n25032);
xnor_4 g20132(new_n14871, new_n14853, n25062);
xnor_4 g20133(new_n17976_1, new_n15420, new_n22482);
xnor_4 g20134(new_n22482, new_n18029, n25083);
xor_4  g20135(new_n11911, new_n11908, n25097);
xnor_4 g20136(new_n16382, new_n16379_1, n25133);
xnor_4 g20137(new_n16986, new_n16968_1, n25155);
xnor_4 g20138(new_n22195, new_n21070, new_n22487);
xnor_4 g20139(new_n22487, new_n22192, n25181);
xnor_4 g20140(new_n19131, new_n19114, n25200);
or_5   g20141(new_n19842, new_n19839, new_n22490);
xnor_4 g20142(new_n19836, new_n22021, new_n22491);
xnor_4 g20143(new_n22491, new_n22490, n25209);
xnor_4 g20144(new_n13875, new_n13874, n25215);
xor_4  g20145(new_n16805, new_n16802, n25244);
xnor_4 g20146(new_n16460_1, new_n16444, n25254);
xor_4  g20147(new_n19314_1, new_n19286, n25256);
and_5  g20148(new_n21613, new_n19916_1, new_n22497);
nor_5  g20149(new_n22497, new_n21621, new_n22498);
xnor_4 g20150(new_n21622, new_n20700_1, new_n22499);
xnor_4 g20151(new_n22499, new_n22498, n25293);
xor_4  g20152(new_n19304, new_n19297, n25328);
xor_4  g20153(new_n10064, new_n3996, n25332);
and_5  g20154(new_n21255, new_n19986, new_n22503);
nor_5  g20155(new_n21278, new_n22503, new_n22504);
nor_5  g20156(new_n21255, new_n19986, new_n22505);
nor_5  g20157(new_n21277, new_n22505, new_n22506);
nor_5  g20158(new_n22506, new_n22504, n25337);
xnor_4 g20159(new_n10391, new_n9868, new_n22508);
xnor_4 g20160(new_n22508, new_n10396, n25356);
xnor_4 g20161(new_n8237, new_n8227, n25362);
xnor_4 g20162(new_n13275, new_n13257, n25412);
xor_4  g20163(new_n14134, new_n14133, n25460);
xnor_4 g20164(new_n6732, new_n6703, n25468);
xnor_4 g20165(new_n13277, new_n13253, n25499);
xnor_4 g20166(new_n18363, new_n18361, n25513);
xnor_4 g20167(new_n11070, new_n11047, n25518);
xnor_4 g20168(new_n12227, new_n12193, n25532);
xnor_4 g20169(new_n18687, new_n18670, n25539);
xnor_4 g20170(new_n15656, new_n15648, n25550);
xnor_4 g20171(new_n19431, new_n19417, n25611);
xor_4  g20172(new_n5004, new_n5001, new_n22521);
xnor_4 g20173(new_n22521, new_n5008, n25614);
xnor_4 g20174(new_n11668, new_n11646, n25619);
and_5  g20175(new_n21506, new_n21372, new_n22524);
nor_5  g20176(new_n21511, new_n22524, new_n22525);
nor_5  g20177(new_n21506, new_n21372, new_n22526);
nor_5  g20178(new_n21510, new_n22526, new_n22527);
nor_5  g20179(new_n22527, new_n22525, n25665);
xnor_4 g20180(new_n8402, new_n8379, n25706);
xnor_4 g20181(new_n21506, new_n18066, new_n22530);
xnor_4 g20182(new_n22530, new_n22157_1, n25719);
xor_4  g20183(new_n8830, new_n8788, n25756);
not_10 g20184(new_n11841_1, new_n22533_1);
nor_5  g20185(new_n11884, new_n22533_1, new_n22534);
nor_5  g20186(new_n11923, new_n22534, new_n22535);
and_5  g20187(new_n11884, new_n22533_1, new_n22536);
nor_5  g20188(new_n11922, new_n22536, new_n22537);
nor_5  g20189(new_n22537, new_n22535, n25758);
xor_4  g20190(new_n13626_1, new_n5312, n25773);
xnor_4 g20191(new_n19223_1, new_n16352, n25784);
xnor_4 g20192(new_n7623, new_n7599, n25792);
xnor_4 g20193(new_n6300, new_n6272, n25816);
xnor_4 g20194(new_n5828, new_n5797, n25826);
xor_4  g20195(new_n11267, new_n11266_1, n25839);
xnor_4 g20196(new_n12886, new_n12846, n25840);
xnor_4 g20197(new_n7447, new_n7420, n25873);
xor_4  g20198(new_n22253_1, new_n22250, n25934);
xnor_4 g20199(new_n19628, new_n19615, n25938);
xnor_4 g20200(new_n19934, new_n19931, n25985);
xor_4  g20201(new_n12709, new_n8229, n25994);
nor_5  g20202(new_n16941, new_n16860, new_n22551);
nor_5  g20203(new_n16998, new_n16942, new_n22552);
or_5   g20204(new_n22552, new_n22551, n26084);
xnor_4 g20205(new_n21274, new_n21261, n26096);
or_5   g20206(new_n10575, new_n21493, new_n22555);
nor_5  g20207(new_n22555, new_n10494, n26111);
xnor_4 g20208(new_n10562, new_n10539, n26113);
xor_4  g20209(new_n18794, new_n18791, n26156);
xnor_4 g20210(new_n15835, new_n15815_1, n26159);
xnor_4 g20211(new_n3512, new_n3471, n26179);
xor_4  g20212(new_n12871_1, new_n12870_1, n26220);
xnor_4 g20213(new_n21312, new_n21309, n26229);
xnor_4 g20214(new_n11602, new_n11574, n26237);
xnor_4 g20215(new_n14522, new_n14508, n26250);
xor_4  g20216(new_n19668, new_n19665, n26274);
xnor_4 g20217(new_n14526, new_n14499, n26287);
xnor_4 g20218(new_n19857, new_n19138, new_n22567);
xnor_4 g20219(new_n22567, new_n22075, n26317);
nor_5  g20220(new_n21824, new_n17249, new_n22569);
nor_5  g20221(new_n22569, new_n17266, new_n22570);
nor_5  g20222(new_n17270, new_n17247, new_n22571);
nor_5  g20223(new_n22571, new_n17265, new_n22572);
nor_5  g20224(new_n22572, new_n22570, n26353);
xnor_4 g20225(new_n18842, new_n18835, n26375);
nor_5  g20226(new_n21646, new_n19972, new_n22575);
nor_5  g20227(new_n21656, new_n21647, new_n22576);
nor_5  g20228(new_n22576, new_n22575, n26396);
xor_4  g20229(new_n5007, new_n5006, n26429);
xnor_4 g20230(new_n13345, new_n13331, n26431);
xnor_4 g20231(new_n6502_1, new_n6448, n26439);
xnor_4 g20232(new_n19065, new_n19064, n26492);
xnor_4 g20233(new_n9253, new_n9252, n26515);
xnor_4 g20234(new_n2517, new_n2494, n26538);
xnor_4 g20235(new_n13812, new_n13798_1, n26590);
xor_4  g20236(new_n18008, new_n15503, n26598);
xnor_4 g20237(new_n21622, new_n19916_1, new_n22586);
xnor_4 g20238(new_n22586, new_n21617, n26605);
xor_4  g20239(new_n21590, new_n21584, new_n22588_1);
xnor_4 g20240(new_n22588_1, new_n21587, n26656);
xnor_4 g20241(new_n10552, new_n10551, n26674);
xnor_4 g20242(new_n8707, new_n8693, n26675);
xnor_4 g20243(new_n19075, new_n19046, n26681);
nor_5  g20244(new_n5242, new_n5070, new_n22593);
nor_5  g20245(new_n5308, new_n22593, new_n22594);
and_5  g20246(new_n5242, new_n5070, new_n22595);
nor_5  g20247(new_n5307, new_n22595, new_n22596);
nor_5  g20248(new_n22596, new_n22594, n26696);
xnor_4 g20249(new_n13586, new_n13568, n26698);
xor_4  g20250(new_n14260, new_n5334, n26707);
xor_4  g20251(new_n22015, new_n22014, n26719);
xnor_4 g20252(new_n8398, new_n8385, n26727);
nor_5  g20253(new_n19986, new_n17855_1, new_n22602);
nor_5  g20254(new_n19990, new_n19987, new_n22603);
nor_5  g20255(new_n22603, new_n22602, n26729);
xor_4  g20256(new_n20011, new_n20008, n26745);
xnor_4 g20257(new_n7192, new_n7162, n26775);
xnor_4 g20258(new_n9570, new_n9553, n26780);
xor_4  g20259(new_n20413, new_n20406, n26794);
xnor_4 g20260(new_n3237, new_n3190, n26795);
xnor_4 g20261(new_n9810, new_n9772, n26801);
xnor_4 g20262(new_n10145, new_n10127, n26815);
xnor_4 g20263(new_n21708, new_n21705, n26847);
xnor_4 g20264(new_n17270, new_n6682, new_n22613);
xnor_4 g20265(new_n22613, new_n21829, n26900);
xor_4  g20266(new_n17411, new_n17410, n26902);
xor_4  g20267(new_n16074, new_n16071, n26905);
xnor_4 g20268(new_n7449, new_n7416, n26921);
xnor_4 g20269(new_n20756, new_n20742, n26923);
xnor_4 g20270(new_n9884, new_n9883, n26929);
xnor_4 g20271(new_n11612, new_n11554, n26930);
xnor_4 g20272(new_n14524, new_n14504, n26943);
xnor_4 g20273(new_n13279, new_n13250, n26970);
xnor_4 g20274(new_n19567, new_n19555, n27004);
xnor_4 g20275(new_n9489, new_n9436, n27011);
xnor_4 g20276(new_n18027, new_n17979, n27019);
xnor_4 g20277(new_n4634, new_n4623, n27031);
xnor_4 g20278(new_n20458, new_n19664_1, new_n22627);
xnor_4 g20279(new_n22627, new_n22228, n27051);
xor_4  g20280(new_n15950, new_n15947_1, n27072);
xnor_4 g20281(new_n14150, new_n14103, n27079);
xor_4  g20282(new_n3997, new_n3996, n27096);
xor_4  g20283(new_n13032, new_n13022, n27110);
xnor_4 g20284(new_n12497, new_n12494, n27112);
xnor_4 g20285(new_n20762, new_n20310, n27130);
xnor_4 g20286(new_n14867, new_n14859, n27145);
and_5  g20287(new_n15302, new_n14733, new_n22636);
nor_5  g20288(new_n20160, new_n20157, new_n22637);
nor_5  g20289(new_n22637, new_n22636, n27158);
xnor_4 g20290(new_n19779, new_n19775, n27163);
xnor_4 g20291(new_n21852, new_n19574, new_n22640);
xnor_4 g20292(new_n22640, new_n21857, n27194);
endmodule


