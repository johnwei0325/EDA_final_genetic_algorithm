// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Thu Jun 27 03:55:57 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533_1, new_n2534,
    new_n2535_1, new_n2536, new_n2537_1, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547_1, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553_1, new_n2554, new_n2555_1, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560_1, new_n2561_1, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2568, new_n2569, new_n2570_1, new_n2571,
    new_n2572, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578_1,
    new_n2579, new_n2580, new_n2581, new_n2582_1, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602_1, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619_1, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826_1, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886_1, new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945, new_n2946,
    new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971_1, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978_1, new_n2979_1, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985_1, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1,
    new_n3019, new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067_1, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076_1, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3163,
    new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235_1,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253_1,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260_1, new_n3261, new_n3262, new_n3263_1, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279_1, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289_1,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301_1,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306_1, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319,
    new_n3320_1, new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332_1, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445,
    new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1,
    new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457,
    new_n3458, new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463,
    new_n3464, new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469,
    new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481,
    new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487,
    new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499,
    new_n3500, new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505,
    new_n3506_1, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511,
    new_n3512, new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3517,
    new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523,
    new_n3524, new_n3525, new_n3526, new_n3527, new_n3528_1, new_n3529,
    new_n3530, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541_1, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555_1, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561_1, new_n3562, new_n3563_1, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570_1, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582_1, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617_1, new_n3618_1, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642_1, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649_1, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665_1, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679_1, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710_1,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725_1, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733_1, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740_1,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755_1, new_n3756, new_n3757, new_n3758_1,
    new_n3759, new_n3760_1, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781_1, new_n3782,
    new_n3783, new_n3784, new_n3785_1, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794_1,
    new_n3795_1, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828_1, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850_1, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866,
    new_n3867, new_n3868, new_n3869_1, new_n3870, new_n3871_1, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891_1,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909_1,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918_1, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925_1, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934_1, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945_1,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952_1, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959_1, new_n3960, new_n3961, new_n3962_1, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971_1, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983_1, new_n3984_1, new_n3985, new_n3986, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000_1, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010_1, new_n4011,
    new_n4012, new_n4013, new_n4014_1, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071_1,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085_1, new_n4086, new_n4087, new_n4088_1, new_n4089_1,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100_1, new_n4101, new_n4102,
    new_n4103_1, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119_1, new_n4120,
    new_n4121, new_n4122, new_n4123_1, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134_1, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146_1, new_n4147, new_n4148, new_n4149, new_n4150_1,
    new_n4151_1, new_n4152_1, new_n4153_1, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165_1, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172_1, new_n4173_1, new_n4174,
    new_n4175, new_n4176_1, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186_1,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204_1,
    new_n4205_1, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215_1, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221_1, new_n4222,
    new_n4223, new_n4224_1, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231_1, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256_1, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266_1, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272_1, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306_1, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319_1,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325_1,
    new_n4326_1, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340_1, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374_1,
    new_n4375, new_n4376_1, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401_1, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409_1, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424_1, new_n4425, new_n4426_1, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432_1, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441_1, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451_1, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476_1,
    new_n4477, new_n4478_1, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4501,
    new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507,
    new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513,
    new_n4514_1, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519,
    new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525,
    new_n4526, new_n4527, new_n4528, new_n4529_1, new_n4530, new_n4531,
    new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537,
    new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543,
    new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549,
    new_n4550, new_n4551, new_n4552_1, new_n4553, new_n4554, new_n4555,
    new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561,
    new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567,
    new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573,
    new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588_1, new_n4589, new_n4590_1, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595_1, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615,
    new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621,
    new_n4622, new_n4623, new_n4624_1, new_n4625, new_n4626, new_n4627,
    new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633,
    new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639,
    new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645,
    new_n4646_1, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651,
    new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657,
    new_n4658, new_n4659, new_n4660, new_n4661, new_n4662, new_n4663,
    new_n4664, new_n4665_1, new_n4666, new_n4667, new_n4668, new_n4669,
    new_n4670, new_n4671, new_n4672, new_n4673, new_n4674_1, new_n4675,
    new_n4676, new_n4677, new_n4678, new_n4679, new_n4680, new_n4681,
    new_n4682, new_n4683, new_n4684, new_n4685, new_n4686, new_n4687,
    new_n4688, new_n4689, new_n4690, new_n4691, new_n4692, new_n4693_1,
    new_n4694, new_n4695, new_n4696, new_n4697, new_n4698, new_n4699,
    new_n4700, new_n4701, new_n4702, new_n4703, new_n4704, new_n4705,
    new_n4706, new_n4707, new_n4708, new_n4709, new_n4710, new_n4711,
    new_n4712, new_n4713, new_n4714, new_n4715, new_n4716, new_n4717,
    new_n4718, new_n4719, new_n4720, new_n4721, new_n4722_1, new_n4723,
    new_n4724, new_n4725, new_n4726, new_n4727, new_n4728, new_n4729,
    new_n4730, new_n4731_1, new_n4732, new_n4733, new_n4734, new_n4735,
    new_n4736, new_n4737, new_n4738, new_n4739, new_n4740, new_n4741,
    new_n4742, new_n4743, new_n4744, new_n4745_1, new_n4746, new_n4747_1,
    new_n4748, new_n4749, new_n4750, new_n4751, new_n4752, new_n4753,
    new_n4754, new_n4755, new_n4756, new_n4757, new_n4758, new_n4759,
    new_n4760, new_n4761, new_n4762, new_n4763, new_n4764, new_n4765,
    new_n4766_1, new_n4767, new_n4768, new_n4769, new_n4770_1, new_n4771,
    new_n4772, new_n4773, new_n4774, new_n4775, new_n4776, new_n4777_1,
    new_n4778, new_n4779, new_n4780, new_n4781, new_n4782, new_n4783,
    new_n4784, new_n4785_1, new_n4786, new_n4787, new_n4788, new_n4789,
    new_n4790, new_n4791, new_n4792, new_n4793, new_n4794, new_n4795,
    new_n4796, new_n4797, new_n4798, new_n4799, new_n4800, new_n4801,
    new_n4802, new_n4803, new_n4804_1, new_n4805, new_n4806, new_n4807,
    new_n4808, new_n4809, new_n4810_1, new_n4811, new_n4812_1, new_n4813,
    new_n4814_1, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819,
    new_n4821, new_n4822, new_n4823, new_n4824, new_n4825, new_n4826,
    new_n4827, new_n4828, new_n4829, new_n4830, new_n4831, new_n4832,
    new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838,
    new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850_1,
    new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858_1, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891_1, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913_1, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925_1, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938, new_n4939_1, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947_1, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952_1,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957_1, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964_1,
    new_n4965, new_n4966_1, new_n4967_1, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972_1, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011_1, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020_1, new_n5021, new_n5022, new_n5023, new_n5024_1, new_n5025_1,
    new_n5026_1, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031_1,
    new_n5032, new_n5033, new_n5034, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046_1, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060_1, new_n5061,
    new_n5062_1, new_n5063, new_n5064_1, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077_1, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082_1, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094, new_n5095, new_n5096, new_n5097,
    new_n5098_1, new_n5099, new_n5100, new_n5101_1, new_n5102, new_n5103,
    new_n5104, new_n5105, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115_1,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120_1, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128_1, new_n5129, new_n5130, new_n5131_1, new_n5132, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140_1, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158_1, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168_1, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184_1, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211_1,
    new_n5212, new_n5213_1, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226_1, new_n5227, new_n5228_1, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255_1, new_n5256_1, new_n5257, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265_1,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273_1, new_n5274_1, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300_1, new_n5301, new_n5302_1,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325_1, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330_1, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337_1, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351_1, new_n5352, new_n5353_1, new_n5354, new_n5356, new_n5357,
    new_n5358, new_n5359, new_n5360, new_n5361, new_n5362, new_n5363,
    new_n5364, new_n5365, new_n5366, new_n5367, new_n5368, new_n5369,
    new_n5370, new_n5371, new_n5372, new_n5373, new_n5374, new_n5375,
    new_n5376_1, new_n5377, new_n5378, new_n5379, new_n5380, new_n5381,
    new_n5382, new_n5383, new_n5384, new_n5385, new_n5386_1, new_n5387,
    new_n5388, new_n5389, new_n5390, new_n5391, new_n5392, new_n5393,
    new_n5394, new_n5395, new_n5396, new_n5397, new_n5398, new_n5399_1,
    new_n5400_1, new_n5401, new_n5402, new_n5403_1, new_n5404, new_n5405,
    new_n5406, new_n5407, new_n5408, new_n5409, new_n5410, new_n5411,
    new_n5412, new_n5413, new_n5414, new_n5415, new_n5416, new_n5417,
    new_n5418, new_n5419, new_n5420, new_n5421, new_n5422, new_n5423,
    new_n5424, new_n5425, new_n5426, new_n5427, new_n5428, new_n5429,
    new_n5430_1, new_n5431, new_n5432, new_n5433, new_n5434, new_n5435,
    new_n5436, new_n5437, new_n5438_1, new_n5439_1, new_n5440, new_n5441,
    new_n5442, new_n5443_1, new_n5444, new_n5445, new_n5446, new_n5447,
    new_n5448, new_n5449, new_n5450, new_n5451_1, new_n5452, new_n5453,
    new_n5454, new_n5455, new_n5456, new_n5457, new_n5458, new_n5459,
    new_n5460, new_n5461, new_n5462, new_n5463, new_n5464, new_n5465,
    new_n5466, new_n5467, new_n5468, new_n5469, new_n5470, new_n5471,
    new_n5472_1, new_n5473, new_n5474, new_n5475, new_n5476, new_n5477,
    new_n5478, new_n5479, new_n5480, new_n5481, new_n5482, new_n5483,
    new_n5484, new_n5485_1, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517_1, new_n5518, new_n5519, new_n5520,
    new_n5521_1, new_n5522, new_n5523, new_n5524_1, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532_1,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564_1, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579_1, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593_1, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603_1, new_n5604,
    new_n5605_1, new_n5606, new_n5607, new_n5608, new_n5609_1, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634_1,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643_1, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680_1, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687_1, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696_1, new_n5697, new_n5698, new_n5699, new_n5700_1,
    new_n5701, new_n5702, new_n5703, new_n5704_1, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732_1, new_n5733, new_n5734, new_n5735, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742_1, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752_1, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765_1, new_n5766, new_n5767,
    new_n5768, new_n5769, new_n5770, new_n5771, new_n5772, new_n5773,
    new_n5774, new_n5775, new_n5776_1, new_n5777, new_n5778, new_n5779,
    new_n5780, new_n5781, new_n5782_1, new_n5783, new_n5784, new_n5785,
    new_n5786, new_n5787, new_n5788, new_n5789, new_n5790, new_n5791,
    new_n5792, new_n5793, new_n5794, new_n5795, new_n5796, new_n5797,
    new_n5798, new_n5799, new_n5800, new_n5801, new_n5802, new_n5803,
    new_n5804, new_n5805, new_n5806, new_n5807, new_n5808, new_n5809,
    new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815,
    new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821,
    new_n5822_1, new_n5823, new_n5824, new_n5825, new_n5826, new_n5827,
    new_n5828, new_n5829, new_n5830, new_n5831, new_n5832, new_n5833_1,
    new_n5834_1, new_n5835, new_n5836, new_n5837, new_n5838, new_n5839,
    new_n5840_1, new_n5841_1, new_n5842_1, new_n5843, new_n5844, new_n5845,
    new_n5846, new_n5847, new_n5848, new_n5849, new_n5850_1, new_n5851,
    new_n5852, new_n5853, new_n5854, new_n5855, new_n5856, new_n5857,
    new_n5858, new_n5859, new_n5860, new_n5861, new_n5862, new_n5863,
    new_n5864, new_n5865, new_n5866, new_n5867, new_n5868, new_n5869,
    new_n5870, new_n5871, new_n5872, new_n5873, new_n5874, new_n5875,
    new_n5876, new_n5877, new_n5878, new_n5879, new_n5880, new_n5881,
    new_n5882_1, new_n5883, new_n5884, new_n5885, new_n5886, new_n5887,
    new_n5888, new_n5889, new_n5890, new_n5891, new_n5892, new_n5893,
    new_n5894, new_n5895, new_n5896, new_n5897, new_n5898, new_n5899,
    new_n5900, new_n5901, new_n5902, new_n5903_1, new_n5904_1, new_n5905,
    new_n5906, new_n5907, new_n5908, new_n5909, new_n5910, new_n5911_1,
    new_n5912, new_n5913, new_n5914, new_n5915, new_n5916, new_n5917,
    new_n5918, new_n5919, new_n5920, new_n5921, new_n5922, new_n5923,
    new_n5924, new_n5925, new_n5926, new_n5927, new_n5928, new_n5929,
    new_n5930, new_n5931, new_n5932, new_n5933, new_n5934, new_n5935,
    new_n5936_1, new_n5937, new_n5938, new_n5939, new_n5940, new_n5941,
    new_n5942, new_n5943_1, new_n5944, new_n5945, new_n5946, new_n5947,
    new_n5948, new_n5949, new_n5950, new_n5951, new_n5952, new_n5953,
    new_n5954, new_n5955, new_n5956, new_n5957, new_n5958, new_n5959,
    new_n5960, new_n5961, new_n5962, new_n5963, new_n5964_1, new_n5965,
    new_n5966, new_n5967, new_n5968, new_n5969, new_n5970, new_n5971,
    new_n5972, new_n5973, new_n5974, new_n5975, new_n5976, new_n5977,
    new_n5978, new_n5979, new_n5980_1, new_n5981, new_n5982, new_n5983,
    new_n5984, new_n5985, new_n5986, new_n5987, new_n5988, new_n5989,
    new_n5990, new_n5991, new_n5992, new_n5993, new_n5994, new_n5995,
    new_n5996, new_n5997, new_n5998, new_n5999, new_n6000, new_n6001,
    new_n6002, new_n6003, new_n6004, new_n6005, new_n6006, new_n6007,
    new_n6008, new_n6009, new_n6010, new_n6011, new_n6012_1, new_n6013,
    new_n6014, new_n6015, new_n6016, new_n6017, new_n6018, new_n6019,
    new_n6020, new_n6021, new_n6022_1, new_n6023, new_n6024, new_n6025,
    new_n6026, new_n6027, new_n6028, new_n6029, new_n6030, new_n6031_1,
    new_n6032, new_n6033, new_n6034, new_n6035, new_n6036, new_n6037,
    new_n6038, new_n6039, new_n6040, new_n6041, new_n6042, new_n6043,
    new_n6044_1, new_n6045, new_n6046_1, new_n6047, new_n6048, new_n6049,
    new_n6050, new_n6051, new_n6052, new_n6053, new_n6054, new_n6055,
    new_n6056, new_n6057, new_n6058, new_n6059, new_n6060, new_n6061,
    new_n6062, new_n6063, new_n6064, new_n6065, new_n6066, new_n6067,
    new_n6068, new_n6069, new_n6070, new_n6071, new_n6072, new_n6073,
    new_n6074, new_n6075, new_n6076, new_n6077, new_n6078, new_n6079,
    new_n6080, new_n6082, new_n6083, new_n6084_1, new_n6085, new_n6086,
    new_n6087, new_n6088, new_n6089, new_n6090, new_n6091, new_n6092,
    new_n6093, new_n6094, new_n6095, new_n6096, new_n6097, new_n6098,
    new_n6099, new_n6100, new_n6101, new_n6102, new_n6103, new_n6104_1,
    new_n6105_1, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160_1, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171_1, new_n6172, new_n6173, new_n6174,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183_1,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189_1,
    new_n6190, new_n6191, new_n6192, new_n6193, new_n6194, new_n6195,
    new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201,
    new_n6202, new_n6203, new_n6204_1, new_n6205, new_n6206, new_n6207,
    new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213,
    new_n6214, new_n6215, new_n6216, new_n6217, new_n6218_1, new_n6219,
    new_n6220, new_n6221, new_n6222, new_n6223_1, new_n6224, new_n6225,
    new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231,
    new_n6232, new_n6233_1, new_n6234, new_n6235, new_n6236, new_n6237,
    new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243,
    new_n6244, new_n6245_1, new_n6246, new_n6247, new_n6248_1, new_n6249,
    new_n6250, new_n6251, new_n6252, new_n6253, new_n6254, new_n6255,
    new_n6256_1, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261,
    new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267,
    new_n6268, new_n6269, new_n6270, new_n6271_1, new_n6272, new_n6273,
    new_n6274, new_n6275, new_n6276_1, new_n6277, new_n6278, new_n6279,
    new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285,
    new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291,
    new_n6292, new_n6293, new_n6294, new_n6295, new_n6296, new_n6297,
    new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303,
    new_n6304, new_n6305, new_n6306, new_n6307, new_n6308_1, new_n6309,
    new_n6310, new_n6311_1, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323_1, new_n6324, new_n6325, new_n6326, new_n6327,
    new_n6328, new_n6329, new_n6330_1, new_n6331, new_n6332, new_n6333,
    new_n6334, new_n6335, new_n6336, new_n6337, new_n6338, new_n6339_1,
    new_n6340, new_n6341, new_n6342, new_n6343, new_n6344, new_n6345,
    new_n6346, new_n6347, new_n6348, new_n6349, new_n6350, new_n6351,
    new_n6352, new_n6353, new_n6354_1, new_n6355, new_n6356_1, new_n6357,
    new_n6358, new_n6359, new_n6360, new_n6361, new_n6362, new_n6363,
    new_n6364, new_n6365, new_n6366, new_n6367, new_n6368, new_n6369_1,
    new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375_1,
    new_n6376, new_n6377, new_n6378, new_n6379_1, new_n6380, new_n6381_1,
    new_n6382, new_n6383_1, new_n6384, new_n6385_1, new_n6386, new_n6387,
    new_n6388, new_n6389, new_n6390, new_n6391, new_n6392, new_n6393,
    new_n6394, new_n6395, new_n6396, new_n6397_1, new_n6398, new_n6399,
    new_n6400, new_n6401, new_n6402, new_n6403, new_n6404, new_n6405,
    new_n6406, new_n6407_1, new_n6408, new_n6409, new_n6410, new_n6411,
    new_n6412, new_n6413, new_n6414, new_n6415, new_n6416, new_n6417,
    new_n6418, new_n6419, new_n6420, new_n6421, new_n6422, new_n6423,
    new_n6424, new_n6425, new_n6426, new_n6427_1, new_n6428, new_n6429,
    new_n6430, new_n6431_1, new_n6432, new_n6433, new_n6434, new_n6435,
    new_n6436, new_n6437_1, new_n6438, new_n6439, new_n6440, new_n6441,
    new_n6442, new_n6443, new_n6444, new_n6445, new_n6446, new_n6447,
    new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453,
    new_n6454, new_n6455, new_n6456_1, new_n6457_1, new_n6458, new_n6459,
    new_n6460, new_n6461, new_n6462, new_n6463, new_n6464, new_n6465_1,
    new_n6466, new_n6467, new_n6468, new_n6469, new_n6470_1, new_n6471,
    new_n6472, new_n6473, new_n6474, new_n6475, new_n6477, new_n6478,
    new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485_1, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502_1,
    new_n6503, new_n6504, new_n6505, new_n6506_1, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513_1, new_n6514_1,
    new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542_1, new_n6543, new_n6544,
    new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550,
    new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556_1,
    new_n6557, new_n6558_1, new_n6559, new_n6560_1, new_n6561, new_n6562,
    new_n6563, new_n6564, new_n6565, new_n6566, new_n6567_1, new_n6568,
    new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574,
    new_n6575, new_n6576_1, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586,
    new_n6587_1, new_n6588, new_n6589, new_n6590_1, new_n6591, new_n6592,
    new_n6593, new_n6594, new_n6595, new_n6596_1, new_n6597, new_n6598,
    new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604,
    new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6610,
    new_n6611_1, new_n6612_1, new_n6613, new_n6614, new_n6615, new_n6616,
    new_n6617, new_n6618, new_n6619, new_n6620, new_n6621, new_n6622,
    new_n6623, new_n6624, new_n6625, new_n6626, new_n6627, new_n6628_1,
    new_n6629, new_n6630_1, new_n6631_1, new_n6632, new_n6633, new_n6634_1,
    new_n6635, new_n6636, new_n6637, new_n6638, new_n6639, new_n6640,
    new_n6641, new_n6642, new_n6643, new_n6644, new_n6645, new_n6646,
    new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652_1,
    new_n6653, new_n6654, new_n6655_1, new_n6656, new_n6657, new_n6658,
    new_n6659_1, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664,
    new_n6665, new_n6666, new_n6667, new_n6668, new_n6669_1, new_n6670,
    new_n6671_1, new_n6672, new_n6673_1, new_n6674_1, new_n6675, new_n6676,
    new_n6677, new_n6678, new_n6679, new_n6680, new_n6681, new_n6682,
    new_n6683, new_n6684_1, new_n6685, new_n6686, new_n6687, new_n6688,
    new_n6689, new_n6690, new_n6691_1, new_n6692, new_n6693, new_n6694,
    new_n6695, new_n6696, new_n6697, new_n6698, new_n6699, new_n6700,
    new_n6701, new_n6702, new_n6703, new_n6704, new_n6705, new_n6706_1,
    new_n6707_1, new_n6708, new_n6709, new_n6710, new_n6711, new_n6712,
    new_n6713, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718,
    new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724,
    new_n6725, new_n6726, new_n6727, new_n6728, new_n6729_1, new_n6730,
    new_n6731, new_n6732, new_n6733, new_n6734, new_n6735, new_n6736_1,
    new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742,
    new_n6743, new_n6744, new_n6745, new_n6746, new_n6747, new_n6748,
    new_n6749, new_n6750, new_n6751, new_n6752, new_n6753, new_n6754,
    new_n6755, new_n6756, new_n6757, new_n6758, new_n6759, new_n6760,
    new_n6761, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773_1,
    new_n6774, new_n6775_1, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785_1,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790_1, new_n6791_1,
    new_n6792, new_n6793, new_n6794_1, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802_1, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814_1, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6826_1, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835_1, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853_1, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6860, new_n6861_1, new_n6862_1, new_n6863_1,
    new_n6864, new_n6865, new_n6866, new_n6867_1, new_n6868, new_n6869,
    new_n6870, new_n6871, new_n6872, new_n6873, new_n6874, new_n6875,
    new_n6876, new_n6877, new_n6878, new_n6879, new_n6880, new_n6881,
    new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887,
    new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893,
    new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899,
    new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905,
    new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911,
    new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6940, new_n6941, new_n6942,
    new_n6944, new_n6945, new_n6946, new_n6947, new_n6948, new_n6949,
    new_n6950, new_n6951, new_n6952, new_n6953, new_n6954, new_n6955,
    new_n6956, new_n6957, new_n6958, new_n6959, new_n6960, new_n6961,
    new_n6962, new_n6963, new_n6964, new_n6965_1, new_n6966, new_n6967_1,
    new_n6968, new_n6969, new_n6970, new_n6971_1, new_n6972, new_n6973,
    new_n6974, new_n6975_1, new_n6976, new_n6977, new_n6978, new_n6979,
    new_n6980, new_n6981, new_n6982, new_n6983_1, new_n6984, new_n6985_1,
    new_n6986, new_n6987, new_n6988, new_n6989, new_n6990, new_n6991,
    new_n6992, new_n6993, new_n6994, new_n6995, new_n6996, new_n6997,
    new_n6998_1, new_n6999, new_n7000, new_n7001, new_n7002, new_n7003,
    new_n7004, new_n7005, new_n7006, new_n7007, new_n7008, new_n7009,
    new_n7010, new_n7011, new_n7012, new_n7013, new_n7014, new_n7015,
    new_n7016, new_n7017, new_n7018, new_n7019, new_n7020, new_n7021,
    new_n7022, new_n7023, new_n7024, new_n7025, new_n7026_1, new_n7027,
    new_n7028, new_n7029, new_n7030, new_n7031, new_n7032_1, new_n7033,
    new_n7034, new_n7036, new_n7037, new_n7038_1, new_n7039, new_n7040,
    new_n7041, new_n7042, new_n7043, new_n7044, new_n7045, new_n7046,
    new_n7047, new_n7048, new_n7049, new_n7050, new_n7051, new_n7052,
    new_n7053, new_n7054, new_n7055, new_n7056, new_n7057_1, new_n7058,
    new_n7059, new_n7060, new_n7061, new_n7062, new_n7063, new_n7064,
    new_n7065, new_n7066, new_n7067, new_n7068, new_n7069, new_n7070,
    new_n7071, new_n7072, new_n7073, new_n7074, new_n7075, new_n7076,
    new_n7077, new_n7078, new_n7079_1, new_n7080, new_n7081, new_n7082,
    new_n7083, new_n7084, new_n7085, new_n7086, new_n7087, new_n7088,
    new_n7089, new_n7090, new_n7091, new_n7092, new_n7093, new_n7094,
    new_n7095, new_n7096, new_n7097, new_n7098, new_n7099_1, new_n7100,
    new_n7101, new_n7102, new_n7103, new_n7104, new_n7105, new_n7106,
    new_n7107, new_n7108, new_n7109, new_n7110, new_n7111, new_n7112,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139_1, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149_1,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190_1, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229_1, new_n7230_1, new_n7231, new_n7232, new_n7233_1,
    new_n7234, new_n7235, new_n7236_1, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253_1, new_n7254, new_n7255, new_n7256_1, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265, new_n7266, new_n7267, new_n7268_1, new_n7269,
    new_n7270, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277_1, new_n7278, new_n7279, new_n7280_1, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294, new_n7295, new_n7296, new_n7297, new_n7298_1, new_n7299,
    new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305_1,
    new_n7306, new_n7307, new_n7308_1, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313_1, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330_1, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335_1,
    new_n7336, new_n7337, new_n7338, new_n7339_1, new_n7340, new_n7341,
    new_n7342, new_n7343, new_n7344, new_n7345, new_n7346_1, new_n7347,
    new_n7348, new_n7349_1, new_n7350, new_n7351, new_n7352, new_n7353,
    new_n7354, new_n7355, new_n7356, new_n7358, new_n7359, new_n7360,
    new_n7361, new_n7362, new_n7363_1, new_n7364, new_n7365, new_n7366,
    new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372,
    new_n7373, new_n7374, new_n7375, new_n7376, new_n7377_1, new_n7378,
    new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384,
    new_n7385, new_n7386, new_n7387, new_n7388, new_n7389, new_n7390_1,
    new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396,
    new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402,
    new_n7403_1, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408_1,
    new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7414,
    new_n7415, new_n7416, new_n7417, new_n7418, new_n7419, new_n7420,
    new_n7421_1, new_n7422, new_n7423, new_n7424, new_n7425, new_n7426,
    new_n7427, new_n7428_1, new_n7429, new_n7430, new_n7431, new_n7432_1,
    new_n7433, new_n7434, new_n7435, new_n7436, new_n7437_1, new_n7438,
    new_n7439, new_n7440, new_n7441, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456,
    new_n7457, new_n7458, new_n7459, new_n7460_1, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475_1, new_n7476, new_n7477_1, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507_1, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514_1, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524_1, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558_1,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566_1, new_n7567, new_n7568, new_n7569_1, new_n7570,
    new_n7571, new_n7572_1, new_n7573, new_n7574, new_n7575_1, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585_1, new_n7586, new_n7587, new_n7588_1,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593_1, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598_1, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607_1, new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616_1, new_n7617, new_n7618,
    new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624,
    new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630_1,
    new_n7631, new_n7632, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7640, new_n7641, new_n7642, new_n7643_1, new_n7644,
    new_n7645, new_n7646, new_n7647_1, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657_1, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670_1, new_n7671, new_n7672, new_n7673, new_n7674_1,
    new_n7675, new_n7676, new_n7677, new_n7678_1, new_n7679_1, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686_1,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692_1,
    new_n7693_1, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698_1,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708_1, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721_1, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731_1, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751_1, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759_1, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769_1, new_n7770,
    new_n7771, new_n7772, new_n7773_1, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780_1, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788_1,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794_1,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811_1, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830_1,
    new_n7831, new_n7832, new_n7833, new_n7834_1, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841_1, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876_1, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884_1,
    new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891,
    new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897,
    new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903,
    new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909,
    new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915,
    new_n7916, new_n7917_1, new_n7918, new_n7919, new_n7920, new_n7921,
    new_n7922, new_n7923, new_n7924, new_n7925, new_n7926, new_n7927,
    new_n7928, new_n7929, new_n7930, new_n7931, new_n7932, new_n7933,
    new_n7934, new_n7935, new_n7936, new_n7937_1, new_n7938, new_n7939,
    new_n7940, new_n7941, new_n7942, new_n7943_1, new_n7944, new_n7945,
    new_n7946, new_n7947, new_n7948, new_n7949_1, new_n7950_1, new_n7951,
    new_n7952, new_n7953, new_n7954, new_n7955, new_n7956, new_n7957,
    new_n7958, new_n7959_1, new_n7960, new_n7961, new_n7962, new_n7963_1,
    new_n7964, new_n7965, new_n7966, new_n7967, new_n7968_1, new_n7969,
    new_n7970, new_n7971, new_n7972, new_n7973, new_n7974, new_n7975,
    new_n7976, new_n7977, new_n7978, new_n7979, new_n7980, new_n7981,
    new_n7982, new_n7983, new_n7984, new_n7985, new_n7986, new_n7987,
    new_n7988, new_n7989, new_n7990, new_n7991, new_n7992_1, new_n7993,
    new_n7994, new_n7995, new_n7996, new_n7997, new_n7998, new_n7999_1,
    new_n8000, new_n8001, new_n8002, new_n8003, new_n8004, new_n8005,
    new_n8006_1, new_n8007, new_n8008, new_n8009, new_n8010, new_n8011,
    new_n8012, new_n8013, new_n8014, new_n8015, new_n8016, new_n8017,
    new_n8018, new_n8019, new_n8020, new_n8021, new_n8022, new_n8023,
    new_n8024, new_n8025, new_n8026, new_n8027_1, new_n8028, new_n8029,
    new_n8030, new_n8031_1, new_n8032, new_n8033, new_n8034, new_n8035,
    new_n8036, new_n8037, new_n8038, new_n8039, new_n8040, new_n8041,
    new_n8042_1, new_n8043, new_n8044, new_n8045, new_n8046, new_n8047,
    new_n8048, new_n8049, new_n8050, new_n8051, new_n8052_1, new_n8053,
    new_n8054, new_n8055, new_n8056, new_n8057, new_n8058, new_n8059,
    new_n8060, new_n8061, new_n8062, new_n8063, new_n8064, new_n8065,
    new_n8066, new_n8067_1, new_n8068, new_n8069, new_n8070, new_n8071,
    new_n8072, new_n8073, new_n8074, new_n8075, new_n8076, new_n8077,
    new_n8078, new_n8079, new_n8080, new_n8081, new_n8082, new_n8083,
    new_n8084, new_n8085, new_n8086, new_n8087, new_n8088, new_n8089,
    new_n8090, new_n8091, new_n8093, new_n8094, new_n8095_1, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103_1, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109_1, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127_1, new_n8128, new_n8129, new_n8130_1, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135_1, new_n8136, new_n8137, new_n8138,
    new_n8139_1, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148_1, new_n8149_1, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159_1, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179_1, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194_1, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215_1, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244_1, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255_1, new_n8256_1, new_n8257, new_n8258,
    new_n8259_1, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267_1, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276_1,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285_1, new_n8286, new_n8287, new_n8288_1,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305_1, new_n8306_1,
    new_n8307, new_n8308, new_n8309_1, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320_1, new_n8321_1, new_n8322, new_n8323, new_n8324_1,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339_1, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363_1, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376_1, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381_1, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399_1, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405_1, new_n8406, new_n8407, new_n8408_1,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8416, new_n8417_1, new_n8418, new_n8419, new_n8420, new_n8421,
    new_n8422, new_n8423, new_n8424, new_n8425, new_n8426, new_n8427,
    new_n8428, new_n8429, new_n8430, new_n8431, new_n8432_1, new_n8433,
    new_n8434, new_n8435, new_n8436, new_n8437, new_n8438, new_n8439_1,
    new_n8440, new_n8441, new_n8442, new_n8443, new_n8444, new_n8445,
    new_n8446, new_n8447, new_n8448, new_n8449, new_n8450, new_n8451,
    new_n8452, new_n8453_1, new_n8454, new_n8455, new_n8456, new_n8457,
    new_n8458, new_n8459, new_n8460, new_n8461, new_n8462, new_n8463,
    new_n8464, new_n8465, new_n8466, new_n8467, new_n8468, new_n8469,
    new_n8470, new_n8471, new_n8472, new_n8473, new_n8474, new_n8475,
    new_n8476, new_n8477, new_n8478, new_n8479, new_n8480_1, new_n8481,
    new_n8482, new_n8483, new_n8484, new_n8485, new_n8486, new_n8487,
    new_n8488, new_n8489_1, new_n8490, new_n8491, new_n8492, new_n8493,
    new_n8494, new_n8495, new_n8496, new_n8497, new_n8498, new_n8499,
    new_n8500, new_n8501, new_n8502, new_n8503, new_n8504, new_n8505_1,
    new_n8506, new_n8507, new_n8508, new_n8509, new_n8510_1, new_n8511,
    new_n8512, new_n8513, new_n8514, new_n8515, new_n8516, new_n8517,
    new_n8518, new_n8519_1, new_n8520, new_n8521, new_n8522, new_n8523,
    new_n8524, new_n8525, new_n8526_1, new_n8527, new_n8528, new_n8529,
    new_n8530, new_n8531, new_n8532, new_n8533, new_n8534, new_n8535_1,
    new_n8536, new_n8537, new_n8538, new_n8539, new_n8540, new_n8541,
    new_n8542, new_n8543, new_n8544, new_n8545, new_n8546, new_n8547,
    new_n8548, new_n8549, new_n8550_1, new_n8551, new_n8552, new_n8553,
    new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559,
    new_n8560, new_n8561, new_n8562, new_n8563_1, new_n8564, new_n8565,
    new_n8566, new_n8567, new_n8568, new_n8569, new_n8570, new_n8571,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8578, new_n8579, new_n8580, new_n8581_1, new_n8582, new_n8583,
    new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589,
    new_n8590, new_n8591, new_n8592, new_n8593, new_n8594_1, new_n8595,
    new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601,
    new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607,
    new_n8608_1, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613,
    new_n8614_1, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619,
    new_n8620_1, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625,
    new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637_1,
    new_n8638_1, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8644, new_n8645, new_n8646, new_n8647, new_n8648, new_n8649,
    new_n8650, new_n8651, new_n8652, new_n8653, new_n8654, new_n8655,
    new_n8656_1, new_n8657, new_n8658, new_n8659, new_n8660, new_n8661,
    new_n8662_1, new_n8663, new_n8664, new_n8665, new_n8666, new_n8667,
    new_n8668, new_n8669, new_n8670, new_n8671, new_n8672, new_n8673,
    new_n8674, new_n8675, new_n8676, new_n8677, new_n8678_1, new_n8679,
    new_n8680, new_n8681, new_n8682, new_n8683, new_n8684, new_n8685,
    new_n8686, new_n8687_1, new_n8688, new_n8689, new_n8690, new_n8691,
    new_n8692, new_n8693, new_n8694_1, new_n8695, new_n8696, new_n8697,
    new_n8698, new_n8699, new_n8700, new_n8701, new_n8702, new_n8703,
    new_n8704, new_n8705, new_n8706, new_n8707, new_n8708, new_n8709,
    new_n8710, new_n8711, new_n8712, new_n8713, new_n8714, new_n8715,
    new_n8716_1, new_n8719, new_n8720, new_n8721_1, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744_1, new_n8745_1, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782_1, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803_1, new_n8804, new_n8805, new_n8806_1, new_n8807,
    new_n8808, new_n8809_1, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819,
    new_n8820, new_n8821_1, new_n8822, new_n8823, new_n8824_1, new_n8825,
    new_n8826, new_n8827_1, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849_1,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856_1, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861_1,
    new_n8862_1, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869_1, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884_1, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909_1,
    new_n8910, new_n8911_1, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8917, new_n8918, new_n8919, new_n8920_1, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943_1, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8958, new_n8959,
    new_n8960, new_n8961, new_n8962, new_n8963, new_n8964_1, new_n8965,
    new_n8966, new_n8967, new_n8968, new_n8969, new_n8970, new_n8971_1,
    new_n8972, new_n8973, new_n8974, new_n8975, new_n8976, new_n8977,
    new_n8978, new_n8979, new_n8980, new_n8981, new_n8982_1, new_n8983,
    new_n8984, new_n8985, new_n8986, new_n8987, new_n8988, new_n8989,
    new_n8990, new_n8991, new_n8992, new_n8993_1, new_n8994, new_n8995,
    new_n8996, new_n8997, new_n8998, new_n8999, new_n9000, new_n9001,
    new_n9002, new_n9003_1, new_n9004, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012_1, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032_1,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042_1, new_n9043, new_n9044,
    new_n9045, new_n9046_1, new_n9047_1, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090_1, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104_1,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9110, new_n9111,
    new_n9112, new_n9113, new_n9114, new_n9115, new_n9116, new_n9117,
    new_n9118, new_n9119, new_n9120, new_n9121, new_n9122, new_n9123,
    new_n9124, new_n9125, new_n9126, new_n9127, new_n9128, new_n9129_1,
    new_n9130, new_n9131, new_n9132, new_n9133, new_n9134, new_n9135,
    new_n9136, new_n9137, new_n9138, new_n9139, new_n9140, new_n9141,
    new_n9142, new_n9143, new_n9144, new_n9145, new_n9146_1, new_n9147,
    new_n9148, new_n9149, new_n9150, new_n9151, new_n9152, new_n9153,
    new_n9154, new_n9155, new_n9156, new_n9157, new_n9158, new_n9159,
    new_n9160, new_n9161, new_n9162, new_n9163, new_n9164_1, new_n9165,
    new_n9166_1, new_n9167, new_n9168, new_n9169, new_n9170, new_n9171,
    new_n9172_1, new_n9173, new_n9174, new_n9175, new_n9176, new_n9177,
    new_n9178, new_n9179, new_n9180, new_n9181, new_n9182_1, new_n9183,
    new_n9184, new_n9185, new_n9186, new_n9187, new_n9188, new_n9189,
    new_n9190, new_n9191_1, new_n9192, new_n9193, new_n9195, new_n9196,
    new_n9197, new_n9198, new_n9199, new_n9200, new_n9201, new_n9202,
    new_n9203, new_n9204, new_n9205, new_n9206, new_n9207, new_n9208,
    new_n9209, new_n9210, new_n9211, new_n9212, new_n9213, new_n9214,
    new_n9215, new_n9216, new_n9217_1, new_n9218, new_n9219, new_n9220_1,
    new_n9221, new_n9222, new_n9223, new_n9224, new_n9225, new_n9226,
    new_n9227, new_n9228, new_n9229, new_n9230, new_n9231, new_n9232,
    new_n9233, new_n9234, new_n9235, new_n9236, new_n9237, new_n9238,
    new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244,
    new_n9245, new_n9246_1, new_n9247, new_n9248, new_n9249, new_n9250,
    new_n9251_1, new_n9252, new_n9253, new_n9254, new_n9255, new_n9256,
    new_n9257, new_n9258, new_n9259_1, new_n9260, new_n9261_1, new_n9262,
    new_n9263, new_n9264, new_n9265, new_n9266, new_n9267, new_n9268,
    new_n9269, new_n9270, new_n9271, new_n9272, new_n9273, new_n9274,
    new_n9275, new_n9276, new_n9277, new_n9278, new_n9279, new_n9280,
    new_n9281, new_n9282, new_n9283, new_n9284, new_n9285, new_n9286,
    new_n9287_1, new_n9288, new_n9289, new_n9290, new_n9291, new_n9292,
    new_n9293, new_n9294, new_n9295, new_n9296, new_n9297, new_n9298,
    new_n9299, new_n9300, new_n9301, new_n9302, new_n9303, new_n9304,
    new_n9305, new_n9306, new_n9307, new_n9308_1, new_n9309, new_n9310,
    new_n9311, new_n9312, new_n9313, new_n9314, new_n9315, new_n9316,
    new_n9317, new_n9318_1, new_n9319, new_n9320, new_n9321, new_n9322,
    new_n9323_1, new_n9324, new_n9325, new_n9326, new_n9327, new_n9328,
    new_n9329, new_n9330, new_n9331, new_n9332, new_n9333, new_n9334,
    new_n9335, new_n9336, new_n9337, new_n9338, new_n9339, new_n9340,
    new_n9341, new_n9342, new_n9343, new_n9344_1, new_n9345, new_n9346,
    new_n9347, new_n9348, new_n9349, new_n9350, new_n9351, new_n9352,
    new_n9353, new_n9354, new_n9355, new_n9356, new_n9357, new_n9358,
    new_n9359, new_n9360, new_n9361, new_n9362, new_n9363, new_n9364_1,
    new_n9365, new_n9366, new_n9367, new_n9368, new_n9369, new_n9370,
    new_n9371_1, new_n9372_1, new_n9373, new_n9374, new_n9375, new_n9376,
    new_n9377, new_n9378, new_n9379, new_n9380_1, new_n9381, new_n9382_1,
    new_n9383, new_n9384, new_n9385, new_n9386, new_n9387, new_n9388,
    new_n9389, new_n9390, new_n9391, new_n9392, new_n9393, new_n9394,
    new_n9395, new_n9396_1, new_n9397, new_n9398, new_n9399_1, new_n9400,
    new_n9401, new_n9402, new_n9403_1, new_n9404, new_n9405, new_n9406,
    new_n9407, new_n9408, new_n9409, new_n9410, new_n9411, new_n9412,
    new_n9413, new_n9414, new_n9415, new_n9416, new_n9417, new_n9418,
    new_n9419_1, new_n9420, new_n9421, new_n9422, new_n9423_1, new_n9424,
    new_n9425, new_n9426, new_n9427, new_n9428, new_n9429, new_n9430_1,
    new_n9431, new_n9432, new_n9433, new_n9434, new_n9435_1, new_n9436,
    new_n9437, new_n9438, new_n9439, new_n9440, new_n9441, new_n9442,
    new_n9443, new_n9444, new_n9445_1, new_n9446, new_n9447, new_n9448,
    new_n9449, new_n9450, new_n9451_1, new_n9452, new_n9453, new_n9454,
    new_n9455, new_n9456, new_n9457, new_n9458_1, new_n9459_1, new_n9460_1,
    new_n9461, new_n9462, new_n9463, new_n9464, new_n9465, new_n9466,
    new_n9467, new_n9468, new_n9469, new_n9470, new_n9471, new_n9472,
    new_n9473, new_n9474, new_n9475, new_n9476, new_n9477, new_n9478,
    new_n9479, new_n9481, new_n9482, new_n9483, new_n9484, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493_1, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507_1, new_n9508_1, new_n9509, new_n9510,
    new_n9511, new_n9512_1, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552_1,
    new_n9553, new_n9554_1, new_n9555, new_n9556_1, new_n9557_1,
    new_n9558_1, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598_1, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616_1, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622_1, new_n9623,
    new_n9624, new_n9625, new_n9626_1, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633_1, new_n9634, new_n9635_1,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646_1, new_n9647,
    new_n9648_1, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689_1, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695_1, new_n9696,
    new_n9697, new_n9698, new_n9699_1, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726_1,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753_1, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761_1, new_n9762,
    new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1, new_n9768,
    new_n9769, new_n9770, new_n9771_1, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778_1, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783_1, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803_1, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832_1, new_n9833_1, new_n9834,
    new_n9835, new_n9836, new_n9841, new_n9842, new_n9843, new_n9844,
    new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850,
    new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856,
    new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862,
    new_n9863, new_n9864, new_n9865, new_n9866, new_n9867_1, new_n9868,
    new_n9869, new_n9870, new_n9871, new_n9872_1, new_n9873, new_n9874,
    new_n9875, new_n9876, new_n9877, new_n9878, new_n9879, new_n9880,
    new_n9881, new_n9882, new_n9883, new_n9884, new_n9885, new_n9886,
    new_n9887, new_n9888, new_n9889, new_n9890_1, new_n9891, new_n9892,
    new_n9893, new_n9894, new_n9895, new_n9896, new_n9897, new_n9898,
    new_n9899, new_n9900, new_n9901, new_n9902, new_n9903, new_n9904,
    new_n9905, new_n9906, new_n9907, new_n9908, new_n9909, new_n9910,
    new_n9911, new_n9912, new_n9913, new_n9914, new_n9915, new_n9916,
    new_n9917_1, new_n9918, new_n9919_1, new_n9920, new_n9921, new_n9922,
    new_n9923, new_n9924, new_n9925, new_n9926_1, new_n9927, new_n9928,
    new_n9929, new_n9930, new_n9931, new_n9932, new_n9933, new_n9934_1,
    new_n9935, new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940,
    new_n9941, new_n9942_1, new_n9943, new_n9944, new_n9945, new_n9946_1,
    new_n9947, new_n9948, new_n9949, new_n9950, new_n9951, new_n9952,
    new_n9953, new_n9954, new_n9955, new_n9956, new_n9957, new_n9958,
    new_n9959, new_n9960, new_n9961, new_n9962, new_n9963, new_n9964,
    new_n9965, new_n9966, new_n9967_1, new_n9968_1, new_n9969, new_n9970,
    new_n9971, new_n9972, new_n9973, new_n9974, new_n9975, new_n9976,
    new_n9977, new_n9978, new_n9979, new_n9980, new_n9981, new_n9982,
    new_n9983, new_n9984, new_n9985, new_n9986, new_n9987, new_n9988,
    new_n9989, new_n9990, new_n9991, new_n9992, new_n9993, new_n9994,
    new_n9995, new_n9996, new_n9997, new_n9998, new_n9999, new_n10000,
    new_n10001, new_n10002, new_n10003, new_n10004, new_n10005, new_n10006,
    new_n10007, new_n10008, new_n10009_1, new_n10010_1, new_n10011,
    new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017_1, new_n10018_1, new_n10019_1, new_n10020, new_n10021_1,
    new_n10022, new_n10023, new_n10025, new_n10026, new_n10027, new_n10028,
    new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034,
    new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10048, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053_1, new_n10054, new_n10055_1, new_n10056, new_n10057_1,
    new_n10058, new_n10059, new_n10060, new_n10061, new_n10062, new_n10063,
    new_n10064, new_n10065, new_n10066, new_n10067, new_n10068, new_n10069,
    new_n10070, new_n10071, new_n10072, new_n10073, new_n10074, new_n10075,
    new_n10076, new_n10077, new_n10078, new_n10079, new_n10080, new_n10081,
    new_n10082, new_n10083, new_n10084, new_n10085, new_n10086, new_n10087,
    new_n10088, new_n10089, new_n10090, new_n10091, new_n10092, new_n10093,
    new_n10094, new_n10095, new_n10096_1, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101_1, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111_1, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117_1, new_n10118, new_n10121,
    new_n10122, new_n10123, new_n10124, new_n10125_1, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158_1, new_n10159, new_n10160, new_n10161,
    new_n10162, new_n10163, new_n10164, new_n10165_1, new_n10166,
    new_n10167, new_n10168, new_n10169, new_n10170, new_n10171, new_n10172,
    new_n10173, new_n10174, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201_1,
    new_n10202, new_n10203, new_n10204, new_n10205, new_n10206, new_n10207,
    new_n10208, new_n10209, new_n10210, new_n10211, new_n10212, new_n10213,
    new_n10214, new_n10215, new_n10216, new_n10217, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236_1, new_n10237,
    new_n10238, new_n10239_1, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244_1, new_n10245, new_n10246, new_n10247,
    new_n10248, new_n10249, new_n10250_1, new_n10251, new_n10252,
    new_n10253, new_n10254, new_n10255, new_n10256, new_n10257, new_n10258,
    new_n10259, new_n10260, new_n10261_1, new_n10262_1, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275_1, new_n10276, new_n10277, new_n10278, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287_1, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295_1,
    new_n10296, new_n10297, new_n10298, new_n10299, new_n10300, new_n10301,
    new_n10302, new_n10303, new_n10304, new_n10305, new_n10306, new_n10307,
    new_n10308, new_n10309, new_n10310, new_n10311, new_n10312, new_n10313,
    new_n10314, new_n10315, new_n10316, new_n10317, new_n10318, new_n10319,
    new_n10320, new_n10321_1, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326_1, new_n10327_1, new_n10328, new_n10329,
    new_n10330_1, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339,
    new_n10340_1, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345_1, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356_1, new_n10357, new_n10358, new_n10359, new_n10360,
    new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366,
    new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372_1, new_n10374, new_n10376, new_n10377, new_n10378,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384,
    new_n10385_1, new_n10386, new_n10387_1, new_n10388_1, new_n10389,
    new_n10390_1, new_n10391, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10400, new_n10402,
    new_n10403, new_n10404_1, new_n10405_1, new_n10406, new_n10407,
    new_n10408, new_n10409_1, new_n10410, new_n10411_1, new_n10412,
    new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418,
    new_n10419, new_n10420_1, new_n10421, new_n10422, new_n10423,
    new_n10424, new_n10425, new_n10426, new_n10427, new_n10428, new_n10429,
    new_n10430, new_n10431, new_n10432_1, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484_1, new_n10485, new_n10486, new_n10487,
    new_n10488, new_n10489_1, new_n10490, new_n10491, new_n10492,
    new_n10493, new_n10494, new_n10495, new_n10496, new_n10497, new_n10498,
    new_n10499, new_n10500, new_n10501, new_n10502, new_n10503, new_n10504,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510,
    new_n10511, new_n10512, new_n10513, new_n10514_1, new_n10515,
    new_n10516, new_n10517, new_n10518, new_n10519, new_n10520, new_n10521,
    new_n10522, new_n10523, new_n10524, new_n10525_1, new_n10526,
    new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540_1, new_n10541, new_n10542, new_n10543,
    new_n10544, new_n10545, new_n10546, new_n10547, new_n10548, new_n10549,
    new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555,
    new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561_1, new_n10562, new_n10563, new_n10564_1, new_n10565,
    new_n10566, new_n10567, new_n10568, new_n10569, new_n10570, new_n10571,
    new_n10572, new_n10573, new_n10574, new_n10575, new_n10576,
    new_n10577_1, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588_1, new_n10589, new_n10590, new_n10591, new_n10592,
    new_n10593_1, new_n10594, new_n10595_1, new_n10596, new_n10597,
    new_n10598, new_n10599, new_n10600, new_n10601, new_n10602, new_n10603,
    new_n10604, new_n10605, new_n10606, new_n10607, new_n10608, new_n10609,
    new_n10610, new_n10611_1, new_n10612, new_n10613, new_n10614_1,
    new_n10615, new_n10616, new_n10617_1, new_n10618, new_n10619,
    new_n10620, new_n10621, new_n10622, new_n10623, new_n10624, new_n10625,
    new_n10626, new_n10627, new_n10628_1, new_n10629, new_n10630,
    new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636,
    new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642,
    new_n10643, new_n10644, new_n10645, new_n10646, new_n10647_1,
    new_n10648, new_n10649, new_n10650_1, new_n10651, new_n10652,
    new_n10653_1, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692_1,
    new_n10693, new_n10694_1, new_n10695, new_n10696, new_n10698,
    new_n10699, new_n10700, new_n10701_1, new_n10702, new_n10703,
    new_n10704, new_n10705, new_n10706, new_n10707, new_n10708, new_n10709,
    new_n10710_1, new_n10711, new_n10712_1, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739_1, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756_1, new_n10757, new_n10758, new_n10759, new_n10760,
    new_n10761, new_n10762, new_n10763_1, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775_1, new_n10776,
    new_n10777, new_n10778, new_n10779, new_n10780_1, new_n10781,
    new_n10782, new_n10783, new_n10784, new_n10785, new_n10786, new_n10787,
    new_n10788, new_n10789, new_n10790, new_n10791, new_n10792_1,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817_1, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834_1, new_n10835, new_n10836, new_n10837, new_n10838,
    new_n10839, new_n10840, new_n10841, new_n10842, new_n10843, new_n10844,
    new_n10845, new_n10846, new_n10847, new_n10848, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874_1, new_n10875, new_n10876, new_n10877, new_n10878,
    new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884,
    new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890,
    new_n10891, new_n10892, new_n10893, new_n10894, new_n10896, new_n10897,
    new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903,
    new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909,
    new_n10910, new_n10911, new_n10912, new_n10913, new_n10914, new_n10915,
    new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921,
    new_n10922, new_n10923, new_n10924_1, new_n10925, new_n10926,
    new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943_1,
    new_n10944, new_n10945, new_n10946, new_n10947, new_n10948, new_n10949,
    new_n10950, new_n10951, new_n10952, new_n10953, new_n10954, new_n10955,
    new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961_1, new_n10962, new_n10963, new_n10964, new_n10965,
    new_n10966, new_n10967, new_n10968, new_n10969, new_n10970, new_n10971,
    new_n10972, new_n10973, new_n10974, new_n10975, new_n10976, new_n10977,
    new_n10978, new_n10979, new_n10980, new_n10981, new_n10982, new_n10983,
    new_n10984, new_n10985, new_n10986, new_n10987, new_n10988, new_n10989,
    new_n10990, new_n10991, new_n10992, new_n10993, new_n10994, new_n10995,
    new_n10996, new_n10997, new_n10998, new_n10999, new_n11000, new_n11001,
    new_n11002, new_n11003, new_n11004, new_n11005_1, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011_1,
    new_n11012, new_n11013, new_n11014, new_n11015, new_n11016, new_n11017,
    new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023_1, new_n11024, new_n11025_1, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044_1,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055,
    new_n11056_1, new_n11057, new_n11058, new_n11059, new_n11060,
    new_n11061, new_n11062, new_n11063_1, new_n11064, new_n11065,
    new_n11066, new_n11067, new_n11068, new_n11069, new_n11070, new_n11071,
    new_n11072, new_n11073, new_n11074, new_n11075, new_n11076, new_n11077,
    new_n11078_1, new_n11079, new_n11080_1, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094_1, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101_1, new_n11102, new_n11103_1,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109,
    new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115,
    new_n11116, new_n11117, new_n11118, new_n11119, new_n11120_1,
    new_n11121_1, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127_1, new_n11128, new_n11129, new_n11130,
    new_n11131, new_n11132_1, new_n11133, new_n11134_1, new_n11135,
    new_n11136, new_n11137, new_n11138_1, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11146,
    new_n11147, new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153, new_n11154, new_n11155, new_n11156, new_n11157, new_n11158,
    new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164,
    new_n11165, new_n11166, new_n11167, new_n11168, new_n11169, new_n11170,
    new_n11171, new_n11173, new_n11174, new_n11175, new_n11176, new_n11177,
    new_n11178, new_n11179, new_n11180, new_n11181, new_n11182_1,
    new_n11183, new_n11184_1, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192_1,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201_1, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216, new_n11217, new_n11218, new_n11219, new_n11220_1,
    new_n11221, new_n11222, new_n11223_1, new_n11224, new_n11225,
    new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231,
    new_n11232, new_n11233, new_n11234_1, new_n11235, new_n11236,
    new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242,
    new_n11243, new_n11244, new_n11245_1, new_n11246, new_n11247,
    new_n11248, new_n11249, new_n11250, new_n11251, new_n11252, new_n11253,
    new_n11254, new_n11255, new_n11256, new_n11257, new_n11258, new_n11259,
    new_n11260, new_n11261_1, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266_1, new_n11267, new_n11268, new_n11269,
    new_n11270, new_n11271, new_n11272, new_n11273_1, new_n11274,
    new_n11275_1, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11281, new_n11282, new_n11283, new_n11284, new_n11285, new_n11286,
    new_n11287, new_n11288, new_n11289, new_n11290_1, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296, new_n11297,
    new_n11298, new_n11299, new_n11300, new_n11301, new_n11302_1,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311, new_n11312, new_n11313_1,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324,
    new_n11325_1, new_n11326_1, new_n11327, new_n11328, new_n11329,
    new_n11330_1, new_n11331, new_n11332, new_n11333, new_n11334,
    new_n11335, new_n11336, new_n11337, new_n11338, new_n11339, new_n11340,
    new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346,
    new_n11347_1, new_n11348_1, new_n11349, new_n11350, new_n11351,
    new_n11352_1, new_n11353, new_n11354, new_n11355, new_n11356_1,
    new_n11357, new_n11358, new_n11359, new_n11360, new_n11361, new_n11362,
    new_n11363, new_n11364, new_n11365, new_n11366, new_n11367, new_n11368,
    new_n11369, new_n11370, new_n11371, new_n11372, new_n11373, new_n11374,
    new_n11375_1, new_n11376, new_n11377, new_n11378, new_n11379_1,
    new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385,
    new_n11386_1, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391_1, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398_1, new_n11399, new_n11400, new_n11401,
    new_n11402, new_n11403_1, new_n11404, new_n11405, new_n11406,
    new_n11407, new_n11408, new_n11409, new_n11410, new_n11411, new_n11412,
    new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418,
    new_n11419_1, new_n11420, new_n11421, new_n11422, new_n11423,
    new_n11424_1, new_n11425, new_n11426, new_n11427, new_n11428,
    new_n11429, new_n11430, new_n11431, new_n11432, new_n11433, new_n11434,
    new_n11435, new_n11436, new_n11437, new_n11438, new_n11439_1,
    new_n11440, new_n11441, new_n11442, new_n11443, new_n11444, new_n11445,
    new_n11446, new_n11447, new_n11448, new_n11449, new_n11450, new_n11451,
    new_n11452, new_n11453, new_n11454, new_n11455_1, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461,
    new_n11462_1, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470_1, new_n11471,
    new_n11472_1, new_n11473_1, new_n11474, new_n11475, new_n11476,
    new_n11477, new_n11478, new_n11479_1, new_n11480, new_n11481_1,
    new_n11482, new_n11483, new_n11484, new_n11485, new_n11486_1,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496_1, new_n11497,
    new_n11498, new_n11499, new_n11500, new_n11501, new_n11502,
    new_n11503_1, new_n11504, new_n11505, new_n11506_1, new_n11507,
    new_n11508, new_n11509, new_n11510, new_n11511, new_n11512, new_n11513,
    new_n11514, new_n11515_1, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535, new_n11536,
    new_n11537, new_n11538_1, new_n11539, new_n11540, new_n11541,
    new_n11542, new_n11543, new_n11544, new_n11545, new_n11546, new_n11547,
    new_n11548_1, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563,
    new_n11564_1, new_n11565, new_n11566_1, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11572, new_n11573, new_n11574, new_n11576,
    new_n11577, new_n11578, new_n11579_1, new_n11580_1, new_n11581,
    new_n11582, new_n11583, new_n11584, new_n11585, new_n11586, new_n11587,
    new_n11588, new_n11589, new_n11590, new_n11591_1, new_n11592,
    new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607_1, new_n11608, new_n11609,
    new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615_1, new_n11616, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627, new_n11628, new_n11629, new_n11630_1,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647_1,
    new_n11648, new_n11649, new_n11650, new_n11651, new_n11652, new_n11653,
    new_n11654, new_n11655, new_n11656, new_n11657, new_n11658, new_n11659,
    new_n11660, new_n11661, new_n11662, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667_1, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682_1,
    new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688,
    new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694,
    new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700,
    new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707, new_n11708, new_n11709, new_n11710_1, new_n11711,
    new_n11712_1, new_n11713, new_n11714, new_n11715, new_n11716,
    new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722,
    new_n11723, new_n11724_1, new_n11725, new_n11726, new_n11727,
    new_n11728, new_n11729, new_n11730, new_n11731, new_n11732, new_n11733,
    new_n11734, new_n11735, new_n11736_1, new_n11737, new_n11738,
    new_n11739, new_n11740, new_n11741_1, new_n11742, new_n11743,
    new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749_1, new_n11750, new_n11751, new_n11752, new_n11753,
    new_n11754, new_n11755, new_n11756, new_n11757, new_n11758, new_n11759,
    new_n11760, new_n11761, new_n11762, new_n11763, new_n11764, new_n11765,
    new_n11766, new_n11767, new_n11768, new_n11769, new_n11770_1,
    new_n11771_1, new_n11772, new_n11773, new_n11774, new_n11775_1,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780, new_n11781,
    new_n11782, new_n11783, new_n11784, new_n11785, new_n11786, new_n11787,
    new_n11788, new_n11789, new_n11790, new_n11791, new_n11792, new_n11793,
    new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799,
    new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805,
    new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811,
    new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818_1, new_n11819, new_n11820, new_n11821, new_n11822,
    new_n11823, new_n11824, new_n11825, new_n11826, new_n11827, new_n11828,
    new_n11829, new_n11830, new_n11831, new_n11832, new_n11833, new_n11834,
    new_n11835, new_n11836, new_n11837_1, new_n11838, new_n11839,
    new_n11840, new_n11841_1, new_n11842_1, new_n11843_1, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897,
    new_n11898_1, new_n11899, new_n11900, new_n11901, new_n11902,
    new_n11903, new_n11904, new_n11905_1, new_n11906, new_n11908,
    new_n11909, new_n11910, new_n11911, new_n11912, new_n11913, new_n11914,
    new_n11915, new_n11916, new_n11917, new_n11918, new_n11919, new_n11920,
    new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926_1, new_n11927, new_n11928, new_n11929, new_n11930,
    new_n11931, new_n11932, new_n11933, new_n11934, new_n11935, new_n11936,
    new_n11937, new_n11938, new_n11939, new_n11940, new_n11941, new_n11942,
    new_n11943, new_n11944, new_n11945, new_n11946, new_n11947, new_n11948,
    new_n11949, new_n11950, new_n11951, new_n11952, new_n11953, new_n11954,
    new_n11955, new_n11956, new_n11957, new_n11958, new_n11959, new_n11960,
    new_n11961, new_n11962, new_n11963, new_n11964, new_n11965_1,
    new_n11966, new_n11967, new_n11968, new_n11969, new_n11971, new_n11972,
    new_n11973, new_n11974, new_n11975, new_n11976, new_n11978, new_n11979,
    new_n11980_1, new_n11981, new_n11982, new_n11983, new_n11984,
    new_n11985, new_n11986, new_n11987, new_n11988, new_n11989, new_n11990,
    new_n11991, new_n11992, new_n11993, new_n11994, new_n11995, new_n11996,
    new_n11997, new_n11998, new_n11999, new_n12000_1, new_n12001,
    new_n12002, new_n12003_1, new_n12004, new_n12005, new_n12006,
    new_n12007, new_n12008, new_n12009, new_n12010, new_n12011_1,
    new_n12012, new_n12013, new_n12014, new_n12015, new_n12016, new_n12017,
    new_n12018, new_n12019, new_n12020, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044, new_n12045, new_n12046, new_n12047,
    new_n12048, new_n12049, new_n12050, new_n12051, new_n12052, new_n12053,
    new_n12054, new_n12055, new_n12056, new_n12057, new_n12058, new_n12059,
    new_n12060, new_n12061, new_n12062, new_n12063, new_n12064, new_n12065,
    new_n12066, new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072_1, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12108, new_n12109, new_n12110,
    new_n12111, new_n12112, new_n12113_1, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120,
    new_n12121_1, new_n12122, new_n12123, new_n12124, new_n12125,
    new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131_1, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142, new_n12143, new_n12144, new_n12145, new_n12146_1,
    new_n12147, new_n12148, new_n12149, new_n12150, new_n12151,
    new_n12152_1, new_n12153_1, new_n12154, new_n12155, new_n12156,
    new_n12157_1, new_n12158_1, new_n12159, new_n12160, new_n12161_1,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173,
    new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179_1, new_n12180, new_n12181, new_n12182, new_n12183,
    new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189,
    new_n12190, new_n12191, new_n12192_1, new_n12193, new_n12194,
    new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200,
    new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206,
    new_n12207, new_n12208, new_n12209_1, new_n12210, new_n12211,
    new_n12212, new_n12213, new_n12214, new_n12215, new_n12216, new_n12217,
    new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223_1, new_n12224, new_n12225_1, new_n12226, new_n12227,
    new_n12228_1, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235_1, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247, new_n12248, new_n12249,
    new_n12250, new_n12251, new_n12252, new_n12253, new_n12254, new_n12255,
    new_n12256, new_n12257, new_n12258, new_n12259, new_n12260, new_n12261,
    new_n12262, new_n12263, new_n12264, new_n12265, new_n12266, new_n12267,
    new_n12268, new_n12269, new_n12270, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299, new_n12300, new_n12301, new_n12302_1, new_n12303,
    new_n12304_1, new_n12305, new_n12306, new_n12307, new_n12308,
    new_n12309, new_n12310, new_n12311, new_n12312, new_n12313, new_n12314,
    new_n12315_1, new_n12316, new_n12317, new_n12318, new_n12319,
    new_n12320, new_n12321, new_n12322, new_n12323, new_n12324_1,
    new_n12325_1, new_n12326, new_n12327, new_n12328, new_n12329_1,
    new_n12330_1, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341_1, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346_1, new_n12347, new_n12348, new_n12349_1, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364_1, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380_1, new_n12381, new_n12382, new_n12383_1, new_n12384_1,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397_1, new_n12398_1, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408_1, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446_1, new_n12447,
    new_n12448, new_n12449_1, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467_1, new_n12468, new_n12469_1, new_n12470, new_n12471,
    new_n12472, new_n12473, new_n12474, new_n12475, new_n12479, new_n12480,
    new_n12481, new_n12482, new_n12483, new_n12484, new_n12485, new_n12486,
    new_n12487, new_n12488, new_n12489, new_n12490, new_n12491, new_n12492,
    new_n12493, new_n12494, new_n12495_1, new_n12496, new_n12497,
    new_n12498, new_n12499, new_n12500, new_n12501, new_n12502, new_n12503,
    new_n12504, new_n12505, new_n12506, new_n12507_1, new_n12508,
    new_n12509, new_n12510, new_n12511, new_n12514, new_n12515_1,
    new_n12516_1, new_n12517, new_n12518, new_n12519, new_n12520,
    new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526,
    new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540_1, new_n12541, new_n12542, new_n12543,
    new_n12544, new_n12545_1, new_n12546_1, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552_1, new_n12553,
    new_n12554, new_n12555, new_n12556, new_n12557, new_n12558, new_n12559,
    new_n12560, new_n12561, new_n12562_1, new_n12563, new_n12564,
    new_n12565, new_n12566_1, new_n12567, new_n12568, new_n12569_1,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587_1, new_n12588, new_n12589, new_n12590, new_n12591,
    new_n12592, new_n12593_1, new_n12594, new_n12595, new_n12596,
    new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602,
    new_n12603, new_n12604, new_n12605, new_n12606, new_n12607_1,
    new_n12608, new_n12609, new_n12610, new_n12611, new_n12612, new_n12613,
    new_n12614, new_n12615, new_n12616, new_n12617, new_n12618, new_n12619,
    new_n12620_1, new_n12621_1, new_n12622, new_n12623, new_n12624,
    new_n12625, new_n12626_1, new_n12627, new_n12628, new_n12629,
    new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635,
    new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641,
    new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648, new_n12649, new_n12650_1, new_n12651, new_n12652,
    new_n12653, new_n12654_1, new_n12655, new_n12656, new_n12657_1,
    new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663,
    new_n12664, new_n12665_1, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670_1, new_n12671, new_n12672, new_n12673,
    new_n12674, new_n12675, new_n12676, new_n12677, new_n12678, new_n12679,
    new_n12680, new_n12681, new_n12682, new_n12683, new_n12684, new_n12685,
    new_n12686, new_n12687, new_n12688, new_n12689, new_n12690, new_n12691,
    new_n12692, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699,
    new_n12700, new_n12701, new_n12702_1, new_n12703, new_n12704,
    new_n12705, new_n12706, new_n12707_1, new_n12708, new_n12709,
    new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715,
    new_n12716, new_n12717, new_n12718, new_n12719, new_n12720, new_n12721,
    new_n12722, new_n12723, new_n12724, new_n12725_1, new_n12726,
    new_n12727_1, new_n12728, new_n12729, new_n12730, new_n12731,
    new_n12732, new_n12733, new_n12734, new_n12735, new_n12736, new_n12737,
    new_n12738, new_n12739, new_n12740_1, new_n12741, new_n12742_1,
    new_n12743, new_n12744, new_n12745, new_n12746_1, new_n12747,
    new_n12748, new_n12749, new_n12750, new_n12751, new_n12752, new_n12753,
    new_n12754, new_n12755, new_n12756_1, new_n12757, new_n12758,
    new_n12759, new_n12760, new_n12761, new_n12762, new_n12763, new_n12764,
    new_n12765, new_n12766, new_n12767, new_n12768, new_n12769, new_n12770,
    new_n12771, new_n12772, new_n12773, new_n12774, new_n12775, new_n12776,
    new_n12777, new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783_1, new_n12784, new_n12785, new_n12786, new_n12787,
    new_n12788, new_n12789, new_n12790, new_n12791, new_n12792, new_n12793,
    new_n12794, new_n12795, new_n12796, new_n12797, new_n12798, new_n12799,
    new_n12800, new_n12801_1, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811_1, new_n12812_1, new_n12813, new_n12814, new_n12815,
    new_n12816_1, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821_1, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12833, new_n12834, new_n12835, new_n12836, new_n12837, new_n12838,
    new_n12839, new_n12840, new_n12841, new_n12842, new_n12843_1,
    new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849,
    new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855,
    new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861_1, new_n12862, new_n12863, new_n12864_1, new_n12865_1,
    new_n12866, new_n12867, new_n12868, new_n12869, new_n12870_1,
    new_n12871_1, new_n12872, new_n12873_1, new_n12874, new_n12875_1,
    new_n12876, new_n12877, new_n12878, new_n12879, new_n12880, new_n12881,
    new_n12882, new_n12883, new_n12884, new_n12885, new_n12886, new_n12887,
    new_n12888, new_n12889, new_n12890, new_n12891, new_n12892_1,
    new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898,
    new_n12899, new_n12900_1, new_n12901, new_n12902, new_n12903,
    new_n12904_1, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917_1, new_n12918, new_n12919,
    new_n12920, new_n12921, new_n12922, new_n12923, new_n12924, new_n12925,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941_1, new_n12942_1,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956_1, new_n12957, new_n12958, new_n12959,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977,
    new_n12978_1, new_n12979, new_n12980_1, new_n12981, new_n12982,
    new_n12983, new_n12984, new_n12985_1, new_n12986, new_n12987_1,
    new_n12988, new_n12989, new_n12990, new_n12991, new_n12992_1,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002, new_n13003, new_n13004, new_n13005_1, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026_1, new_n13027, new_n13028, new_n13029,
    new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043_1, new_n13044_1, new_n13045, new_n13046,
    new_n13047, new_n13048_1, new_n13049, new_n13050, new_n13051,
    new_n13052, new_n13053, new_n13054_1, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13072, new_n13073, new_n13074_1, new_n13075,
    new_n13076, new_n13077, new_n13078, new_n13079, new_n13080, new_n13081,
    new_n13082_1, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096_1, new_n13097,
    new_n13098, new_n13099, new_n13100, new_n13101, new_n13102, new_n13103,
    new_n13104, new_n13105, new_n13106, new_n13107, new_n13108, new_n13109,
    new_n13110_1, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116_1, new_n13117, new_n13118, new_n13119,
    new_n13120, new_n13121, new_n13122_1, new_n13123, new_n13124,
    new_n13125, new_n13126, new_n13127, new_n13128, new_n13129, new_n13130,
    new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137_1, new_n13138, new_n13139, new_n13140, new_n13141_1,
    new_n13142, new_n13143, new_n13144_1, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168_1, new_n13169,
    new_n13170, new_n13171, new_n13172, new_n13173, new_n13174, new_n13175,
    new_n13176, new_n13177, new_n13178, new_n13179, new_n13180, new_n13181,
    new_n13182, new_n13183, new_n13184, new_n13185, new_n13186, new_n13187,
    new_n13188, new_n13189, new_n13190_1, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197,
    new_n13198_1, new_n13199_1, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13204_1, new_n13205, new_n13206, new_n13207,
    new_n13208, new_n13209_1, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263_1, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270_1,
    new_n13271, new_n13272, new_n13273_1, new_n13274, new_n13275,
    new_n13276, new_n13277, new_n13278, new_n13279, new_n13280, new_n13281,
    new_n13282, new_n13283, new_n13284, new_n13285_1, new_n13286,
    new_n13287, new_n13288, new_n13289, new_n13290, new_n13291, new_n13292,
    new_n13293, new_n13294, new_n13295, new_n13296, new_n13297, new_n13298,
    new_n13299, new_n13300, new_n13301, new_n13302, new_n13303, new_n13304,
    new_n13305, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312,
    new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318,
    new_n13319_1, new_n13320, new_n13321, new_n13322, new_n13323,
    new_n13324, new_n13325, new_n13326, new_n13327, new_n13328, new_n13329,
    new_n13330, new_n13331, new_n13332, new_n13333_1, new_n13334,
    new_n13335, new_n13336, new_n13337, new_n13338_1, new_n13339,
    new_n13340, new_n13341, new_n13343, new_n13344, new_n13345, new_n13346,
    new_n13347, new_n13348, new_n13349, new_n13350, new_n13351, new_n13352,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367_1, new_n13368, new_n13369,
    new_n13370, new_n13371, new_n13372, new_n13373, new_n13374, new_n13375,
    new_n13376, new_n13377, new_n13378, new_n13379, new_n13380, new_n13381,
    new_n13382, new_n13383, new_n13384, new_n13385, new_n13386, new_n13387,
    new_n13388, new_n13389, new_n13390, new_n13391, new_n13392, new_n13393,
    new_n13394, new_n13395, new_n13396, new_n13397, new_n13398, new_n13399,
    new_n13400, new_n13401, new_n13402, new_n13403, new_n13404, new_n13405,
    new_n13406, new_n13407_1, new_n13408, new_n13409_1, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419_1, new_n13420, new_n13421,
    new_n13422, new_n13423, new_n13424_1, new_n13425, new_n13426,
    new_n13427, new_n13428, new_n13429, new_n13430, new_n13431, new_n13432,
    new_n13433, new_n13434, new_n13435, new_n13436, new_n13437, new_n13438,
    new_n13439, new_n13440, new_n13441, new_n13442, new_n13443, new_n13444,
    new_n13445, new_n13446, new_n13447, new_n13448, new_n13449, new_n13450,
    new_n13451, new_n13452, new_n13453_1, new_n13454, new_n13455,
    new_n13456_1, new_n13457_1, new_n13458, new_n13459, new_n13460_1,
    new_n13461, new_n13462, new_n13463, new_n13464, new_n13465, new_n13466,
    new_n13467, new_n13468, new_n13469, new_n13470, new_n13471, new_n13472,
    new_n13473, new_n13474, new_n13475, new_n13476, new_n13477_1,
    new_n13478, new_n13479, new_n13480, new_n13481, new_n13482, new_n13483,
    new_n13484_1, new_n13485, new_n13486_1, new_n13487_1, new_n13488,
    new_n13489, new_n13490_1, new_n13491, new_n13492, new_n13493,
    new_n13494_1, new_n13495, new_n13496, new_n13497, new_n13498,
    new_n13499, new_n13500_1, new_n13501_1, new_n13502, new_n13503,
    new_n13504, new_n13505, new_n13506_1, new_n13507, new_n13508,
    new_n13509, new_n13510, new_n13511, new_n13512, new_n13513, new_n13514,
    new_n13515, new_n13516, new_n13517, new_n13518, new_n13519, new_n13520,
    new_n13521, new_n13522, new_n13523, new_n13524, new_n13525, new_n13526,
    new_n13527, new_n13528, new_n13529, new_n13530, new_n13531, new_n13532,
    new_n13533, new_n13534, new_n13535, new_n13536, new_n13537, new_n13538,
    new_n13539, new_n13540, new_n13541, new_n13542, new_n13543, new_n13544,
    new_n13545, new_n13546, new_n13547, new_n13548_1, new_n13549_1,
    new_n13550, new_n13551_1, new_n13552, new_n13553, new_n13554,
    new_n13555, new_n13556, new_n13557, new_n13558, new_n13559, new_n13560,
    new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566,
    new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572,
    new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578,
    new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584,
    new_n13585, new_n13586, new_n13587, new_n13588, new_n13589, new_n13590,
    new_n13591, new_n13592, new_n13593, new_n13594, new_n13595, new_n13596,
    new_n13597, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602_1, new_n13603, new_n13604, new_n13605, new_n13606,
    new_n13607, new_n13608, new_n13609, new_n13610, new_n13611, new_n13612,
    new_n13613, new_n13614, new_n13615, new_n13616, new_n13617, new_n13618,
    new_n13619, new_n13620, new_n13621, new_n13622, new_n13623, new_n13624,
    new_n13625, new_n13626_1, new_n13627, new_n13628, new_n13629,
    new_n13630, new_n13631, new_n13632, new_n13633, new_n13634, new_n13635,
    new_n13636, new_n13637, new_n13638, new_n13639, new_n13640, new_n13641,
    new_n13642, new_n13643, new_n13644, new_n13645, new_n13646, new_n13647,
    new_n13648, new_n13649, new_n13650, new_n13651, new_n13652, new_n13653,
    new_n13654, new_n13655, new_n13656, new_n13657, new_n13658, new_n13659,
    new_n13660, new_n13661, new_n13662, new_n13663, new_n13664, new_n13665,
    new_n13666, new_n13667, new_n13668_1, new_n13669, new_n13670,
    new_n13671, new_n13672, new_n13673, new_n13674, new_n13675, new_n13676,
    new_n13679, new_n13680, new_n13681, new_n13682, new_n13683_1,
    new_n13684, new_n13685, new_n13686, new_n13687, new_n13688, new_n13689,
    new_n13690, new_n13691, new_n13692, new_n13693, new_n13694, new_n13695,
    new_n13696, new_n13697, new_n13698, new_n13699, new_n13700, new_n13701,
    new_n13702, new_n13703, new_n13704, new_n13705, new_n13706, new_n13707,
    new_n13708_1, new_n13709, new_n13710_1, new_n13711, new_n13712,
    new_n13713, new_n13714_1, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719_1, new_n13720, new_n13721, new_n13722_1,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13756,
    new_n13757, new_n13758, new_n13759, new_n13760, new_n13761, new_n13762,
    new_n13763, new_n13764_1, new_n13765, new_n13766, new_n13767,
    new_n13768, new_n13769, new_n13770, new_n13771, new_n13772, new_n13773,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781_1,
    new_n13782, new_n13783_1, new_n13784, new_n13785, new_n13786,
    new_n13787, new_n13788, new_n13789, new_n13790, new_n13791, new_n13792,
    new_n13793, new_n13794, new_n13795, new_n13796, new_n13797,
    new_n13798_1, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13806, new_n13807, new_n13808, new_n13809, new_n13810, new_n13811,
    new_n13812, new_n13813, new_n13814, new_n13815, new_n13816, new_n13817,
    new_n13818, new_n13819, new_n13820, new_n13821, new_n13822, new_n13823,
    new_n13824, new_n13825, new_n13826, new_n13827, new_n13828, new_n13829,
    new_n13830, new_n13831, new_n13832, new_n13833, new_n13834,
    new_n13835_1, new_n13836, new_n13837, new_n13838, new_n13839,
    new_n13840, new_n13841, new_n13842, new_n13843, new_n13844, new_n13845,
    new_n13847, new_n13848, new_n13849, new_n13850_1, new_n13851_1,
    new_n13852, new_n13853, new_n13854, new_n13855, new_n13856, new_n13857,
    new_n13858, new_n13859, new_n13860, new_n13861, new_n13862, new_n13863,
    new_n13864, new_n13865, new_n13866, new_n13867, new_n13868, new_n13869,
    new_n13870, new_n13871, new_n13872, new_n13873, new_n13874, new_n13875,
    new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884,
    new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890,
    new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13911, new_n13912_1, new_n13913,
    new_n13914_1, new_n13915, new_n13916, new_n13917, new_n13918,
    new_n13919, new_n13920, new_n13921, new_n13922_1, new_n13923_1,
    new_n13924, new_n13925, new_n13926, new_n13927, new_n13928, new_n13929,
    new_n13932, new_n13933, new_n13934, new_n13935, new_n13936, new_n13937,
    new_n13938, new_n13939, new_n13940, new_n13941, new_n13942, new_n13943,
    new_n13944, new_n13945, new_n13946, new_n13947, new_n13948, new_n13949,
    new_n13950, new_n13951_1, new_n13952, new_n13953, new_n13954,
    new_n13955, new_n13956, new_n13957, new_n13958, new_n13959, new_n13960,
    new_n13961, new_n13962, new_n13963, new_n13964, new_n13965, new_n13966,
    new_n13967, new_n13968, new_n13969, new_n13970, new_n13971, new_n13972,
    new_n13973, new_n13974, new_n13975, new_n13976, new_n13977, new_n13978,
    new_n13979, new_n13980, new_n13981, new_n13982, new_n13983, new_n13984,
    new_n13985, new_n13986, new_n13987, new_n13988, new_n13989, new_n13990,
    new_n13991, new_n13992, new_n13993, new_n13994, new_n13995, new_n13996,
    new_n13997, new_n13998, new_n13999, new_n14000, new_n14001, new_n14002,
    new_n14003, new_n14004_1, new_n14005, new_n14006, new_n14007,
    new_n14008, new_n14009, new_n14010, new_n14011, new_n14012, new_n14013,
    new_n14014, new_n14015, new_n14016, new_n14017, new_n14018, new_n14019,
    new_n14020, new_n14021, new_n14022, new_n14023, new_n14024, new_n14025,
    new_n14026, new_n14027, new_n14028, new_n14029, new_n14030, new_n14031,
    new_n14032, new_n14033, new_n14034, new_n14035, new_n14036_1,
    new_n14037, new_n14038, new_n14039, new_n14040, new_n14041, new_n14042,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059_1, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071_1,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081_1, new_n14082,
    new_n14083, new_n14084, new_n14085, new_n14086, new_n14087, new_n14088,
    new_n14089, new_n14090_1, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095_1, new_n14096, new_n14097, new_n14098,
    new_n14099, new_n14100, new_n14101, new_n14102, new_n14103, new_n14104,
    new_n14105, new_n14106, new_n14107_1, new_n14108, new_n14109,
    new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121_1, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126_1, new_n14127, new_n14128, new_n14129, new_n14130_1,
    new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136_1, new_n14137, new_n14138, new_n14139, new_n14140,
    new_n14141, new_n14142, new_n14143, new_n14144, new_n14145, new_n14146,
    new_n14147_1, new_n14148_1, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14168, new_n14169, new_n14170,
    new_n14171, new_n14172, new_n14173, new_n14174_1, new_n14175,
    new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181,
    new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187,
    new_n14188, new_n14189, new_n14190_1, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211_1, new_n14212, new_n14213, new_n14214, new_n14215,
    new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221,
    new_n14222_1, new_n14223, new_n14226, new_n14227, new_n14228,
    new_n14229, new_n14230_1, new_n14231, new_n14232, new_n14233,
    new_n14234, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267_1, new_n14268, new_n14269,
    new_n14270, new_n14271_1, new_n14272, new_n14273, new_n14274,
    new_n14275_1, new_n14276, new_n14277_1, new_n14278, new_n14279,
    new_n14280, new_n14281, new_n14282, new_n14283, new_n14284, new_n14285,
    new_n14286, new_n14287, new_n14288, new_n14289, new_n14290, new_n14291,
    new_n14292, new_n14293, new_n14294_1, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310_1, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14320, new_n14321, new_n14322, new_n14323_1, new_n14324,
    new_n14325, new_n14326_1, new_n14327, new_n14328, new_n14329,
    new_n14330, new_n14331, new_n14332, new_n14333, new_n14334, new_n14335,
    new_n14336, new_n14337, new_n14338, new_n14339, new_n14340, new_n14341,
    new_n14342_1, new_n14343, new_n14344, new_n14345_1, new_n14346,
    new_n14347, new_n14348, new_n14349, new_n14350, new_n14351, new_n14352,
    new_n14353_1, new_n14354, new_n14355, new_n14356, new_n14357,
    new_n14358, new_n14359, new_n14360, new_n14361, new_n14362, new_n14363,
    new_n14364_1, new_n14365, new_n14366, new_n14367, new_n14368,
    new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374,
    new_n14375_1, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385,
    new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391,
    new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397,
    new_n14398, new_n14399, new_n14400, new_n14401, new_n14402, new_n14403,
    new_n14404, new_n14405, new_n14406, new_n14407, new_n14408, new_n14409,
    new_n14410, new_n14411, new_n14412_1, new_n14413, new_n14414_1,
    new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420,
    new_n14421, new_n14422, new_n14423, new_n14424, new_n14427, new_n14428,
    new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440_1, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457_1, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464_1, new_n14465, new_n14466,
    new_n14467, new_n14468, new_n14469, new_n14470, new_n14471_1,
    new_n14472, new_n14473, new_n14474, new_n14475_1, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510_1, new_n14512,
    new_n14513, new_n14514, new_n14515, new_n14516, new_n14517, new_n14518,
    new_n14519, new_n14522, new_n14523, new_n14524, new_n14525, new_n14526,
    new_n14527, new_n14528, new_n14529, new_n14530, new_n14531, new_n14532,
    new_n14533, new_n14534, new_n14535, new_n14536, new_n14537, new_n14538,
    new_n14539, new_n14540, new_n14541_1, new_n14542, new_n14543,
    new_n14544, new_n14545, new_n14546_1, new_n14547_1, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570_1, new_n14571,
    new_n14572, new_n14573, new_n14574, new_n14575_1, new_n14576_1,
    new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582,
    new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588,
    new_n14589, new_n14590, new_n14591, new_n14592, new_n14593_1,
    new_n14594, new_n14595, new_n14596, new_n14597, new_n14598, new_n14599,
    new_n14600, new_n14601, new_n14602, new_n14603_1, new_n14604,
    new_n14605, new_n14606, new_n14607, new_n14608, new_n14609, new_n14610,
    new_n14611, new_n14612, new_n14613, new_n14614, new_n14616, new_n14617,
    new_n14618, new_n14619, new_n14620, new_n14621, new_n14622, new_n14623,
    new_n14624, new_n14625, new_n14626, new_n14627, new_n14628, new_n14629,
    new_n14630, new_n14631, new_n14632, new_n14633_1, new_n14634,
    new_n14635, new_n14636_1, new_n14637, new_n14638, new_n14639,
    new_n14640, new_n14641, new_n14642, new_n14643, new_n14644, new_n14645,
    new_n14646, new_n14647, new_n14648, new_n14649, new_n14650, new_n14651,
    new_n14652, new_n14653, new_n14654, new_n14655, new_n14656, new_n14657,
    new_n14658, new_n14659, new_n14660, new_n14661, new_n14662, new_n14663,
    new_n14664, new_n14665, new_n14666, new_n14667, new_n14668, new_n14669,
    new_n14670, new_n14671, new_n14672, new_n14673, new_n14674, new_n14675,
    new_n14676, new_n14677, new_n14678, new_n14679, new_n14680_1,
    new_n14681, new_n14682, new_n14683, new_n14684_1, new_n14685,
    new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692_1, new_n14693, new_n14694, new_n14695, new_n14696,
    new_n14697, new_n14698, new_n14699, new_n14700, new_n14701_1,
    new_n14702_1, new_n14703, new_n14704_1, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730,
    new_n14731, new_n14732, new_n14733, new_n14734_1, new_n14735,
    new_n14736, new_n14737, new_n14738, new_n14739, new_n14740, new_n14741,
    new_n14742, new_n14743, new_n14744, new_n14745, new_n14746_1,
    new_n14747, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754,
    new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760,
    new_n14761, new_n14762, new_n14763_1, new_n14764, new_n14765,
    new_n14766, new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772_1, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790_1, new_n14791, new_n14792, new_n14793,
    new_n14794, new_n14795, new_n14796, new_n14797, new_n14798,
    new_n14801_1, new_n14802, new_n14803, new_n14804, new_n14805,
    new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819_1, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826_1, new_n14827_1,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839_1, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14848,
    new_n14849_1, new_n14850, new_n14851, new_n14852, new_n14853,
    new_n14854, new_n14855, new_n14856, new_n14857, new_n14858, new_n14859,
    new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865,
    new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871,
    new_n14872, new_n14873, new_n14874, new_n14875, new_n14876, new_n14877,
    new_n14878, new_n14879, new_n14880, new_n14881, new_n14882, new_n14883,
    new_n14884, new_n14885, new_n14886, new_n14887, new_n14888, new_n14889,
    new_n14890, new_n14891_1, new_n14892, new_n14893, new_n14894,
    new_n14895, new_n14896, new_n14897, new_n14898, new_n14899_1,
    new_n14900, new_n14901, new_n14902, new_n14903, new_n14904, new_n14905,
    new_n14906, new_n14907, new_n14908, new_n14909, new_n14910, new_n14911,
    new_n14912, new_n14913, new_n14914, new_n14915, new_n14916, new_n14917,
    new_n14918, new_n14919, new_n14920, new_n14921, new_n14922, new_n14923,
    new_n14924, new_n14925, new_n14926, new_n14927, new_n14928, new_n14929,
    new_n14930, new_n14931_1, new_n14932, new_n14933, new_n14934,
    new_n14935, new_n14936, new_n14937, new_n14938, new_n14939, new_n14940,
    new_n14941, new_n14942, new_n14943, new_n14944_1, new_n14945,
    new_n14946, new_n14947, new_n14948, new_n14949, new_n14950, new_n14952,
    new_n14953, new_n14954_1, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977_1, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14985, new_n14986, new_n14987,
    new_n14988, new_n14989_1, new_n14990, new_n14991, new_n14992,
    new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998,
    new_n14999, new_n15000, new_n15001, new_n15002_1, new_n15003,
    new_n15004_1, new_n15005, new_n15006, new_n15007, new_n15008,
    new_n15009, new_n15010, new_n15011_1, new_n15012, new_n15013,
    new_n15014, new_n15015, new_n15016, new_n15017, new_n15018,
    new_n15019_1, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031_1, new_n15032, new_n15033_1, new_n15034,
    new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040,
    new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046,
    new_n15047, new_n15048, new_n15049, new_n15050, new_n15051,
    new_n15052_1, new_n15053_1, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077_1, new_n15078, new_n15079,
    new_n15080, new_n15081, new_n15082_1, new_n15083, new_n15084,
    new_n15085, new_n15086, new_n15087, new_n15088, new_n15089, new_n15090,
    new_n15091, new_n15092, new_n15093, new_n15094_1, new_n15095,
    new_n15096, new_n15097, new_n15098, new_n15099, new_n15100, new_n15101,
    new_n15102, new_n15103, new_n15104, new_n15105, new_n15106, new_n15107,
    new_n15108, new_n15109, new_n15110, new_n15111, new_n15112, new_n15113,
    new_n15114, new_n15115, new_n15116, new_n15117, new_n15118_1,
    new_n15119, new_n15120, new_n15121, new_n15122, new_n15123, new_n15124,
    new_n15125, new_n15126, new_n15127, new_n15128_1, new_n15129,
    new_n15130, new_n15131, new_n15132, new_n15133, new_n15134, new_n15135,
    new_n15136, new_n15137, new_n15138, new_n15139_1, new_n15140,
    new_n15141, new_n15142, new_n15143, new_n15144, new_n15145_1,
    new_n15146_1, new_n15147, new_n15148, new_n15149, new_n15150,
    new_n15151, new_n15152, new_n15153, new_n15154, new_n15155, new_n15156,
    new_n15157, new_n15158, new_n15159, new_n15160, new_n15161, new_n15162,
    new_n15163, new_n15164, new_n15165_1, new_n15166, new_n15167_1,
    new_n15168, new_n15169, new_n15170, new_n15171, new_n15172, new_n15173,
    new_n15174, new_n15175, new_n15176_1, new_n15177, new_n15178,
    new_n15179, new_n15180_1, new_n15181, new_n15182_1, new_n15183,
    new_n15184, new_n15185, new_n15186, new_n15187, new_n15188, new_n15189,
    new_n15190, new_n15191, new_n15192, new_n15193, new_n15194, new_n15195,
    new_n15196, new_n15197, new_n15198, new_n15199, new_n15200, new_n15202,
    new_n15203, new_n15204, new_n15205_1, new_n15206, new_n15207,
    new_n15208, new_n15209, new_n15210, new_n15211, new_n15212, new_n15213,
    new_n15214, new_n15215, new_n15216, new_n15217, new_n15218, new_n15219,
    new_n15220, new_n15221, new_n15222, new_n15223, new_n15224, new_n15225,
    new_n15226, new_n15227, new_n15228, new_n15229, new_n15230_1,
    new_n15231, new_n15232, new_n15233, new_n15234, new_n15235, new_n15236,
    new_n15237, new_n15238, new_n15239, new_n15240, new_n15241_1,
    new_n15242, new_n15243, new_n15244, new_n15245, new_n15246, new_n15247,
    new_n15248, new_n15249, new_n15250, new_n15251, new_n15252, new_n15253,
    new_n15254, new_n15255_1, new_n15256, new_n15257, new_n15258_1,
    new_n15259, new_n15260, new_n15261, new_n15262, new_n15263, new_n15264,
    new_n15265, new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271_1, new_n15272, new_n15273, new_n15274, new_n15275_1,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289_1, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300_1, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307_1, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327_1, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332_1, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342,
    new_n15343, new_n15344, new_n15345_1, new_n15346, new_n15347,
    new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353_1, new_n15354, new_n15355, new_n15356, new_n15357,
    new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363,
    new_n15364, new_n15365, new_n15366_1, new_n15367, new_n15368,
    new_n15369, new_n15370, new_n15371, new_n15373, new_n15374, new_n15375,
    new_n15376, new_n15377, new_n15378_1, new_n15379, new_n15380,
    new_n15381, new_n15382_1, new_n15383, new_n15384, new_n15385,
    new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391,
    new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397,
    new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403,
    new_n15404, new_n15405, new_n15406, new_n15407_1, new_n15408,
    new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414,
    new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420,
    new_n15421, new_n15422, new_n15423, new_n15424_1, new_n15425,
    new_n15426, new_n15427, new_n15428_1, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435_1,
    new_n15436, new_n15437, new_n15438_1, new_n15439, new_n15440,
    new_n15441, new_n15442, new_n15443, new_n15444, new_n15445, new_n15446,
    new_n15447, new_n15448, new_n15449, new_n15450, new_n15451, new_n15452,
    new_n15453, new_n15454, new_n15455, new_n15456, new_n15457, new_n15458,
    new_n15459, new_n15460, new_n15461, new_n15462, new_n15463, new_n15464,
    new_n15465_1, new_n15466, new_n15467_1, new_n15468, new_n15469,
    new_n15470_1, new_n15471, new_n15472, new_n15473, new_n15474,
    new_n15475, new_n15476, new_n15477_1, new_n15478, new_n15479,
    new_n15480, new_n15481_1, new_n15482, new_n15483, new_n15484,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489,
    new_n15490_1, new_n15491, new_n15492, new_n15493, new_n15494,
    new_n15495, new_n15496_1, new_n15497, new_n15498, new_n15499,
    new_n15500, new_n15501_1, new_n15502, new_n15503, new_n15504,
    new_n15505, new_n15506_1, new_n15507, new_n15508_1, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15526, new_n15527, new_n15528,
    new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534,
    new_n15535, new_n15536, new_n15537, new_n15538, new_n15539_1,
    new_n15540, new_n15541, new_n15542, new_n15543, new_n15544, new_n15545,
    new_n15546_1, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555_1,
    new_n15556, new_n15557, new_n15558_1, new_n15559_1, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570_1, new_n15571,
    new_n15572, new_n15573_1, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588_1, new_n15589, new_n15590_1, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598_1, new_n15599, new_n15600, new_n15601, new_n15602_1,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613,
    new_n15614_1, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635,
    new_n15636_1, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15645, new_n15646, new_n15647,
    new_n15648, new_n15649, new_n15650, new_n15651, new_n15652_1,
    new_n15653, new_n15654, new_n15655, new_n15656, new_n15657, new_n15658,
    new_n15659, new_n15660, new_n15661, new_n15662_1, new_n15663,
    new_n15664, new_n15665, new_n15666, new_n15667, new_n15668, new_n15669,
    new_n15670, new_n15671, new_n15672, new_n15673, new_n15674, new_n15675,
    new_n15676, new_n15677, new_n15678, new_n15679, new_n15680, new_n15681,
    new_n15682, new_n15683, new_n15684, new_n15685, new_n15686, new_n15687,
    new_n15688, new_n15689, new_n15690, new_n15691, new_n15692, new_n15693,
    new_n15694, new_n15695, new_n15696, new_n15697, new_n15698, new_n15699,
    new_n15700, new_n15701, new_n15702, new_n15703, new_n15704, new_n15705,
    new_n15706, new_n15707, new_n15708, new_n15711, new_n15712, new_n15713,
    new_n15714, new_n15715, new_n15716_1, new_n15717, new_n15718,
    new_n15719, new_n15720, new_n15721, new_n15722, new_n15723, new_n15724,
    new_n15725, new_n15726, new_n15727, new_n15728, new_n15729, new_n15730,
    new_n15731, new_n15732, new_n15733, new_n15734, new_n15735, new_n15736,
    new_n15737, new_n15738, new_n15739, new_n15740, new_n15741, new_n15742,
    new_n15743_1, new_n15744, new_n15745, new_n15746, new_n15747,
    new_n15748, new_n15749_1, new_n15750, new_n15751, new_n15752,
    new_n15753, new_n15754, new_n15755, new_n15756, new_n15757, new_n15758,
    new_n15759, new_n15760, new_n15761_1, new_n15762_1, new_n15763,
    new_n15764, new_n15765, new_n15766_1, new_n15767, new_n15768,
    new_n15769, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774,
    new_n15775, new_n15776, new_n15777, new_n15778, new_n15779,
    new_n15780_1, new_n15781, new_n15782, new_n15783, new_n15784,
    new_n15785, new_n15786, new_n15787, new_n15788, new_n15789, new_n15790,
    new_n15791, new_n15792, new_n15793_1, new_n15794, new_n15795,
    new_n15796, new_n15797, new_n15798, new_n15799, new_n15800, new_n15801,
    new_n15802, new_n15803, new_n15804, new_n15805, new_n15806, new_n15807,
    new_n15808, new_n15809, new_n15810, new_n15811, new_n15812_1,
    new_n15813, new_n15814, new_n15815_1, new_n15816_1, new_n15817,
    new_n15818, new_n15819, new_n15820, new_n15821, new_n15822, new_n15823,
    new_n15824, new_n15825, new_n15826, new_n15827, new_n15828, new_n15829,
    new_n15830, new_n15831_1, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15845,
    new_n15846_1, new_n15847, new_n15848, new_n15849, new_n15850,
    new_n15851, new_n15852, new_n15853, new_n15854, new_n15855, new_n15856,
    new_n15858, new_n15859_1, new_n15860, new_n15861, new_n15862,
    new_n15863, new_n15864, new_n15865, new_n15866, new_n15867, new_n15868,
    new_n15869_1, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884_1,
    new_n15885_1, new_n15886, new_n15887, new_n15888, new_n15889_1,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917_1, new_n15918_1,
    new_n15919, new_n15920, new_n15921, new_n15922_1, new_n15923,
    new_n15924, new_n15925, new_n15926, new_n15927, new_n15928, new_n15929,
    new_n15930, new_n15931, new_n15932, new_n15933, new_n15934, new_n15935,
    new_n15936_1, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947_1, new_n15948, new_n15949, new_n15950, new_n15951,
    new_n15952, new_n15953, new_n15954, new_n15955, new_n15956_1,
    new_n15957, new_n15958_1, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967_1, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15979_1, new_n15982, new_n15983,
    new_n15984, new_n15986_1, new_n15987, new_n15988, new_n15989,
    new_n15990, new_n15991, new_n15992, new_n15993, new_n15994, new_n15995,
    new_n15996, new_n15997, new_n15998, new_n15999, new_n16000, new_n16001,
    new_n16002, new_n16003, new_n16004, new_n16005, new_n16006, new_n16007,
    new_n16008, new_n16009, new_n16010, new_n16011, new_n16012,
    new_n16013_1, new_n16014, new_n16015, new_n16016, new_n16017,
    new_n16018, new_n16019, new_n16022, new_n16023, new_n16024, new_n16025,
    new_n16026, new_n16027, new_n16028, new_n16029_1, new_n16030,
    new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036,
    new_n16037, new_n16038, new_n16039, new_n16040, new_n16041, new_n16042,
    new_n16043, new_n16044, new_n16045, new_n16046, new_n16047, new_n16048,
    new_n16049, new_n16050, new_n16051, new_n16052, new_n16053, new_n16054,
    new_n16055, new_n16056, new_n16057, new_n16058, new_n16059,
    new_n16060_1, new_n16061, new_n16062_1, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068_1, new_n16069,
    new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075,
    new_n16076, new_n16077, new_n16078, new_n16079, new_n16080_1,
    new_n16081, new_n16082, new_n16083, new_n16084, new_n16085, new_n16086,
    new_n16087, new_n16088, new_n16089, new_n16090, new_n16091, new_n16092,
    new_n16098_1, new_n16099, new_n16100, new_n16101, new_n16102,
    new_n16103, new_n16104, new_n16105, new_n16106, new_n16107, new_n16108,
    new_n16109, new_n16110_1, new_n16111, new_n16112, new_n16113,
    new_n16114, new_n16115, new_n16116, new_n16117, new_n16118, new_n16119,
    new_n16120, new_n16121, new_n16122, new_n16123, new_n16124, new_n16125,
    new_n16126, new_n16127, new_n16128, new_n16129, new_n16130, new_n16131,
    new_n16132, new_n16133, new_n16134, new_n16135, new_n16136, new_n16137,
    new_n16138, new_n16139, new_n16140, new_n16141, new_n16142_1,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158_1, new_n16159,
    new_n16160, new_n16161, new_n16162, new_n16163, new_n16164, new_n16165,
    new_n16166, new_n16167_1, new_n16168, new_n16169, new_n16170,
    new_n16171, new_n16172, new_n16173, new_n16174, new_n16175, new_n16176,
    new_n16177, new_n16178, new_n16179, new_n16180, new_n16181, new_n16182,
    new_n16183, new_n16184, new_n16185_1, new_n16186, new_n16187,
    new_n16188, new_n16189, new_n16190, new_n16191, new_n16192, new_n16193,
    new_n16194, new_n16195, new_n16196_1, new_n16197, new_n16198,
    new_n16199, new_n16200, new_n16201, new_n16202, new_n16203, new_n16204,
    new_n16205, new_n16206_1, new_n16207, new_n16208, new_n16209,
    new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215_1, new_n16216, new_n16217_1, new_n16218_1, new_n16219_1,
    new_n16220, new_n16221, new_n16222, new_n16223_1, new_n16224,
    new_n16225, new_n16226, new_n16227, new_n16228, new_n16229,
    new_n16230_1, new_n16231, new_n16232, new_n16233, new_n16234,
    new_n16237, new_n16238, new_n16239, new_n16240, new_n16241, new_n16242,
    new_n16243_1, new_n16244, new_n16245, new_n16246, new_n16247_1,
    new_n16248, new_n16249, new_n16250, new_n16251, new_n16252, new_n16253,
    new_n16254, new_n16255, new_n16256, new_n16257, new_n16258, new_n16259,
    new_n16260, new_n16261, new_n16262, new_n16263, new_n16264, new_n16265,
    new_n16266, new_n16267, new_n16268, new_n16269, new_n16270, new_n16271,
    new_n16272, new_n16273, new_n16274, new_n16275_1, new_n16276,
    new_n16277, new_n16278, new_n16279_1, new_n16280, new_n16281,
    new_n16282, new_n16283, new_n16284, new_n16285, new_n16286, new_n16287,
    new_n16288, new_n16289, new_n16290, new_n16291, new_n16292, new_n16293,
    new_n16294, new_n16295, new_n16296, new_n16297, new_n16298, new_n16299,
    new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305,
    new_n16306, new_n16308, new_n16309, new_n16310, new_n16311, new_n16312,
    new_n16313, new_n16314, new_n16315, new_n16316, new_n16317, new_n16318,
    new_n16319, new_n16320, new_n16321, new_n16322_1, new_n16323,
    new_n16324, new_n16325, new_n16326, new_n16327_1, new_n16328,
    new_n16329, new_n16330, new_n16331, new_n16332, new_n16333, new_n16334,
    new_n16335, new_n16336, new_n16337, new_n16338, new_n16339, new_n16342,
    new_n16343, new_n16344, new_n16345, new_n16346, new_n16347, new_n16348,
    new_n16349, new_n16350_1, new_n16351, new_n16352, new_n16353,
    new_n16354, new_n16355, new_n16356, new_n16357, new_n16358, new_n16359,
    new_n16360, new_n16361, new_n16362, new_n16363, new_n16364, new_n16365,
    new_n16366, new_n16367_1, new_n16368, new_n16369, new_n16370,
    new_n16371, new_n16372, new_n16373, new_n16374, new_n16375,
    new_n16376_1, new_n16377, new_n16378, new_n16379_1, new_n16380,
    new_n16381, new_n16382, new_n16383, new_n16384, new_n16385, new_n16386,
    new_n16387, new_n16389, new_n16390, new_n16391, new_n16392, new_n16393,
    new_n16394, new_n16395, new_n16396_1, new_n16397, new_n16398_1,
    new_n16399, new_n16400, new_n16401, new_n16402, new_n16403, new_n16404,
    new_n16405, new_n16406_1, new_n16407_1, new_n16408, new_n16409,
    new_n16410, new_n16411, new_n16412, new_n16413, new_n16414, new_n16415,
    new_n16416, new_n16417, new_n16418, new_n16419_1, new_n16420,
    new_n16421, new_n16422, new_n16423, new_n16424_1, new_n16425,
    new_n16426, new_n16427, new_n16428_1, new_n16429, new_n16430,
    new_n16431, new_n16432, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439_1, new_n16440_1, new_n16441, new_n16442,
    new_n16443, new_n16444, new_n16445_1, new_n16446, new_n16447,
    new_n16448, new_n16449, new_n16450, new_n16451, new_n16452, new_n16453,
    new_n16454, new_n16455, new_n16456, new_n16457, new_n16458, new_n16459,
    new_n16460_1, new_n16461, new_n16462, new_n16463, new_n16464,
    new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470,
    new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476_1, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481_1, new_n16482_1, new_n16483, new_n16484, new_n16485,
    new_n16486, new_n16487, new_n16488, new_n16489, new_n16490, new_n16491,
    new_n16492, new_n16493_1, new_n16494, new_n16495, new_n16496,
    new_n16497, new_n16498, new_n16499, new_n16500, new_n16501,
    new_n16502_1, new_n16503, new_n16504, new_n16505, new_n16506_1,
    new_n16507_1, new_n16508, new_n16509, new_n16510, new_n16511,
    new_n16512, new_n16513, new_n16514, new_n16515, new_n16516_1,
    new_n16517_1, new_n16518, new_n16519, new_n16520, new_n16521_1,
    new_n16522, new_n16523, new_n16524_1, new_n16525, new_n16526,
    new_n16527_1, new_n16528, new_n16529, new_n16530, new_n16531,
    new_n16532, new_n16533, new_n16534, new_n16535, new_n16536, new_n16537,
    new_n16538, new_n16539, new_n16540, new_n16541, new_n16542, new_n16543,
    new_n16544_1, new_n16545, new_n16546, new_n16547, new_n16548,
    new_n16549, new_n16550, new_n16551, new_n16552, new_n16553,
    new_n16554_1, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583_1, new_n16584_1, new_n16585, new_n16586, new_n16587,
    new_n16588, new_n16589_1, new_n16590, new_n16591, new_n16592,
    new_n16593, new_n16594, new_n16595, new_n16596_1, new_n16597,
    new_n16598, new_n16599, new_n16600, new_n16601, new_n16602, new_n16603,
    new_n16604, new_n16605, new_n16606, new_n16607, new_n16608_1,
    new_n16609, new_n16610, new_n16611, new_n16612, new_n16613, new_n16614,
    new_n16615, new_n16616, new_n16617_1, new_n16618, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16632, new_n16633, new_n16634, new_n16635,
    new_n16636, new_n16637, new_n16638, new_n16639, new_n16640_1,
    new_n16641, new_n16642, new_n16643, new_n16644, new_n16645, new_n16646,
    new_n16647, new_n16650, new_n16651, new_n16652, new_n16653, new_n16654,
    new_n16655, new_n16656_1, new_n16657, new_n16658, new_n16659,
    new_n16660, new_n16661, new_n16662, new_n16663, new_n16664, new_n16665,
    new_n16666, new_n16667, new_n16668, new_n16669, new_n16670, new_n16671,
    new_n16672, new_n16673, new_n16674_1, new_n16675, new_n16676,
    new_n16677, new_n16678, new_n16679, new_n16680, new_n16681,
    new_n16682_1, new_n16683, new_n16684_1, new_n16685, new_n16686,
    new_n16687, new_n16688_1, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722_1, new_n16723, new_n16724, new_n16725, new_n16726,
    new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732,
    new_n16733_1, new_n16734, new_n16735, new_n16736, new_n16737,
    new_n16738, new_n16739, new_n16740, new_n16741, new_n16742,
    new_n16743_1, new_n16744, new_n16745, new_n16746, new_n16747,
    new_n16748, new_n16749, new_n16750, new_n16751, new_n16752, new_n16753,
    new_n16754, new_n16755, new_n16756, new_n16757, new_n16758, new_n16759,
    new_n16762, new_n16763, new_n16764, new_n16765, new_n16766, new_n16767,
    new_n16768, new_n16769, new_n16770, new_n16771, new_n16772, new_n16773,
    new_n16774, new_n16775, new_n16776, new_n16777, new_n16778, new_n16779,
    new_n16780, new_n16781, new_n16782, new_n16783, new_n16784, new_n16785,
    new_n16786, new_n16787, new_n16788, new_n16789, new_n16790, new_n16792,
    new_n16793, new_n16794, new_n16795, new_n16796, new_n16797,
    new_n16798_1, new_n16799, new_n16800, new_n16801, new_n16802,
    new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812_1, new_n16815,
    new_n16816, new_n16817, new_n16818_1, new_n16819, new_n16820,
    new_n16821, new_n16822, new_n16823, new_n16824_1, new_n16825,
    new_n16826, new_n16827, new_n16828, new_n16829, new_n16830, new_n16831,
    new_n16832, new_n16833, new_n16834_1, new_n16835, new_n16836,
    new_n16837_1, new_n16838, new_n16839, new_n16840, new_n16841_1,
    new_n16842, new_n16843, new_n16844, new_n16845, new_n16846, new_n16847,
    new_n16848, new_n16849, new_n16850, new_n16851, new_n16852, new_n16853,
    new_n16854, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860,
    new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866,
    new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872,
    new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878,
    new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885_1, new_n16886, new_n16887, new_n16888, new_n16889,
    new_n16890, new_n16891, new_n16892, new_n16893, new_n16894, new_n16895,
    new_n16896, new_n16897, new_n16898, new_n16899, new_n16900, new_n16901,
    new_n16902, new_n16903, new_n16904, new_n16905_1, new_n16906,
    new_n16907, new_n16908, new_n16909, new_n16910, new_n16911_1,
    new_n16912, new_n16913, new_n16914, new_n16915, new_n16916, new_n16917,
    new_n16918, new_n16919, new_n16920, new_n16921, new_n16922, new_n16923,
    new_n16924, new_n16925, new_n16926, new_n16927, new_n16928, new_n16929,
    new_n16930, new_n16931, new_n16932, new_n16933, new_n16934, new_n16935,
    new_n16936, new_n16937, new_n16938, new_n16939, new_n16940, new_n16941,
    new_n16942, new_n16943, new_n16944, new_n16945, new_n16946, new_n16947,
    new_n16948, new_n16949, new_n16950, new_n16951_1, new_n16952,
    new_n16953, new_n16954_1, new_n16955, new_n16956, new_n16957,
    new_n16958, new_n16959, new_n16960, new_n16961, new_n16962, new_n16963,
    new_n16964, new_n16965, new_n16966, new_n16967, new_n16968_1,
    new_n16969, new_n16970, new_n16971_1, new_n16972, new_n16973,
    new_n16974, new_n16975, new_n16976, new_n16977, new_n16978, new_n16979,
    new_n16980, new_n16981, new_n16982, new_n16983, new_n16984, new_n16985,
    new_n16986, new_n16987, new_n16988_1, new_n16989_1, new_n16990,
    new_n16991, new_n16992, new_n16993, new_n16994_1, new_n16995,
    new_n16996, new_n16997, new_n16998, new_n16999, new_n17000, new_n17001,
    new_n17002, new_n17003, new_n17004, new_n17005, new_n17006_1,
    new_n17007, new_n17008, new_n17009, new_n17010, new_n17011, new_n17012,
    new_n17013, new_n17014, new_n17015, new_n17016, new_n17017, new_n17018,
    new_n17019, new_n17020, new_n17021, new_n17022, new_n17023, new_n17024,
    new_n17025, new_n17026, new_n17027, new_n17028, new_n17029, new_n17030,
    new_n17031, new_n17032, new_n17033, new_n17034, new_n17035_1,
    new_n17036, new_n17037_1, new_n17038, new_n17039, new_n17040,
    new_n17041, new_n17042, new_n17043, new_n17044, new_n17045, new_n17046,
    new_n17047, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052,
    new_n17053, new_n17054, new_n17055, new_n17056, new_n17057, new_n17059,
    new_n17060, new_n17061, new_n17062, new_n17063, new_n17064, new_n17065,
    new_n17066, new_n17067, new_n17068_1, new_n17069_1, new_n17070_1,
    new_n17071, new_n17072, new_n17073, new_n17074, new_n17075_1,
    new_n17076, new_n17077_1, new_n17078, new_n17079, new_n17080,
    new_n17081, new_n17082, new_n17083, new_n17084_1, new_n17085,
    new_n17086, new_n17087, new_n17088, new_n17089, new_n17090_1,
    new_n17091, new_n17092, new_n17093, new_n17094, new_n17095_1,
    new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101,
    new_n17102, new_n17103, new_n17104_1, new_n17105, new_n17106_1,
    new_n17107, new_n17108, new_n17109, new_n17110, new_n17111, new_n17112,
    new_n17113, new_n17114, new_n17115, new_n17116, new_n17117, new_n17118,
    new_n17119_1, new_n17120, new_n17121, new_n17122, new_n17123,
    new_n17124, new_n17125, new_n17126, new_n17127, new_n17128, new_n17129,
    new_n17130_1, new_n17131, new_n17132, new_n17133, new_n17134,
    new_n17135, new_n17136, new_n17137, new_n17138_1, new_n17139,
    new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17147, new_n17148, new_n17149, new_n17150, new_n17151,
    new_n17152, new_n17153, new_n17154, new_n17155, new_n17156, new_n17157,
    new_n17158, new_n17159, new_n17160, new_n17161, new_n17162,
    new_n17163_1, new_n17164, new_n17165, new_n17166, new_n17169,
    new_n17170, new_n17171, new_n17172, new_n17173, new_n17174, new_n17175,
    new_n17176, new_n17177, new_n17178, new_n17179, new_n17180, new_n17181,
    new_n17182, new_n17183, new_n17184, new_n17185, new_n17186, new_n17187,
    new_n17188, new_n17189, new_n17190, new_n17191, new_n17192, new_n17193,
    new_n17194, new_n17195, new_n17196, new_n17197, new_n17198, new_n17199,
    new_n17200, new_n17201, new_n17202_1, new_n17203, new_n17204,
    new_n17205, new_n17206, new_n17207, new_n17208, new_n17209, new_n17210,
    new_n17211, new_n17212, new_n17213, new_n17214, new_n17215, new_n17216,
    new_n17217, new_n17218, new_n17219_1, new_n17220, new_n17221,
    new_n17222, new_n17223, new_n17224, new_n17225, new_n17226, new_n17227,
    new_n17228, new_n17229, new_n17230, new_n17231, new_n17232_1,
    new_n17233, new_n17234, new_n17235, new_n17236_1, new_n17237,
    new_n17238, new_n17239, new_n17240, new_n17241, new_n17242,
    new_n17243_1, new_n17244, new_n17245, new_n17246, new_n17247,
    new_n17248, new_n17249, new_n17250_1, new_n17251_1, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263_1,
    new_n17264, new_n17265, new_n17266, new_n17267, new_n17268, new_n17269,
    new_n17270, new_n17271, new_n17272, new_n17273, new_n17274, new_n17275,
    new_n17276, new_n17277, new_n17278, new_n17279, new_n17281, new_n17282,
    new_n17283, new_n17284, new_n17285_1, new_n17286, new_n17287,
    new_n17288, new_n17289, new_n17290, new_n17291, new_n17292, new_n17293,
    new_n17294, new_n17295, new_n17296, new_n17297, new_n17298, new_n17299,
    new_n17300, new_n17301, new_n17302_1, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320_1, new_n17321,
    new_n17322, new_n17323, new_n17324, new_n17325, new_n17326, new_n17327,
    new_n17328, new_n17329, new_n17330, new_n17331, new_n17332, new_n17333,
    new_n17334, new_n17335, new_n17336, new_n17337_1, new_n17338,
    new_n17340, new_n17341, new_n17342, new_n17343, new_n17344_1,
    new_n17345, new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351_1, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359_1, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17368,
    new_n17369, new_n17370, new_n17371, new_n17372, new_n17373, new_n17374,
    new_n17375, new_n17376, new_n17377, new_n17378, new_n17379, new_n17380,
    new_n17381, new_n17382, new_n17383, new_n17384, new_n17385, new_n17386,
    new_n17387_1, new_n17388, new_n17389, new_n17390, new_n17391_1,
    new_n17392_1, new_n17393, new_n17394, new_n17395, new_n17396,
    new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402,
    new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408,
    new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414,
    new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420,
    new_n17421_1, new_n17422, new_n17423, new_n17424, new_n17425,
    new_n17426, new_n17427, new_n17428, new_n17429, new_n17430, new_n17431,
    new_n17432_1, new_n17433, new_n17434, new_n17435, new_n17436_1,
    new_n17437, new_n17438, new_n17439, new_n17440_1, new_n17441,
    new_n17442, new_n17443, new_n17444, new_n17445, new_n17446, new_n17447,
    new_n17448, new_n17449, new_n17450_1, new_n17451, new_n17452,
    new_n17453, new_n17454, new_n17455, new_n17456, new_n17457,
    new_n17458_1, new_n17462, new_n17463, new_n17464, new_n17465,
    new_n17466_1, new_n17467, new_n17468, new_n17469, new_n17470,
    new_n17471, new_n17472, new_n17473, new_n17474, new_n17478, new_n17479,
    new_n17480, new_n17481, new_n17482, new_n17483, new_n17484, new_n17485,
    new_n17486, new_n17487, new_n17488, new_n17489, new_n17490, new_n17491,
    new_n17492, new_n17493_1, new_n17494, new_n17495, new_n17496,
    new_n17497, new_n17498, new_n17499, new_n17500_1, new_n17501,
    new_n17502, new_n17503, new_n17504, new_n17505, new_n17506, new_n17507,
    new_n17508, new_n17511, new_n17512, new_n17513, new_n17514, new_n17515,
    new_n17516, new_n17517, new_n17518, new_n17519, new_n17520, new_n17521,
    new_n17522, new_n17523, new_n17524_1, new_n17525, new_n17526,
    new_n17527, new_n17528, new_n17529_1, new_n17530, new_n17531,
    new_n17532, new_n17533, new_n17534, new_n17535, new_n17536, new_n17537,
    new_n17538, new_n17539, new_n17540, new_n17541, new_n17542, new_n17543,
    new_n17544, new_n17545, new_n17546, new_n17547, new_n17548, new_n17549,
    new_n17550, new_n17551, new_n17552, new_n17553, new_n17554, new_n17555,
    new_n17556, new_n17557_1, new_n17558, new_n17559, new_n17560,
    new_n17561, new_n17562, new_n17563, new_n17564, new_n17565, new_n17566,
    new_n17567, new_n17568, new_n17569, new_n17570, new_n17571, new_n17572,
    new_n17573, new_n17574, new_n17575, new_n17576, new_n17577, new_n17578,
    new_n17579, new_n17580, new_n17581, new_n17582, new_n17583_1,
    new_n17584, new_n17585, new_n17586, new_n17587, new_n17588, new_n17589,
    new_n17590, new_n17591, new_n17592_1, new_n17593, new_n17594,
    new_n17595, new_n17596, new_n17597, new_n17598, new_n17599, new_n17600,
    new_n17601, new_n17602, new_n17603, new_n17604, new_n17605, new_n17606,
    new_n17607, new_n17608, new_n17609, new_n17610, new_n17611, new_n17612,
    new_n17613, new_n17614, new_n17615, new_n17616, new_n17617, new_n17618,
    new_n17619, new_n17620, new_n17624, new_n17625, new_n17626, new_n17627,
    new_n17628, new_n17629, new_n17630, new_n17631, new_n17632, new_n17633,
    new_n17634, new_n17635, new_n17636, new_n17637, new_n17638_1,
    new_n17639, new_n17640, new_n17641, new_n17642, new_n17643, new_n17644,
    new_n17645, new_n17646, new_n17647, new_n17648, new_n17649, new_n17650,
    new_n17651, new_n17652, new_n17653, new_n17654, new_n17655, new_n17656,
    new_n17657, new_n17658, new_n17659, new_n17660, new_n17661, new_n17662,
    new_n17663, new_n17664_1, new_n17665, new_n17666, new_n17667,
    new_n17668, new_n17669, new_n17670, new_n17671, new_n17672, new_n17673,
    new_n17674, new_n17675, new_n17676, new_n17677, new_n17678, new_n17679,
    new_n17680, new_n17681, new_n17682, new_n17683, new_n17684, new_n17685,
    new_n17686, new_n17687_1, new_n17688, new_n17689, new_n17690,
    new_n17691, new_n17692, new_n17693, new_n17694, new_n17695, new_n17696,
    new_n17697, new_n17698, new_n17699, new_n17700, new_n17701, new_n17702,
    new_n17703, new_n17704, new_n17705, new_n17706, new_n17707, new_n17708,
    new_n17709, new_n17710, new_n17711, new_n17712, new_n17713, new_n17714,
    new_n17715, new_n17716, new_n17717, new_n17718, new_n17719, new_n17720,
    new_n17721_1, new_n17722, new_n17723, new_n17724, new_n17725,
    new_n17726, new_n17727, new_n17728, new_n17729, new_n17730, new_n17731,
    new_n17732, new_n17733, new_n17734, new_n17735_1, new_n17736,
    new_n17737, new_n17738_1, new_n17739, new_n17740, new_n17741,
    new_n17742, new_n17743, new_n17744, new_n17745, new_n17746_1,
    new_n17747, new_n17748, new_n17749_1, new_n17750, new_n17751,
    new_n17752, new_n17753, new_n17754, new_n17755, new_n17756, new_n17757,
    new_n17758, new_n17759, new_n17760, new_n17762, new_n17763, new_n17764,
    new_n17765, new_n17766, new_n17767, new_n17768, new_n17769, new_n17770,
    new_n17771, new_n17772, new_n17773, new_n17775, new_n17776, new_n17777,
    new_n17778, new_n17779, new_n17780, new_n17781, new_n17782, new_n17783,
    new_n17784_1, new_n17785, new_n17786, new_n17787, new_n17788,
    new_n17789, new_n17790, new_n17791, new_n17792, new_n17793, new_n17794,
    new_n17795, new_n17796, new_n17797, new_n17798, new_n17799, new_n17800,
    new_n17801, new_n17802, new_n17803, new_n17804, new_n17805, new_n17806,
    new_n17807, new_n17808, new_n17809, new_n17810, new_n17811, new_n17812,
    new_n17813, new_n17814, new_n17815, new_n17816, new_n17817, new_n17818,
    new_n17820_1, new_n17821, new_n17822, new_n17823, new_n17824,
    new_n17825, new_n17826, new_n17827, new_n17828, new_n17829, new_n17830,
    new_n17831, new_n17832, new_n17833, new_n17834, new_n17835, new_n17836,
    new_n17837, new_n17838, new_n17839, new_n17840, new_n17841, new_n17842,
    new_n17843, new_n17844, new_n17845, new_n17846, new_n17847, new_n17848,
    new_n17849, new_n17850, new_n17851, new_n17852, new_n17853, new_n17854,
    new_n17855_1, new_n17856, new_n17857, new_n17858, new_n17860,
    new_n17861, new_n17862, new_n17863, new_n17864, new_n17865, new_n17866,
    new_n17867, new_n17868, new_n17869, new_n17870, new_n17871, new_n17872,
    new_n17873, new_n17874, new_n17875, new_n17876, new_n17877_1,
    new_n17878, new_n17879, new_n17880, new_n17881, new_n17882, new_n17883,
    new_n17884, new_n17885, new_n17886, new_n17887, new_n17888, new_n17891,
    new_n17892, new_n17893, new_n17894, new_n17895, new_n17896, new_n17897,
    new_n17898, new_n17899, new_n17900, new_n17901, new_n17902, new_n17903,
    new_n17904, new_n17905, new_n17906, new_n17907, new_n17908, new_n17909,
    new_n17910, new_n17911_1, new_n17912_1, new_n17913, new_n17914,
    new_n17915, new_n17916, new_n17918, new_n17919, new_n17920, new_n17921,
    new_n17922, new_n17923, new_n17924, new_n17925, new_n17926,
    new_n17927_1, new_n17928, new_n17929, new_n17930, new_n17931_1,
    new_n17932, new_n17933, new_n17934, new_n17935, new_n17936, new_n17937,
    new_n17938, new_n17939, new_n17940, new_n17941, new_n17942, new_n17943,
    new_n17944, new_n17945, new_n17946, new_n17947, new_n17948_1,
    new_n17949, new_n17950, new_n17951, new_n17952, new_n17953,
    new_n17954_1, new_n17955, new_n17956_1, new_n17957, new_n17958,
    new_n17959_1, new_n17960, new_n17961, new_n17962, new_n17963_1,
    new_n17964, new_n17965, new_n17966, new_n17967, new_n17968_1,
    new_n17969, new_n17970, new_n17971, new_n17972, new_n17973, new_n17974,
    new_n17975, new_n17976_1, new_n17977, new_n17978, new_n17979,
    new_n17980, new_n17981, new_n17982, new_n17983, new_n17984, new_n17985,
    new_n17986, new_n17987, new_n17988, new_n17989, new_n17990, new_n17991,
    new_n17992, new_n17993, new_n17994, new_n17996, new_n17997,
    new_n17998_1, new_n17999, new_n18000, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020,
    new_n18021, new_n18022, new_n18023, new_n18024, new_n18025_1,
    new_n18026, new_n18027, new_n18028, new_n18029, new_n18030, new_n18031,
    new_n18032, new_n18033, new_n18034, new_n18035_1, new_n18036,
    new_n18037, new_n18038, new_n18039, new_n18040, new_n18041, new_n18042,
    new_n18043_1, new_n18044, new_n18045_1, new_n18046, new_n18047,
    new_n18048, new_n18049, new_n18050, new_n18051, new_n18052, new_n18053,
    new_n18054, new_n18055, new_n18056, new_n18057, new_n18058,
    new_n18059_1, new_n18060, new_n18061_1, new_n18062, new_n18063,
    new_n18064, new_n18065, new_n18066, new_n18067, new_n18068, new_n18069,
    new_n18070, new_n18071_1, new_n18072, new_n18073, new_n18074,
    new_n18075, new_n18076, new_n18077, new_n18078, new_n18079, new_n18080,
    new_n18081, new_n18082, new_n18083, new_n18084, new_n18085, new_n18086,
    new_n18087, new_n18088, new_n18089, new_n18090, new_n18091, new_n18092,
    new_n18093, new_n18094, new_n18095, new_n18096, new_n18097, new_n18098,
    new_n18099, new_n18100, new_n18101, new_n18102, new_n18103, new_n18104,
    new_n18105_1, new_n18106, new_n18107, new_n18108, new_n18109,
    new_n18110, new_n18111, new_n18112, new_n18113, new_n18114, new_n18115,
    new_n18116, new_n18117, new_n18118, new_n18119, new_n18120, new_n18121,
    new_n18122, new_n18123, new_n18124, new_n18125, new_n18126, new_n18127,
    new_n18128, new_n18129, new_n18130, new_n18131, new_n18132, new_n18133,
    new_n18134, new_n18135, new_n18136, new_n18137, new_n18138, new_n18139,
    new_n18140, new_n18141, new_n18142, new_n18143_1, new_n18144,
    new_n18145_1, new_n18146, new_n18147, new_n18148, new_n18149,
    new_n18150, new_n18151_1, new_n18152_1, new_n18153, new_n18154,
    new_n18155, new_n18156, new_n18157_1, new_n18158, new_n18159,
    new_n18160, new_n18161, new_n18162, new_n18163, new_n18164, new_n18165,
    new_n18166, new_n18167, new_n18168, new_n18169, new_n18170,
    new_n18171_1, new_n18172, new_n18174, new_n18175, new_n18176,
    new_n18177, new_n18178, new_n18179, new_n18180, new_n18181, new_n18182,
    new_n18183, new_n18184, new_n18185, new_n18186, new_n18187, new_n18188,
    new_n18189, new_n18190, new_n18191, new_n18194, new_n18195, new_n18196,
    new_n18197, new_n18198, new_n18199, new_n18200, new_n18201, new_n18202,
    new_n18203, new_n18204, new_n18205, new_n18206, new_n18207, new_n18212,
    new_n18213, new_n18214, new_n18215, new_n18216, new_n18217, new_n18218,
    new_n18219, new_n18220, new_n18221, new_n18222, new_n18223, new_n18224,
    new_n18231, new_n18232_1, new_n18233, new_n18234, new_n18235,
    new_n18236, new_n18237, new_n18238_1, new_n18239, new_n18240,
    new_n18241_1, new_n18242, new_n18243, new_n18244, new_n18245,
    new_n18246, new_n18247, new_n18248, new_n18249, new_n18250, new_n18251,
    new_n18252, new_n18253, new_n18254_1, new_n18255, new_n18256,
    new_n18257, new_n18258, new_n18259, new_n18260, new_n18261, new_n18262,
    new_n18263, new_n18264, new_n18265, new_n18266, new_n18267, new_n18268,
    new_n18269, new_n18270, new_n18271, new_n18272, new_n18273,
    new_n18274_1, new_n18275, new_n18276, new_n18277, new_n18278,
    new_n18279, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284,
    new_n18285, new_n18286, new_n18287, new_n18288_1, new_n18289,
    new_n18290_1, new_n18291, new_n18292, new_n18293, new_n18294,
    new_n18295_1, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301_1, new_n18302, new_n18303, new_n18304_1,
    new_n18305, new_n18306, new_n18307, new_n18308, new_n18309,
    new_n18310_1, new_n18311_1, new_n18312, new_n18313, new_n18314,
    new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320,
    new_n18321, new_n18322, new_n18323_1, new_n18324, new_n18325,
    new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332_1, new_n18334, new_n18335, new_n18336, new_n18337,
    new_n18338, new_n18339, new_n18340, new_n18341, new_n18342,
    new_n18343_1, new_n18344, new_n18345_1, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350_1, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362_1, new_n18363,
    new_n18364, new_n18365, new_n18366, new_n18367, new_n18368, new_n18369,
    new_n18370, new_n18371, new_n18372, new_n18373, new_n18374, new_n18375,
    new_n18376, new_n18377_1, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386,
    new_n18387, new_n18388, new_n18389, new_n18391, new_n18392, new_n18393,
    new_n18394, new_n18395, new_n18396, new_n18397, new_n18398, new_n18399,
    new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405_1, new_n18406, new_n18407, new_n18408, new_n18409_1,
    new_n18410, new_n18411, new_n18412, new_n18413, new_n18414_1,
    new_n18415, new_n18416, new_n18417, new_n18418_1, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437_1, new_n18438, new_n18439_1, new_n18440, new_n18441,
    new_n18442, new_n18443, new_n18444_1, new_n18445_1, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451,
    new_n18452_1, new_n18453, new_n18454, new_n18455, new_n18456,
    new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462,
    new_n18463, new_n18464, new_n18465, new_n18466, new_n18467_1,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482_1, new_n18483_1, new_n18484,
    new_n18485, new_n18486, new_n18487, new_n18488, new_n18489, new_n18490,
    new_n18491, new_n18492, new_n18493, new_n18494, new_n18495,
    new_n18496_1, new_n18497, new_n18498, new_n18499, new_n18500,
    new_n18501, new_n18502, new_n18503, new_n18504, new_n18505, new_n18506,
    new_n18507, new_n18508, new_n18509_1, new_n18510, new_n18511,
    new_n18512, new_n18513_1, new_n18514, new_n18515_1, new_n18516,
    new_n18517, new_n18518, new_n18519, new_n18520, new_n18521, new_n18522,
    new_n18523, new_n18524, new_n18525, new_n18526, new_n18527, new_n18528,
    new_n18529, new_n18530, new_n18531, new_n18532, new_n18533, new_n18534,
    new_n18535, new_n18536, new_n18537_1, new_n18538, new_n18539,
    new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545,
    new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551,
    new_n18552, new_n18553, new_n18555, new_n18556, new_n18557,
    new_n18558_1, new_n18559, new_n18560, new_n18561, new_n18562,
    new_n18563, new_n18564, new_n18565, new_n18566, new_n18567, new_n18568,
    new_n18569, new_n18570, new_n18571, new_n18572_1, new_n18573,
    new_n18574_1, new_n18575, new_n18576_1, new_n18577, new_n18578_1,
    new_n18579, new_n18580, new_n18581, new_n18582_1, new_n18583_1,
    new_n18584_1, new_n18585, new_n18586, new_n18587, new_n18588,
    new_n18589, new_n18590, new_n18591, new_n18592, new_n18593, new_n18594,
    new_n18595, new_n18596, new_n18597, new_n18598, new_n18599, new_n18600,
    new_n18601, new_n18602, new_n18603, new_n18604, new_n18605, new_n18608,
    new_n18609, new_n18610_1, new_n18611, new_n18612, new_n18613,
    new_n18614, new_n18615, new_n18616, new_n18617, new_n18618, new_n18619,
    new_n18620, new_n18621, new_n18624, new_n18625, new_n18626, new_n18627,
    new_n18628, new_n18629, new_n18630, new_n18631, new_n18632, new_n18633,
    new_n18637, new_n18638, new_n18639, new_n18640, new_n18641, new_n18642,
    new_n18643, new_n18644, new_n18645, new_n18646, new_n18647, new_n18648,
    new_n18649_1, new_n18650, new_n18651, new_n18652, new_n18653_1,
    new_n18654, new_n18655, new_n18656, new_n18657, new_n18658, new_n18659,
    new_n18660, new_n18661, new_n18662, new_n18663, new_n18664, new_n18665,
    new_n18666, new_n18667, new_n18668, new_n18669, new_n18670, new_n18671,
    new_n18672, new_n18673, new_n18674, new_n18675, new_n18676, new_n18677,
    new_n18678, new_n18679_1, new_n18680, new_n18681, new_n18682,
    new_n18683, new_n18686, new_n18687, new_n18688, new_n18689,
    new_n18690_1, new_n18691, new_n18692, new_n18693_1, new_n18694,
    new_n18695, new_n18696, new_n18697, new_n18698, new_n18699, new_n18700,
    new_n18701, new_n18702, new_n18703, new_n18704, new_n18705, new_n18706,
    new_n18707, new_n18708_1, new_n18709, new_n18710, new_n18711,
    new_n18712, new_n18713, new_n18714, new_n18715, new_n18716, new_n18717,
    new_n18718, new_n18719, new_n18720, new_n18721_1, new_n18722,
    new_n18723, new_n18724, new_n18725_1, new_n18726, new_n18727,
    new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733,
    new_n18734, new_n18735, new_n18736, new_n18737_1, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745_1, new_n18746, new_n18747, new_n18748, new_n18749,
    new_n18750, new_n18751_1, new_n18752, new_n18753, new_n18754,
    new_n18755, new_n18756, new_n18757, new_n18758, new_n18759, new_n18760,
    new_n18761, new_n18762, new_n18763, new_n18764, new_n18765, new_n18766,
    new_n18767, new_n18768, new_n18769, new_n18770, new_n18771, new_n18772,
    new_n18773, new_n18774, new_n18775, new_n18776, new_n18778, new_n18779,
    new_n18780_1, new_n18781, new_n18782_1, new_n18783, new_n18784,
    new_n18785, new_n18786, new_n18787, new_n18788, new_n18789, new_n18790,
    new_n18791, new_n18792, new_n18793, new_n18794, new_n18795, new_n18796,
    new_n18797, new_n18798, new_n18799, new_n18800, new_n18801,
    new_n18802_1, new_n18803, new_n18804, new_n18805, new_n18806,
    new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812,
    new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818,
    new_n18819, new_n18820, new_n18822, new_n18823, new_n18824, new_n18825,
    new_n18826, new_n18827, new_n18828, new_n18829, new_n18830_1,
    new_n18831_1, new_n18832, new_n18833, new_n18834, new_n18835,
    new_n18836, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841,
    new_n18842, new_n18843_1, new_n18844, new_n18845, new_n18846,
    new_n18847, new_n18848, new_n18849, new_n18850, new_n18851, new_n18852,
    new_n18853, new_n18854, new_n18855, new_n18856, new_n18857,
    new_n18858_1, new_n18859_1, new_n18860, new_n18861, new_n18862,
    new_n18863, new_n18864_1, new_n18865_1, new_n18866, new_n18867,
    new_n18868, new_n18869, new_n18870, new_n18871, new_n18872, new_n18873,
    new_n18874, new_n18875, new_n18876, new_n18877, new_n18878, new_n18879,
    new_n18880_1, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901_1, new_n18902, new_n18903, new_n18904, new_n18905,
    new_n18906, new_n18907_1, new_n18908, new_n18909, new_n18910,
    new_n18911, new_n18912, new_n18913, new_n18914, new_n18915, new_n18916,
    new_n18917, new_n18918, new_n18919_1, new_n18920, new_n18921,
    new_n18922, new_n18923, new_n18924, new_n18925, new_n18926_1,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940_1, new_n18941, new_n18942, new_n18943,
    new_n18944, new_n18945_1, new_n18946, new_n18947, new_n18948,
    new_n18949, new_n18950, new_n18951, new_n18952, new_n18953, new_n18954,
    new_n18955, new_n18956, new_n18957, new_n18958, new_n18959, new_n18960,
    new_n18961, new_n18962_1, new_n18963, new_n18964, new_n18965,
    new_n18966, new_n18969, new_n18970_1, new_n18971, new_n18972,
    new_n18973, new_n18974, new_n18975, new_n18976, new_n18977_1,
    new_n18978, new_n18979, new_n18980, new_n18981, new_n18982_1,
    new_n18983, new_n18984, new_n18985, new_n18986, new_n18987, new_n18988,
    new_n18989, new_n18990, new_n18991, new_n18992, new_n18993, new_n18994,
    new_n18995, new_n18996, new_n18997, new_n18998, new_n18999_1,
    new_n19000, new_n19003, new_n19004, new_n19005_1, new_n19006,
    new_n19007, new_n19008, new_n19009, new_n19010, new_n19011, new_n19012,
    new_n19013, new_n19014, new_n19015, new_n19016, new_n19017, new_n19018,
    new_n19019, new_n19020, new_n19021, new_n19023, new_n19028, new_n19029,
    new_n19030, new_n19031, new_n19032, new_n19033_1, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042_1, new_n19043, new_n19044_1, new_n19045,
    new_n19046, new_n19047, new_n19048, new_n19049, new_n19050, new_n19051,
    new_n19052, new_n19053, new_n19054, new_n19055, new_n19056, new_n19057,
    new_n19058, new_n19059, new_n19060, new_n19061, new_n19062, new_n19063,
    new_n19064, new_n19065, new_n19066, new_n19067, new_n19068, new_n19069,
    new_n19070, new_n19071, new_n19072, new_n19073, new_n19074, new_n19075,
    new_n19076, new_n19077, new_n19078, new_n19079, new_n19080,
    new_n19081_1, new_n19082, new_n19083, new_n19084, new_n19085,
    new_n19086, new_n19087, new_n19088, new_n19089, new_n19090, new_n19091,
    new_n19092, new_n19093, new_n19094, new_n19095, new_n19096, new_n19097,
    new_n19098, new_n19099, new_n19100, new_n19101, new_n19102, new_n19103,
    new_n19104, new_n19105, new_n19106, new_n19107_1, new_n19108,
    new_n19109, new_n19110, new_n19111, new_n19112, new_n19113, new_n19114,
    new_n19115, new_n19116_1, new_n19117, new_n19118, new_n19119,
    new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125_1, new_n19126, new_n19127, new_n19128, new_n19129,
    new_n19130, new_n19131, new_n19132, new_n19133, new_n19134, new_n19135,
    new_n19136, new_n19137, new_n19138, new_n19139, new_n19140,
    new_n19141_1, new_n19142, new_n19143, new_n19144_1, new_n19145,
    new_n19146, new_n19147, new_n19148, new_n19152, new_n19153, new_n19154,
    new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160,
    new_n19161, new_n19162, new_n19163_1, new_n19164_1, new_n19165,
    new_n19166, new_n19167, new_n19168, new_n19169, new_n19170, new_n19171,
    new_n19172, new_n19173, new_n19174_1, new_n19175, new_n19176_1,
    new_n19177, new_n19178, new_n19179, new_n19180, new_n19181, new_n19188,
    new_n19189, new_n19190, new_n19191, new_n19192, new_n19193, new_n19194,
    new_n19195, new_n19196_1, new_n19197, new_n19198, new_n19199,
    new_n19200, new_n19201, new_n19202_1, new_n19203, new_n19204,
    new_n19205, new_n19206, new_n19207, new_n19208, new_n19209, new_n19210,
    new_n19211, new_n19212, new_n19213, new_n19214, new_n19215, new_n19216,
    new_n19217, new_n19218, new_n19219, new_n19220_1, new_n19221_1,
    new_n19222, new_n19223_1, new_n19224_1, new_n19225, new_n19226,
    new_n19227, new_n19228_1, new_n19229, new_n19230, new_n19231,
    new_n19232, new_n19233_1, new_n19234_1, new_n19235, new_n19236,
    new_n19237, new_n19238, new_n19239, new_n19240, new_n19241, new_n19242,
    new_n19243, new_n19244_1, new_n19245, new_n19246, new_n19247,
    new_n19248, new_n19249, new_n19250, new_n19251, new_n19252, new_n19253,
    new_n19254, new_n19255, new_n19256, new_n19257, new_n19258, new_n19259,
    new_n19260, new_n19261, new_n19262, new_n19263, new_n19264, new_n19265,
    new_n19266, new_n19267, new_n19268, new_n19269, new_n19270_1,
    new_n19271, new_n19274, new_n19275, new_n19276, new_n19277, new_n19278,
    new_n19279, new_n19280, new_n19281, new_n19282_1, new_n19283,
    new_n19284, new_n19285, new_n19286, new_n19287, new_n19288, new_n19289,
    new_n19290, new_n19291, new_n19292, new_n19293, new_n19294, new_n19295,
    new_n19296, new_n19297, new_n19298, new_n19299, new_n19300, new_n19301,
    new_n19302, new_n19303, new_n19304, new_n19305, new_n19306, new_n19307,
    new_n19308, new_n19309, new_n19310, new_n19311, new_n19312, new_n19313,
    new_n19314_1, new_n19315_1, new_n19316, new_n19317, new_n19318,
    new_n19319, new_n19320, new_n19321, new_n19322, new_n19323_1,
    new_n19324, new_n19325, new_n19326, new_n19327_1, new_n19328,
    new_n19329, new_n19330, new_n19331, new_n19332, new_n19333_1,
    new_n19334, new_n19335, new_n19336, new_n19337, new_n19338, new_n19339,
    new_n19340, new_n19341, new_n19342, new_n19343, new_n19344, new_n19345,
    new_n19346, new_n19347, new_n19348_1, new_n19349, new_n19350,
    new_n19351, new_n19352, new_n19353, new_n19354_1, new_n19356,
    new_n19357_1, new_n19358, new_n19359, new_n19360, new_n19361_1,
    new_n19362, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367_1, new_n19368, new_n19369, new_n19370, new_n19371,
    new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377,
    new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383,
    new_n19384, new_n19385_1, new_n19386, new_n19387, new_n19388,
    new_n19389_1, new_n19390, new_n19391, new_n19392, new_n19393,
    new_n19394, new_n19395, new_n19396, new_n19397, new_n19398, new_n19399,
    new_n19400, new_n19401_1, new_n19402, new_n19403, new_n19404,
    new_n19405, new_n19406, new_n19407, new_n19408, new_n19409, new_n19410,
    new_n19411, new_n19412, new_n19413, new_n19415, new_n19416, new_n19417,
    new_n19418, new_n19419, new_n19420, new_n19421, new_n19422, new_n19423,
    new_n19424_1, new_n19425, new_n19426, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19442, new_n19443, new_n19444, new_n19445, new_n19446,
    new_n19447, new_n19448, new_n19449, new_n19450_1, new_n19451,
    new_n19452, new_n19453, new_n19454_1, new_n19455, new_n19456,
    new_n19457, new_n19458_1, new_n19459, new_n19460, new_n19461,
    new_n19466, new_n19467_1, new_n19468, new_n19469, new_n19470,
    new_n19471, new_n19472_1, new_n19473, new_n19474, new_n19475,
    new_n19476, new_n19477_1, new_n19478, new_n19479, new_n19480,
    new_n19485, new_n19486, new_n19487, new_n19488, new_n19489, new_n19490,
    new_n19491, new_n19492, new_n19493, new_n19494_1, new_n19495,
    new_n19496_1, new_n19497, new_n19498, new_n19499, new_n19500,
    new_n19501, new_n19502, new_n19503, new_n19504, new_n19505, new_n19506,
    new_n19507, new_n19508, new_n19509, new_n19510, new_n19511, new_n19512,
    new_n19513, new_n19514_1, new_n19515_1, new_n19516, new_n19517,
    new_n19518, new_n19519, new_n19520, new_n19521, new_n19522,
    new_n19523_1, new_n19524, new_n19525, new_n19526, new_n19527,
    new_n19528, new_n19529, new_n19530, new_n19531_1, new_n19532,
    new_n19533, new_n19534, new_n19535, new_n19536, new_n19537, new_n19538,
    new_n19539_1, new_n19541, new_n19542, new_n19543, new_n19544,
    new_n19545, new_n19546, new_n19548, new_n19549, new_n19550, new_n19551,
    new_n19552, new_n19553, new_n19554, new_n19555, new_n19556, new_n19557,
    new_n19558, new_n19559, new_n19563, new_n19564, new_n19565, new_n19566,
    new_n19567, new_n19568, new_n19569, new_n19570_1, new_n19571,
    new_n19572, new_n19573, new_n19574, new_n19575_1, new_n19576,
    new_n19577, new_n19578, new_n19579, new_n19580, new_n19581, new_n19582,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641_1, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648_1,
    new_n19649, new_n19650, new_n19652_1, new_n19653, new_n19654,
    new_n19655, new_n19656, new_n19657, new_n19658, new_n19659, new_n19660,
    new_n19661, new_n19663, new_n19664_1, new_n19665, new_n19666,
    new_n19667, new_n19668, new_n19669, new_n19670, new_n19671, new_n19672,
    new_n19673, new_n19674, new_n19675, new_n19676, new_n19677, new_n19678,
    new_n19679, new_n19680_1, new_n19681, new_n19682, new_n19683,
    new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689,
    new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695,
    new_n19696, new_n19697, new_n19698, new_n19699, new_n19700,
    new_n19701_1, new_n19702, new_n19703, new_n19704, new_n19705,
    new_n19706, new_n19707, new_n19708, new_n19709, new_n19710, new_n19711,
    new_n19712, new_n19713, new_n19714, new_n19715, new_n19716, new_n19717,
    new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723,
    new_n19724, new_n19725, new_n19726, new_n19727, new_n19728, new_n19729,
    new_n19730, new_n19731, new_n19732, new_n19733, new_n19734, new_n19735,
    new_n19736_1, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749_1, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756_1,
    new_n19757, new_n19758, new_n19759, new_n19760, new_n19761, new_n19762,
    new_n19763, new_n19764, new_n19765, new_n19766, new_n19767_1,
    new_n19768, new_n19769, new_n19770_1, new_n19771, new_n19772,
    new_n19773, new_n19774, new_n19775, new_n19776, new_n19777, new_n19778,
    new_n19779, new_n19780_1, new_n19781, new_n19782, new_n19783,
    new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789_1, new_n19790, new_n19791, new_n19792_1, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798_1,
    new_n19799, new_n19800, new_n19801, new_n19802, new_n19803_1,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19866, new_n19867, new_n19868, new_n19869,
    new_n19870, new_n19871, new_n19872, new_n19873_1, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19880,
    new_n19881, new_n19882, new_n19883, new_n19884, new_n19885, new_n19886,
    new_n19887, new_n19888, new_n19890, new_n19892, new_n19893, new_n19894,
    new_n19895, new_n19896, new_n19897, new_n19898, new_n19899, new_n19900,
    new_n19901, new_n19902, new_n19903, new_n19904, new_n19905_1,
    new_n19906, new_n19907, new_n19908, new_n19909_1, new_n19910,
    new_n19911_1, new_n19912, new_n19913, new_n19914, new_n19915,
    new_n19916_1, new_n19917, new_n19918, new_n19919, new_n19920,
    new_n19921, new_n19922_1, new_n19924, new_n19925, new_n19926,
    new_n19927, new_n19928, new_n19929, new_n19930_1, new_n19931,
    new_n19932, new_n19933, new_n19934, new_n19935, new_n19936, new_n19937,
    new_n19938, new_n19939, new_n19940, new_n19941_1, new_n19942,
    new_n19943, new_n19946, new_n19947, new_n19948, new_n19949, new_n19950,
    new_n19951, new_n19952, new_n19953, new_n19954, new_n19959, new_n19960,
    new_n19961, new_n19962, new_n19963, new_n19964, new_n19965, new_n19966,
    new_n19967, new_n19968_1, new_n19969, new_n19970, new_n19971,
    new_n19972, new_n19973, new_n19974, new_n19975, new_n19976, new_n19977,
    new_n19978, new_n19979, new_n19980, new_n19981, new_n19982, new_n19983,
    new_n19984, new_n19985, new_n19986, new_n19987, new_n19988_1,
    new_n19989, new_n19990, new_n19991, new_n19992, new_n19993, new_n19994,
    new_n19995, new_n19996, new_n19997, new_n19998, new_n19999, new_n20000,
    new_n20001, new_n20002, new_n20003, new_n20004_1, new_n20005,
    new_n20006, new_n20007, new_n20008, new_n20009, new_n20010, new_n20011,
    new_n20012, new_n20013_1, new_n20014, new_n20015, new_n20016,
    new_n20017_1, new_n20018, new_n20019, new_n20020, new_n20021,
    new_n20022, new_n20023, new_n20024, new_n20025, new_n20026, new_n20027,
    new_n20028, new_n20029, new_n20030, new_n20031, new_n20032,
    new_n20033_1, new_n20034, new_n20035, new_n20036_1, new_n20037,
    new_n20038, new_n20039, new_n20040_1, new_n20041, new_n20042,
    new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061_1, new_n20062, new_n20063, new_n20064, new_n20065,
    new_n20066, new_n20067, new_n20068, new_n20069_1, new_n20070,
    new_n20071, new_n20072, new_n20073, new_n20074, new_n20075, new_n20076,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086_1, new_n20087, new_n20088, new_n20089,
    new_n20090, new_n20091, new_n20092, new_n20093, new_n20094, new_n20095,
    new_n20096_1, new_n20097, new_n20099, new_n20100, new_n20101,
    new_n20102, new_n20103_1, new_n20104, new_n20105, new_n20106,
    new_n20107, new_n20108, new_n20109, new_n20110, new_n20111, new_n20112,
    new_n20113, new_n20114, new_n20115, new_n20116, new_n20117, new_n20118,
    new_n20119, new_n20120, new_n20121, new_n20122, new_n20123, new_n20124,
    new_n20125, new_n20126_1, new_n20127, new_n20128, new_n20129,
    new_n20130, new_n20131, new_n20132, new_n20133, new_n20134, new_n20135,
    new_n20136, new_n20137, new_n20138_1, new_n20139, new_n20140,
    new_n20141, new_n20142, new_n20143, new_n20144, new_n20145, new_n20146,
    new_n20147, new_n20148, new_n20149_1, new_n20150, new_n20151_1,
    new_n20152, new_n20153, new_n20154, new_n20155, new_n20156, new_n20157,
    new_n20158, new_n20159, new_n20162, new_n20163, new_n20164, new_n20165,
    new_n20166, new_n20167, new_n20168, new_n20169_1, new_n20170,
    new_n20171, new_n20172, new_n20173, new_n20174, new_n20175, new_n20176,
    new_n20177, new_n20178, new_n20179_1, new_n20180, new_n20181,
    new_n20182, new_n20183, new_n20184, new_n20185, new_n20186,
    new_n20187_1, new_n20188, new_n20189, new_n20190, new_n20191,
    new_n20192, new_n20193, new_n20194, new_n20195, new_n20196, new_n20198,
    new_n20199, new_n20200, new_n20201, new_n20202, new_n20203, new_n20204,
    new_n20205, new_n20206, new_n20207, new_n20208, new_n20209, new_n20210,
    new_n20211, new_n20212, new_n20213_1, new_n20214, new_n20215,
    new_n20216, new_n20217, new_n20218, new_n20219, new_n20220, new_n20221,
    new_n20222, new_n20223, new_n20224, new_n20225, new_n20226, new_n20227,
    new_n20228, new_n20229, new_n20230, new_n20231, new_n20232, new_n20233,
    new_n20234, new_n20235_1, new_n20236, new_n20240, new_n20242,
    new_n20243, new_n20244, new_n20245, new_n20246, new_n20247, new_n20248,
    new_n20249, new_n20250_1, new_n20251, new_n20252, new_n20253,
    new_n20254, new_n20255, new_n20256, new_n20257, new_n20258,
    new_n20259_1, new_n20260, new_n20261, new_n20262, new_n20263,
    new_n20264, new_n20269, new_n20270, new_n20271, new_n20272, new_n20273,
    new_n20274, new_n20275, new_n20276, new_n20277, new_n20278,
    new_n20279_1, new_n20280, new_n20281, new_n20282, new_n20283,
    new_n20284, new_n20285, new_n20286, new_n20287_1, new_n20288,
    new_n20289, new_n20290, new_n20291, new_n20292, new_n20293, new_n20294,
    new_n20295, new_n20296, new_n20297, new_n20298, new_n20299, new_n20300,
    new_n20301_1, new_n20302, new_n20303, new_n20304, new_n20305,
    new_n20306, new_n20307, new_n20308, new_n20309, new_n20310, new_n20311,
    new_n20312, new_n20313, new_n20314, new_n20315, new_n20316, new_n20317,
    new_n20318, new_n20319, new_n20320, new_n20321, new_n20322, new_n20323,
    new_n20324, new_n20325, new_n20326, new_n20327, new_n20328, new_n20329,
    new_n20330_1, new_n20331, new_n20332, new_n20333_1, new_n20334,
    new_n20335, new_n20336, new_n20337, new_n20338, new_n20339, new_n20340,
    new_n20341, new_n20342, new_n20343, new_n20344, new_n20345, new_n20346,
    new_n20347, new_n20348, new_n20349_1, new_n20350, new_n20351,
    new_n20352, new_n20353, new_n20354, new_n20355_1, new_n20356,
    new_n20357, new_n20363, new_n20364, new_n20365, new_n20366_1,
    new_n20367, new_n20368, new_n20369, new_n20370, new_n20371, new_n20372,
    new_n20373, new_n20374, new_n20375, new_n20376, new_n20377, new_n20378,
    new_n20379, new_n20380, new_n20382, new_n20383, new_n20384,
    new_n20385_1, new_n20386, new_n20387, new_n20388_1, new_n20389,
    new_n20390, new_n20391, new_n20392, new_n20393, new_n20394, new_n20395,
    new_n20396, new_n20397, new_n20398, new_n20399, new_n20400, new_n20401,
    new_n20402_1, new_n20403_1, new_n20404, new_n20405, new_n20406,
    new_n20407, new_n20408, new_n20409_1, new_n20410, new_n20411_1,
    new_n20412, new_n20413, new_n20414, new_n20415, new_n20416, new_n20417,
    new_n20418, new_n20419, new_n20420, new_n20421, new_n20422, new_n20423,
    new_n20424_1, new_n20425, new_n20426, new_n20427, new_n20428,
    new_n20429_1, new_n20430, new_n20431, new_n20432, new_n20433,
    new_n20434, new_n20435, new_n20436_1, new_n20437, new_n20438,
    new_n20439, new_n20440, new_n20441_1, new_n20442, new_n20443,
    new_n20444, new_n20445_1, new_n20446, new_n20447, new_n20448,
    new_n20449, new_n20450_1, new_n20451, new_n20452, new_n20453,
    new_n20454, new_n20455_1, new_n20456, new_n20457, new_n20458,
    new_n20459, new_n20460, new_n20461, new_n20462, new_n20467, new_n20468,
    new_n20469, new_n20470_1, new_n20471, new_n20472, new_n20473,
    new_n20474, new_n20475, new_n20476, new_n20477, new_n20478_1,
    new_n20479, new_n20480, new_n20481, new_n20482, new_n20483, new_n20484,
    new_n20485, new_n20486, new_n20487, new_n20488, new_n20489_1,
    new_n20490_1, new_n20491, new_n20492, new_n20493, new_n20494,
    new_n20495_1, new_n20496, new_n20497, new_n20498, new_n20499,
    new_n20500, new_n20501, new_n20502, new_n20503, new_n20504, new_n20505,
    new_n20506, new_n20507, new_n20508, new_n20509, new_n20510, new_n20511,
    new_n20512, new_n20513, new_n20514, new_n20515_1, new_n20516,
    new_n20517, new_n20518, new_n20519, new_n20520, new_n20521, new_n20522,
    new_n20523, new_n20524, new_n20525, new_n20526, new_n20527, new_n20528,
    new_n20529, new_n20530, new_n20531, new_n20532, new_n20533_1,
    new_n20534, new_n20535, new_n20536, new_n20537, new_n20538, new_n20539,
    new_n20540, new_n20541, new_n20542, new_n20543, new_n20544, new_n20545,
    new_n20546, new_n20547, new_n20548, new_n20549, new_n20550, new_n20551,
    new_n20552, new_n20553, new_n20554, new_n20557, new_n20558, new_n20559,
    new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571,
    new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582_1,
    new_n20583, new_n20584, new_n20585, new_n20586, new_n20587, new_n20588,
    new_n20589, new_n20590_1, new_n20591, new_n20592, new_n20593,
    new_n20594, new_n20595, new_n20596, new_n20597, new_n20598, new_n20599,
    new_n20600, new_n20601, new_n20602_1, new_n20603, new_n20604_1,
    new_n20605, new_n20606, new_n20607, new_n20608, new_n20609_1,
    new_n20610, new_n20611, new_n20612, new_n20613, new_n20614, new_n20615,
    new_n20616, new_n20617, new_n20618, new_n20619, new_n20620, new_n20621,
    new_n20622, new_n20623_1, new_n20624, new_n20625, new_n20626,
    new_n20627, new_n20628, new_n20629_1, new_n20630, new_n20631,
    new_n20632, new_n20635, new_n20636, new_n20637, new_n20638, new_n20639,
    new_n20640, new_n20641, new_n20642, new_n20643, new_n20644, new_n20645,
    new_n20646, new_n20647, new_n20648, new_n20649, new_n20650, new_n20651,
    new_n20652, new_n20654, new_n20655, new_n20656, new_n20657,
    new_n20658_1, new_n20659, new_n20660, new_n20661_1, new_n20662,
    new_n20663, new_n20664, new_n20665, new_n20666, new_n20667, new_n20668,
    new_n20669, new_n20670, new_n20671, new_n20672, new_n20673_1,
    new_n20674, new_n20675, new_n20676, new_n20677, new_n20679,
    new_n20680_1, new_n20681, new_n20682, new_n20683, new_n20684,
    new_n20685_1, new_n20686, new_n20687, new_n20688, new_n20689,
    new_n20690, new_n20691_1, new_n20692, new_n20693, new_n20694,
    new_n20695, new_n20696_1, new_n20697, new_n20698, new_n20699,
    new_n20700_1, new_n20701, new_n20702, new_n20703, new_n20704_1,
    new_n20705_1, new_n20706, new_n20707, new_n20708, new_n20709_1,
    new_n20710, new_n20711, new_n20712, new_n20713_1, new_n20714,
    new_n20715, new_n20716, new_n20717, new_n20718, new_n20719, new_n20720,
    new_n20721, new_n20722_1, new_n20723_1, new_n20724, new_n20725,
    new_n20726, new_n20727, new_n20729, new_n20732, new_n20733, new_n20734,
    new_n20735, new_n20736, new_n20737, new_n20738, new_n20739, new_n20740,
    new_n20741, new_n20742, new_n20743, new_n20744, new_n20745, new_n20746,
    new_n20747, new_n20748_1, new_n20749, new_n20750, new_n20751,
    new_n20752, new_n20753, new_n20754, new_n20755, new_n20756, new_n20757,
    new_n20758, new_n20759, new_n20760, new_n20761_1, new_n20762,
    new_n20763, new_n20764, new_n20765, new_n20766, new_n20767, new_n20768,
    new_n20769, new_n20770, new_n20771, new_n20772, new_n20773,
    new_n20774_1, new_n20775, new_n20776, new_n20777, new_n20778,
    new_n20779, new_n20780, new_n20781, new_n20782, new_n20783, new_n20784,
    new_n20786, new_n20787, new_n20788_1, new_n20789, new_n20790,
    new_n20791, new_n20792, new_n20793, new_n20794_1, new_n20795_1,
    new_n20796, new_n20797, new_n20798, new_n20799, new_n20800, new_n20801,
    new_n20802, new_n20803_1, new_n20804, new_n20805, new_n20806,
    new_n20807, new_n20808, new_n20809, new_n20810, new_n20811, new_n20812,
    new_n20813, new_n20814, new_n20815, new_n20816, new_n20817, new_n20818,
    new_n20820, new_n20821, new_n20822, new_n20823, new_n20824, new_n20825,
    new_n20826_1, new_n20827, new_n20828, new_n20829, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20836,
    new_n20837, new_n20838, new_n20843, new_n20844, new_n20845, new_n20846,
    new_n20847, new_n20848, new_n20849, new_n20850, new_n20851, new_n20854,
    new_n20855, new_n20856, new_n20857, new_n20858, new_n20859, new_n20860,
    new_n20861, new_n20862, new_n20863, new_n20864, new_n20865, new_n20866,
    new_n20867, new_n20868, new_n20869_1, new_n20870, new_n20871,
    new_n20872, new_n20873, new_n20874, new_n20875, new_n20876, new_n20877,
    new_n20878, new_n20879_1, new_n20880, new_n20881, new_n20882,
    new_n20883, new_n20884, new_n20885, new_n20886, new_n20887, new_n20888,
    new_n20889, new_n20890, new_n20891, new_n20892, new_n20893, new_n20894,
    new_n20895, new_n20896, new_n20897, new_n20898, new_n20899, new_n20900,
    new_n20901, new_n20902, new_n20903, new_n20904, new_n20905, new_n20906,
    new_n20907, new_n20908, new_n20909, new_n20910, new_n20911, new_n20912,
    new_n20913, new_n20914, new_n20915_1, new_n20916, new_n20917,
    new_n20918, new_n20919, new_n20920, new_n20921, new_n20922, new_n20927,
    new_n20928, new_n20929_1, new_n20930, new_n20931, new_n20932,
    new_n20933, new_n20934, new_n20935_1, new_n20936_1, new_n20937,
    new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943,
    new_n20944, new_n20945, new_n20946_1, new_n20947, new_n20948,
    new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20957,
    new_n20958, new_n20959, new_n20960, new_n20961, new_n20962, new_n20963,
    new_n20964, new_n20965, new_n20966, new_n20967, new_n20968, new_n20969,
    new_n20970, new_n20971, new_n20972, new_n20973, new_n20974, new_n20975,
    new_n20976, new_n20977, new_n20978, new_n20979, new_n20980, new_n20981,
    new_n20982, new_n20983, new_n20984, new_n20985, new_n20986_1,
    new_n20987, new_n20988, new_n20989, new_n20990, new_n20991, new_n20992,
    new_n20993, new_n20994, new_n20995, new_n20996, new_n20997, new_n20998,
    new_n20999, new_n21000, new_n21001, new_n21002, new_n21003, new_n21004,
    new_n21005, new_n21006, new_n21007, new_n21008_1, new_n21009,
    new_n21010, new_n21011, new_n21012, new_n21013, new_n21014, new_n21015,
    new_n21016, new_n21017_1, new_n21018, new_n21019, new_n21020,
    new_n21021, new_n21022, new_n21023, new_n21024, new_n21025, new_n21026,
    new_n21027, new_n21028, new_n21029, new_n21030, new_n21031, new_n21032,
    new_n21033, new_n21034_1, new_n21035, new_n21036, new_n21037,
    new_n21038, new_n21039, new_n21040, new_n21041, new_n21042, new_n21043,
    new_n21044, new_n21045, new_n21046_1, new_n21047, new_n21048,
    new_n21049, new_n21050, new_n21051, new_n21052, new_n21053, new_n21054,
    new_n21055, new_n21056, new_n21057, new_n21058, new_n21059, new_n21060,
    new_n21061, new_n21062_1, new_n21063, new_n21064, new_n21065,
    new_n21066, new_n21067, new_n21068, new_n21069, new_n21077,
    new_n21078_1, new_n21079, new_n21080, new_n21081, new_n21082,
    new_n21083, new_n21084, new_n21085, new_n21086, new_n21087, new_n21088,
    new_n21089, new_n21090, new_n21091, new_n21092, new_n21093_1,
    new_n21094_1, new_n21095_1, new_n21096, new_n21097, new_n21098,
    new_n21099, new_n21100, new_n21101, new_n21102, new_n21103, new_n21104,
    new_n21105, new_n21106, new_n21107, new_n21108, new_n21109, new_n21110,
    new_n21111, new_n21112, new_n21113, new_n21114, new_n21115, new_n21116,
    new_n21117, new_n21118, new_n21122, new_n21123_1, new_n21124,
    new_n21125, new_n21126, new_n21127, new_n21128, new_n21129, new_n21130,
    new_n21131, new_n21132, new_n21133, new_n21134_1, new_n21135,
    new_n21136, new_n21137, new_n21138_1, new_n21139, new_n21140,
    new_n21141, new_n21142, new_n21143, new_n21144, new_n21145, new_n21146,
    new_n21147, new_n21148, new_n21149, new_n21150, new_n21151, new_n21152,
    new_n21153, new_n21154_1, new_n21155, new_n21156, new_n21157_1,
    new_n21158, new_n21159, new_n21160, new_n21161, new_n21162, new_n21163,
    new_n21164, new_n21165, new_n21166, new_n21167, new_n21168_1,
    new_n21169, new_n21170, new_n21171, new_n21172, new_n21173_1,
    new_n21174, new_n21175, new_n21176_1, new_n21177, new_n21178,
    new_n21179, new_n21180, new_n21181, new_n21182_1, new_n21183,
    new_n21184, new_n21185, new_n21186, new_n21187, new_n21188, new_n21189,
    new_n21190, new_n21191, new_n21192, new_n21193_1, new_n21194,
    new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200,
    new_n21201, new_n21202, new_n21203_1, new_n21204, new_n21205,
    new_n21206, new_n21207, new_n21208, new_n21209, new_n21210, new_n21211,
    new_n21212, new_n21213, new_n21214, new_n21215, new_n21216, new_n21217,
    new_n21218, new_n21219, new_n21220, new_n21221, new_n21222_1,
    new_n21223, new_n21224, new_n21225_1, new_n21226_1, new_n21227,
    new_n21228, new_n21229, new_n21230, new_n21231, new_n21232, new_n21234,
    new_n21235, new_n21236, new_n21237, new_n21238_1, new_n21239,
    new_n21240, new_n21241, new_n21242, new_n21243, new_n21244, new_n21245,
    new_n21246, new_n21250, new_n21251, new_n21252, new_n21253,
    new_n21254_1, new_n21255, new_n21256, new_n21257, new_n21258,
    new_n21259, new_n21260, new_n21261, new_n21262, new_n21263, new_n21264,
    new_n21265, new_n21266, new_n21267, new_n21268, new_n21269, new_n21270,
    new_n21271, new_n21272, new_n21273, new_n21274, new_n21275,
    new_n21276_1, new_n21277, new_n21278, new_n21280, new_n21281,
    new_n21282, new_n21283, new_n21284, new_n21285, new_n21286,
    new_n21287_1, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298_1, new_n21299, new_n21300, new_n21301, new_n21302_1,
    new_n21303, new_n21304, new_n21305, new_n21306, new_n21307, new_n21308,
    new_n21309, new_n21310, new_n21311, new_n21312, new_n21313, new_n21314,
    new_n21315, new_n21316, new_n21317_1, new_n21318, new_n21319,
    new_n21320, new_n21321, new_n21322, new_n21323, new_n21324, new_n21325,
    new_n21326, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331,
    new_n21332, new_n21333, new_n21334, new_n21335, new_n21336, new_n21337,
    new_n21338, new_n21339, new_n21340, new_n21341, new_n21342, new_n21343,
    new_n21344, new_n21345, new_n21346, new_n21347, new_n21348,
    new_n21349_1, new_n21350, new_n21351, new_n21352, new_n21353,
    new_n21355, new_n21358, new_n21359, new_n21360, new_n21361, new_n21362,
    new_n21363, new_n21364, new_n21365_1, new_n21366, new_n21367_1,
    new_n21368, new_n21369, new_n21370, new_n21371, new_n21372, new_n21373,
    new_n21374, new_n21375, new_n21376, new_n21377, new_n21378, new_n21379,
    new_n21380, new_n21381, new_n21382, new_n21383, new_n21384, new_n21385,
    new_n21386, new_n21387, new_n21388, new_n21389, new_n21390, new_n21391,
    new_n21392, new_n21393, new_n21394, new_n21395, new_n21396_1,
    new_n21397, new_n21398_1, new_n21399_1, new_n21400, new_n21401,
    new_n21402, new_n21403, new_n21404_1, new_n21405, new_n21406,
    new_n21407, new_n21408, new_n21409, new_n21410, new_n21411, new_n21412,
    new_n21413, new_n21414, new_n21415, new_n21416, new_n21417, new_n21418,
    new_n21419, new_n21420, new_n21421, new_n21422, new_n21423, new_n21424,
    new_n21425, new_n21426, new_n21427, new_n21428, new_n21429, new_n21430,
    new_n21431, new_n21432, new_n21433, new_n21434, new_n21435, new_n21436,
    new_n21437, new_n21438, new_n21439, new_n21440, new_n21441, new_n21442,
    new_n21443, new_n21444, new_n21445, new_n21446_1, new_n21447,
    new_n21448, new_n21449, new_n21450, new_n21451, new_n21452, new_n21453,
    new_n21454, new_n21455, new_n21456, new_n21457, new_n21458, new_n21459,
    new_n21460, new_n21461, new_n21462, new_n21463, new_n21464, new_n21465,
    new_n21466, new_n21467, new_n21468, new_n21469, new_n21470,
    new_n21471_1, new_n21472_1, new_n21473, new_n21474, new_n21475,
    new_n21476, new_n21477, new_n21478, new_n21479, new_n21482, new_n21483,
    new_n21484, new_n21485, new_n21486, new_n21487, new_n21488,
    new_n21489_1, new_n21490, new_n21491, new_n21492, new_n21493,
    new_n21494, new_n21495, new_n21496, new_n21497, new_n21498, new_n21499,
    new_n21500, new_n21501, new_n21502, new_n21503, new_n21504, new_n21505,
    new_n21506, new_n21507, new_n21508, new_n21509, new_n21510, new_n21511,
    new_n21512, new_n21513, new_n21514, new_n21515, new_n21516, new_n21517,
    new_n21518, new_n21519, new_n21520, new_n21521, new_n21522, new_n21523,
    new_n21524, new_n21525_1, new_n21526, new_n21527, new_n21528,
    new_n21529, new_n21530, new_n21531, new_n21532, new_n21533, new_n21534,
    new_n21535, new_n21536, new_n21537, new_n21538_1, new_n21539,
    new_n21540, new_n21541, new_n21542, new_n21543, new_n21544, new_n21545,
    new_n21546, new_n21547, new_n21548, new_n21549_1, new_n21550,
    new_n21551, new_n21552, new_n21553, new_n21554, new_n21555, new_n21556,
    new_n21557, new_n21558, new_n21559, new_n21560, new_n21561, new_n21568,
    new_n21569, new_n21570, new_n21571, new_n21575, new_n21576, new_n21577,
    new_n21578, new_n21579, new_n21580, new_n21581, new_n21582, new_n21583,
    new_n21584, new_n21585, new_n21586, new_n21587, new_n21588, new_n21589,
    new_n21590, new_n21591, new_n21592, new_n21593, new_n21594, new_n21595,
    new_n21596, new_n21597, new_n21598, new_n21599_1, new_n21600,
    new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606,
    new_n21607, new_n21608, new_n21609, new_n21610, new_n21611, new_n21612,
    new_n21613, new_n21614, new_n21615_1, new_n21616, new_n21617,
    new_n21618, new_n21619, new_n21620, new_n21621, new_n21622, new_n21623,
    new_n21624, new_n21625, new_n21626, new_n21627, new_n21628_1,
    new_n21629, new_n21630, new_n21631, new_n21632, new_n21633, new_n21634,
    new_n21635, new_n21636, new_n21637_1, new_n21638, new_n21639,
    new_n21640, new_n21641, new_n21642, new_n21643, new_n21644,
    new_n21645_1, new_n21646, new_n21647, new_n21648, new_n21649_1,
    new_n21650, new_n21651, new_n21652, new_n21653, new_n21654_1,
    new_n21655, new_n21656, new_n21657, new_n21658, new_n21659, new_n21660,
    new_n21661, new_n21662, new_n21663, new_n21664, new_n21665_1,
    new_n21666, new_n21667, new_n21668, new_n21669, new_n21670, new_n21671,
    new_n21672, new_n21673, new_n21674_1, new_n21675, new_n21676,
    new_n21677, new_n21678, new_n21679, new_n21680_1, new_n21681,
    new_n21682, new_n21683, new_n21684, new_n21685_1, new_n21686,
    new_n21687_1, new_n21688, new_n21689, new_n21690, new_n21691,
    new_n21692, new_n21693, new_n21694, new_n21695, new_n21696, new_n21697,
    new_n21698, new_n21699, new_n21700, new_n21701, new_n21702, new_n21703,
    new_n21704, new_n21705, new_n21706, new_n21707, new_n21708, new_n21709,
    new_n21710, new_n21711, new_n21712, new_n21713, new_n21714, new_n21715,
    new_n21716, new_n21717_1, new_n21718, new_n21719_1, new_n21720,
    new_n21721, new_n21722, new_n21723, new_n21724, new_n21727, new_n21728,
    new_n21729, new_n21730, new_n21731, new_n21732, new_n21733, new_n21734,
    new_n21735_1, new_n21736, new_n21737, new_n21738, new_n21739,
    new_n21740, new_n21741, new_n21742, new_n21743, new_n21744, new_n21745,
    new_n21746, new_n21747, new_n21748, new_n21749_1, new_n21750_1,
    new_n21751, new_n21752, new_n21753_1, new_n21754, new_n21755,
    new_n21756, new_n21757, new_n21758, new_n21759, new_n21760, new_n21761,
    new_n21762, new_n21763, new_n21764, new_n21765_1, new_n21766,
    new_n21767, new_n21768, new_n21769, new_n21770, new_n21771, new_n21772,
    new_n21773, new_n21774, new_n21775, new_n21776, new_n21777, new_n21778,
    new_n21779_1, new_n21780, new_n21781, new_n21782, new_n21783,
    new_n21784_1, new_n21785, new_n21786, new_n21787, new_n21788,
    new_n21789, new_n21790, new_n21791, new_n21792, new_n21793, new_n21794,
    new_n21795, new_n21796, new_n21797, new_n21798, new_n21799,
    new_n21800_1, new_n21801, new_n21802, new_n21803, new_n21804,
    new_n21805, new_n21806, new_n21807, new_n21808, new_n21809, new_n21810,
    new_n21811, new_n21812, new_n21813, new_n21814, new_n21815, new_n21816,
    new_n21817, new_n21818, new_n21819, new_n21820_1, new_n21821,
    new_n21822, new_n21827, new_n21828, new_n21829, new_n21830, new_n21831,
    new_n21832_1, new_n21833, new_n21834, new_n21835, new_n21836,
    new_n21837, new_n21838, new_n21839_1, new_n21840, new_n21841,
    new_n21842, new_n21843, new_n21844, new_n21845, new_n21846, new_n21847,
    new_n21848, new_n21849, new_n21850, new_n21851, new_n21852, new_n21853,
    new_n21854, new_n21855, new_n21856, new_n21857, new_n21858, new_n21859,
    new_n21860, new_n21861, new_n21862, new_n21863, new_n21864, new_n21865,
    new_n21866, new_n21867, new_n21868, new_n21869, new_n21870, new_n21871,
    new_n21872, new_n21873, new_n21874_1, new_n21875, new_n21876,
    new_n21877, new_n21878, new_n21879, new_n21880, new_n21881, new_n21882,
    new_n21883, new_n21884, new_n21885, new_n21886, new_n21887, new_n21888,
    new_n21889, new_n21890, new_n21891, new_n21892, new_n21893, new_n21894,
    new_n21895, new_n21896, new_n21897, new_n21898_1, new_n21899,
    new_n21900, new_n21901, new_n21902, new_n21903, new_n21904,
    new_n21905_1, new_n21906, new_n21907, new_n21908, new_n21909,
    new_n21910, new_n21911, new_n21912, new_n21913, new_n21914,
    new_n21915_1, new_n21916, new_n21917, new_n21918, new_n21919,
    new_n21920, new_n21921, new_n21922, new_n21923, new_n21924, new_n21925,
    new_n21926, new_n21927, new_n21928, new_n21929, new_n21930, new_n21931,
    new_n21932, new_n21933, new_n21935, new_n21936, new_n21937, new_n21938,
    new_n21939, new_n21940, new_n21941, new_n21942, new_n21943_1,
    new_n21945, new_n21946, new_n21947, new_n21948, new_n21949, new_n21950,
    new_n21951, new_n21952, new_n21953, new_n21954, new_n21955, new_n21956,
    new_n21957_1, new_n21958, new_n21959, new_n21960_1, new_n21961,
    new_n21962, new_n21963, new_n21964, new_n21965, new_n21966, new_n21967,
    new_n21968, new_n21969, new_n21970, new_n21971, new_n21972, new_n21973,
    new_n21974, new_n21975, new_n21982, new_n21983, new_n21984, new_n21985,
    new_n21986_1, new_n21987, new_n21988, new_n21989, new_n21990,
    new_n21991, new_n21992, new_n21993_1, new_n21994, new_n21995,
    new_n21996, new_n21997_1, new_n21998, new_n21999, new_n22011,
    new_n22012, new_n22013, new_n22014, new_n22015, new_n22016_1,
    new_n22017, new_n22018, new_n22019, new_n22020, new_n22021, new_n22022,
    new_n22023, new_n22024, new_n22025, new_n22026, new_n22027_1,
    new_n22028, new_n22029, new_n22030, new_n22031, new_n22032, new_n22033,
    new_n22034, new_n22035, new_n22036, new_n22037, new_n22038, new_n22039,
    new_n22040, new_n22041, new_n22042, new_n22043_1, new_n22044,
    new_n22045, new_n22046, new_n22047, new_n22048, new_n22049,
    new_n22050_1, new_n22051, new_n22052, new_n22053, new_n22054,
    new_n22055, new_n22056, new_n22057, new_n22058, new_n22059, new_n22061,
    new_n22062, new_n22063_1, new_n22064, new_n22065, new_n22066,
    new_n22067, new_n22068_1, new_n22069, new_n22070, new_n22071,
    new_n22072_1, new_n22073, new_n22074, new_n22075, new_n22076_1,
    new_n22077, new_n22078, new_n22079, new_n22080, new_n22081, new_n22082,
    new_n22083, new_n22084, new_n22085, new_n22086, new_n22087, new_n22088,
    new_n22089, new_n22090_1, new_n22092, new_n22093, new_n22094,
    new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100,
    new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106,
    new_n22107_1, new_n22108, new_n22109, new_n22110, new_n22111,
    new_n22112, new_n22113_1, new_n22114, new_n22115, new_n22116,
    new_n22117, new_n22118, new_n22119, new_n22120, new_n22121, new_n22122,
    new_n22123, new_n22124_1, new_n22125, new_n22126_1, new_n22127,
    new_n22128, new_n22129, new_n22130_1, new_n22131, new_n22132,
    new_n22133, new_n22134, new_n22135, new_n22136, new_n22137, new_n22138,
    new_n22139, new_n22140, new_n22141, new_n22142, new_n22143,
    new_n22144_1, new_n22145, new_n22146, new_n22147, new_n22148,
    new_n22149, new_n22150_1, new_n22151, new_n22152, new_n22153,
    new_n22154, new_n22155, new_n22156, new_n22157_1, new_n22158,
    new_n22159, new_n22160, new_n22161, new_n22162, new_n22163, new_n22164,
    new_n22165, new_n22166, new_n22167, new_n22168, new_n22169, new_n22170,
    new_n22171, new_n22172, new_n22173_1, new_n22174, new_n22175,
    new_n22176, new_n22177, new_n22178, new_n22179, new_n22180, new_n22181,
    new_n22182, new_n22183, new_n22184, new_n22185, new_n22186, new_n22187,
    new_n22188, new_n22189, new_n22190, new_n22191, new_n22192, new_n22193,
    new_n22194, new_n22195, new_n22196, new_n22197, new_n22198_1,
    new_n22199, new_n22200, new_n22201_1, new_n22202, new_n22203,
    new_n22204, new_n22205, new_n22206, new_n22207, new_n22208, new_n22209,
    new_n22210, new_n22211, new_n22212, new_n22213_1, new_n22214,
    new_n22215, new_n22216, new_n22217, new_n22218, new_n22219, new_n22220,
    new_n22221, new_n22222, new_n22223, new_n22224, new_n22225, new_n22226,
    new_n22227, new_n22228, new_n22229, new_n22230, new_n22231, new_n22232,
    new_n22233, new_n22234, new_n22235, new_n22236, new_n22237, new_n22238,
    new_n22239, new_n22240, new_n22241, new_n22242, new_n22243, new_n22244,
    new_n22245, new_n22246, new_n22247, new_n22248, new_n22249, new_n22250,
    new_n22251, new_n22252, new_n22253_1, new_n22254, new_n22255,
    new_n22256, new_n22257, new_n22258, new_n22259, new_n22260, new_n22265,
    new_n22266, new_n22267, new_n22268, new_n22269, new_n22270_1,
    new_n22271, new_n22272, new_n22273, new_n22274_1, new_n22275,
    new_n22276, new_n22277, new_n22278, new_n22279, new_n22280, new_n22281,
    new_n22282, new_n22283_1, new_n22284, new_n22285, new_n22286,
    new_n22287, new_n22290_1, new_n22291, new_n22292, new_n22293,
    new_n22294, new_n22295, new_n22296, new_n22297, new_n22298, new_n22299,
    new_n22300, new_n22301, new_n22302, new_n22303, new_n22304, new_n22305,
    new_n22306, new_n22307, new_n22308, new_n22309_1, new_n22310,
    new_n22313, new_n22314, new_n22315, new_n22316, new_n22317_1,
    new_n22318, new_n22319, new_n22320, new_n22325, new_n22326, new_n22330,
    new_n22331, new_n22332_1, new_n22333, new_n22334, new_n22335_1,
    new_n22336, new_n22337, new_n22338, new_n22339, new_n22340,
    new_n22341_1, new_n22342, new_n22343, new_n22344, new_n22345,
    new_n22346, new_n22350, new_n22351, new_n22352, new_n22353_1,
    new_n22354, new_n22355, new_n22356, new_n22357, new_n22358_1,
    new_n22359_1, new_n22360, new_n22362, new_n22363, new_n22364,
    new_n22365, new_n22366, new_n22367, new_n22368, new_n22369, new_n22370,
    new_n22371, new_n22372, new_n22373, new_n22374, new_n22375, new_n22376,
    new_n22377, new_n22378, new_n22379_1, new_n22380, new_n22381,
    new_n22383, new_n22384, new_n22385, new_n22386, new_n22387, new_n22388,
    new_n22389, new_n22390, new_n22391, new_n22392, new_n22393, new_n22394,
    new_n22395, new_n22396, new_n22397, new_n22398, new_n22399, new_n22400,
    new_n22401, new_n22402, new_n22403, new_n22404, new_n22405, new_n22406,
    new_n22407, new_n22408, new_n22409, new_n22410, new_n22411, new_n22412,
    new_n22413, new_n22414, new_n22415, new_n22416, new_n22417, new_n22418,
    new_n22419, new_n22420, new_n22421, new_n22423, new_n22424, new_n22425,
    new_n22426, new_n22427, new_n22428, new_n22429, new_n22430, new_n22431,
    new_n22432, new_n22433_1, new_n22434, new_n22435, new_n22436,
    new_n22437, new_n22438, new_n22439, new_n22440, new_n22441,
    new_n22442_1, new_n22443, new_n22444_1, new_n22445, new_n22446,
    new_n22447, new_n22448, new_n22449, new_n22450, new_n22451, new_n22452,
    new_n22453, new_n22454, new_n22455, new_n22456, new_n22457, new_n22458,
    new_n22459, new_n22460, new_n22461, new_n22462, new_n22463, new_n22464,
    new_n22465, new_n22466, new_n22467_1, new_n22468, new_n22469,
    new_n22470_1, new_n22471, new_n22472, new_n22473, new_n22474,
    new_n22475, new_n22476, new_n22477, new_n22478, new_n22479, new_n22480,
    new_n22481, new_n22482, new_n22483, new_n22484_1, new_n22485,
    new_n22486, new_n22487, new_n22488, new_n22489_1, new_n22490,
    new_n22491, new_n22492_1, new_n22493, new_n22494_1, new_n22495,
    new_n22496, new_n22497, new_n22498, new_n22499, new_n22500, new_n22501,
    new_n22502, new_n22503, new_n22504, new_n22505, new_n22506, new_n22507,
    new_n22508, new_n22513, new_n22514, new_n22515, new_n22516, new_n22517,
    new_n22518, new_n22519, new_n22520, new_n22521, new_n22522, new_n22523,
    new_n22524, new_n22525, new_n22526, new_n22527, new_n22528, new_n22529,
    new_n22530, new_n22531, new_n22532, new_n22533_1, new_n22534,
    new_n22535, new_n22536, new_n22537, new_n22538, new_n22539, new_n22540,
    new_n22541, new_n22542, new_n22543, new_n22544, new_n22545, new_n22546,
    new_n22547, new_n22548, new_n22549, new_n22550, new_n22551, new_n22552,
    new_n22553, new_n22554_1, new_n22555, new_n22556, new_n22557,
    new_n22558, new_n22559, new_n22560, new_n22561, new_n22562, new_n22563,
    new_n22564, new_n22565, new_n22566, new_n22567, new_n22568, new_n22569,
    new_n22570, new_n22571, new_n22572, new_n22573, new_n22574, new_n22575,
    new_n22576, new_n22577, new_n22578, new_n22579, new_n22580, new_n22581,
    new_n22582, new_n22583, new_n22584_1, new_n22585, new_n22586,
    new_n22587, new_n22588_1, new_n22589_1, new_n22590, new_n22591_1,
    new_n22592, new_n22593, new_n22594, new_n22595, new_n22596,
    new_n22597_1, new_n22598, new_n22599, new_n22600, new_n22601,
    new_n22602, new_n22603, new_n22604, new_n22605, new_n22606, new_n22607,
    new_n22608, new_n22609, new_n22610, new_n22611, new_n22612, new_n22613,
    new_n22614, new_n22615, new_n22616, new_n22617, new_n22618,
    new_n22619_1, new_n22620_1, new_n22621, new_n22622, new_n22623_1,
    new_n22624, new_n22625, new_n22626_1, new_n22627, new_n22628,
    new_n22629, new_n22630, new_n22631_1, new_n22632, new_n22633,
    new_n22634, new_n22635, new_n22636, new_n22637, new_n22638, new_n22639,
    new_n22640, new_n22641, new_n22642, new_n22643, new_n22644, new_n22646,
    new_n22647, new_n22648, new_n22653, new_n22656, new_n22657, new_n22658,
    new_n22659, new_n22660_1, new_n22661, new_n22662, new_n22663,
    new_n22664, new_n22665, new_n22666, new_n22667, new_n22668, new_n22669,
    new_n22670, new_n22671, new_n22672, new_n22673, new_n22674, new_n22675,
    new_n22676, new_n22677, new_n22678, new_n22679, new_n22680, new_n22681,
    new_n22682, new_n22683, new_n22684, new_n22685, new_n22686, new_n22687,
    new_n22688, new_n22689, new_n22690, new_n22691, new_n22692, new_n22694,
    new_n22695, new_n22696, new_n22697_1, new_n22698, new_n22699,
    new_n22700, new_n22701, new_n22702, new_n22703, new_n22704, new_n22705,
    new_n22706, new_n22707, new_n22708, new_n22709, new_n22710, new_n22711,
    new_n22712, new_n22713, new_n22714_1, new_n22715, new_n22716,
    new_n22717, new_n22718, new_n22719, new_n22720, new_n22721, new_n22722,
    new_n22723, new_n22724, new_n22725, new_n22726, new_n22727, new_n22728,
    new_n22729, new_n22738, new_n22739, new_n22740, new_n22741, new_n22742,
    new_n22743, new_n22744, new_n22745, new_n22746, new_n22747, new_n22748,
    new_n22749, new_n22750, new_n22751, new_n22755, new_n22756, new_n22757,
    new_n22758, new_n22759, new_n22760, new_n22761_1, new_n22762,
    new_n22763, new_n22764_1, new_n22765, new_n22766, new_n22767,
    new_n22768, new_n22769, new_n22770, new_n22771, new_n22772, new_n22773,
    new_n22774, new_n22775, new_n22776, new_n22777, new_n22778,
    new_n22779_1, new_n22780, new_n22781, new_n22782, new_n22783,
    new_n22784, new_n22785, new_n22786, new_n22787_1, new_n22788,
    new_n22789, new_n22792, new_n22793_1, new_n22794, new_n22795,
    new_n22796, new_n22797, new_n22798, new_n22799, new_n22800, new_n22801,
    new_n22802, new_n22803, new_n22804, new_n22805, new_n22806, new_n22807,
    new_n22808, new_n22809, new_n22810, new_n22811, new_n22812, new_n22813,
    new_n22814, new_n22815, new_n22816, new_n22817, new_n22818,
    new_n22819_1, new_n22820, new_n22821, new_n22822, new_n22823,
    new_n22824, new_n22825, new_n22826, new_n22827, new_n22828, new_n22829,
    new_n22830, new_n22831, new_n22832, new_n22833, new_n22834, new_n22835,
    new_n22836, new_n22837, new_n22838, new_n22839, new_n22840, new_n22841,
    new_n22842, new_n22843_1, new_n22844, new_n22845, new_n22846,
    new_n22847, new_n22848, new_n22849, new_n22850, new_n22851, new_n22852,
    new_n22853, new_n22854, new_n22855, new_n22856, new_n22857,
    new_n22858_1, new_n22859, new_n22860, new_n22861, new_n22862,
    new_n22863, new_n22864, new_n22865, new_n22866, new_n22867, new_n22869,
    new_n22870_1, new_n22871_1, new_n22872, new_n22873, new_n22874,
    new_n22875, new_n22876, new_n22877, new_n22878, new_n22879_1,
    new_n22880, new_n22881, new_n22882, new_n22883, new_n22884, new_n22885,
    new_n22886, new_n22887, new_n22888, new_n22889, new_n22890,
    new_n22891_1, new_n22892, new_n22893, new_n22894, new_n22895,
    new_n22896, new_n22897_1, new_n22898, new_n22899, new_n22900,
    new_n22901, new_n22902, new_n22903_1, new_n22904, new_n22905,
    new_n22907_1, new_n22908, new_n22909, new_n22911, new_n22912,
    new_n22913, new_n22914_1, new_n22915, new_n22916, new_n22917,
    new_n22918_1, new_n22919, new_n22920, new_n22921, new_n22922,
    new_n22923, new_n22924, new_n22925, new_n22926, new_n22927, new_n22928,
    new_n22929, new_n22930, new_n22931, new_n22932, new_n22933, new_n22934,
    new_n22935, new_n22936, new_n22937, new_n22938, new_n22939_1,
    new_n22940, new_n22941, new_n22942, new_n22943, new_n22944, new_n22945,
    new_n22946, new_n22947, new_n22948, new_n22951, new_n22952, new_n22953,
    new_n22956, new_n22957, new_n22958, new_n22959, new_n22960, new_n22961,
    new_n22962, new_n22963, new_n22964, new_n22965, new_n22966, new_n22967,
    new_n22968, new_n22969, new_n22970, new_n22971, new_n22972, new_n22973,
    new_n22974, new_n22975, new_n22976, new_n22977, new_n22978, new_n22979,
    new_n22980, new_n22981, new_n22982, new_n22983, new_n22984, new_n22985,
    new_n22986, new_n22987, new_n22988, new_n22989, new_n22990, new_n22991,
    new_n22992, new_n22993, new_n22994, new_n22997, new_n22998_1,
    new_n22999, new_n23000, new_n23001, new_n23002, new_n23003, new_n23004,
    new_n23005, new_n23006_1, new_n23007_1, new_n23008, new_n23009_1,
    new_n23010, new_n23011, new_n23012, new_n23013, new_n23014_1,
    new_n23015, new_n23016, new_n23017, new_n23018, new_n23026, new_n23027,
    new_n23028, new_n23029, new_n23030, new_n23031, new_n23032, new_n23033,
    new_n23034, new_n23035_1, new_n23036, new_n23037, new_n23038,
    new_n23039_1, new_n23040, new_n23041, new_n23042, new_n23043,
    new_n23044, new_n23045, new_n23046, new_n23047_1, new_n23048,
    new_n23049, new_n23050, new_n23051, new_n23052, new_n23053, new_n23054,
    new_n23055, new_n23056, new_n23057, new_n23058_1, new_n23059,
    new_n23060, new_n23061, new_n23062, new_n23063, new_n23064,
    new_n23065_1, new_n23066_1, new_n23067_1, new_n23068_1, new_n23069,
    new_n23070, new_n23071, new_n23072, new_n23073, new_n23074, new_n23075,
    new_n23076, new_n23077, new_n23078, new_n23079, new_n23080, new_n23081,
    new_n23082, new_n23083, new_n23084, new_n23092, new_n23095, new_n23096,
    new_n23097, new_n23098, new_n23099, new_n23100, new_n23101, new_n23102,
    new_n23103, new_n23104, new_n23105, new_n23106, new_n23118, new_n23123,
    new_n23125, new_n23126, new_n23127, new_n23128, new_n23129, new_n23130,
    new_n23131, new_n23132, new_n23133, new_n23134, new_n23135, new_n23136,
    new_n23137, new_n23138, new_n23139, new_n23140, new_n23141, new_n23142,
    new_n23143, new_n23144, new_n23145, new_n23146_1, new_n23148,
    new_n23149, new_n23150, new_n23151, new_n23152, new_n23153, new_n23154,
    new_n23155, new_n23156, new_n23157, new_n23158, new_n23159,
    new_n23160_1, new_n23161, new_n23162, new_n23163, new_n23164,
    new_n23165, new_n23166_1, new_n23167, new_n23168, new_n23169,
    new_n23171, new_n23172, new_n23173, new_n23174, new_n23175, new_n23176,
    new_n23177, new_n23178, new_n23179, new_n23180, new_n23181, new_n23182,
    new_n23183, new_n23184, new_n23185, new_n23186, new_n23191, new_n23192,
    new_n23193, new_n23194, new_n23195, new_n23196, new_n23197, new_n23198,
    new_n23199, new_n23200_1, new_n23201, new_n23202, new_n23203,
    new_n23204, new_n23205, new_n23206, new_n23207, new_n23208, new_n23209,
    new_n23210, new_n23211, new_n23212, new_n23213, new_n23214, new_n23223,
    new_n23224, new_n23225, new_n23226, new_n23227, new_n23228, new_n23229,
    new_n23230, new_n23231, new_n23232, new_n23238_1, new_n23239,
    new_n23240, new_n23241, new_n23242, new_n23243, new_n23244, new_n23245,
    new_n23246, new_n23247_1, new_n23248_1, new_n23253, new_n23259,
    new_n23260, new_n23261, new_n23262, new_n23263, new_n23264, new_n23265,
    new_n23266, new_n23267, new_n23268, new_n23269, new_n23270_1,
    new_n23271, new_n23272_1, new_n23273, new_n23274, new_n23275,
    new_n23276, new_n23277, new_n23282, new_n23283, new_n23284, new_n23285,
    new_n23286, new_n23287, new_n23288, new_n23289_1, new_n23290,
    new_n23291, new_n23298, new_n23299, new_n23300, new_n23301, new_n23302,
    new_n23303, new_n23304_1, new_n23305_1, new_n23306, new_n23307,
    new_n23308, new_n23309, new_n23310, new_n23311, new_n23312, new_n23313,
    new_n23314, new_n23315, new_n23316, new_n23317, new_n23318, new_n23319,
    new_n23320, new_n23321, new_n23322, new_n23323, new_n23324, new_n23325,
    new_n23326, new_n23327, new_n23328, new_n23329, new_n23330, new_n23331,
    new_n23332, new_n23333_1, new_n23334, new_n23335, new_n23336,
    new_n23337, new_n23338, new_n23339, new_n23340, new_n23341_1,
    new_n23342_1, new_n23343, new_n23344, new_n23345, new_n23346,
    new_n23347, new_n23348, new_n23349, new_n23350, new_n23351, new_n23352,
    new_n23355_1, new_n23356, new_n23357, new_n23358, new_n23359,
    new_n23360, new_n23361, new_n23362, new_n23363, new_n23364, new_n23366,
    new_n23367, new_n23368, new_n23369_1, new_n23370, new_n23371_1,
    new_n23372, new_n23373, new_n23374, new_n23375, new_n23376, new_n23377,
    new_n23378, new_n23379, new_n23380, new_n23381, new_n23382, new_n23383,
    new_n23384, new_n23394, new_n23395, new_n23396, new_n23397, new_n23398,
    new_n23399, new_n23400, new_n23401_1, new_n23402, new_n23403,
    new_n23404, new_n23405, new_n23406, new_n23407, new_n23408, new_n23409,
    new_n23410, new_n23411, new_n23412, new_n23413, new_n23414_1,
    new_n23415, new_n23416, new_n23417, new_n23418, new_n23419, new_n23420,
    new_n23421, new_n23422, new_n23423, new_n23424, new_n23425, new_n23426,
    new_n23427, new_n23428, new_n23429_1, new_n23435, new_n23436,
    new_n23437, new_n23438, new_n23448, new_n23449, new_n23450_1,
    new_n23451, new_n23452, new_n23453, new_n23454, new_n23455, new_n23456,
    new_n23457, new_n23458, new_n23459, new_n23460, new_n23461, new_n23462,
    new_n23463_1, new_n23464, new_n23465, new_n23466, new_n23467,
    new_n23468, new_n23469, new_n23470, new_n23471_1, new_n23472,
    new_n23473, new_n23474, new_n23475, new_n23476, new_n23477, new_n23478,
    new_n23479, new_n23480_1, new_n23481, new_n23482, new_n23483,
    new_n23484, new_n23485, new_n23486, new_n23487, new_n23488, new_n23489,
    new_n23490, new_n23491, new_n23492, new_n23493_1, new_n23494,
    new_n23495, new_n23496, new_n23497, new_n23498, new_n23499, new_n23500,
    new_n23501, new_n23502, new_n23503, new_n23504, new_n23505, new_n23506,
    new_n23507, new_n23508, new_n23509, new_n23510, new_n23511, new_n23512,
    new_n23513_1, new_n23514, new_n23515, new_n23516, new_n23517,
    new_n23518, new_n23519, new_n23520, new_n23521, new_n23522, new_n23523,
    new_n23524, new_n23525, new_n23526, new_n23527, new_n23528,
    new_n23529_1, new_n23530, new_n23531, new_n23532, new_n23534,
    new_n23535, new_n23536, new_n23537, new_n23538, new_n23539, new_n23540,
    new_n23541_1, new_n23542, new_n23543, new_n23544, new_n23545,
    new_n23546_1, new_n23547, new_n23548, new_n23549, new_n23550_1,
    new_n23551, new_n23552, new_n23553, new_n23554, new_n23555, new_n23556,
    new_n23557, new_n23558, new_n23559, new_n23560, new_n23561, new_n23562,
    new_n23563, new_n23564, new_n23565, new_n23566, new_n23567, new_n23568,
    new_n23569, new_n23570, new_n23571, new_n23572, new_n23573, new_n23574,
    new_n23575, new_n23576, new_n23577, new_n23578, new_n23579, new_n23580,
    new_n23581, new_n23582, new_n23583, new_n23584, new_n23585_1,
    new_n23586_1, new_n23587, new_n23588_1, new_n23589, new_n23590,
    new_n23591, new_n23592, new_n23593, new_n23594, new_n23595, new_n23596,
    new_n23597, new_n23598, new_n23599, new_n23600, new_n23601, new_n23602,
    new_n23603, new_n23604, new_n23605, new_n23606, new_n23607, new_n23608,
    new_n23609, new_n23610, new_n23611, new_n23614, new_n23615, new_n23616,
    new_n23617, new_n23618, new_n23619_1, new_n23620, new_n23621,
    new_n23622, new_n23623, new_n23624_1, new_n23625, new_n23626,
    new_n23627, new_n23628_1, new_n23629, new_n23630, new_n23632,
    new_n23637_1, new_n23638, new_n23639, new_n23640, new_n23641,
    new_n23642, new_n23643, new_n23644, new_n23645, new_n23646, new_n23647,
    new_n23648, new_n23649, new_n23650, new_n23651, new_n23652, new_n23653,
    new_n23654, new_n23655, new_n23656, new_n23657_1, new_n23658,
    new_n23659, new_n23660, new_n23661, new_n23662, new_n23663_1,
    new_n23664, new_n23665, new_n23666, new_n23667, new_n23668,
    new_n23669_1, new_n23670, new_n23671, new_n23672, new_n23673,
    new_n23674, new_n23675, new_n23676, new_n23677, new_n23678, new_n23679,
    new_n23680, new_n23681, new_n23682, new_n23683, new_n23684_1,
    new_n23685, new_n23686, new_n23687, new_n23688, new_n23689,
    new_n23690_1, new_n23691, new_n23692, new_n23693, new_n23694,
    new_n23695, new_n23696, new_n23697_1, new_n23698, new_n23699,
    new_n23700, new_n23701, new_n23702, new_n23703, new_n23704, new_n23705,
    new_n23706, new_n23707, new_n23708, new_n23709, new_n23710, new_n23711,
    new_n23712, new_n23713, new_n23714_1, new_n23715, new_n23716,
    new_n23717_1, new_n23718, new_n23719_1, new_n23720, new_n23721,
    new_n23722, new_n23723, new_n23724, new_n23725, new_n23726, new_n23727,
    new_n23728, new_n23729, new_n23730, new_n23731, new_n23732, new_n23734,
    new_n23735, new_n23736, new_n23737, new_n23738, new_n23739, new_n23740,
    new_n23741, new_n23742, new_n23743, new_n23744, new_n23745,
    new_n23748_1, new_n23749, new_n23750, new_n23751, new_n23752,
    new_n23753, new_n23754, new_n23755_1, new_n23756, new_n23757,
    new_n23758, new_n23759, new_n23765, new_n23766, new_n23767, new_n23768,
    new_n23769, new_n23770, new_n23771, new_n23772, new_n23773, new_n23774,
    new_n23775_1, new_n23776, new_n23777, new_n23778, new_n23779,
    new_n23780, new_n23781, new_n23782, new_n23783, new_n23784, new_n23785,
    new_n23786, new_n23787, new_n23788, new_n23789, new_n23790, new_n23791,
    new_n23792, new_n23793, new_n23794, new_n23795, new_n23796, new_n23797,
    new_n23798, new_n23799, new_n23800, new_n23801, new_n23802, new_n23803,
    new_n23804, new_n23805, new_n23806, new_n23807, new_n23808, new_n23809,
    new_n23810, new_n23811, new_n23812, new_n23813, new_n23814, new_n23815,
    new_n23816, new_n23817, new_n23818, new_n23819, new_n23820, new_n23821,
    new_n23822, new_n23823, new_n23824, new_n23825, new_n23826, new_n23827,
    new_n23828, new_n23829, new_n23830, new_n23831_1, new_n23832,
    new_n23833, new_n23834, new_n23835, new_n23836, new_n23837, new_n23838,
    new_n23839, new_n23840, new_n23841, new_n23842_1, new_n23843,
    new_n23844, new_n23845, new_n23846, new_n23847, new_n23848,
    new_n23849_1, new_n23850, new_n23857, new_n23859, new_n23860,
    new_n23861, new_n23862, new_n23863, new_n23864, new_n23869, new_n23872,
    new_n23874, new_n23875, new_n23876, new_n23877, new_n23878, new_n23879,
    new_n23880, new_n23881, new_n23882, new_n23883_1, new_n23884,
    new_n23885, new_n23886, new_n23887, new_n23888_1, new_n23889,
    new_n23890, new_n23891, new_n23892, new_n23893, new_n23894,
    new_n23895_1, new_n23896, new_n23897, new_n23898, new_n23899_1,
    new_n23900, new_n23901, new_n23902, new_n23903_1, new_n23904,
    new_n23905, new_n23906, new_n23907, new_n23908, new_n23909, new_n23910,
    new_n23911, new_n23912_1, new_n23913_1, new_n23914, new_n23915,
    new_n23916, new_n23917, new_n23918, new_n23919, new_n23920, new_n23921,
    new_n23922, new_n23923_1, new_n23924_1, new_n23925, new_n23926,
    new_n23927, new_n23928, new_n23929, new_n23930, new_n23931, new_n23934,
    new_n23935_1, new_n23936, new_n23937, new_n23938, new_n23946,
    new_n23947, new_n23948, new_n23949, new_n23950, new_n23951, new_n23952,
    new_n23953, new_n23954_1, new_n23955, new_n23956, new_n23960,
    new_n23968, new_n23969, new_n23970, new_n23971, new_n23972, new_n23973,
    new_n23974_1, new_n23975, new_n23976, new_n23977, new_n23978,
    new_n23979, new_n23980, new_n23981, new_n23982, new_n23983, new_n23984,
    new_n23985, new_n23986_1, new_n23988, new_n23989, new_n23990,
    new_n23991, new_n23992, new_n23993, new_n23994, new_n23995, new_n23996,
    new_n23997, new_n23998, new_n23999, new_n24000, new_n24001,
    new_n24002_1, new_n24003, new_n24004_1, new_n24005, new_n24006,
    new_n24007, new_n24013, new_n24014, new_n24015, new_n24016, new_n24017,
    new_n24018, new_n24019, new_n24020, new_n24021, new_n24022, new_n24023,
    new_n24024, new_n24025, new_n24026, new_n24027, new_n24028, new_n24029,
    new_n24030, new_n24031, new_n24032_1, new_n24033, new_n24034,
    new_n24035, new_n24036, new_n24037, new_n24038, new_n24039_1,
    new_n24040, new_n24043, new_n24044, new_n24045, new_n24046, new_n24047,
    new_n24048_1, new_n24049, new_n24050, new_n24051, new_n24052_1,
    new_n24053, new_n24054, new_n24055, new_n24056, new_n24057, new_n24058,
    new_n24059, new_n24060, new_n24061, new_n24062, new_n24063, new_n24064,
    new_n24065, new_n24066, new_n24067, new_n24068, new_n24070, new_n24071,
    new_n24072, new_n24073, new_n24074, new_n24075, new_n24076, new_n24077,
    new_n24078, new_n24079, new_n24080, new_n24081, new_n24082, new_n24086,
    new_n24088, new_n24089, new_n24090, new_n24095, new_n24096_1,
    new_n24097_1, new_n24098, new_n24099, new_n24100, new_n24101,
    new_n24102, new_n24103, new_n24104, new_n24105_1, new_n24106,
    new_n24107, new_n24108, new_n24109, new_n24110, new_n24111, new_n24112,
    new_n24113, new_n24114, new_n24115, new_n24116, new_n24117, new_n24118,
    new_n24119_1, new_n24120, new_n24121, new_n24122, new_n24123,
    new_n24124, new_n24125, new_n24126, new_n24127, new_n24128,
    new_n24129_1, new_n24130, new_n24131, new_n24132, new_n24133_1,
    new_n24134, new_n24135, new_n24136, new_n24137, new_n24138, new_n24139,
    new_n24140, new_n24141_1, new_n24142, new_n24143, new_n24145_1,
    new_n24146_1, new_n24147, new_n24148, new_n24149, new_n24150_1,
    new_n24151, new_n24152, new_n24153, new_n24154, new_n24155_1,
    new_n24156, new_n24157, new_n24158, new_n24159, new_n24160_1,
    new_n24161, new_n24162, new_n24163, new_n24164, new_n24165, new_n24166,
    new_n24167_1, new_n24168, new_n24169, new_n24170_1, new_n24171,
    new_n24172_1, new_n24173, new_n24174, new_n24175, new_n24176,
    new_n24177_1, new_n24178, new_n24179, new_n24180, new_n24181,
    new_n24182, new_n24183, new_n24184, new_n24185, new_n24186, new_n24187,
    new_n24188, new_n24189, new_n24190, new_n24191, new_n24192, new_n24193,
    new_n24194, new_n24195, new_n24196_1, new_n24197, new_n24198,
    new_n24204, new_n24213, new_n24214, new_n24215, new_n24216, new_n24217,
    new_n24221, new_n24224, new_n24231, new_n24232, new_n24233, new_n24234,
    new_n24235, new_n24236, new_n24237, new_n24238, new_n24239, new_n24240,
    new_n24241, new_n24242, new_n24243, new_n24244, new_n24245, new_n24246,
    new_n24247, new_n24248, new_n24249, new_n24250, new_n24251, new_n24252,
    new_n24253, new_n24254, new_n24255, new_n24256, new_n24257,
    new_n24258_1, new_n24259, new_n24260_1, new_n24261, new_n24262,
    new_n24263, new_n24264, new_n24265, new_n24266, new_n24267, new_n24268,
    new_n24269, new_n24270, new_n24272, new_n24274, new_n24275, new_n24276,
    new_n24277, new_n24278_1, new_n24279, new_n24280, new_n24281,
    new_n24282, new_n24283, new_n24284, new_n24285, new_n24286, new_n24293,
    new_n24294, new_n24295, new_n24296, new_n24297_1, new_n24298,
    new_n24299, new_n24300, new_n24301, new_n24302, new_n24303, new_n24304,
    new_n24305, new_n24306, new_n24307_1, new_n24308, new_n24309,
    new_n24310, new_n24311, new_n24312, new_n24313, new_n24314, new_n24315,
    new_n24316, new_n24317, new_n24318, new_n24319_1, new_n24320,
    new_n24321, new_n24322, new_n24323_1, new_n24324, new_n24325,
    new_n24326, new_n24327_1, new_n24328, new_n24329, new_n24330,
    new_n24331, new_n24332, new_n24333, new_n24334, new_n24335, new_n24336,
    new_n24337, new_n24338, new_n24339, new_n24340, new_n24341,
    new_n24342_1, new_n24343, new_n24344, new_n24345_1, new_n24346,
    new_n24347_1, new_n24348, new_n24349, new_n24350, new_n24351,
    new_n24352, new_n24353, new_n24354, new_n24355, new_n24356, new_n24357,
    new_n24358, new_n24359, new_n24360, new_n24361, new_n24362, new_n24363,
    new_n24364, new_n24365, new_n24366, new_n24367, new_n24368, new_n24369,
    new_n24370, new_n24371, new_n24372, new_n24373_1, new_n24374_1,
    new_n24375, new_n24376, new_n24377, new_n24378, new_n24379, new_n24380,
    new_n24381, new_n24382, new_n24383, new_n24384, new_n24385, new_n24386,
    new_n24387, new_n24388, new_n24389, new_n24390, new_n24391, new_n24392,
    new_n24393, new_n24394, new_n24395, new_n24396, new_n24397, new_n24398,
    new_n24399, new_n24400, new_n24401, new_n24402, new_n24403, new_n24404,
    new_n24405, new_n24406_1, new_n24407, new_n24408, new_n24409,
    new_n24410, new_n24411, new_n24412, new_n24413, new_n24414,
    new_n24415_1, new_n24416, new_n24417, new_n24418, new_n24419,
    new_n24420, new_n24421_1, new_n24422, new_n24423, new_n24424,
    new_n24425, new_n24426, new_n24427, new_n24428, new_n24429, new_n24430,
    new_n24431_1, new_n24432, new_n24433, new_n24434, new_n24435,
    new_n24436, new_n24440, new_n24443, new_n24444, new_n24445, new_n24446,
    new_n24447, new_n24448, new_n24449, new_n24450, new_n24451, new_n24452,
    new_n24453, new_n24454, new_n24455, new_n24456, new_n24457, new_n24458,
    new_n24459, new_n24464, new_n24465, new_n24466, new_n24467, new_n24468,
    new_n24469, new_n24470, new_n24471, new_n24472_1, new_n24473,
    new_n24474, new_n24475, new_n24476_1, new_n24477, new_n24478,
    new_n24479, new_n24480, new_n24481, new_n24482, new_n24483_1,
    new_n24484, new_n24485_1, new_n24486, new_n24487, new_n24488,
    new_n24489, new_n24490, new_n24492, new_n24493, new_n24494, new_n24495,
    new_n24496, new_n24497, new_n24498, new_n24499, new_n24503, new_n24504,
    new_n24505, new_n24506, new_n24516, new_n24517, new_n24518, new_n24519,
    new_n24520, new_n24521, new_n24522, new_n24523, new_n24524, new_n24525,
    new_n24526, new_n24527, new_n24528, new_n24529, new_n24530, new_n24531,
    new_n24532, new_n24533, new_n24534, new_n24535, new_n24536, new_n24537,
    new_n24538, new_n24539, new_n24540, new_n24541, new_n24542, new_n24552,
    new_n24564, new_n24565, new_n24566, new_n24567, new_n24568, new_n24569,
    new_n24570, new_n24571, new_n24572, new_n24573, new_n24574, new_n24575,
    new_n24576_1, new_n24577, new_n24578, new_n24579_1, new_n24580,
    new_n24581, new_n24582, new_n24583, new_n24584, new_n24585, new_n24586,
    new_n24587, new_n24588, new_n24589, new_n24590, new_n24591, new_n24592,
    new_n24593, new_n24594, new_n24595, new_n24596, new_n24597, new_n24598,
    new_n24599, new_n24600, new_n24601, new_n24602_1, new_n24603,
    new_n24604_1, new_n24605, new_n24613, new_n24614, new_n24615,
    new_n24616, new_n24617, new_n24618_1, new_n24619, new_n24620_1,
    new_n24621, new_n24622, new_n24623, new_n24624, new_n24625,
    new_n24626_1, new_n24627, new_n24628, new_n24632, new_n24633,
    new_n24634, new_n24637, new_n24638_1, new_n24639, new_n24640,
    new_n24641, new_n24642, new_n24643, new_n24644, new_n24645, new_n24647,
    new_n24649, new_n24650, new_n24651, new_n24652, new_n24653, new_n24654,
    new_n24655, new_n24656, new_n24657, new_n24658, new_n24659, new_n24660,
    new_n24661, new_n24662, new_n24663, new_n24664, new_n24665, new_n24666,
    new_n24667, new_n24668, new_n24669, new_n24670, new_n24673, new_n24674,
    new_n24675, new_n24676, new_n24677, new_n24678, new_n24679, new_n24680,
    new_n24681, new_n24682, new_n24683, new_n24684, new_n24685, new_n24686,
    new_n24687, new_n24688, new_n24689, new_n24690, new_n24691, new_n24692,
    new_n24693, new_n24694, new_n24695, new_n24696, new_n24697, new_n24698,
    new_n24699, new_n24700, new_n24701, new_n24702, new_n24703, new_n24704,
    new_n24705, new_n24706, new_n24707, new_n24708, new_n24709, new_n24710,
    new_n24711, new_n24712, new_n24713, new_n24734, new_n24738, new_n24739,
    new_n24740, new_n24741, new_n24742, new_n24743, new_n24744, new_n24745,
    new_n24746, new_n24747, new_n24748, new_n24749_1, new_n24750,
    new_n24751, new_n24752, new_n24755, new_n24756, new_n24757,
    new_n24758_1, new_n24759, new_n24760, new_n24761, new_n24762,
    new_n24763, new_n24764, new_n24765, new_n24766, new_n24767,
    new_n24768_1, new_n24769, new_n24770, new_n24771, new_n24772,
    new_n24773, new_n24774, new_n24775, new_n24776, new_n24777, new_n24778,
    new_n24779, new_n24783, new_n24784_1, new_n24785, new_n24786_1,
    new_n24787, new_n24788, new_n24789, new_n24790, new_n24794, new_n24799,
    new_n24800, new_n24801, new_n24802, new_n24803, new_n24804, new_n24805,
    new_n24806, new_n24808, new_n24809, new_n24810, new_n24811, new_n24812,
    new_n24813, new_n24814, new_n24815, new_n24816, new_n24817, new_n24818,
    new_n24819, new_n24820, new_n24821, new_n24822, new_n24823, new_n24824,
    new_n24825, new_n24846, new_n24849, new_n24850, new_n24851, new_n24852,
    new_n24853_1, new_n24854, new_n24855, new_n24856, new_n24857_1,
    new_n24858, new_n24859, new_n24860, new_n24861, new_n24862, new_n24863,
    new_n24864, new_n24865, new_n24866, new_n24867, new_n24868, new_n24869,
    new_n24870, new_n24871, new_n24872, new_n24873, new_n24874, new_n24875,
    new_n24880, new_n24881, new_n24882, new_n24883, new_n24884, new_n24896,
    new_n24899, new_n24914, new_n24915, new_n24916, new_n24917, new_n24918,
    new_n24919, new_n24933, new_n24934_1, new_n24935, new_n24936,
    new_n24937_1, new_n24938, new_n24939, new_n24940, new_n24941,
    new_n24945, new_n24946, new_n24947, new_n24948, new_n24949, new_n24950,
    new_n24951, new_n24952, new_n24953, new_n24958, new_n24959, new_n24960,
    new_n24961, new_n24962, new_n24963, new_n24964, new_n24965, new_n24966,
    new_n24967, new_n24968, new_n24971, new_n24972, new_n24973, new_n24988,
    new_n24989, new_n24990, new_n24991, new_n24994, new_n24995, new_n24996,
    new_n24997, new_n24998_1, new_n25005, new_n25007, new_n25008,
    new_n25009, new_n25015, new_n25019, new_n25029, new_n25030, new_n25031,
    new_n25032_1, new_n25033, new_n25034, new_n25035, new_n25036,
    new_n25037, new_n25038, new_n25039, new_n25048, new_n25049, new_n25050,
    new_n25051, new_n25052, new_n25053, new_n25054, new_n25055, new_n25056,
    new_n25057, new_n25058, new_n25059, new_n25060, new_n25061, new_n25063,
    new_n25064, new_n25065, new_n25066, new_n25067, new_n25068_1,
    new_n25069, new_n25070, new_n25071, new_n25082, new_n25083_1,
    new_n25085, new_n25086, new_n25087, new_n25088, new_n25089, new_n25090,
    new_n25091, new_n25092, new_n25093, new_n25094_1, new_n25095,
    new_n25096, new_n25097_1, new_n25098, new_n25099, new_n25100,
    new_n25101, new_n25102, new_n25120_1, new_n25121, new_n25122,
    new_n25123, new_n25124, new_n25125, new_n25126_1, new_n25127,
    new_n25128, new_n25129, new_n25130, new_n25131, new_n25132,
    new_n25133_1, new_n25134, new_n25135, new_n25136, new_n25139,
    new_n25140, new_n25141, new_n25142, new_n25147, new_n25148, new_n25149,
    new_n25150, new_n25151, new_n25152, new_n25153, new_n25154, new_n25157,
    new_n25158, new_n25159, new_n25160, new_n25161, new_n25162, new_n25163,
    new_n25164, new_n25167, new_n25168_1, new_n25169, new_n25170,
    new_n25171, new_n25172, new_n25173, new_n25175, new_n25176, new_n25177,
    new_n25178, new_n25179, new_n25180, new_n25181_1, new_n25182,
    new_n25183, new_n25184, new_n25185, new_n25186, new_n25187, new_n25188,
    new_n25189, new_n25190, new_n25191, new_n25192, new_n25193, new_n25194,
    new_n25195, new_n25196, new_n25197, new_n25198, new_n25202, new_n25203,
    new_n25204, new_n25205, new_n25206, new_n25207, new_n25208, new_n25222,
    new_n25223, new_n25234, new_n25241, new_n25242, new_n25243,
    new_n25244_1, new_n25245, new_n25246, new_n25247, new_n25255,
    new_n25258, new_n25275, new_n25295, new_n25298, new_n25299, new_n25300,
    new_n25314, new_n25315, new_n25316_1, new_n25317, new_n25318,
    new_n25319, new_n25320, new_n25321, new_n25322, new_n25323, new_n25324,
    new_n25326, new_n25332_1, new_n25340, new_n25341, new_n25342,
    new_n25343, new_n25344, new_n25345_1, new_n25346, new_n25347,
    new_n25348, new_n25349, new_n25350, new_n25351, new_n25352, new_n25353,
    new_n25354, new_n25360, new_n25361, new_n25362_1, new_n25363,
    new_n25364, new_n25365_1, new_n25366, new_n25367, new_n25368,
    new_n25369, new_n25370_1, new_n25373, new_n25374, new_n25375,
    new_n25376, new_n25377, new_n25383, new_n25384, new_n25385, new_n25386,
    new_n25388, new_n25389, new_n25390, new_n25391, new_n25392, new_n25393,
    new_n25394, new_n25395, new_n25396, new_n25397, new_n25398, new_n25399,
    new_n25400, new_n25401, new_n25402, new_n25403, new_n25404, new_n25405,
    new_n25417, new_n25418, new_n25419, new_n25420, new_n25421, new_n25422,
    new_n25423, new_n25424, new_n25425, new_n25453, new_n25454, new_n25455,
    new_n25456, new_n25457, new_n25468_1, new_n25474, new_n25475_1,
    new_n25476, new_n25477, new_n25478, new_n25479, new_n25492, new_n25495,
    new_n25502, new_n25503, new_n25504, new_n25505, new_n25506, new_n25507,
    new_n25508, new_n25509, new_n25510, new_n25511, new_n25517, new_n25527,
    new_n25528, new_n25529, new_n25530, new_n25531, new_n25532_1,
    new_n25533, new_n25534, new_n25535, new_n25536, new_n25541, new_n25544,
    new_n25548, new_n25549, new_n25550_1, new_n25551, new_n25552,
    new_n25553, new_n25554, new_n25555, new_n25556, new_n25557, new_n25558,
    new_n25562, new_n25572, new_n25573, new_n25574, new_n25575, new_n25579,
    new_n25584, new_n25585, new_n25586_1, new_n25587, new_n25594,
    new_n25595, new_n25596, new_n25597, new_n25598, new_n25599, new_n25600,
    new_n25601, new_n25607, new_n25608, new_n25616, new_n25617, new_n25618,
    new_n25619_1, new_n25620, new_n25621, new_n25622, new_n25625,
    new_n25626, new_n25627, new_n25630, new_n25631, new_n25632, new_n25633,
    new_n25634, new_n25635, new_n25636, new_n25637, new_n25638, new_n25651,
    new_n25652, new_n25653, new_n25654, new_n25655, new_n25657, new_n25658,
    new_n25669, new_n25670, new_n25671, new_n25672, new_n25673, new_n25676,
    new_n25684, new_n25685, new_n25686, new_n25687, new_n25688, new_n25689,
    new_n25690, new_n25691, new_n25692, new_n25694_1, new_n25699,
    new_n25700, new_n25701, new_n25702, new_n25704, new_n25705,
    new_n25706_1, new_n25707, new_n25712, new_n25713, new_n25714,
    new_n25715, new_n25716, new_n25717, new_n25718, new_n25719_1,
    new_n25720, new_n25721, new_n25722, new_n25723, new_n25724, new_n25725,
    new_n25726, new_n25727, new_n25728, new_n25729, new_n25730, new_n25731,
    new_n25732, new_n25733, new_n25734, new_n25735, new_n25736, new_n25737,
    new_n25738_1, new_n25739, new_n25740, new_n25745, new_n25746,
    new_n25747, new_n25748, new_n25749_1, new_n25753, new_n25763,
    new_n25764, new_n25765, new_n25766, new_n25767, new_n25768, new_n25769,
    new_n25782, new_n25789, new_n25790, new_n25791, new_n25792_1,
    new_n25793, new_n25794, new_n25795, new_n25797_1, new_n25798,
    new_n25799, new_n25800, new_n25801, new_n25802, new_n25803, new_n25814,
    new_n25826_1, new_n25827, new_n25828, new_n25832, new_n25833,
    new_n25834, new_n25835, new_n25836, new_n25838, new_n25839_1,
    new_n25840_1, new_n25841, new_n25843, new_n25853, new_n25854,
    new_n25855, new_n25856, new_n25857, new_n25858, new_n25859, new_n25860,
    new_n25861, new_n25870, new_n25871, new_n25882, new_n25891, new_n25899,
    new_n25901, new_n25902, new_n25912, new_n25913, new_n25914, new_n25915,
    new_n25916, new_n25922, new_n25923_1, new_n25924, new_n25925,
    new_n25928, new_n25929, new_n25930, new_n25931, new_n25932, new_n25949,
    new_n25954, new_n25974_1, new_n25984, new_n25985_1, new_n25986,
    new_n26000, new_n26001, new_n26016, new_n26032, new_n26037, new_n26040,
    new_n26041, new_n26047, new_n26048, new_n26049, new_n26053_1,
    new_n26054_1, new_n26055, new_n26056, new_n26057, new_n26059,
    new_n26072, new_n26075, new_n26076, new_n26077, new_n26078, new_n26079,
    new_n26082, new_n26085, new_n26086, new_n26087, new_n26088, new_n26089,
    new_n26090, new_n26104, new_n26105, new_n26106, new_n26109, new_n26119,
    new_n26122, new_n26124, new_n26125, new_n26126, new_n26127, new_n26128,
    new_n26131, new_n26132, new_n26133, new_n26134, new_n26144, new_n26146,
    new_n26151, new_n26152, new_n26153, new_n26154, new_n26160, new_n26161,
    new_n26162, new_n26164, new_n26173, new_n26187, new_n26196, new_n26197,
    new_n26198, new_n26201;
xnor_4 g00000(n10739, n9942, new_n2349);
not_8  g00001(n21753, new_n2350);
or_5   g00002(n25643, new_n2350, new_n2351);
xnor_4 g00003(n25643, n21753, new_n2352);
not_8  g00004(n21832, new_n2353);
nor_5  g00005(new_n2353, n9557, new_n2354);
xnor_4 g00006(n21832, n9557, new_n2355_1);
not_8  g00007(n26913, new_n2356);
nor_5  g00008(new_n2356, n3136, new_n2357);
not_8  g00009(new_n2357, new_n2358);
xnor_4 g00010(n26913, n3136, new_n2359);
not_8  g00011(n6385, new_n2360);
nor_5  g00012(n16223, new_n2360, new_n2361_1);
not_8  g00013(n16223, new_n2362);
nor_5  g00014(new_n2362, n6385, new_n2363_1);
not_8  g00015(n20138, new_n2364);
nor_5  g00016(new_n2364, n19494, new_n2365);
not_8  g00017(n19494, new_n2366);
nor_5  g00018(n20138, new_n2366, new_n2367);
not_8  g00019(n2387, new_n2368);
nand_5 g00020(n9251, new_n2368, new_n2369);
nor_5  g00021(new_n2369, new_n2367, new_n2370);
nor_5  g00022(new_n2370, new_n2365, new_n2371);
nor_5  g00023(new_n2371, new_n2363_1, new_n2372);
nor_5  g00024(new_n2372, new_n2361_1, new_n2373);
nand_5 g00025(new_n2373, new_n2359, new_n2374_1);
nand_5 g00026(new_n2374_1, new_n2358, new_n2375);
and_5  g00027(new_n2375, new_n2355_1, new_n2376);
nor_5  g00028(new_n2376, new_n2354, new_n2377);
not_8  g00029(new_n2377, new_n2378);
nand_5 g00030(new_n2378, new_n2352, new_n2379);
nand_5 g00031(new_n2379, new_n2351, new_n2380);
xnor_4 g00032(new_n2380, new_n2349, new_n2381);
xnor_4 g00033(n13781, n5704, new_n2382);
not_8  g00034(new_n2382, new_n2383);
nand_5 g00035(n13781, n5704, new_n2384);
not_8  g00036(new_n2384, new_n2385);
xnor_4 g00037(n18409, n11486, new_n2386);
xnor_4 g00038(new_n2386, new_n2385, new_n2387_1);
nor_5  g00039(new_n2387_1, new_n2383, new_n2388_1);
not_8  g00040(new_n2388_1, new_n2389);
not_8  g00041(n13708, new_n2390);
xnor_4 g00042(n16722, new_n2390, new_n2391);
nor_5  g00043(n18409, n11486, new_n2392);
nor_5  g00044(new_n2386, new_n2385, new_n2393);
nor_5  g00045(new_n2393, new_n2392, new_n2394);
xnor_4 g00046(new_n2394, new_n2391, new_n2395);
not_8  g00047(new_n2395, new_n2396);
nor_5  g00048(new_n2396, new_n2389, new_n2397);
not_8  g00049(n3480, new_n2398);
xnor_4 g00050(n19911, new_n2398, new_n2399);
nor_5  g00051(n16722, n13708, new_n2400);
not_8  g00052(new_n2391, new_n2401);
nor_5  g00053(new_n2394, new_n2401, new_n2402);
nor_5  g00054(new_n2402, new_n2400, new_n2403);
xnor_4 g00055(new_n2403, new_n2399, new_n2404);
nand_5 g00056(new_n2404, new_n2397, new_n2405);
not_8  g00057(n2731, new_n2406);
xnor_4 g00058(n3018, new_n2406, new_n2407);
not_8  g00059(new_n2407, new_n2408);
nor_5  g00060(n19911, n3480, new_n2409_1);
not_8  g00061(new_n2399, new_n2410);
nor_5  g00062(new_n2403, new_n2410, new_n2411);
nor_5  g00063(new_n2411, new_n2409_1, new_n2412);
xnor_4 g00064(new_n2412, new_n2408, new_n2413);
nor_5  g00065(new_n2413, new_n2405, new_n2414);
not_8  g00066(n18907, new_n2415);
xnor_4 g00067(n26660, new_n2415, new_n2416_1);
nor_5  g00068(n3018, n2731, new_n2417);
nor_5  g00069(new_n2412, new_n2408, new_n2418);
nor_5  g00070(new_n2418, new_n2417, new_n2419);
xnor_4 g00071(new_n2419, new_n2416_1, new_n2420_1);
nand_5 g00072(new_n2420_1, new_n2414, new_n2421_1);
not_8  g00073(n13783, new_n2422);
xnor_4 g00074(n22332, new_n2422, new_n2423);
nor_5  g00075(n26660, n18907, new_n2424);
not_8  g00076(new_n2416_1, new_n2425);
nor_5  g00077(new_n2419, new_n2425, new_n2426);
nor_5  g00078(new_n2426, new_n2424, new_n2427);
xnor_4 g00079(new_n2427, new_n2423, new_n2428);
xnor_4 g00080(new_n2428, new_n2421_1, new_n2429);
not_8  g00081(n7751, new_n2430);
xnor_4 g00082(n13490, new_n2430, new_n2431);
not_8  g00083(new_n2431, new_n2432);
not_8  g00084(n22660, new_n2433);
not_8  g00085(n26823, new_n2434);
nand_5 g00086(new_n2434, new_n2433, new_n2435);
xnor_4 g00087(n26823, new_n2433, new_n2436);
not_8  g00088(n1777, new_n2437);
not_8  g00089(n4812, new_n2438);
nand_5 g00090(new_n2438, new_n2437, new_n2439);
xnor_4 g00091(n4812, new_n2437, new_n2440_1);
not_8  g00092(n8745, new_n2441);
not_8  g00093(n24278, new_n2442);
nand_5 g00094(new_n2442, new_n2441, new_n2443);
xnor_4 g00095(n24278, new_n2441, new_n2444_1);
not_8  g00096(n15636, new_n2445);
not_8  g00097(n24618, new_n2446);
nand_5 g00098(new_n2446, new_n2445, new_n2447);
xnor_4 g00099(n24618, n15636, new_n2448);
not_8  g00100(new_n2448, new_n2449);
nand_5 g00101(n20077, n3952, new_n2450);
not_8  g00102(new_n2450, new_n2451);
nor_5  g00103(n20077, n3952, new_n2452);
nand_5 g00104(n12315, n6794, new_n2453);
nor_5  g00105(new_n2453, new_n2452, new_n2454);
nor_5  g00106(new_n2454, new_n2451, new_n2455);
nand_5 g00107(new_n2455, new_n2449, new_n2456);
nand_5 g00108(new_n2456, new_n2447, new_n2457);
nand_5 g00109(new_n2457, new_n2444_1, new_n2458);
nand_5 g00110(new_n2458, new_n2443, new_n2459);
nand_5 g00111(new_n2459, new_n2440_1, new_n2460);
nand_5 g00112(new_n2460, new_n2439, new_n2461);
nand_5 g00113(new_n2461, new_n2436, new_n2462);
nand_5 g00114(new_n2462, new_n2435, new_n2463);
xnor_4 g00115(new_n2463, new_n2432, new_n2464);
xnor_4 g00116(new_n2464, new_n2429, new_n2465);
not_8  g00117(new_n2420_1, new_n2466);
xnor_4 g00118(new_n2466, new_n2414, new_n2467);
not_8  g00119(new_n2467, new_n2468);
not_8  g00120(new_n2436, new_n2469);
xnor_4 g00121(new_n2461, new_n2469, new_n2470);
nand_5 g00122(new_n2470, new_n2468, new_n2471);
not_8  g00123(new_n2413, new_n2472);
xnor_4 g00124(new_n2472, new_n2405, new_n2473);
not_8  g00125(new_n2473, new_n2474);
not_8  g00126(new_n2440_1, new_n2475);
xnor_4 g00127(new_n2459, new_n2475, new_n2476);
nand_5 g00128(new_n2476, new_n2474, new_n2477);
xnor_4 g00129(new_n2476, new_n2473, new_n2478);
xnor_4 g00130(new_n2404, new_n2397, new_n2479_1);
not_8  g00131(new_n2444_1, new_n2480);
xnor_4 g00132(new_n2457, new_n2480, new_n2481);
nand_5 g00133(new_n2481, new_n2479_1, new_n2482);
not_8  g00134(new_n2482, new_n2483);
xnor_4 g00135(new_n2395, new_n2388_1, new_n2484);
xnor_4 g00136(new_n2455, new_n2448, new_n2485);
nand_5 g00137(new_n2485, new_n2484, new_n2486);
not_8  g00138(new_n2486, new_n2487);
xnor_4 g00139(new_n2485, new_n2484, new_n2488);
xnor_4 g00140(n12315, n6794, new_n2489);
nor_5  g00141(new_n2489, new_n2382, new_n2490);
xnor_4 g00142(n20077, n3952, new_n2491);
xnor_4 g00143(new_n2491, new_n2453, new_n2492);
not_8  g00144(new_n2492, new_n2493);
nor_5  g00145(new_n2493, new_n2490, new_n2494);
nor_5  g00146(n13781, n5704, new_n2495);
not_8  g00147(new_n2393, new_n2496);
nor_5  g00148(new_n2496, new_n2495, new_n2497);
nor_5  g00149(new_n2497, new_n2388_1, new_n2498);
not_8  g00150(new_n2491, new_n2499);
nand_5 g00151(new_n2499, new_n2490, new_n2500);
not_8  g00152(new_n2500, new_n2501);
nor_5  g00153(new_n2501, new_n2494, new_n2502);
not_8  g00154(new_n2502, new_n2503);
nor_5  g00155(new_n2503, new_n2498, new_n2504);
nor_5  g00156(new_n2504, new_n2494, new_n2505);
nor_5  g00157(new_n2505, new_n2488, new_n2506);
nor_5  g00158(new_n2506, new_n2487, new_n2507);
xnor_4 g00159(new_n2481, new_n2479_1, new_n2508);
nor_5  g00160(new_n2508, new_n2507, new_n2509);
nor_5  g00161(new_n2509, new_n2483, new_n2510);
not_8  g00162(new_n2510, new_n2511);
nand_5 g00163(new_n2511, new_n2478, new_n2512);
nand_5 g00164(new_n2512, new_n2477, new_n2513_1);
xnor_4 g00165(new_n2470, new_n2467, new_n2514);
nand_5 g00166(new_n2514, new_n2513_1, new_n2515_1);
nand_5 g00167(new_n2515_1, new_n2471, new_n2516);
xnor_4 g00168(new_n2516, new_n2465, new_n2517);
not_8  g00169(new_n2517, new_n2518);
xnor_4 g00170(new_n2518, new_n2381, new_n2519);
xnor_4 g00171(new_n2377, new_n2352, new_n2520);
not_8  g00172(new_n2520, new_n2521);
not_8  g00173(new_n2514, new_n2522);
xnor_4 g00174(new_n2522, new_n2513_1, new_n2523);
nand_5 g00175(new_n2523, new_n2521, new_n2524);
xnor_4 g00176(new_n2523, new_n2520, new_n2525);
not_8  g00177(new_n2355_1, new_n2526);
xnor_4 g00178(new_n2375, new_n2526, new_n2527);
not_8  g00179(new_n2527, new_n2528);
xnor_4 g00180(new_n2510, new_n2478, new_n2529);
nand_5 g00181(new_n2529, new_n2528, new_n2530);
xnor_4 g00182(new_n2529, new_n2527, new_n2531);
xnor_4 g00183(new_n2373, new_n2359, new_n2532);
not_8  g00184(new_n2532, new_n2533_1);
xnor_4 g00185(new_n2508, new_n2507, new_n2534);
nor_5  g00186(new_n2534, new_n2533_1, new_n2535_1);
not_8  g00187(new_n2535_1, new_n2536);
xnor_4 g00188(new_n2534, new_n2532, new_n2537_1);
xnor_4 g00189(new_n2505, new_n2488, new_n2538);
xnor_4 g00190(n16223, n6385, new_n2539);
xnor_4 g00191(new_n2539, new_n2371, new_n2540);
not_8  g00192(new_n2540, new_n2541);
nor_5  g00193(new_n2541, new_n2538, new_n2542);
not_8  g00194(new_n2542, new_n2543);
xnor_4 g00195(new_n2540, new_n2538, new_n2544);
xnor_4 g00196(n9251, n2387, new_n2545);
not_8  g00197(new_n2489, new_n2546);
xnor_4 g00198(new_n2546, new_n2382, new_n2547_1);
not_8  g00199(new_n2547_1, new_n2548);
nor_5  g00200(new_n2548, new_n2545, new_n2549);
xnor_4 g00201(n20138, n19494, new_n2550);
xnor_4 g00202(new_n2550, new_n2369, new_n2551);
not_8  g00203(new_n2551, new_n2552);
nor_5  g00204(new_n2552, new_n2549, new_n2553_1);
not_8  g00205(new_n2553_1, new_n2554);
xnor_4 g00206(new_n2502, new_n2498, new_n2555_1);
xnor_4 g00207(new_n2551, new_n2549, new_n2556);
nand_5 g00208(new_n2556, new_n2555_1, new_n2557);
nand_5 g00209(new_n2557, new_n2554, new_n2558);
nand_5 g00210(new_n2558, new_n2544, new_n2559);
nand_5 g00211(new_n2559, new_n2543, new_n2560_1);
nand_5 g00212(new_n2560_1, new_n2537_1, new_n2561_1);
nand_5 g00213(new_n2561_1, new_n2536, new_n2562);
nand_5 g00214(new_n2562, new_n2531, new_n2563);
nand_5 g00215(new_n2563, new_n2530, new_n2564);
nand_5 g00216(new_n2564, new_n2525, new_n2565);
nand_5 g00217(new_n2565, new_n2524, new_n2566);
xor_4  g00218(new_n2566, new_n2519, n7);
not_8  g00219(n1681, new_n2568);
xnor_4 g00220(n3618, new_n2568, new_n2569);
xnor_4 g00221(new_n2569, n4588, new_n2570_1);
xnor_4 g00222(n22843, n583, new_n2571);
xnor_4 g00223(new_n2571, n22201, new_n2572);
xnor_4 g00224(new_n2572, new_n2570_1, n50);
not_8  g00225(n21687, new_n2574);
not_8  g00226(n6773, new_n2575);
xnor_4 g00227(n19922, new_n2575, new_n2576);
xnor_4 g00228(new_n2576, new_n2574, new_n2577);
not_8  g00229(new_n2577, new_n2578_1);
not_8  g00230(n25926, new_n2579);
not_8  g00231(n14090, new_n2580);
xnor_4 g00232(n21398, new_n2580, new_n2581);
xnor_4 g00233(new_n2581, new_n2579, new_n2582_1);
xnor_4 g00234(new_n2582_1, new_n2578_1, n55);
not_8  g00235(n9396, new_n2584);
xnor_4 g00236(n20040, new_n2584, new_n2585);
not_8  g00237(new_n2585, new_n2586);
or_5   g00238(n19531, n1999, new_n2587);
not_8  g00239(n1999, new_n2588);
xnor_4 g00240(n19531, new_n2588, new_n2589);
or_5   g00241(n25168, n18345, new_n2590);
not_8  g00242(n18345, new_n2591);
xnor_4 g00243(n25168, new_n2591, new_n2592);
nor_5  g00244(n13190, n9318, new_n2593);
not_8  g00245(new_n2593, new_n2594);
not_8  g00246(n9318, new_n2595);
xnor_4 g00247(n13190, new_n2595, new_n2596);
nor_5  g00248(n19477, n3460, new_n2597);
not_8  g00249(new_n2597, new_n2598);
not_8  g00250(n3460, new_n2599);
xnor_4 g00251(n19477, new_n2599, new_n2600);
nor_5  g00252(n11223, n5226, new_n2601);
not_8  g00253(new_n2601, new_n2602_1);
not_8  g00254(n5226, new_n2603);
xnor_4 g00255(n11223, new_n2603, new_n2604);
nor_5  g00256(n17664, n5115, new_n2605);
not_8  g00257(n5115, new_n2606);
xnor_4 g00258(n17664, new_n2606, new_n2607);
not_8  g00259(new_n2607, new_n2608);
nor_5  g00260(n26572, n23369, new_n2609);
not_8  g00261(n23369, new_n2610);
xnor_4 g00262(n26572, new_n2610, new_n2611);
not_8  g00263(new_n2611, new_n2612);
nor_5  g00264(n11667, n1136, new_n2613);
nand_5 g00265(n21398, n19234, new_n2614);
not_8  g00266(new_n2614, new_n2615);
xnor_4 g00267(n11667, n1136, new_n2616);
nor_5  g00268(new_n2616, new_n2615, new_n2617);
nor_5  g00269(new_n2617, new_n2613, new_n2618);
nor_5  g00270(new_n2618, new_n2612, new_n2619_1);
nor_5  g00271(new_n2619_1, new_n2609, new_n2620);
nor_5  g00272(new_n2620, new_n2608, new_n2621);
nor_5  g00273(new_n2621, new_n2605, new_n2622);
not_8  g00274(new_n2622, new_n2623);
nand_5 g00275(new_n2623, new_n2604, new_n2624);
nand_5 g00276(new_n2624, new_n2602_1, new_n2625);
nand_5 g00277(new_n2625, new_n2600, new_n2626);
nand_5 g00278(new_n2626, new_n2598, new_n2627);
nand_5 g00279(new_n2627, new_n2596, new_n2628);
nand_5 g00280(new_n2628, new_n2594, new_n2629);
nand_5 g00281(new_n2629, new_n2592, new_n2630);
nand_5 g00282(new_n2630, new_n2590, new_n2631);
nand_5 g00283(new_n2631, new_n2589, new_n2632);
nand_5 g00284(new_n2632, new_n2587, new_n2633);
xnor_4 g00285(new_n2633, new_n2586, new_n2634);
xnor_4 g00286(new_n2634, n25365, new_n2635);
not_8  g00287(n14704, new_n2636);
not_8  g00288(new_n2589, new_n2637);
xnor_4 g00289(new_n2631, new_n2637, new_n2638);
nor_5  g00290(new_n2638, new_n2636, new_n2639);
xnor_4 g00291(new_n2638, n14704, new_n2640);
not_8  g00292(new_n2640, new_n2641);
not_8  g00293(n19270, new_n2642);
not_8  g00294(new_n2592, new_n2643);
xnor_4 g00295(new_n2629, new_n2643, new_n2644);
nor_5  g00296(new_n2644, new_n2642, new_n2645);
xnor_4 g00297(new_n2644, new_n2642, new_n2646_1);
not_8  g00298(n8687, new_n2647);
not_8  g00299(new_n2596, new_n2648);
xnor_4 g00300(new_n2627, new_n2648, new_n2649);
nor_5  g00301(new_n2649, new_n2647, new_n2650);
not_8  g00302(new_n2604, new_n2651);
nor_5  g00303(new_n2622, new_n2651, new_n2652);
nor_5  g00304(new_n2652, new_n2601, new_n2653);
xnor_4 g00305(new_n2653, new_n2600, new_n2654);
not_8  g00306(new_n2654, new_n2655);
nor_5  g00307(new_n2655, n24768, new_n2656);
not_8  g00308(new_n2656, new_n2657);
xnor_4 g00309(new_n2654, n24768, new_n2658);
xnor_4 g00310(new_n2622, new_n2604, new_n2659_1);
not_8  g00311(new_n2659_1, new_n2660);
nor_5  g00312(new_n2660, n26483, new_n2661_1);
not_8  g00313(new_n2661_1, new_n2662);
xnor_4 g00314(new_n2659_1, n26483, new_n2663);
not_8  g00315(n15979, new_n2664);
xnor_4 g00316(new_n2620, new_n2607, new_n2665);
nor_5  g00317(new_n2665, new_n2664, new_n2666);
xnor_4 g00318(new_n2665, n15979, new_n2667);
not_8  g00319(new_n2667, new_n2668);
not_8  g00320(n8638, new_n2669);
xnor_4 g00321(new_n2618, new_n2611, new_n2670);
nor_5  g00322(new_n2670, new_n2669, new_n2671);
xnor_4 g00323(new_n2616, new_n2614, new_n2672);
not_8  g00324(new_n2672, new_n2673);
nor_5  g00325(new_n2673, n16247, new_n2674);
not_8  g00326(new_n2674, new_n2675);
not_8  g00327(n23541, new_n2676);
xnor_4 g00328(n21398, n19234, new_n2677);
nor_5  g00329(new_n2677, new_n2676, new_n2678);
not_8  g00330(new_n2678, new_n2679);
xnor_4 g00331(new_n2672, n16247, new_n2680_1);
nand_5 g00332(new_n2680_1, new_n2679, new_n2681);
nand_5 g00333(new_n2681, new_n2675, new_n2682);
xnor_4 g00334(new_n2670, n8638, new_n2683);
not_8  g00335(new_n2683, new_n2684);
nor_5  g00336(new_n2684, new_n2682, new_n2685);
nor_5  g00337(new_n2685, new_n2671, new_n2686);
nor_5  g00338(new_n2686, new_n2668, new_n2687);
nor_5  g00339(new_n2687, new_n2666, new_n2688);
nand_5 g00340(new_n2688, new_n2663, new_n2689);
nand_5 g00341(new_n2689, new_n2662, new_n2690);
nand_5 g00342(new_n2690, new_n2658, new_n2691);
nand_5 g00343(new_n2691, new_n2657, new_n2692);
xnor_4 g00344(new_n2649, n8687, new_n2693_1);
not_8  g00345(new_n2693_1, new_n2694);
nor_5  g00346(new_n2694, new_n2692, new_n2695);
nor_5  g00347(new_n2695, new_n2650, new_n2696);
nor_5  g00348(new_n2696, new_n2646_1, new_n2697);
nor_5  g00349(new_n2697, new_n2645, new_n2698);
nor_5  g00350(new_n2698, new_n2641, new_n2699);
nor_5  g00351(new_n2699, new_n2639, new_n2700);
xnor_4 g00352(new_n2700, new_n2635, new_n2701);
not_8  g00353(new_n2701, new_n2702);
not_8  g00354(n25523, new_n2703_1);
not_8  g00355(n23430, new_n2704);
not_8  g00356(n16971, new_n2705);
nor_5  g00357(n18151, n11503, new_n2706_1);
nand_5 g00358(new_n2706_1, new_n2705, new_n2707);
nor_5  g00359(new_n2707, n10411, new_n2708);
nand_5 g00360(new_n2708, new_n2704, new_n2709);
nor_5  g00361(new_n2709, n5579, new_n2710);
nand_5 g00362(new_n2710, new_n2703_1, new_n2711_1);
nor_5  g00363(new_n2711_1, n8439, new_n2712);
not_8  g00364(new_n2712, new_n2713);
nor_5  g00365(new_n2713, n22793, new_n2714);
xnor_4 g00366(new_n2714, n13951, new_n2715);
not_8  g00367(new_n2715, new_n2716);
not_8  g00368(n2944, new_n2717);
xnor_4 g00369(n22270, new_n2717, new_n2718);
or_5   g00370(n8806, n767, new_n2719);
not_8  g00371(n767, new_n2720);
xnor_4 g00372(n8806, new_n2720, new_n2721);
or_5   g00373(n7330, n2479, new_n2722);
not_8  g00374(n7330, new_n2723);
xnor_4 g00375(new_n2723, n2479, new_n2724);
nor_5  g00376(n22492, n9372, new_n2725);
not_8  g00377(n22492, new_n2726);
xnor_4 g00378(new_n2726, n9372, new_n2727);
not_8  g00379(new_n2727, new_n2728);
nor_5  g00380(n12821, n6596, new_n2729);
not_8  g00381(n6596, new_n2730);
xnor_4 g00382(n12821, new_n2730, new_n2731_1);
not_8  g00383(new_n2731_1, new_n2732);
nor_5  g00384(n15289, n3468, new_n2733);
not_8  g00385(n3468, new_n2734);
xnor_4 g00386(n15289, new_n2734, new_n2735);
not_8  g00387(new_n2735, new_n2736);
nor_5  g00388(n18558, n6556, new_n2737);
not_8  g00389(n6556, new_n2738);
xnor_4 g00390(n18558, new_n2738, new_n2739);
not_8  g00391(new_n2739, new_n2740);
nor_5  g00392(n22871, n7149, new_n2741);
not_8  g00393(n7149, new_n2742);
xnor_4 g00394(n22871, new_n2742, new_n2743_1);
not_8  g00395(new_n2743_1, new_n2744);
nor_5  g00396(n14275, n14148, new_n2745);
nand_5 g00397(n25023, n1152, new_n2746);
not_8  g00398(new_n2746, new_n2747);
xnor_4 g00399(n14275, n14148, new_n2748);
nor_5  g00400(new_n2748, new_n2747, new_n2749);
nor_5  g00401(new_n2749, new_n2745, new_n2750);
nor_5  g00402(new_n2750, new_n2744, new_n2751);
nor_5  g00403(new_n2751, new_n2741, new_n2752);
nor_5  g00404(new_n2752, new_n2740, new_n2753);
nor_5  g00405(new_n2753, new_n2737, new_n2754);
nor_5  g00406(new_n2754, new_n2736, new_n2755);
nor_5  g00407(new_n2755, new_n2733, new_n2756);
nor_5  g00408(new_n2756, new_n2732, new_n2757);
nor_5  g00409(new_n2757, new_n2729, new_n2758);
nor_5  g00410(new_n2758, new_n2728, new_n2759);
nor_5  g00411(new_n2759, new_n2725, new_n2760);
not_8  g00412(new_n2760, new_n2761_1);
nand_5 g00413(new_n2761_1, new_n2724, new_n2762);
nand_5 g00414(new_n2762, new_n2722, new_n2763);
nand_5 g00415(new_n2763, new_n2721, new_n2764);
nand_5 g00416(new_n2764, new_n2719, new_n2765);
xnor_4 g00417(new_n2765, new_n2718, new_n2766);
xnor_4 g00418(new_n2766, new_n2716, new_n2767);
not_8  g00419(new_n2767, new_n2768);
xnor_4 g00420(new_n2712, n22793, new_n2769);
not_8  g00421(new_n2769, new_n2770);
xnor_4 g00422(new_n2763, new_n2721, new_n2771);
nor_5  g00423(new_n2771, new_n2770, new_n2772);
xnor_4 g00424(new_n2771, new_n2770, new_n2773);
xnor_4 g00425(new_n2711_1, n8439, new_n2774_1);
xnor_4 g00426(new_n2760, new_n2724, new_n2775);
not_8  g00427(new_n2775, new_n2776);
nand_5 g00428(new_n2776, new_n2774_1, new_n2777);
xnor_4 g00429(new_n2775, new_n2774_1, new_n2778);
xnor_4 g00430(new_n2710, new_n2703_1, new_n2779_1);
xnor_4 g00431(new_n2758, new_n2727, new_n2780);
not_8  g00432(new_n2780, new_n2781);
nand_5 g00433(new_n2781, new_n2779_1, new_n2782);
xnor_4 g00434(new_n2780, new_n2779_1, new_n2783_1);
xnor_4 g00435(new_n2709, n5579, new_n2784);
xnor_4 g00436(new_n2756, new_n2731_1, new_n2785);
not_8  g00437(new_n2785, new_n2786);
nand_5 g00438(new_n2786, new_n2784, new_n2787);
xnor_4 g00439(new_n2785, new_n2784, new_n2788);
xnor_4 g00440(new_n2708, n23430, new_n2789);
xnor_4 g00441(new_n2754, new_n2735, new_n2790);
nor_5  g00442(new_n2790, new_n2789, new_n2791);
not_8  g00443(n10411, new_n2792);
xnor_4 g00444(new_n2707, new_n2792, new_n2793);
xnor_4 g00445(new_n2752, new_n2739, new_n2794);
nor_5  g00446(new_n2794, new_n2793, new_n2795);
xnor_4 g00447(new_n2794, new_n2793, new_n2796);
xnor_4 g00448(new_n2706_1, n16971, new_n2797);
xnor_4 g00449(new_n2750, new_n2743_1, new_n2798);
nor_5  g00450(new_n2798, new_n2797, new_n2799);
xnor_4 g00451(new_n2798, new_n2797, new_n2800);
not_8  g00452(n11503, new_n2801);
xnor_4 g00453(n18151, new_n2801, new_n2802);
xnor_4 g00454(new_n2748, new_n2746, new_n2803);
nor_5  g00455(new_n2803, new_n2802, new_n2804);
not_8  g00456(n1152, new_n2805);
xnor_4 g00457(n25023, new_n2805, new_n2806);
not_8  g00458(new_n2806, new_n2807);
nor_5  g00459(new_n2807, n18151, new_n2808);
not_8  g00460(new_n2808, new_n2809_1);
xnor_4 g00461(new_n2803, new_n2802, new_n2810);
nor_5  g00462(new_n2810, new_n2809_1, new_n2811);
nor_5  g00463(new_n2811, new_n2804, new_n2812);
nor_5  g00464(new_n2812, new_n2800, new_n2813);
nor_5  g00465(new_n2813, new_n2799, new_n2814);
nor_5  g00466(new_n2814, new_n2796, new_n2815);
nor_5  g00467(new_n2815, new_n2795, new_n2816_1);
xnor_4 g00468(new_n2790, new_n2789, new_n2817);
nor_5  g00469(new_n2817, new_n2816_1, new_n2818);
nor_5  g00470(new_n2818, new_n2791, new_n2819);
not_8  g00471(new_n2819, new_n2820);
nand_5 g00472(new_n2820, new_n2788, new_n2821);
nand_5 g00473(new_n2821, new_n2787, new_n2822);
nand_5 g00474(new_n2822, new_n2783_1, new_n2823);
nand_5 g00475(new_n2823, new_n2782, new_n2824);
nand_5 g00476(new_n2824, new_n2778, new_n2825);
nand_5 g00477(new_n2825, new_n2777, new_n2826_1);
nor_5  g00478(new_n2826_1, new_n2773, new_n2827);
nor_5  g00479(new_n2827, new_n2772, new_n2828);
xnor_4 g00480(new_n2828, new_n2768, new_n2829);
xnor_4 g00481(new_n2829, new_n2702, new_n2830);
xnor_4 g00482(new_n2698, new_n2640, new_n2831);
not_8  g00483(new_n2831, new_n2832);
xnor_4 g00484(new_n2826_1, new_n2773, new_n2833);
nor_5  g00485(new_n2833, new_n2832, new_n2834);
xnor_4 g00486(new_n2833, new_n2831, new_n2835);
not_8  g00487(new_n2835, new_n2836);
xnor_4 g00488(new_n2696, new_n2646_1, new_n2837);
not_8  g00489(new_n2837, new_n2838);
xnor_4 g00490(new_n2824, new_n2778, new_n2839);
nor_5  g00491(new_n2839, new_n2838, new_n2840);
not_8  g00492(new_n2840, new_n2841);
xnor_4 g00493(new_n2839, new_n2837, new_n2842);
xnor_4 g00494(new_n2693_1, new_n2692, new_n2843);
xnor_4 g00495(new_n2822, new_n2783_1, new_n2844);
nor_5  g00496(new_n2844, new_n2843, new_n2845);
not_8  g00497(new_n2845, new_n2846);
not_8  g00498(new_n2843, new_n2847);
xnor_4 g00499(new_n2844, new_n2847, new_n2848);
not_8  g00500(new_n2658, new_n2849);
xnor_4 g00501(new_n2690, new_n2849, new_n2850);
xnor_4 g00502(new_n2819, new_n2788, new_n2851);
nor_5  g00503(new_n2851, new_n2850, new_n2852);
xnor_4 g00504(new_n2851, new_n2850, new_n2853_1);
xnor_4 g00505(new_n2688, new_n2663, new_n2854);
xnor_4 g00506(new_n2817, new_n2816_1, new_n2855);
nor_5  g00507(new_n2855, new_n2854, new_n2856);
not_8  g00508(new_n2856, new_n2857);
not_8  g00509(new_n2854, new_n2858_1);
xnor_4 g00510(new_n2855, new_n2858_1, new_n2859);
xnor_4 g00511(new_n2814, new_n2796, new_n2860_1);
xnor_4 g00512(new_n2686, new_n2667, new_n2861);
nor_5  g00513(new_n2861, new_n2860_1, new_n2862);
not_8  g00514(new_n2862, new_n2863);
not_8  g00515(new_n2861, new_n2864);
xnor_4 g00516(new_n2864, new_n2860_1, new_n2865);
xnor_4 g00517(new_n2812, new_n2800, new_n2866);
xnor_4 g00518(new_n2683, new_n2682, new_n2867);
and_5  g00519(new_n2867, new_n2866, new_n2868);
not_8  g00520(new_n2867, new_n2869);
xnor_4 g00521(new_n2869, new_n2866, new_n2870);
not_8  g00522(new_n2870, new_n2871);
xnor_4 g00523(new_n2810, new_n2808, new_n2872);
xnor_4 g00524(new_n2680_1, new_n2678, new_n2873);
nand_5 g00525(new_n2873, new_n2872, new_n2874);
xnor_4 g00526(new_n2677, n23541, new_n2875);
not_8  g00527(new_n2875, new_n2876);
xnor_4 g00528(new_n2806, n18151, new_n2877);
nor_5  g00529(new_n2877, new_n2876, new_n2878);
not_8  g00530(new_n2878, new_n2879);
not_8  g00531(new_n2873, new_n2880);
xnor_4 g00532(new_n2880, new_n2872, new_n2881);
nand_5 g00533(new_n2881, new_n2879, new_n2882);
nand_5 g00534(new_n2882, new_n2874, new_n2883);
nor_5  g00535(new_n2883, new_n2871, new_n2884);
nor_5  g00536(new_n2884, new_n2868, new_n2885);
nand_5 g00537(new_n2885, new_n2865, new_n2886_1);
nand_5 g00538(new_n2886_1, new_n2863, new_n2887_1);
nand_5 g00539(new_n2887_1, new_n2859, new_n2888);
nand_5 g00540(new_n2888, new_n2857, new_n2889);
nor_5  g00541(new_n2889, new_n2853_1, new_n2890);
nor_5  g00542(new_n2890, new_n2852, new_n2891);
nand_5 g00543(new_n2891, new_n2848, new_n2892);
nand_5 g00544(new_n2892, new_n2846, new_n2893);
nand_5 g00545(new_n2893, new_n2842, new_n2894);
nand_5 g00546(new_n2894, new_n2841, new_n2895);
nor_5  g00547(new_n2895, new_n2836, new_n2896);
nor_5  g00548(new_n2896, new_n2834, new_n2897);
xnor_4 g00549(new_n2897, new_n2830, n108);
xnor_4 g00550(n22379, n767, new_n2899);
not_8  g00551(n1662, new_n2900);
or_5   g00552(n7330, new_n2900, new_n2901);
xnor_4 g00553(n7330, n1662, new_n2902);
not_8  g00554(n12875, new_n2903);
or_5   g00555(n22492, new_n2903, new_n2904);
xnor_4 g00556(n22492, n12875, new_n2905);
not_8  g00557(n2035, new_n2906);
or_5   g00558(n12821, new_n2906, new_n2907);
xnor_4 g00559(n12821, n2035, new_n2908);
not_8  g00560(n5213, new_n2909);
nor_5  g00561(new_n2909, n3468, new_n2910);
xnor_4 g00562(n5213, n3468, new_n2911);
not_8  g00563(n4665, new_n2912);
nor_5  g00564(n18558, new_n2912, new_n2913);
not_8  g00565(new_n2913, new_n2914);
xnor_4 g00566(n18558, n4665, new_n2915);
nor_5  g00567(n19005, new_n2742, new_n2916);
not_8  g00568(n19005, new_n2917);
nor_5  g00569(new_n2917, n7149, new_n2918);
not_8  g00570(n14148, new_n2919);
nor_5  g00571(new_n2919, n4326, new_n2920);
not_8  g00572(n4326, new_n2921);
nor_5  g00573(n14148, new_n2921, new_n2922);
nor_5  g00574(n5438, new_n2805, new_n2923);
not_8  g00575(new_n2923, new_n2924);
nor_5  g00576(new_n2924, new_n2922, new_n2925);
nor_5  g00577(new_n2925, new_n2920, new_n2926);
nor_5  g00578(new_n2926, new_n2918, new_n2927);
nor_5  g00579(new_n2927, new_n2916, new_n2928);
nand_5 g00580(new_n2928, new_n2915, new_n2929_1);
nand_5 g00581(new_n2929_1, new_n2914, new_n2930);
and_5  g00582(new_n2930, new_n2911, new_n2931);
nor_5  g00583(new_n2931, new_n2910, new_n2932);
not_8  g00584(new_n2932, new_n2933);
nand_5 g00585(new_n2933, new_n2908, new_n2934);
nand_5 g00586(new_n2934, new_n2907, new_n2935);
nand_5 g00587(new_n2935, new_n2905, new_n2936);
nand_5 g00588(new_n2936, new_n2904, new_n2937);
nand_5 g00589(new_n2937, new_n2902, new_n2938);
nand_5 g00590(new_n2938, new_n2901, new_n2939);
xnor_4 g00591(new_n2939, new_n2899, new_n2940);
not_8  g00592(n6814, new_n2941);
xnor_4 g00593(n10763, new_n2941, new_n2942);
or_5   g00594(n19701, n7437, new_n2943);
not_8  g00595(n7437, new_n2944_1);
xnor_4 g00596(n19701, new_n2944_1, new_n2945);
nor_5  g00597(n23529, n20700, new_n2946);
not_8  g00598(n20700, new_n2947);
xnor_4 g00599(n23529, new_n2947, new_n2948_1);
not_8  g00600(new_n2948_1, new_n2949);
nor_5  g00601(n24620, n7099, new_n2950);
not_8  g00602(n7099, new_n2951);
xnor_4 g00603(n24620, new_n2951, new_n2952);
not_8  g00604(new_n2952, new_n2953);
nor_5  g00605(n12811, n5211, new_n2954);
not_8  g00606(n5211, new_n2955);
xnor_4 g00607(n12811, new_n2955, new_n2956);
not_8  g00608(new_n2956, new_n2957);
nor_5  g00609(n12956, n1118, new_n2958);
not_8  g00610(n1118, new_n2959);
xnor_4 g00611(n12956, new_n2959, new_n2960);
not_8  g00612(new_n2960, new_n2961_1);
nor_5  g00613(n25974, n18295, new_n2962);
not_8  g00614(n18295, new_n2963);
xnor_4 g00615(n25974, new_n2963, new_n2964);
not_8  g00616(new_n2964, new_n2965);
nor_5  g00617(n6502, n1630, new_n2966);
nand_5 g00618(n15780, n1451, new_n2967);
not_8  g00619(new_n2967, new_n2968);
xnor_4 g00620(n6502, n1630, new_n2969);
nor_5  g00621(new_n2969, new_n2968, new_n2970);
nor_5  g00622(new_n2970, new_n2966, new_n2971_1);
nor_5  g00623(new_n2971_1, new_n2965, new_n2972);
nor_5  g00624(new_n2972, new_n2962, new_n2973);
nor_5  g00625(new_n2973, new_n2961_1, new_n2974);
nor_5  g00626(new_n2974, new_n2958, new_n2975);
nor_5  g00627(new_n2975, new_n2957, new_n2976);
nor_5  g00628(new_n2976, new_n2954, new_n2977);
nor_5  g00629(new_n2977, new_n2953, new_n2978_1);
nor_5  g00630(new_n2978_1, new_n2950, new_n2979_1);
nor_5  g00631(new_n2979_1, new_n2949, new_n2980);
nor_5  g00632(new_n2980, new_n2946, new_n2981);
not_8  g00633(new_n2981, new_n2982);
nand_5 g00634(new_n2982, new_n2945, new_n2983);
nand_5 g00635(new_n2983, new_n2943, new_n2984);
xnor_4 g00636(new_n2984, new_n2942, new_n2985_1);
not_8  g00637(n12657, new_n2986);
xnor_4 g00638(n27089, new_n2986, new_n2987);
not_8  g00639(new_n2987, new_n2988);
or_5   g00640(n17077, n11841, new_n2989);
not_8  g00641(n11841, new_n2990);
xnor_4 g00642(n17077, new_n2990, new_n2991);
nor_5  g00643(n26510, n10710, new_n2992);
not_8  g00644(new_n2992, new_n2993);
not_8  g00645(n10710, new_n2994);
xnor_4 g00646(n26510, new_n2994, new_n2995);
nor_5  g00647(n23068, n20929, new_n2996);
not_8  g00648(new_n2996, new_n2997);
not_8  g00649(n20929, new_n2998);
xnor_4 g00650(n23068, new_n2998, new_n2999_1);
nor_5  g00651(n19514, n8006, new_n3000);
not_8  g00652(new_n3000, new_n3001);
not_8  g00653(n8006, new_n3002);
xnor_4 g00654(n19514, new_n3002, new_n3003);
nor_5  g00655(n25074, n10053, new_n3004);
not_8  g00656(new_n3004, new_n3005);
not_8  g00657(n10053, new_n3006);
xnor_4 g00658(n25074, new_n3006, new_n3007);
nor_5  g00659(n16396, n8399, new_n3008);
not_8  g00660(n8399, new_n3009);
xnor_4 g00661(n16396, new_n3009, new_n3010_1);
not_8  g00662(new_n3010_1, new_n3011);
nor_5  g00663(n9507, n9399, new_n3012);
nand_5 g00664(n26979, n2088, new_n3013);
not_8  g00665(new_n3013, new_n3014);
xnor_4 g00666(n9507, n9399, new_n3015);
nor_5  g00667(new_n3015, new_n3014, new_n3016);
nor_5  g00668(new_n3016, new_n3012, new_n3017_1);
nor_5  g00669(new_n3017_1, new_n3011, new_n3018_1);
nor_5  g00670(new_n3018_1, new_n3008, new_n3019);
not_8  g00671(new_n3019, new_n3020_1);
nand_5 g00672(new_n3020_1, new_n3007, new_n3021);
nand_5 g00673(new_n3021, new_n3005, new_n3022);
nand_5 g00674(new_n3022, new_n3003, new_n3023);
nand_5 g00675(new_n3023, new_n3001, new_n3024);
nand_5 g00676(new_n3024, new_n2999_1, new_n3025);
nand_5 g00677(new_n3025, new_n2997, new_n3026);
nand_5 g00678(new_n3026, new_n2995, new_n3027);
nand_5 g00679(new_n3027, new_n2993, new_n3028);
nand_5 g00680(new_n3028, new_n2991, new_n3029);
nand_5 g00681(new_n3029, new_n2989, new_n3030_1);
xnor_4 g00682(new_n3030_1, new_n2988, new_n3031);
not_8  g00683(new_n3031, new_n3032);
xnor_4 g00684(new_n3032, new_n2985_1, new_n3033);
xnor_4 g00685(new_n2981, new_n2945, new_n3034);
xnor_4 g00686(new_n3028, new_n2991, new_n3035);
nor_5  g00687(new_n3035, new_n3034, new_n3036);
not_8  g00688(new_n3035, new_n3037);
xnor_4 g00689(new_n3037, new_n3034, new_n3038);
not_8  g00690(new_n3038, new_n3039);
xnor_4 g00691(new_n2979_1, new_n2948_1, new_n3040);
not_8  g00692(new_n3040, new_n3041);
xnor_4 g00693(new_n3026, new_n2995, new_n3042);
not_8  g00694(new_n3042, new_n3043);
nor_5  g00695(new_n3043, new_n3041, new_n3044);
not_8  g00696(new_n3044, new_n3045);
xnor_4 g00697(new_n3043, new_n3040, new_n3046);
xnor_4 g00698(new_n2977, new_n2952, new_n3047);
not_8  g00699(new_n3047, new_n3048);
xnor_4 g00700(new_n3024, new_n2999_1, new_n3049);
not_8  g00701(new_n3049, new_n3050);
nor_5  g00702(new_n3050, new_n3048, new_n3051);
not_8  g00703(new_n3051, new_n3052);
xnor_4 g00704(new_n3049, new_n3048, new_n3053);
xnor_4 g00705(new_n2975, new_n2956, new_n3054);
not_8  g00706(new_n3054, new_n3055);
xnor_4 g00707(new_n3022, new_n3003, new_n3056);
not_8  g00708(new_n3056, new_n3057);
nor_5  g00709(new_n3057, new_n3055, new_n3058);
xnor_4 g00710(new_n3056, new_n3055, new_n3059);
not_8  g00711(new_n3059, new_n3060);
xnor_4 g00712(new_n2973, new_n2960, new_n3061);
not_8  g00713(new_n3061, new_n3062);
xnor_4 g00714(new_n3019, new_n3007, new_n3063);
nor_5  g00715(new_n3063, new_n3062, new_n3064);
xnor_4 g00716(new_n3063, new_n3061, new_n3065);
not_8  g00717(new_n3065, new_n3066);
xnor_4 g00718(new_n2971_1, new_n2964, new_n3067_1);
xnor_4 g00719(new_n3017_1, new_n3010_1, new_n3068);
not_8  g00720(new_n3068, new_n3069);
nor_5  g00721(new_n3069, new_n3067_1, new_n3070);
not_8  g00722(new_n3070, new_n3071);
xnor_4 g00723(new_n3068, new_n3067_1, new_n3072);
xnor_4 g00724(new_n2969, new_n2968, new_n3073);
xnor_4 g00725(new_n3015, new_n3013, new_n3074);
nor_5  g00726(new_n3074, new_n3073, new_n3075);
xnor_4 g00727(n15780, n1451, new_n3076_1);
not_8  g00728(new_n3076_1, new_n3077);
not_8  g00729(n2088, new_n3078);
xnor_4 g00730(n26979, new_n3078, new_n3079);
not_8  g00731(new_n3079, new_n3080);
nor_5  g00732(new_n3080, new_n3077, new_n3081);
not_8  g00733(new_n3073, new_n3082);
xnor_4 g00734(new_n3074, new_n3082, new_n3083);
nand_5 g00735(new_n3083, new_n3081, new_n3084);
not_8  g00736(new_n3084, new_n3085);
nor_5  g00737(new_n3085, new_n3075, new_n3086);
nand_5 g00738(new_n3086, new_n3072, new_n3087);
nand_5 g00739(new_n3087, new_n3071, new_n3088);
nor_5  g00740(new_n3088, new_n3066, new_n3089_1);
nor_5  g00741(new_n3089_1, new_n3064, new_n3090);
nor_5  g00742(new_n3090, new_n3060, new_n3091);
nor_5  g00743(new_n3091, new_n3058, new_n3092);
not_8  g00744(new_n3092, new_n3093);
nand_5 g00745(new_n3093, new_n3053, new_n3094);
nand_5 g00746(new_n3094, new_n3052, new_n3095);
nand_5 g00747(new_n3095, new_n3046, new_n3096);
nand_5 g00748(new_n3096, new_n3045, new_n3097);
nor_5  g00749(new_n3097, new_n3039, new_n3098);
nor_5  g00750(new_n3098, new_n3036, new_n3099);
xnor_4 g00751(new_n3099, new_n3033, new_n3100);
xnor_4 g00752(new_n3100, new_n2940, new_n3101);
xnor_4 g00753(new_n2937, new_n2902, new_n3102);
xnor_4 g00754(new_n3097, new_n3038, new_n3103);
not_8  g00755(new_n3103, new_n3104);
nand_5 g00756(new_n3104, new_n3102, new_n3105);
xnor_4 g00757(new_n3103, new_n3102, new_n3106);
xnor_4 g00758(new_n2935, new_n2905, new_n3107);
xnor_4 g00759(new_n3095, new_n3046, new_n3108);
not_8  g00760(new_n3108, new_n3109);
nand_5 g00761(new_n3109, new_n3107, new_n3110);
xnor_4 g00762(new_n3108, new_n3107, new_n3111);
xnor_4 g00763(new_n2932, new_n2908, new_n3112);
not_8  g00764(new_n3112, new_n3113);
xnor_4 g00765(new_n3092, new_n3053, new_n3114);
nand_5 g00766(new_n3114, new_n3113, new_n3115);
xnor_4 g00767(new_n3114, new_n3112, new_n3116);
xnor_4 g00768(new_n2930, new_n2911, new_n3117);
xnor_4 g00769(new_n3090, new_n3059, new_n3118);
nand_5 g00770(new_n3118, new_n3117, new_n3119);
not_8  g00771(new_n3118, new_n3120);
xnor_4 g00772(new_n3120, new_n3117, new_n3121);
xnor_4 g00773(new_n3088, new_n3065, new_n3122);
not_8  g00774(new_n3122, new_n3123);
xnor_4 g00775(new_n2928, new_n2915, new_n3124);
not_8  g00776(new_n3124, new_n3125_1);
nor_5  g00777(new_n3125_1, new_n3123, new_n3126_1);
xnor_4 g00778(new_n3125_1, new_n3122, new_n3127);
not_8  g00779(new_n3127, new_n3128);
xnor_4 g00780(new_n3086, new_n3072, new_n3129);
not_8  g00781(new_n3129, new_n3130);
xnor_4 g00782(n19005, n7149, new_n3131);
xnor_4 g00783(new_n3131, new_n2926, new_n3132);
not_8  g00784(new_n3132, new_n3133);
nor_5  g00785(new_n3133, new_n3130, new_n3134);
xnor_4 g00786(new_n3133, new_n3129, new_n3135);
not_8  g00787(new_n3135, new_n3136_1);
xnor_4 g00788(n5438, n1152, new_n3137);
xnor_4 g00789(new_n3079, new_n3077, new_n3138);
nor_5  g00790(new_n3138, new_n3137, new_n3139);
xnor_4 g00791(n14148, n4326, new_n3140);
xnor_4 g00792(new_n3140, new_n2924, new_n3141);
not_8  g00793(new_n3141, new_n3142);
nor_5  g00794(new_n3142, new_n3139, new_n3143);
xnor_4 g00795(new_n3083, new_n3081, new_n3144);
xnor_4 g00796(new_n3141, new_n3139, new_n3145);
not_8  g00797(new_n3145, new_n3146);
nor_5  g00798(new_n3146, new_n3144, new_n3147);
nor_5  g00799(new_n3147, new_n3143, new_n3148);
nor_5  g00800(new_n3148, new_n3136_1, new_n3149);
nor_5  g00801(new_n3149, new_n3134, new_n3150);
nor_5  g00802(new_n3150, new_n3128, new_n3151);
nor_5  g00803(new_n3151, new_n3126_1, new_n3152);
not_8  g00804(new_n3152, new_n3153);
nand_5 g00805(new_n3153, new_n3121, new_n3154);
nand_5 g00806(new_n3154, new_n3119, new_n3155);
nand_5 g00807(new_n3155, new_n3116, new_n3156);
nand_5 g00808(new_n3156, new_n3115, new_n3157);
nand_5 g00809(new_n3157, new_n3111, new_n3158);
nand_5 g00810(new_n3158, new_n3110, new_n3159);
nand_5 g00811(new_n3159, new_n3106, new_n3160);
nand_5 g00812(new_n3160, new_n3105, new_n3161_1);
xnor_4 g00813(new_n3161_1, new_n3101, n142);
not_8  g00814(n5025, new_n3163);
not_8  g00815(n4319, new_n3164_1);
xnor_4 g00816(n7335, new_n3164_1, new_n3165);
not_8  g00817(new_n3165, new_n3166);
or_5   g00818(n23463, n5696, new_n3167);
not_8  g00819(n5696, new_n3168);
xnor_4 g00820(n23463, new_n3168, new_n3169);
or_5   g00821(n13367, n13074, new_n3170);
not_8  g00822(n13074, new_n3171);
xnor_4 g00823(n13367, new_n3171, new_n3172);
nor_5  g00824(n10739, n932, new_n3173);
not_8  g00825(new_n3173, new_n3174);
not_8  g00826(n932, new_n3175);
xnor_4 g00827(n10739, new_n3175, new_n3176);
nor_5  g00828(n21753, n6691, new_n3177);
not_8  g00829(new_n3177, new_n3178);
not_8  g00830(n6691, new_n3179);
xnor_4 g00831(n21753, new_n3179, new_n3180);
nor_5  g00832(n21832, n3260, new_n3181);
not_8  g00833(new_n3181, new_n3182);
not_8  g00834(n3260, new_n3183);
xnor_4 g00835(n21832, new_n3183, new_n3184);
nor_5  g00836(n26913, n20489, new_n3185);
not_8  g00837(new_n3185, new_n3186);
not_8  g00838(n20489, new_n3187);
xnor_4 g00839(n26913, new_n3187, new_n3188);
nor_5  g00840(n16223, n2355, new_n3189);
not_8  g00841(new_n3189, new_n3190);
not_8  g00842(n2355, new_n3191);
xnor_4 g00843(n16223, new_n3191, new_n3192);
nor_5  g00844(n19494, n11121, new_n3193);
not_8  g00845(new_n3193, new_n3194);
nand_5 g00846(n16217, n2387, new_n3195);
not_8  g00847(new_n3195, new_n3196);
xnor_4 g00848(n19494, n11121, new_n3197);
nor_5  g00849(new_n3197, new_n3196, new_n3198);
not_8  g00850(new_n3198, new_n3199);
nand_5 g00851(new_n3199, new_n3194, new_n3200);
nand_5 g00852(new_n3200, new_n3192, new_n3201);
nand_5 g00853(new_n3201, new_n3190, new_n3202);
nand_5 g00854(new_n3202, new_n3188, new_n3203);
nand_5 g00855(new_n3203, new_n3186, new_n3204);
nand_5 g00856(new_n3204, new_n3184, new_n3205);
nand_5 g00857(new_n3205, new_n3182, new_n3206);
nand_5 g00858(new_n3206, new_n3180, new_n3207);
nand_5 g00859(new_n3207, new_n3178, new_n3208_1);
nand_5 g00860(new_n3208_1, new_n3176, new_n3209);
nand_5 g00861(new_n3209, new_n3174, new_n3210);
nand_5 g00862(new_n3210, new_n3172, new_n3211);
nand_5 g00863(new_n3211, new_n3170, new_n3212);
nand_5 g00864(new_n3212, new_n3169, new_n3213);
nand_5 g00865(new_n3213, new_n3167, new_n3214);
xnor_4 g00866(new_n3214, new_n3166, new_n3215);
not_8  g00867(new_n3215, new_n3216);
nand_5 g00868(new_n3216, new_n3163, new_n3217);
xnor_4 g00869(new_n3215, new_n3163, new_n3218);
not_8  g00870(n6485, new_n3219_1);
not_8  g00871(new_n3169, new_n3220);
xnor_4 g00872(new_n3212, new_n3220, new_n3221);
not_8  g00873(new_n3221, new_n3222);
nand_5 g00874(new_n3222, new_n3219_1, new_n3223);
xnor_4 g00875(new_n3221, new_n3219_1, new_n3224);
not_8  g00876(n26036, new_n3225);
not_8  g00877(new_n3172, new_n3226);
xnor_4 g00878(new_n3210, new_n3226, new_n3227);
not_8  g00879(new_n3227, new_n3228_1);
nand_5 g00880(new_n3228_1, new_n3225, new_n3229);
xnor_4 g00881(new_n3227, new_n3225, new_n3230);
not_8  g00882(n19770, new_n3231);
not_8  g00883(new_n3176, new_n3232);
xnor_4 g00884(new_n3208_1, new_n3232, new_n3233);
not_8  g00885(new_n3233, new_n3234);
nand_5 g00886(new_n3234, new_n3231, new_n3235_1);
xnor_4 g00887(new_n3233, new_n3231, new_n3236);
not_8  g00888(n8782, new_n3237);
xnor_4 g00889(new_n3206, new_n3180, new_n3238);
nand_5 g00890(new_n3238, new_n3237, new_n3239);
xnor_4 g00891(new_n3238, n8782, new_n3240);
not_8  g00892(n8678, new_n3241);
not_8  g00893(new_n3184, new_n3242);
not_8  g00894(new_n3188, new_n3243);
not_8  g00895(new_n3192, new_n3244_1);
nor_5  g00896(new_n3198, new_n3193, new_n3245);
nor_5  g00897(new_n3245, new_n3244_1, new_n3246);
nor_5  g00898(new_n3246, new_n3189, new_n3247);
nor_5  g00899(new_n3247, new_n3243, new_n3248);
nor_5  g00900(new_n3248, new_n3185, new_n3249);
xnor_4 g00901(new_n3249, new_n3242, new_n3250);
nand_5 g00902(new_n3250, new_n3241, new_n3251);
xnor_4 g00903(new_n3250, n8678, new_n3252);
not_8  g00904(n1432, new_n3253_1);
xnor_4 g00905(new_n3247, new_n3188, new_n3254);
not_8  g00906(new_n3254, new_n3255);
nand_5 g00907(new_n3255, new_n3253_1, new_n3256);
xnor_4 g00908(new_n3254, new_n3253_1, new_n3257);
not_8  g00909(n21599, new_n3258);
xnor_4 g00910(new_n3245, new_n3192, new_n3259);
not_8  g00911(new_n3259, new_n3260_1);
nand_5 g00912(new_n3260_1, new_n3258, new_n3261);
xnor_4 g00913(new_n3259, new_n3258, new_n3262);
not_8  g00914(n25336, new_n3263_1);
xnor_4 g00915(n16217, n2387, new_n3264);
nor_5  g00916(new_n3264, n11424, new_n3265);
nand_5 g00917(new_n3265, new_n3263_1, new_n3266);
xnor_4 g00918(new_n3265, n25336, new_n3267);
xnor_4 g00919(new_n3197, new_n3195, new_n3268);
not_8  g00920(new_n3268, new_n3269);
nand_5 g00921(new_n3269, new_n3267, new_n3270);
nand_5 g00922(new_n3270, new_n3266, new_n3271);
nand_5 g00923(new_n3271, new_n3262, new_n3272);
nand_5 g00924(new_n3272, new_n3261, new_n3273);
nand_5 g00925(new_n3273, new_n3257, new_n3274);
nand_5 g00926(new_n3274, new_n3256, new_n3275);
nand_5 g00927(new_n3275, new_n3252, new_n3276);
nand_5 g00928(new_n3276, new_n3251, new_n3277);
nand_5 g00929(new_n3277, new_n3240, new_n3278);
nand_5 g00930(new_n3278, new_n3239, new_n3279_1);
nand_5 g00931(new_n3279_1, new_n3236, new_n3280);
nand_5 g00932(new_n3280, new_n3235_1, new_n3281);
nand_5 g00933(new_n3281, new_n3230, new_n3282);
nand_5 g00934(new_n3282, new_n3229, new_n3283);
nand_5 g00935(new_n3283, new_n3224, new_n3284);
nand_5 g00936(new_n3284, new_n3223, new_n3285);
nand_5 g00937(new_n3285, new_n3218, new_n3286);
nand_5 g00938(new_n3286, new_n3217, new_n3287);
or_5   g00939(n7335, n4319, new_n3288);
nand_5 g00940(new_n3214, new_n3165, new_n3289_1);
nand_5 g00941(new_n3289_1, new_n3288, new_n3290);
not_8  g00942(new_n3290, new_n3291);
nor_5  g00943(new_n3291, new_n3287, new_n3292);
not_8  g00944(new_n3292, new_n3293);
not_8  g00945(n3425, new_n3294);
not_8  g00946(n9967, new_n3295);
nor_5  g00947(n12315, n3952, new_n3296);
nand_5 g00948(new_n3296, new_n2446, new_n3297);
nor_5  g00949(new_n3297, n24278, new_n3298);
nand_5 g00950(new_n3298, new_n2438, new_n3299);
nor_5  g00951(new_n3299, n26823, new_n3300);
nand_5 g00952(new_n3300, new_n2430, new_n3301_1);
nor_5  g00953(new_n3301_1, n20946, new_n3302);
nand_5 g00954(new_n3302, new_n3295, new_n3303);
xnor_4 g00955(new_n3303, new_n3294, new_n3304);
not_8  g00956(new_n3304, new_n3305);
xnor_4 g00957(new_n3285, new_n3218, new_n3306_1);
not_8  g00958(new_n3306_1, new_n3307);
nor_5  g00959(new_n3307, new_n3305, new_n3308);
nor_5  g00960(new_n3303, n3425, new_n3309);
not_8  g00961(new_n3309, new_n3310);
xnor_4 g00962(new_n3306_1, new_n3305, new_n3311);
xnor_4 g00963(new_n3302, n9967, new_n3312);
xnor_4 g00964(new_n3283, new_n3224, new_n3313);
nand_5 g00965(new_n3313, new_n3312, new_n3314);
not_8  g00966(new_n3312, new_n3315);
xnor_4 g00967(new_n3313, new_n3315, new_n3316_1);
not_8  g00968(n20946, new_n3317);
xnor_4 g00969(new_n3301_1, new_n3317, new_n3318);
xnor_4 g00970(new_n3281, new_n3230, new_n3319);
nand_5 g00971(new_n3319, new_n3318, new_n3320_1);
not_8  g00972(new_n3318, new_n3321);
xnor_4 g00973(new_n3319, new_n3321, new_n3322);
xnor_4 g00974(new_n3300, n7751, new_n3323);
xnor_4 g00975(new_n3279_1, new_n3236, new_n3324_1);
nand_5 g00976(new_n3324_1, new_n3323, new_n3325);
not_8  g00977(new_n3323, new_n3326);
xnor_4 g00978(new_n3324_1, new_n3326, new_n3327);
xnor_4 g00979(new_n3299, new_n2434, new_n3328);
xnor_4 g00980(new_n3277, new_n3240, new_n3329);
nand_5 g00981(new_n3329, new_n3328, new_n3330);
not_8  g00982(new_n3328, new_n3331);
xnor_4 g00983(new_n3329, new_n3331, new_n3332_1);
xnor_4 g00984(new_n3298, n4812, new_n3333);
xnor_4 g00985(new_n3275, new_n3252, new_n3334);
nand_5 g00986(new_n3334, new_n3333, new_n3335);
not_8  g00987(new_n3333, new_n3336);
xnor_4 g00988(new_n3334, new_n3336, new_n3337);
xnor_4 g00989(new_n3297, new_n2442, new_n3338);
xnor_4 g00990(new_n3273, new_n3257, new_n3339);
nand_5 g00991(new_n3339, new_n3338, new_n3340_1);
not_8  g00992(new_n3338, new_n3341);
xnor_4 g00993(new_n3339, new_n3341, new_n3342);
xnor_4 g00994(new_n3296, n24618, new_n3343_1);
xnor_4 g00995(new_n3271, new_n3262, new_n3344);
nand_5 g00996(new_n3344, new_n3343_1, new_n3345);
not_8  g00997(new_n3343_1, new_n3346);
xnor_4 g00998(new_n3344, new_n3346, new_n3347);
not_8  g00999(n3952, new_n3348);
not_8  g01000(n12315, new_n3349_1);
not_8  g01001(n11424, new_n3350);
xnor_4 g01002(new_n3264, new_n3350, new_n3351);
nor_5  g01003(new_n3351, new_n3349_1, new_n3352);
nand_5 g01004(new_n3352, new_n3348, new_n3353);
not_8  g01005(new_n3353, new_n3354);
xnor_4 g01006(new_n3268, new_n3267, new_n3355);
xnor_4 g01007(n12315, new_n3348, new_n3356);
nor_5  g01008(new_n3356, new_n3352, new_n3357);
not_8  g01009(new_n3357, new_n3358);
nand_5 g01010(new_n3358, new_n3353, new_n3359);
nor_5  g01011(new_n3359, new_n3355, new_n3360);
nor_5  g01012(new_n3360, new_n3354, new_n3361);
not_8  g01013(new_n3361, new_n3362);
nand_5 g01014(new_n3362, new_n3347, new_n3363);
nand_5 g01015(new_n3363, new_n3345, new_n3364);
nand_5 g01016(new_n3364, new_n3342, new_n3365);
nand_5 g01017(new_n3365, new_n3340_1, new_n3366_1);
nand_5 g01018(new_n3366_1, new_n3337, new_n3367);
nand_5 g01019(new_n3367, new_n3335, new_n3368);
nand_5 g01020(new_n3368, new_n3332_1, new_n3369);
nand_5 g01021(new_n3369, new_n3330, new_n3370);
nand_5 g01022(new_n3370, new_n3327, new_n3371);
nand_5 g01023(new_n3371, new_n3325, new_n3372);
nand_5 g01024(new_n3372, new_n3322, new_n3373);
nand_5 g01025(new_n3373, new_n3320_1, new_n3374);
nand_5 g01026(new_n3374, new_n3316_1, new_n3375);
nand_5 g01027(new_n3375, new_n3314, new_n3376);
nand_5 g01028(new_n3376, new_n3311, new_n3377);
nand_5 g01029(new_n3377, new_n3310, new_n3378);
nor_5  g01030(new_n3378, new_n3308, new_n3379);
not_8  g01031(new_n3379, new_n3380);
nor_5  g01032(new_n3380, new_n3293, new_n3381);
not_8  g01033(new_n3381, new_n3382);
or_5   g01034(n7593, n5101, new_n3383);
not_8  g01035(n5101, new_n3384);
xnor_4 g01036(n7593, new_n3384, new_n3385);
or_5   g01037(n16507, n337, new_n3386);
not_8  g01038(n337, new_n3387);
xnor_4 g01039(n16507, new_n3387, new_n3388);
or_5   g01040(n22470, n3228, new_n3389);
not_8  g01041(n3228, new_n3390_1);
xnor_4 g01042(n22470, new_n3390_1, new_n3391);
nor_5  g01043(n19116, n5302, new_n3392);
not_8  g01044(n5302, new_n3393);
xnor_4 g01045(n19116, new_n3393, new_n3394);
not_8  g01046(new_n3394, new_n3395);
nor_5  g01047(n25738, n6861, new_n3396);
not_8  g01048(n6861, new_n3397);
xnor_4 g01049(n25738, new_n3397, new_n3398);
not_8  g01050(new_n3398, new_n3399);
nor_5  g01051(n21471, n19357, new_n3400);
not_8  g01052(n19357, new_n3401);
xnor_4 g01053(n21471, new_n3401, new_n3402);
not_8  g01054(new_n3402, new_n3403);
nor_5  g01055(n18737, n2328, new_n3404);
not_8  g01056(n2328, new_n3405);
xnor_4 g01057(n18737, new_n3405, new_n3406);
not_8  g01058(new_n3406, new_n3407);
nor_5  g01059(n15053, n14603, new_n3408);
not_8  g01060(n14603, new_n3409);
xnor_4 g01061(n15053, new_n3409, new_n3410);
not_8  g01062(new_n3410, new_n3411);
nor_5  g01063(n25471, n20794, new_n3412);
nand_5 g01064(n23333, n16502, new_n3413);
not_8  g01065(new_n3413, new_n3414);
not_8  g01066(n20794, new_n3415);
xnor_4 g01067(n25471, new_n3415, new_n3416);
not_8  g01068(new_n3416, new_n3417);
nor_5  g01069(new_n3417, new_n3414, new_n3418);
nor_5  g01070(new_n3418, new_n3412, new_n3419);
nor_5  g01071(new_n3419, new_n3411, new_n3420);
nor_5  g01072(new_n3420, new_n3408, new_n3421);
nor_5  g01073(new_n3421, new_n3407, new_n3422);
nor_5  g01074(new_n3422, new_n3404, new_n3423);
nor_5  g01075(new_n3423, new_n3403, new_n3424);
nor_5  g01076(new_n3424, new_n3400, new_n3425_1);
nor_5  g01077(new_n3425_1, new_n3399, new_n3426_1);
nor_5  g01078(new_n3426_1, new_n3396, new_n3427);
nor_5  g01079(new_n3427, new_n3395, new_n3428);
nor_5  g01080(new_n3428, new_n3392, new_n3429);
not_8  g01081(new_n3429, new_n3430);
nand_5 g01082(new_n3430, new_n3391, new_n3431);
nand_5 g01083(new_n3431, new_n3389, new_n3432);
nand_5 g01084(new_n3432, new_n3388, new_n3433);
nand_5 g01085(new_n3433, new_n3386, new_n3434);
nand_5 g01086(new_n3434, new_n3385, new_n3435);
nand_5 g01087(new_n3435, new_n3383, new_n3436);
xnor_4 g01088(new_n3290, new_n3287, new_n3437);
not_8  g01089(new_n3437, new_n3438);
xnor_4 g01090(new_n3438, new_n3379, new_n3439);
not_8  g01091(new_n3439, new_n3440);
nor_5  g01092(new_n3440, new_n3436, new_n3441);
not_8  g01093(new_n3436, new_n3442);
nor_5  g01094(new_n3439, new_n3442, new_n3443);
xnor_4 g01095(new_n3376, new_n3311, new_n3444);
xnor_4 g01096(new_n3434, new_n3385, new_n3445);
not_8  g01097(new_n3445, new_n3446);
nand_5 g01098(new_n3446, new_n3444, new_n3447);
xnor_4 g01099(new_n3445, new_n3444, new_n3448);
xnor_4 g01100(new_n3374, new_n3316_1, new_n3449);
xnor_4 g01101(new_n3432, new_n3388, new_n3450);
not_8  g01102(new_n3450, new_n3451_1);
nand_5 g01103(new_n3451_1, new_n3449, new_n3452);
xnor_4 g01104(new_n3450, new_n3449, new_n3453);
xnor_4 g01105(new_n3372, new_n3322, new_n3454);
xnor_4 g01106(new_n3429, new_n3391, new_n3455);
nand_5 g01107(new_n3455, new_n3454, new_n3456);
not_8  g01108(new_n3455, new_n3457);
xnor_4 g01109(new_n3457, new_n3454, new_n3458);
xnor_4 g01110(new_n3370, new_n3327, new_n3459_1);
xnor_4 g01111(new_n3427, new_n3394, new_n3460_1);
nand_5 g01112(new_n3460_1, new_n3459_1, new_n3461);
not_8  g01113(new_n3460_1, new_n3462);
xnor_4 g01114(new_n3462, new_n3459_1, new_n3463);
xnor_4 g01115(new_n3329, new_n3328, new_n3464);
xnor_4 g01116(new_n3368, new_n3464, new_n3465);
not_8  g01117(new_n3465, new_n3466);
xnor_4 g01118(new_n3425_1, new_n3398, new_n3467);
nand_5 g01119(new_n3467, new_n3466, new_n3468_1);
xnor_4 g01120(new_n3467, new_n3465, new_n3469);
xnor_4 g01121(new_n3366_1, new_n3337, new_n3470);
xnor_4 g01122(new_n3423, new_n3402, new_n3471);
nand_5 g01123(new_n3471, new_n3470, new_n3472);
not_8  g01124(new_n3471, new_n3473);
xnor_4 g01125(new_n3473, new_n3470, new_n3474);
xnor_4 g01126(new_n3339, new_n3338, new_n3475);
xnor_4 g01127(new_n3364, new_n3475, new_n3476);
not_8  g01128(new_n3476, new_n3477);
xnor_4 g01129(new_n3421, new_n3406, new_n3478);
nand_5 g01130(new_n3478, new_n3477, new_n3479);
xnor_4 g01131(new_n3478, new_n3476, new_n3480_1);
xnor_4 g01132(new_n3362, new_n3347, new_n3481);
xnor_4 g01133(new_n3419, new_n3410, new_n3482);
nand_5 g01134(new_n3482, new_n3481, new_n3483);
not_8  g01135(new_n3482, new_n3484);
xnor_4 g01136(new_n3484, new_n3481, new_n3485);
not_8  g01137(n16502, new_n3486);
xnor_4 g01138(n23333, new_n3486, new_n3487);
not_8  g01139(new_n3487, new_n3488);
xnor_4 g01140(new_n3351, n12315, new_n3489);
not_8  g01141(new_n3489, new_n3490);
nor_5  g01142(new_n3490, new_n3488, new_n3491);
xnor_4 g01143(new_n3416, new_n3414, new_n3492);
not_8  g01144(new_n3492, new_n3493);
nor_5  g01145(new_n3493, new_n3491, new_n3494);
not_8  g01146(new_n3355, new_n3495);
xnor_4 g01147(new_n3359, new_n3495, new_n3496);
not_8  g01148(new_n3491, new_n3497);
nor_5  g01149(new_n3497, new_n3417, new_n3498);
nor_5  g01150(new_n3498, new_n3494, new_n3499);
not_8  g01151(new_n3499, new_n3500);
nor_5  g01152(new_n3500, new_n3496, new_n3501);
nor_5  g01153(new_n3501, new_n3494, new_n3502_1);
not_8  g01154(new_n3502_1, new_n3503);
nand_5 g01155(new_n3503, new_n3485, new_n3504);
nand_5 g01156(new_n3504, new_n3483, new_n3505);
nand_5 g01157(new_n3505, new_n3480_1, new_n3506_1);
nand_5 g01158(new_n3506_1, new_n3479, new_n3507);
nand_5 g01159(new_n3507, new_n3474, new_n3508);
nand_5 g01160(new_n3508, new_n3472, new_n3509);
nand_5 g01161(new_n3509, new_n3469, new_n3510);
nand_5 g01162(new_n3510, new_n3468_1, new_n3511);
nand_5 g01163(new_n3511, new_n3463, new_n3512);
nand_5 g01164(new_n3512, new_n3461, new_n3513);
nand_5 g01165(new_n3513, new_n3458, new_n3514);
nand_5 g01166(new_n3514, new_n3456, new_n3515);
nand_5 g01167(new_n3515, new_n3453, new_n3516_1);
nand_5 g01168(new_n3516_1, new_n3452, new_n3517);
nand_5 g01169(new_n3517, new_n3448, new_n3518);
nand_5 g01170(new_n3518, new_n3447, new_n3519);
nor_5  g01171(new_n3519, new_n3443, new_n3520);
nor_5  g01172(new_n3520, new_n3441, new_n3521);
nor_5  g01173(new_n3521, new_n3382, new_n3522);
nor_5  g01174(new_n3379, new_n3293, new_n3523);
not_8  g01175(new_n3523, new_n3524);
nand_5 g01176(new_n3291, new_n3287, new_n3525);
not_8  g01177(new_n3525, new_n3526);
nand_5 g01178(new_n3526, new_n3379, new_n3527);
nand_5 g01179(new_n3527, new_n3524, new_n3528_1);
nor_5  g01180(new_n3528_1, new_n3521, new_n3529);
nor_5  g01181(new_n3529, new_n3381, new_n3530);
nor_5  g01182(new_n3530, new_n3522, n175);
not_8  g01183(n26180, new_n3532);
not_8  g01184(n8856, new_n3533);
not_8  g01185(n14130, new_n3534);
not_8  g01186(n9942, new_n3535);
not_8  g01187(n9557, new_n3536);
nor_5  g01188(n20138, n9251, new_n3537);
nand_5 g01189(new_n3537, new_n2360, new_n3538);
nor_5  g01190(new_n3538, n3136, new_n3539);
nand_5 g01191(new_n3539, new_n3536, new_n3540);
nor_5  g01192(new_n3540, n25643, new_n3541_1);
nand_5 g01193(new_n3541_1, new_n3535, new_n3542);
nor_5  g01194(new_n3542, n16482, new_n3543);
nand_5 g01195(new_n3543, new_n3534, new_n3544);
xnor_4 g01196(new_n3544, new_n3533, new_n3545);
xnor_4 g01197(new_n3545, n25494, new_n3546);
not_8  g01198(new_n3546, new_n3547);
not_8  g01199(n10117, new_n3548);
xnor_4 g01200(new_n3543, n14130, new_n3549);
not_8  g01201(new_n3549, new_n3550);
nand_5 g01202(new_n3550, new_n3548, new_n3551);
xnor_4 g01203(new_n3549, new_n3548, new_n3552);
not_8  g01204(n13460, new_n3553);
not_8  g01205(n16482, new_n3554);
xnor_4 g01206(new_n3542, new_n3554, new_n3555_1);
not_8  g01207(new_n3555_1, new_n3556);
nand_5 g01208(new_n3556, new_n3553, new_n3557);
xnor_4 g01209(new_n3555_1, new_n3553, new_n3558);
not_8  g01210(n6104, new_n3559);
xnor_4 g01211(new_n3541_1, n9942, new_n3560);
not_8  g01212(new_n3560, new_n3561_1);
nand_5 g01213(new_n3561_1, new_n3559, new_n3562);
xnor_4 g01214(new_n3560, new_n3559, new_n3563_1);
not_8  g01215(n4119, new_n3564);
not_8  g01216(n25643, new_n3565);
xnor_4 g01217(new_n3540, new_n3565, new_n3566);
not_8  g01218(new_n3566, new_n3567);
nand_5 g01219(new_n3567, new_n3564, new_n3568);
xnor_4 g01220(new_n3566, new_n3564, new_n3569);
not_8  g01221(n14510, new_n3570_1);
xnor_4 g01222(new_n3539, n9557, new_n3571);
not_8  g01223(new_n3571, new_n3572);
nand_5 g01224(new_n3572, new_n3570_1, new_n3573);
xnor_4 g01225(new_n3571, new_n3570_1, new_n3574);
not_8  g01226(n13263, new_n3575);
not_8  g01227(n3136, new_n3576);
xnor_4 g01228(new_n3538, new_n3576, new_n3577);
not_8  g01229(new_n3577, new_n3578);
nand_5 g01230(new_n3578, new_n3575, new_n3579);
not_8  g01231(n20455, new_n3580);
xnor_4 g01232(new_n3537, n6385, new_n3581);
not_8  g01233(new_n3581, new_n3582_1);
nand_5 g01234(new_n3582_1, new_n3580, new_n3583);
xnor_4 g01235(new_n3581, new_n3580, new_n3584);
not_8  g01236(n1639, new_n3585);
xnor_4 g01237(n20138, n9251, new_n3586);
nand_5 g01238(new_n3586, new_n3585, new_n3587);
nand_5 g01239(n16968, n9251, new_n3588);
xnor_4 g01240(new_n3586, n1639, new_n3589);
nand_5 g01241(new_n3589, new_n3588, new_n3590);
nand_5 g01242(new_n3590, new_n3587, new_n3591);
nand_5 g01243(new_n3591, new_n3584, new_n3592);
nand_5 g01244(new_n3592, new_n3583, new_n3593);
xnor_4 g01245(new_n3577, new_n3575, new_n3594);
nand_5 g01246(new_n3594, new_n3593, new_n3595);
nand_5 g01247(new_n3595, new_n3579, new_n3596);
nand_5 g01248(new_n3596, new_n3574, new_n3597);
nand_5 g01249(new_n3597, new_n3573, new_n3598);
nand_5 g01250(new_n3598, new_n3569, new_n3599);
nand_5 g01251(new_n3599, new_n3568, new_n3600);
nand_5 g01252(new_n3600, new_n3563_1, new_n3601);
nand_5 g01253(new_n3601, new_n3562, new_n3602);
nand_5 g01254(new_n3602, new_n3558, new_n3603);
nand_5 g01255(new_n3603, new_n3557, new_n3604);
nand_5 g01256(new_n3604, new_n3552, new_n3605);
nand_5 g01257(new_n3605, new_n3551, new_n3606);
xnor_4 g01258(new_n3606, new_n3547, new_n3607);
xnor_4 g01259(new_n3607, new_n3532, new_n3608);
not_8  g01260(n24004, new_n3609);
xnor_4 g01261(new_n3604, new_n3552, new_n3610);
not_8  g01262(new_n3610, new_n3611);
nand_5 g01263(new_n3611, new_n3609, new_n3612);
xnor_4 g01264(new_n3610, new_n3609, new_n3613);
not_8  g01265(n12871, new_n3614);
xnor_4 g01266(new_n3602, new_n3558, new_n3615);
not_8  g01267(new_n3615, new_n3616);
nand_5 g01268(new_n3616, new_n3614, new_n3617_1);
xnor_4 g01269(new_n3615, new_n3614, new_n3618_1);
not_8  g01270(n23304, new_n3619);
xnor_4 g01271(new_n3600, new_n3563_1, new_n3620);
not_8  g01272(new_n3620, new_n3621);
nand_5 g01273(new_n3621, new_n3619, new_n3622);
xnor_4 g01274(new_n3620, new_n3619, new_n3623);
not_8  g01275(n19361, new_n3624);
xnor_4 g01276(new_n3598, new_n3569, new_n3625);
not_8  g01277(new_n3625, new_n3626);
nand_5 g01278(new_n3626, new_n3624, new_n3627);
xnor_4 g01279(new_n3625, new_n3624, new_n3628);
not_8  g01280(n1437, new_n3629);
xnor_4 g01281(new_n3596, new_n3574, new_n3630);
not_8  g01282(new_n3630, new_n3631);
nand_5 g01283(new_n3631, new_n3629, new_n3632);
xnor_4 g01284(new_n3630, new_n3629, new_n3633);
xnor_4 g01285(new_n3594, new_n3593, new_n3634);
nor_5  g01286(new_n3634, n4722, new_n3635);
not_8  g01287(new_n3635, new_n3636);
not_8  g01288(n4722, new_n3637);
xnor_4 g01289(new_n3634, new_n3637, new_n3638);
not_8  g01290(n14633, new_n3639);
xnor_4 g01291(new_n3591, new_n3584, new_n3640);
not_8  g01292(new_n3640, new_n3641);
nor_5  g01293(new_n3641, new_n3639, new_n3642_1);
xnor_4 g01294(new_n3640, new_n3639, new_n3643);
not_8  g01295(new_n3643, new_n3644);
not_8  g01296(n8721, new_n3645);
xnor_4 g01297(new_n3589, new_n3588, new_n3646);
not_8  g01298(new_n3646, new_n3647);
nor_5  g01299(new_n3647, new_n3645, new_n3648);
not_8  g01300(n18578, new_n3649_1);
not_8  g01301(n9251, new_n3650);
xnor_4 g01302(n16968, new_n3650, new_n3651);
not_8  g01303(new_n3651, new_n3652);
nor_5  g01304(new_n3652, new_n3649_1, new_n3653);
not_8  g01305(new_n3653, new_n3654);
xnor_4 g01306(new_n3646, n8721, new_n3655);
nor_5  g01307(new_n3655, new_n3654, new_n3656);
nor_5  g01308(new_n3656, new_n3648, new_n3657);
nor_5  g01309(new_n3657, new_n3644, new_n3658);
nor_5  g01310(new_n3658, new_n3642_1, new_n3659);
nand_5 g01311(new_n3659, new_n3638, new_n3660);
nand_5 g01312(new_n3660, new_n3636, new_n3661);
nand_5 g01313(new_n3661, new_n3633, new_n3662);
nand_5 g01314(new_n3662, new_n3632, new_n3663);
nand_5 g01315(new_n3663, new_n3628, new_n3664);
nand_5 g01316(new_n3664, new_n3627, new_n3665_1);
nand_5 g01317(new_n3665_1, new_n3623, new_n3666);
nand_5 g01318(new_n3666, new_n3622, new_n3667);
nand_5 g01319(new_n3667, new_n3618_1, new_n3668);
nand_5 g01320(new_n3668, new_n3617_1, new_n3669);
nand_5 g01321(new_n3669, new_n3613, new_n3670);
nand_5 g01322(new_n3670, new_n3612, new_n3671);
xnor_4 g01323(new_n3671, new_n3608, new_n3672);
not_8  g01324(new_n3672, new_n3673);
xnor_4 g01325(n3506, n2743, new_n3674);
not_8  g01326(n7026, new_n3675);
or_5   g01327(n14899, new_n3675, new_n3676);
xnor_4 g01328(n14899, n7026, new_n3677);
not_8  g01329(n13719, new_n3678);
or_5   g01330(n18444, new_n3678, new_n3679_1);
xnor_4 g01331(n18444, n13719, new_n3680);
not_8  g01332(n442, new_n3681);
or_5   g01333(n24638, new_n3681, new_n3682);
xnor_4 g01334(n24638, n442, new_n3683);
not_8  g01335(n9172, new_n3684);
or_5   g01336(n21674, new_n3684, new_n3685);
xnor_4 g01337(n21674, n9172, new_n3686);
not_8  g01338(n4913, new_n3687);
nor_5  g01339(n17251, new_n3687, new_n3688);
not_8  g01340(new_n3688, new_n3689);
xnor_4 g01341(n17251, n4913, new_n3690);
not_8  g01342(n604, new_n3691);
nor_5  g01343(n14790, new_n3691, new_n3692);
xnor_4 g01344(n14790, n604, new_n3693);
not_8  g01345(n10096, new_n3694);
nor_5  g01346(n16824, new_n3694, new_n3695);
not_8  g01347(n16824, new_n3696);
nor_5  g01348(new_n3696, n10096, new_n3697);
not_8  g01349(n16994, new_n3698);
nor_5  g01350(new_n3698, n16521, new_n3699);
not_8  g01351(n16521, new_n3700);
nor_5  g01352(n16994, new_n3700, new_n3701);
not_8  g01353(n7139, new_n3702);
nand_5 g01354(n9246, new_n3702, new_n3703);
nor_5  g01355(new_n3703, new_n3701, new_n3704);
nor_5  g01356(new_n3704, new_n3699, new_n3705);
nor_5  g01357(new_n3705, new_n3697, new_n3706);
nor_5  g01358(new_n3706, new_n3695, new_n3707);
nand_5 g01359(new_n3707, new_n3693, new_n3708);
not_8  g01360(new_n3708, new_n3709);
nor_5  g01361(new_n3709, new_n3692, new_n3710_1);
not_8  g01362(new_n3710_1, new_n3711);
nand_5 g01363(new_n3711, new_n3690, new_n3712);
nand_5 g01364(new_n3712, new_n3689, new_n3713);
nand_5 g01365(new_n3713, new_n3686, new_n3714);
nand_5 g01366(new_n3714, new_n3685, new_n3715);
nand_5 g01367(new_n3715, new_n3683, new_n3716);
nand_5 g01368(new_n3716, new_n3682, new_n3717);
nand_5 g01369(new_n3717, new_n3680, new_n3718);
nand_5 g01370(new_n3718, new_n3679_1, new_n3719);
nand_5 g01371(new_n3719, new_n3677, new_n3720);
nand_5 g01372(new_n3720, new_n3676, new_n3721);
xnor_4 g01373(new_n3721, new_n3674, new_n3722);
not_8  g01374(n9259, new_n3723);
not_8  g01375(n21489, new_n3724);
not_8  g01376(n13912, new_n3725_1);
not_8  g01377(n9598, new_n3726);
not_8  g01378(n11273, new_n3727);
nor_5  g01379(n25565, n21993, new_n3728);
nand_5 g01380(new_n3728, new_n3727, new_n3729);
nor_5  g01381(new_n3729, n22290, new_n3730);
nand_5 g01382(new_n3730, new_n3726, new_n3731);
nor_5  g01383(new_n3731, n7670, new_n3732);
nand_5 g01384(new_n3732, new_n3725_1, new_n3733_1);
nor_5  g01385(new_n3733_1, n20213, new_n3734);
nand_5 g01386(new_n3734, new_n3724, new_n3735);
xnor_4 g01387(new_n3735, new_n3723, new_n3736);
xnor_4 g01388(new_n3736, new_n3722, new_n3737);
not_8  g01389(new_n3677, new_n3738);
xnor_4 g01390(new_n3719, new_n3738, new_n3739);
not_8  g01391(new_n3739, new_n3740_1);
xnor_4 g01392(new_n3734, n21489, new_n3741);
not_8  g01393(new_n3741, new_n3742);
nor_5  g01394(new_n3742, new_n3740_1, new_n3743);
xnor_4 g01395(new_n3741, new_n3739, new_n3744);
xnor_4 g01396(new_n3717, new_n3680, new_n3745);
not_8  g01397(n20213, new_n3746);
xnor_4 g01398(new_n3733_1, new_n3746, new_n3747);
not_8  g01399(new_n3747, new_n3748);
nand_5 g01400(new_n3748, new_n3745, new_n3749);
xnor_4 g01401(new_n3747, new_n3745, new_n3750);
xnor_4 g01402(new_n3715, new_n3683, new_n3751);
xnor_4 g01403(new_n3732, n13912, new_n3752);
not_8  g01404(new_n3752, new_n3753);
nand_5 g01405(new_n3753, new_n3751, new_n3754);
xnor_4 g01406(new_n3752, new_n3751, new_n3755_1);
xnor_4 g01407(new_n3713, new_n3686, new_n3756);
not_8  g01408(n7670, new_n3757);
xnor_4 g01409(new_n3731, new_n3757, new_n3758_1);
not_8  g01410(new_n3758_1, new_n3759);
nand_5 g01411(new_n3759, new_n3756, new_n3760_1);
xnor_4 g01412(new_n3758_1, new_n3756, new_n3761);
xnor_4 g01413(new_n3730, n9598, new_n3762);
not_8  g01414(new_n3762, new_n3763);
xnor_4 g01415(new_n3710_1, new_n3690, new_n3764);
not_8  g01416(new_n3764, new_n3765);
nand_5 g01417(new_n3765, new_n3763, new_n3766);
xnor_4 g01418(new_n3764, new_n3763, new_n3767);
not_8  g01419(n22290, new_n3768);
xnor_4 g01420(new_n3729, new_n3768, new_n3769);
not_8  g01421(new_n3769, new_n3770);
xnor_4 g01422(new_n3707, new_n3693, new_n3771);
nand_5 g01423(new_n3771, new_n3770, new_n3772);
xnor_4 g01424(new_n3728, n11273, new_n3773);
not_8  g01425(new_n3773, new_n3774);
xnor_4 g01426(n16824, n10096, new_n3775);
xnor_4 g01427(new_n3775, new_n3705, new_n3776);
nand_5 g01428(new_n3776, new_n3774, new_n3777);
xnor_4 g01429(new_n3776, new_n3773, new_n3778);
not_8  g01430(n21993, new_n3779);
xnor_4 g01431(n25565, new_n3779, new_n3780);
not_8  g01432(new_n3780, new_n3781_1);
xnor_4 g01433(n16994, n16521, new_n3782);
xnor_4 g01434(new_n3782, new_n3703, new_n3783);
and_5  g01435(new_n3783, new_n3781_1, new_n3784);
xnor_4 g01436(n9246, n7139, new_n3785_1);
nor_5  g01437(new_n3785_1, new_n3779, new_n3786);
xnor_4 g01438(new_n3783, new_n3780, new_n3787);
not_8  g01439(new_n3787, new_n3788);
nor_5  g01440(new_n3788, new_n3786, new_n3789);
nor_5  g01441(new_n3789, new_n3784, new_n3790);
not_8  g01442(new_n3790, new_n3791);
nand_5 g01443(new_n3791, new_n3778, new_n3792);
nand_5 g01444(new_n3792, new_n3777, new_n3793);
xnor_4 g01445(new_n3771, new_n3769, new_n3794_1);
nand_5 g01446(new_n3794_1, new_n3793, new_n3795_1);
nand_5 g01447(new_n3795_1, new_n3772, new_n3796);
nand_5 g01448(new_n3796, new_n3767, new_n3797);
nand_5 g01449(new_n3797, new_n3766, new_n3798);
nand_5 g01450(new_n3798, new_n3761, new_n3799);
nand_5 g01451(new_n3799, new_n3760_1, new_n3800);
nand_5 g01452(new_n3800, new_n3755_1, new_n3801);
nand_5 g01453(new_n3801, new_n3754, new_n3802);
nand_5 g01454(new_n3802, new_n3750, new_n3803);
nand_5 g01455(new_n3803, new_n3749, new_n3804);
nor_5  g01456(new_n3804, new_n3744, new_n3805);
nor_5  g01457(new_n3805, new_n3743, new_n3806);
xnor_4 g01458(new_n3806, new_n3737, new_n3807);
xnor_4 g01459(new_n3807, new_n3673, new_n3808);
xnor_4 g01460(new_n3669, new_n3613, new_n3809);
not_8  g01461(new_n3809, new_n3810);
not_8  g01462(new_n3744, new_n3811);
xnor_4 g01463(new_n3804, new_n3811, new_n3812);
not_8  g01464(new_n3812, new_n3813);
nand_5 g01465(new_n3813, new_n3810, new_n3814);
xnor_4 g01466(new_n3812, new_n3810, new_n3815);
xnor_4 g01467(new_n3667, new_n3618_1, new_n3816);
not_8  g01468(new_n3816, new_n3817);
xnor_4 g01469(new_n3802, new_n3750, new_n3818);
not_8  g01470(new_n3818, new_n3819);
nand_5 g01471(new_n3819, new_n3817, new_n3820);
xnor_4 g01472(new_n3818, new_n3817, new_n3821);
xnor_4 g01473(new_n3665_1, new_n3623, new_n3822);
not_8  g01474(new_n3822, new_n3823);
xnor_4 g01475(new_n3800, new_n3755_1, new_n3824);
not_8  g01476(new_n3824, new_n3825);
nand_5 g01477(new_n3825, new_n3823, new_n3826);
xnor_4 g01478(new_n3824, new_n3823, new_n3827);
xnor_4 g01479(new_n3663, new_n3628, new_n3828_1);
not_8  g01480(new_n3828_1, new_n3829);
not_8  g01481(new_n3761, new_n3830);
xnor_4 g01482(new_n3798, new_n3830, new_n3831);
nand_5 g01483(new_n3831, new_n3829, new_n3832);
xnor_4 g01484(new_n3831, new_n3828_1, new_n3833);
xnor_4 g01485(new_n3661, new_n3633, new_n3834);
not_8  g01486(new_n3834, new_n3835);
xnor_4 g01487(new_n3796, new_n3767, new_n3836);
not_8  g01488(new_n3836, new_n3837);
nand_5 g01489(new_n3837, new_n3835, new_n3838);
xnor_4 g01490(new_n3836, new_n3835, new_n3839);
not_8  g01491(new_n3638, new_n3840);
xnor_4 g01492(new_n3659, new_n3840, new_n3841);
xnor_4 g01493(new_n3794_1, new_n3793, new_n3842_1);
not_8  g01494(new_n3842_1, new_n3843);
nand_5 g01495(new_n3843, new_n3841, new_n3844);
xnor_4 g01496(new_n3842_1, new_n3841, new_n3845);
xnor_4 g01497(new_n3657, new_n3643, new_n3846);
not_8  g01498(new_n3846, new_n3847);
xnor_4 g01499(new_n3790, new_n3778, new_n3848);
nand_5 g01500(new_n3848, new_n3847, new_n3849);
xnor_4 g01501(new_n3848, new_n3846, new_n3850_1);
xnor_4 g01502(new_n3787, new_n3786, new_n3851);
xnor_4 g01503(new_n3655, new_n3654, new_n3852);
nand_5 g01504(new_n3852, new_n3851, new_n3853);
xnor_4 g01505(new_n3651, new_n3649_1, new_n3854);
xnor_4 g01506(new_n3785_1, n21993, new_n3855);
and_5  g01507(new_n3855, new_n3854, new_n3856);
not_8  g01508(new_n3856, new_n3857);
not_8  g01509(new_n3852, new_n3858);
xnor_4 g01510(new_n3858, new_n3851, new_n3859);
nand_5 g01511(new_n3859, new_n3857, new_n3860);
nand_5 g01512(new_n3860, new_n3853, new_n3861);
nand_5 g01513(new_n3861, new_n3850_1, new_n3862);
nand_5 g01514(new_n3862, new_n3849, new_n3863);
nand_5 g01515(new_n3863, new_n3845, new_n3864);
nand_5 g01516(new_n3864, new_n3844, new_n3865);
nand_5 g01517(new_n3865, new_n3839, new_n3866);
nand_5 g01518(new_n3866, new_n3838, new_n3867);
nand_5 g01519(new_n3867, new_n3833, new_n3868);
nand_5 g01520(new_n3868, new_n3832, new_n3869_1);
nand_5 g01521(new_n3869_1, new_n3827, new_n3870);
nand_5 g01522(new_n3870, new_n3826, new_n3871_1);
nand_5 g01523(new_n3871_1, new_n3821, new_n3872);
nand_5 g01524(new_n3872, new_n3820, new_n3873);
nand_5 g01525(new_n3873, new_n3815, new_n3874);
nand_5 g01526(new_n3874, new_n3814, new_n3875);
xnor_4 g01527(new_n3875, new_n3808, n235);
not_8  g01528(n25749, new_n3877);
not_8  g01529(n19327, new_n3878);
not_8  g01530(n6369, new_n3879);
not_8  g01531(n15967, new_n3880);
nor_5  g01532(n25435, n13319, new_n3881);
nand_5 g01533(new_n3881, new_n3880, new_n3882);
nor_5  g01534(new_n3882, n25797, new_n3883);
nand_5 g01535(new_n3883, new_n3879, new_n3884);
nor_5  g01536(new_n3884, n21134, new_n3885);
xnor_4 g01537(new_n3885, n2113, new_n3886);
xnor_4 g01538(new_n3886, new_n3878, new_n3887);
not_8  g01539(n22597, new_n3888);
not_8  g01540(n21134, new_n3889);
xnor_4 g01541(new_n3884, new_n3889, new_n3890);
not_8  g01542(new_n3890, new_n3891_1);
nand_5 g01543(new_n3891_1, new_n3888, new_n3892);
xnor_4 g01544(new_n3890, new_n3888, new_n3893);
not_8  g01545(n26107, new_n3894);
xnor_4 g01546(new_n3883, n6369, new_n3895);
not_8  g01547(new_n3895, new_n3896);
nand_5 g01548(new_n3896, new_n3894, new_n3897);
xnor_4 g01549(new_n3895, new_n3894, new_n3898);
not_8  g01550(n342, new_n3899);
not_8  g01551(n25797, new_n3900);
xnor_4 g01552(new_n3882, new_n3900, new_n3901);
not_8  g01553(new_n3901, new_n3902);
nand_5 g01554(new_n3902, new_n3899, new_n3903);
not_8  g01555(n26553, new_n3904);
xnor_4 g01556(new_n3881, n15967, new_n3905);
not_8  g01557(new_n3905, new_n3906);
nand_5 g01558(new_n3906, new_n3904, new_n3907);
xnor_4 g01559(new_n3905, new_n3904, new_n3908);
not_8  g01560(n4964, new_n3909_1);
xnor_4 g01561(n25435, n13319, new_n3910);
nand_5 g01562(new_n3910, new_n3909_1, new_n3911);
nand_5 g01563(n25435, n7876, new_n3912);
xnor_4 g01564(new_n3910, n4964, new_n3913);
nand_5 g01565(new_n3913, new_n3912, new_n3914);
nand_5 g01566(new_n3914, new_n3911, new_n3915);
nand_5 g01567(new_n3915, new_n3908, new_n3916);
nand_5 g01568(new_n3916, new_n3907, new_n3917);
xnor_4 g01569(new_n3901, new_n3899, new_n3918_1);
nand_5 g01570(new_n3918_1, new_n3917, new_n3919);
nand_5 g01571(new_n3919, new_n3903, new_n3920);
nand_5 g01572(new_n3920, new_n3898, new_n3921);
nand_5 g01573(new_n3921, new_n3897, new_n3922);
nand_5 g01574(new_n3922, new_n3893, new_n3923);
nand_5 g01575(new_n3923, new_n3892, new_n3924);
xnor_4 g01576(new_n3924, new_n3887, new_n3925_1);
xnor_4 g01577(new_n3925_1, new_n3877, new_n3926);
xnor_4 g01578(new_n3922, new_n3893, new_n3927);
nand_5 g01579(new_n3927, n3161, new_n3928);
not_8  g01580(n3161, new_n3929);
xnor_4 g01581(new_n3927, new_n3929, new_n3930);
xnor_4 g01582(new_n3920, new_n3898, new_n3931);
nand_5 g01583(new_n3931, n9003, new_n3932_1);
not_8  g01584(n9003, new_n3933);
xnor_4 g01585(new_n3931, new_n3933, new_n3934_1);
xnor_4 g01586(new_n3918_1, new_n3917, new_n3935);
nand_5 g01587(new_n3935, n4957, new_n3936);
not_8  g01588(n4957, new_n3937);
xnor_4 g01589(new_n3935, new_n3937, new_n3938);
xnor_4 g01590(new_n3915, new_n3908, new_n3939);
nand_5 g01591(new_n3939, n7524, new_n3940);
not_8  g01592(n7524, new_n3941);
xnor_4 g01593(new_n3939, new_n3941, new_n3942);
xnor_4 g01594(new_n3913, new_n3912, new_n3943);
nand_5 g01595(new_n3943, n15743, new_n3944);
not_8  g01596(n20658, new_n3945_1);
not_8  g01597(n7876, new_n3946);
xnor_4 g01598(n25435, new_n3946, new_n3947);
not_8  g01599(new_n3947, new_n3948);
nor_5  g01600(new_n3948, new_n3945_1, new_n3949);
not_8  g01601(n15743, new_n3950);
xnor_4 g01602(new_n3943, new_n3950, new_n3951);
nand_5 g01603(new_n3951, new_n3949, new_n3952_1);
nand_5 g01604(new_n3952_1, new_n3944, new_n3953);
nand_5 g01605(new_n3953, new_n3942, new_n3954);
nand_5 g01606(new_n3954, new_n3940, new_n3955);
nand_5 g01607(new_n3955, new_n3938, new_n3956);
nand_5 g01608(new_n3956, new_n3936, new_n3957);
nand_5 g01609(new_n3957, new_n3934_1, new_n3958);
nand_5 g01610(new_n3958, new_n3932_1, new_n3959_1);
nand_5 g01611(new_n3959_1, new_n3930, new_n3960);
nand_5 g01612(new_n3960, new_n3928, new_n3961);
xnor_4 g01613(new_n3961, new_n3926, new_n3962_1);
xnor_4 g01614(n26510, n22332, new_n3963);
or_5   g01615(n23068, new_n2415, new_n3964);
xnor_4 g01616(n23068, n18907, new_n3965);
nor_5  g01617(n19514, new_n2406, new_n3966);
not_8  g01618(new_n3966, new_n3967);
xnor_4 g01619(n19514, n2731, new_n3968);
not_8  g01620(n19911, new_n3969);
nor_5  g01621(new_n3969, n10053, new_n3970);
not_8  g01622(new_n3970, new_n3971_1);
xnor_4 g01623(n19911, n10053, new_n3972);
nor_5  g01624(n13708, new_n3009, new_n3973);
nor_5  g01625(new_n2390, n8399, new_n3974);
not_8  g01626(n9507, new_n3975);
nor_5  g01627(n18409, new_n3975, new_n3976);
not_8  g01628(n18409, new_n3977);
nor_5  g01629(new_n3977, n9507, new_n3978);
not_8  g01630(n26979, new_n3979);
nor_5  g01631(new_n3979, n5704, new_n3980);
not_8  g01632(new_n3980, new_n3981);
nor_5  g01633(new_n3981, new_n3978, new_n3982);
nor_5  g01634(new_n3982, new_n3976, new_n3983_1);
nor_5  g01635(new_n3983_1, new_n3974, new_n3984_1);
nor_5  g01636(new_n3984_1, new_n3973, new_n3985);
nand_5 g01637(new_n3985, new_n3972, new_n3986);
nand_5 g01638(new_n3986, new_n3971_1, new_n3987);
nand_5 g01639(new_n3987, new_n3968, new_n3988);
nand_5 g01640(new_n3988, new_n3967, new_n3989);
nand_5 g01641(new_n3989, new_n3965, new_n3990);
nand_5 g01642(new_n3990, new_n3964, new_n3991);
xnor_4 g01643(new_n3991, new_n3963, new_n3992);
not_8  g01644(n626, new_n3993);
not_8  g01645(n19618, new_n3994);
nor_5  g01646(n22043, n12121, new_n3995);
nand_5 g01647(new_n3995, new_n3994, new_n3996);
nor_5  g01648(new_n3996, n1204, new_n3997);
nand_5 g01649(new_n3997, new_n3993, new_n3998);
nor_5  g01650(new_n3998, n5337, new_n3999);
xnor_4 g01651(new_n3999, n4325, new_n4000_1);
xnor_4 g01652(new_n4000_1, new_n3992, new_n4001);
xnor_4 g01653(new_n3989, new_n3965, new_n4002);
not_8  g01654(n5337, new_n4003);
xnor_4 g01655(new_n3998, new_n4003, new_n4004);
not_8  g01656(new_n4004, new_n4005);
nand_5 g01657(new_n4005, new_n4002, new_n4006);
xnor_4 g01658(new_n4004, new_n4002, new_n4007);
not_8  g01659(new_n3968, new_n4008);
xnor_4 g01660(new_n3987, new_n4008, new_n4009);
not_8  g01661(new_n4009, new_n4010_1);
xnor_4 g01662(new_n3997, n626, new_n4011);
not_8  g01663(new_n4011, new_n4012);
nand_5 g01664(new_n4012, new_n4010_1, new_n4013);
xnor_4 g01665(new_n4012, new_n4009, new_n4014_1);
not_8  g01666(n1204, new_n4015);
xnor_4 g01667(new_n3996, new_n4015, new_n4016);
not_8  g01668(new_n4016, new_n4017);
not_8  g01669(new_n3972, new_n4018);
xnor_4 g01670(new_n3985, new_n4018, new_n4019);
not_8  g01671(new_n4019, new_n4020);
nand_5 g01672(new_n4020, new_n4017, new_n4021);
xnor_4 g01673(new_n4019, new_n4017, new_n4022);
xnor_4 g01674(new_n3995, n19618, new_n4023);
not_8  g01675(new_n4023, new_n4024);
xnor_4 g01676(n13708, n8399, new_n4025);
not_8  g01677(new_n4025, new_n4026);
xnor_4 g01678(new_n4026, new_n3983_1, new_n4027);
not_8  g01679(new_n4027, new_n4028);
nand_5 g01680(new_n4028, new_n4024, new_n4029);
xnor_4 g01681(new_n4027, new_n4024, new_n4030);
not_8  g01682(n12121, new_n4031);
xnor_4 g01683(n22043, new_n4031, new_n4032);
not_8  g01684(new_n4032, new_n4033);
xnor_4 g01685(n18409, n9507, new_n4034);
xnor_4 g01686(new_n4034, new_n3980, new_n4035);
not_8  g01687(new_n4035, new_n4036);
nor_5  g01688(new_n4036, new_n4033, new_n4037);
xnor_4 g01689(n26979, n5704, new_n4038);
nor_5  g01690(new_n4038, new_n4031, new_n4039);
not_8  g01691(new_n4039, new_n4040);
xnor_4 g01692(new_n4035, new_n4033, new_n4041);
not_8  g01693(new_n4041, new_n4042);
nor_5  g01694(new_n4042, new_n4040, new_n4043);
nor_5  g01695(new_n4043, new_n4037, new_n4044);
nand_5 g01696(new_n4044, new_n4030, new_n4045);
nand_5 g01697(new_n4045, new_n4029, new_n4046);
nand_5 g01698(new_n4046, new_n4022, new_n4047);
nand_5 g01699(new_n4047, new_n4021, new_n4048);
nand_5 g01700(new_n4048, new_n4014_1, new_n4049);
nand_5 g01701(new_n4049, new_n4013, new_n4050);
nand_5 g01702(new_n4050, new_n4007, new_n4051);
nand_5 g01703(new_n4051, new_n4006, new_n4052);
xnor_4 g01704(new_n4052, new_n4001, new_n4053);
xnor_4 g01705(new_n4053, new_n3962_1, new_n4054);
xnor_4 g01706(new_n4050, new_n4007, new_n4055);
not_8  g01707(new_n4055, new_n4056);
xnor_4 g01708(new_n3959_1, new_n3930, new_n4057);
nand_5 g01709(new_n4057, new_n4056, new_n4058);
xnor_4 g01710(new_n4057, new_n4055, new_n4059);
xnor_4 g01711(new_n4048, new_n4014_1, new_n4060);
not_8  g01712(new_n4060, new_n4061);
xnor_4 g01713(new_n3957, new_n3934_1, new_n4062);
nand_5 g01714(new_n4062, new_n4061, new_n4063);
xnor_4 g01715(new_n4062, new_n4060, new_n4064);
xnor_4 g01716(new_n4046, new_n4022, new_n4065);
not_8  g01717(new_n4065, new_n4066);
xnor_4 g01718(new_n3955, new_n3938, new_n4067);
nand_5 g01719(new_n4067, new_n4066, new_n4068);
xnor_4 g01720(new_n4067, new_n4065, new_n4069);
xnor_4 g01721(new_n4044, new_n4030, new_n4070);
not_8  g01722(new_n4070, new_n4071_1);
xnor_4 g01723(new_n3953, new_n3942, new_n4072);
nand_5 g01724(new_n4072, new_n4071_1, new_n4073);
xnor_4 g01725(new_n4072, new_n4070, new_n4074);
xnor_4 g01726(new_n4041, new_n4040, new_n4075);
not_8  g01727(new_n4075, new_n4076);
xnor_4 g01728(new_n3951, new_n3949, new_n4077);
nand_5 g01729(new_n4077, new_n4076, new_n4078);
xnor_4 g01730(new_n3947, new_n3945_1, new_n4079);
xnor_4 g01731(new_n4038, n12121, new_n4080);
and_5  g01732(new_n4080, new_n4079, new_n4081);
not_8  g01733(new_n4081, new_n4082);
xnor_4 g01734(new_n4077, new_n4075, new_n4083);
nand_5 g01735(new_n4083, new_n4082, new_n4084);
nand_5 g01736(new_n4084, new_n4078, new_n4085_1);
nand_5 g01737(new_n4085_1, new_n4074, new_n4086);
nand_5 g01738(new_n4086, new_n4073, new_n4087);
nand_5 g01739(new_n4087, new_n4069, new_n4088_1);
nand_5 g01740(new_n4088_1, new_n4068, new_n4089_1);
nand_5 g01741(new_n4089_1, new_n4064, new_n4090);
nand_5 g01742(new_n4090, new_n4063, new_n4091);
nand_5 g01743(new_n4091, new_n4059, new_n4092);
nand_5 g01744(new_n4092, new_n4058, new_n4093);
xnor_4 g01745(new_n4093, new_n4054, n242);
not_8  g01746(n13677, new_n4095);
not_8  g01747(n11223, new_n4096);
not_8  g01748(n26572, new_n4097);
nor_5  g01749(n21398, n11667, new_n4098);
nand_5 g01750(new_n4098, new_n4097, new_n4099);
nor_5  g01751(new_n4099, n5115, new_n4100_1);
nand_5 g01752(new_n4100_1, new_n4096, new_n4101);
xnor_4 g01753(new_n4101, n19477, new_n4102);
xnor_4 g01754(new_n4102, n11011, new_n4103_1);
not_8  g01755(n16029, new_n4104);
xnor_4 g01756(new_n4100_1, n11223, new_n4105);
not_8  g01757(new_n4105, new_n4106);
nand_5 g01758(new_n4106, new_n4104, new_n4107);
xnor_4 g01759(new_n4105, new_n4104, new_n4108);
not_8  g01760(n16476, new_n4109);
xnor_4 g01761(new_n4099, new_n2606, new_n4110);
not_8  g01762(new_n4110, new_n4111);
nor_5  g01763(new_n4111, new_n4109, new_n4112);
xnor_4 g01764(new_n4110, new_n4109, new_n4113);
not_8  g01765(new_n4113, new_n4114);
not_8  g01766(n11615, new_n4115);
xnor_4 g01767(new_n4098, n26572, new_n4116);
not_8  g01768(new_n4116, new_n4117);
nand_5 g01769(new_n4117, new_n4115, new_n4118);
xnor_4 g01770(new_n4116, new_n4115, new_n4119_1);
not_8  g01771(n22433, new_n4120);
xnor_4 g01772(n21398, n11667, new_n4121);
nand_5 g01773(new_n4121, new_n4120, new_n4122);
nand_5 g01774(n21398, n14090, new_n4123_1);
xnor_4 g01775(new_n4121, n22433, new_n4124);
nand_5 g01776(new_n4124, new_n4123_1, new_n4125);
nand_5 g01777(new_n4125, new_n4122, new_n4126);
nand_5 g01778(new_n4126, new_n4119_1, new_n4127);
nand_5 g01779(new_n4127, new_n4118, new_n4128);
nor_5  g01780(new_n4128, new_n4114, new_n4129);
nor_5  g01781(new_n4129, new_n4112, new_n4130);
nand_5 g01782(new_n4130, new_n4108, new_n4131);
nand_5 g01783(new_n4131, new_n4107, new_n4132);
xnor_4 g01784(new_n4132, new_n4103_1, new_n4133);
xnor_4 g01785(new_n4133, new_n4095, new_n4134_1);
xnor_4 g01786(new_n4130, new_n4108, new_n4135);
nor_5  g01787(new_n4135, n18926, new_n4136);
not_8  g01788(new_n4136, new_n4137);
not_8  g01789(n5451, new_n4138);
xnor_4 g01790(new_n4128, new_n4113, new_n4139);
not_8  g01791(new_n4139, new_n4140);
nor_5  g01792(new_n4140, new_n4138, new_n4141);
xnor_4 g01793(new_n4139, new_n4138, new_n4142);
not_8  g01794(new_n4142, new_n4143);
not_8  g01795(n5330, new_n4144);
xnor_4 g01796(new_n4126, new_n4119_1, new_n4145);
not_8  g01797(new_n4145, new_n4146_1);
nor_5  g01798(new_n4146_1, new_n4144, new_n4147);
xnor_4 g01799(new_n4145, new_n4144, new_n4148);
not_8  g01800(new_n4148, new_n4149);
not_8  g01801(n7657, new_n4150_1);
xnor_4 g01802(new_n4124, new_n4123_1, new_n4151_1);
not_8  g01803(new_n4151_1, new_n4152_1);
nor_5  g01804(new_n4152_1, new_n4150_1, new_n4153_1);
not_8  g01805(new_n2581, new_n4154);
nor_5  g01806(new_n4154, new_n2579, new_n4155);
xnor_4 g01807(new_n4151_1, new_n4150_1, new_n4156);
nand_5 g01808(new_n4156, new_n4155, new_n4157);
not_8  g01809(new_n4157, new_n4158);
nor_5  g01810(new_n4158, new_n4153_1, new_n4159);
nor_5  g01811(new_n4159, new_n4149, new_n4160);
nor_5  g01812(new_n4160, new_n4147, new_n4161);
nor_5  g01813(new_n4161, new_n4143, new_n4162);
nor_5  g01814(new_n4162, new_n4141, new_n4163);
not_8  g01815(n18926, new_n4164);
xnor_4 g01816(new_n4135, new_n4164, new_n4165_1);
nand_5 g01817(new_n4165_1, new_n4163, new_n4166);
nand_5 g01818(new_n4166, new_n4137, new_n4167);
xnor_4 g01819(new_n4167, new_n4134_1, new_n4168);
not_8  g01820(n12398, new_n4169);
not_8  g01821(n19789, new_n4170);
not_8  g01822(n8285, new_n4171);
nor_5  g01823(n21687, n6729, new_n4172_1);
nand_5 g01824(new_n4172_1, new_n4171, new_n4173_1);
nor_5  g01825(new_n4173_1, n20169, new_n4174);
nand_5 g01826(new_n4174, new_n4170, new_n4175);
xnor_4 g01827(new_n4175, new_n4169, new_n4176_1);
not_8  g01828(n15424, new_n4177);
not_8  g01829(n9323, new_n4178);
nor_5  g01830(n19922, n10792, new_n4179);
nand_5 g01831(new_n4179, new_n4178, new_n4180);
nor_5  g01832(new_n4180, n1949, new_n4181);
nand_5 g01833(new_n4181, new_n4177, new_n4182);
xnor_4 g01834(new_n4182, n25694, new_n4183);
xnor_4 g01835(new_n4183, n20151, new_n4184);
not_8  g01836(n7693, new_n4185);
xnor_4 g01837(new_n4181, n15424, new_n4186_1);
not_8  g01838(new_n4186_1, new_n4187);
nor_5  g01839(new_n4187, new_n4185, new_n4188);
not_8  g01840(n10405, new_n4189);
not_8  g01841(n1949, new_n4190);
xnor_4 g01842(new_n4180, new_n4190, new_n4191);
not_8  g01843(new_n4191, new_n4192);
nor_5  g01844(new_n4192, new_n4189, new_n4193);
xnor_4 g01845(new_n4191, new_n4189, new_n4194);
not_8  g01846(new_n4194, new_n4195);
xnor_4 g01847(new_n4179, n9323, new_n4196);
nor_5  g01848(new_n4196, n11302, new_n4197);
not_8  g01849(new_n4197, new_n4198);
not_8  g01850(n11302, new_n4199);
xnor_4 g01851(new_n4196, new_n4199, new_n4200);
not_8  g01852(n17090, new_n4201);
xnor_4 g01853(n19922, n10792, new_n4202);
nand_5 g01854(new_n4202, new_n4201, new_n4203);
nand_5 g01855(n19922, n6773, new_n4204_1);
xnor_4 g01856(new_n4202, n17090, new_n4205_1);
nand_5 g01857(new_n4205_1, new_n4204_1, new_n4206);
nand_5 g01858(new_n4206, new_n4203, new_n4207);
nand_5 g01859(new_n4207, new_n4200, new_n4208);
nand_5 g01860(new_n4208, new_n4198, new_n4209);
nor_5  g01861(new_n4209, new_n4195, new_n4210);
nor_5  g01862(new_n4210, new_n4193, new_n4211);
xnor_4 g01863(new_n4186_1, new_n4185, new_n4212);
not_8  g01864(new_n4212, new_n4213);
nor_5  g01865(new_n4213, new_n4211, new_n4214);
nor_5  g01866(new_n4214, new_n4188, new_n4215_1);
not_8  g01867(new_n4215_1, new_n4216);
xnor_4 g01868(new_n4216, new_n4184, new_n4217);
xnor_4 g01869(new_n4217, new_n4176_1, new_n4218);
xnor_4 g01870(new_n4174, n19789, new_n4219);
not_8  g01871(new_n4219, new_n4220);
xnor_4 g01872(new_n4212, new_n4211, new_n4221_1);
not_8  g01873(new_n4221_1, new_n4222);
nor_5  g01874(new_n4222, new_n4220, new_n4223);
not_8  g01875(new_n4223, new_n4224_1);
xnor_4 g01876(new_n4221_1, new_n4220, new_n4225);
xnor_4 g01877(new_n4209, new_n4194, new_n4226);
not_8  g01878(n20169, new_n4227);
xnor_4 g01879(new_n4173_1, new_n4227, new_n4228);
nor_5  g01880(new_n4228, new_n4226, new_n4229);
xnor_4 g01881(new_n4228, new_n4226, new_n4230);
xnor_4 g01882(new_n4207, new_n4200, new_n4231_1);
not_8  g01883(new_n4231_1, new_n4232);
xnor_4 g01884(new_n4172_1, n8285, new_n4233);
not_8  g01885(new_n4233, new_n4234);
nor_5  g01886(new_n4234, new_n4232, new_n4235);
not_8  g01887(new_n4235, new_n4236);
xnor_4 g01888(new_n4234, new_n4231_1, new_n4237);
not_8  g01889(n6729, new_n4238);
xnor_4 g01890(n21687, new_n4238, new_n4239);
not_8  g01891(new_n4239, new_n4240);
xnor_4 g01892(new_n4205_1, new_n4204_1, new_n4241);
not_8  g01893(new_n4241, new_n4242);
nor_5  g01894(new_n4242, new_n4240, new_n4243);
not_8  g01895(new_n4243, new_n4244);
not_8  g01896(new_n2576, new_n4245);
nor_5  g01897(new_n4245, new_n2574, new_n4246);
xnor_4 g01898(new_n4241, new_n4240, new_n4247);
nand_5 g01899(new_n4247, new_n4246, new_n4248);
nand_5 g01900(new_n4248, new_n4244, new_n4249);
nand_5 g01901(new_n4249, new_n4237, new_n4250);
nand_5 g01902(new_n4250, new_n4236, new_n4251);
nor_5  g01903(new_n4251, new_n4230, new_n4252);
nor_5  g01904(new_n4252, new_n4229, new_n4253);
nand_5 g01905(new_n4253, new_n4225, new_n4254);
nand_5 g01906(new_n4254, new_n4224_1, new_n4255);
xnor_4 g01907(new_n4255, new_n4218, new_n4256_1);
xnor_4 g01908(new_n4256_1, new_n4168, new_n4257);
xnor_4 g01909(new_n4253, new_n4225, new_n4258);
xnor_4 g01910(new_n4165_1, new_n4163, new_n4259);
not_8  g01911(new_n4259, new_n4260);
nand_5 g01912(new_n4260, new_n4258, new_n4261);
xnor_4 g01913(new_n4259, new_n4258, new_n4262);
not_8  g01914(new_n4251, new_n4263);
xnor_4 g01915(new_n4263, new_n4230, new_n4264);
xnor_4 g01916(new_n4161, new_n4142, new_n4265);
not_8  g01917(new_n4265, new_n4266_1);
nand_5 g01918(new_n4266_1, new_n4264, new_n4267);
xnor_4 g01919(new_n4265, new_n4264, new_n4268);
xnor_4 g01920(new_n4159, new_n4148, new_n4269);
not_8  g01921(new_n4269, new_n4270);
xnor_4 g01922(new_n4249, new_n4237, new_n4271);
nand_5 g01923(new_n4271, new_n4270, new_n4272_1);
xnor_4 g01924(new_n4271, new_n4269, new_n4273);
xnor_4 g01925(new_n4247, new_n4246, new_n4274);
not_8  g01926(new_n4274, new_n4275);
xnor_4 g01927(new_n4156, new_n4155, new_n4276);
not_8  g01928(new_n4276, new_n4277);
nor_5  g01929(new_n4277, new_n4275, new_n4278);
not_8  g01930(new_n4278, new_n4279);
not_8  g01931(new_n2582_1, new_n4280);
nor_5  g01932(new_n4280, new_n2578_1, new_n4281);
not_8  g01933(new_n4281, new_n4282);
xnor_4 g01934(new_n4276, new_n4275, new_n4283);
nand_5 g01935(new_n4283, new_n4282, new_n4284);
nand_5 g01936(new_n4284, new_n4279, new_n4285);
nand_5 g01937(new_n4285, new_n4273, new_n4286);
nand_5 g01938(new_n4286, new_n4272_1, new_n4287);
nand_5 g01939(new_n4287, new_n4268, new_n4288);
nand_5 g01940(new_n4288, new_n4267, new_n4289);
nand_5 g01941(new_n4289, new_n4262, new_n4290);
nand_5 g01942(new_n4290, new_n4261, new_n4291);
xnor_4 g01943(new_n4291, new_n4257, n243);
xnor_4 g01944(n24786, new_n4199, new_n4293);
nor_5  g01945(n27120, n17090, new_n4294);
nand_5 g01946(n23065, n6773, new_n4295);
not_8  g01947(new_n4295, new_n4296);
xnor_4 g01948(n27120, n17090, new_n4297);
nor_5  g01949(new_n4297, new_n4296, new_n4298);
nor_5  g01950(new_n4298, new_n4294, new_n4299);
xnor_4 g01951(new_n4299, new_n4293, new_n4300);
not_8  g01952(n1689, new_n4301);
xnor_4 g01953(n20036, new_n4301, new_n4302);
not_8  g01954(n22274, new_n4303);
nor_5  g01955(new_n4303, n11192, new_n4304);
not_8  g01956(n11192, new_n4305);
nor_5  g01957(n22274, new_n4305, new_n4306_1);
not_8  g01958(n9380, new_n4307);
nand_5 g01959(n24129, new_n4307, new_n4308);
nor_5  g01960(new_n4308, new_n4306_1, new_n4309);
nor_5  g01961(new_n4309, new_n4304, new_n4310);
xnor_4 g01962(new_n4310, new_n4302, new_n4311);
xnor_4 g01963(new_n4311, new_n4300, new_n4312);
xnor_4 g01964(new_n4297, new_n4295, new_n4313);
xnor_4 g01965(n22274, n11192, new_n4314);
xnor_4 g01966(new_n4314, new_n4308, new_n4315);
nor_5  g01967(new_n4315, new_n4313, new_n4316);
xnor_4 g01968(n23065, n6773, new_n4317);
not_8  g01969(new_n4317, new_n4318);
xnor_4 g01970(n24129, n9380, new_n4319_1);
not_8  g01971(new_n4319_1, new_n4320);
nand_5 g01972(new_n4320, new_n4318, new_n4321);
xnor_4 g01973(new_n4315, new_n4313, new_n4322);
nor_5  g01974(new_n4322, new_n4321, new_n4323);
nor_5  g01975(new_n4323, new_n4316, new_n4324);
xnor_4 g01976(new_n4324, new_n4312, new_n4325_1);
not_8  g01977(new_n4325_1, new_n4326_1);
not_8  g01978(n919, new_n4327);
xnor_4 g01979(n5330, new_n4327, new_n4328);
nor_5  g01980(n25316, n7657, new_n4329);
nand_5 g01981(n25926, n20385, new_n4330);
xnor_4 g01982(n25316, new_n4150_1, new_n4331);
and_5  g01983(new_n4331, new_n4330, new_n4332);
nor_5  g01984(new_n4332, new_n4329, new_n4333);
xnor_4 g01985(new_n4333, new_n4328, new_n4334);
xnor_4 g01986(new_n4334, new_n4326_1, new_n4335);
not_8  g01987(new_n4335, new_n4336);
xnor_4 g01988(new_n4322, new_n4321, new_n4337);
not_8  g01989(new_n4330, new_n4338);
xnor_4 g01990(new_n4331, new_n4338, new_n4339);
not_8  g01991(new_n4339, new_n4340_1);
and_5  g01992(new_n4340_1, new_n4337, new_n4341);
not_8  g01993(n20385, new_n4342);
xnor_4 g01994(n25926, new_n4342, new_n4343);
not_8  g01995(new_n4343, new_n4344);
xnor_4 g01996(new_n4319_1, new_n4318, new_n4345);
nor_5  g01997(new_n4345, new_n4344, new_n4346);
not_8  g01998(new_n4346, new_n4347);
xnor_4 g01999(new_n4339, new_n4337, new_n4348);
not_8  g02000(new_n4348, new_n4349);
nor_5  g02001(new_n4349, new_n4347, new_n4350);
nor_5  g02002(new_n4350, new_n4341, new_n4351);
xnor_4 g02003(new_n4351, new_n4336, n248);
not_8  g02004(n14684, new_n4353);
nor_5  g02005(n24732, n6631, new_n4354);
nand_5 g02006(new_n4354, new_n4353, new_n4355);
nor_5  g02007(new_n4355, n17035, new_n4356);
xnor_4 g02008(new_n4356, n19905, new_n4357);
xnor_4 g02009(new_n4357, new_n3879, new_n4358);
not_8  g02010(n17035, new_n4359);
xnor_4 g02011(new_n4355, new_n4359, new_n4360);
and_5  g02012(new_n4360, n25797, new_n4361);
xnor_4 g02013(new_n4360, new_n3900, new_n4362);
not_8  g02014(new_n4362, new_n4363);
xnor_4 g02015(new_n4354, n14684, new_n4364);
not_8  g02016(new_n4364, new_n4365);
nand_5 g02017(new_n4365, new_n3880, new_n4366);
xnor_4 g02018(new_n4364, new_n3880, new_n4367);
not_8  g02019(n13319, new_n4368);
xnor_4 g02020(n24732, n6631, new_n4369);
nand_5 g02021(new_n4369, new_n4368, new_n4370);
not_8  g02022(new_n4370, new_n4371);
nand_5 g02023(n25435, n24732, new_n4372);
not_8  g02024(new_n4372, new_n4373);
xnor_4 g02025(new_n4369, n13319, new_n4374_1);
not_8  g02026(new_n4374_1, new_n4375);
nor_5  g02027(new_n4375, new_n4373, new_n4376_1);
nor_5  g02028(new_n4376_1, new_n4371, new_n4377);
not_8  g02029(new_n4377, new_n4378);
nand_5 g02030(new_n4378, new_n4367, new_n4379);
nand_5 g02031(new_n4379, new_n4366, new_n4380);
nor_5  g02032(new_n4380, new_n4363, new_n4381);
nor_5  g02033(new_n4381, new_n4361, new_n4382);
xnor_4 g02034(new_n4382, new_n4358, new_n4383);
nor_5  g02035(n14148, n1152, new_n4384);
nand_5 g02036(new_n4384, new_n2742, new_n4385);
nor_5  g02037(new_n4385, n18558, new_n4386);
xnor_4 g02038(new_n4386, n3468, new_n4387);
not_8  g02039(new_n4387, new_n4388);
xnor_4 g02040(new_n4388, n19514, new_n4389);
not_8  g02041(n18558, new_n4390);
xnor_4 g02042(new_n4385, new_n4390, new_n4391);
nand_5 g02043(new_n4391, n10053, new_n4392);
xnor_4 g02044(new_n4391, new_n3006, new_n4393);
xnor_4 g02045(new_n4384, n7149, new_n4394);
nand_5 g02046(new_n4394, n8399, new_n4395);
xnor_4 g02047(new_n4394, new_n3009, new_n4396);
xnor_4 g02048(n14148, n1152, new_n4397);
nor_5  g02049(new_n4397, new_n3975, new_n4398);
not_8  g02050(new_n4398, new_n4399);
nand_5 g02051(n26979, n1152, new_n4400);
not_8  g02052(new_n4400, new_n4401_1);
xnor_4 g02053(new_n4397, n9507, new_n4402);
nand_5 g02054(new_n4402, new_n4401_1, new_n4403);
nand_5 g02055(new_n4403, new_n4399, new_n4404);
nand_5 g02056(new_n4404, new_n4396, new_n4405);
nand_5 g02057(new_n4405, new_n4395, new_n4406);
nand_5 g02058(new_n4406, new_n4393, new_n4407);
nand_5 g02059(new_n4407, new_n4392, new_n4408);
xnor_4 g02060(new_n4408, new_n4389, new_n4409_1);
not_8  g02061(new_n4409_1, new_n4410);
not_8  g02062(n26748, new_n4411);
nor_5  g02063(n10057, n8920, new_n4412);
nand_5 g02064(new_n4412, new_n4411, new_n4413);
nor_5  g02065(new_n4413, n21276, new_n4414);
xnor_4 g02066(new_n4414, n13668, new_n4415);
xnor_4 g02067(new_n4415, new_n3993, new_n4416);
not_8  g02068(n21276, new_n4417);
xnor_4 g02069(new_n4413, new_n4417, new_n4418);
nand_5 g02070(new_n4418, n1204, new_n4419);
xnor_4 g02071(new_n4418, new_n4015, new_n4420);
xnor_4 g02072(new_n4412, n26748, new_n4421);
nand_5 g02073(new_n4421, n19618, new_n4422);
xnor_4 g02074(new_n4421, new_n3994, new_n4423);
not_8  g02075(n22043, new_n4424_1);
xnor_4 g02076(n10057, n8920, new_n4425);
nand_5 g02077(new_n4425, new_n4424_1, new_n4426_1);
not_8  g02078(new_n4426_1, new_n4427);
nand_5 g02079(n12121, n8920, new_n4428);
not_8  g02080(new_n4428, new_n4429);
xnor_4 g02081(new_n4425, n22043, new_n4430);
not_8  g02082(new_n4430, new_n4431);
nor_5  g02083(new_n4431, new_n4429, new_n4432_1);
nor_5  g02084(new_n4432_1, new_n4427, new_n4433);
nand_5 g02085(new_n4433, new_n4423, new_n4434);
nand_5 g02086(new_n4434, new_n4422, new_n4435);
nand_5 g02087(new_n4435, new_n4420, new_n4436);
nand_5 g02088(new_n4436, new_n4419, new_n4437);
xnor_4 g02089(new_n4437, new_n4416, new_n4438);
xnor_4 g02090(new_n4438, new_n4410, new_n4439);
xnor_4 g02091(new_n4406, new_n4393, new_n4440);
not_8  g02092(new_n4440, new_n4441_1);
xnor_4 g02093(new_n4435, new_n4420, new_n4442);
not_8  g02094(new_n4442, new_n4443);
nand_5 g02095(new_n4443, new_n4441_1, new_n4444);
xnor_4 g02096(new_n4442, new_n4441_1, new_n4445);
xnor_4 g02097(new_n4433, new_n4423, new_n4446);
not_8  g02098(new_n4446, new_n4447);
xnor_4 g02099(new_n4402, new_n4400, new_n4448);
xnor_4 g02100(new_n4430, new_n4429, new_n4449);
not_8  g02101(new_n4449, new_n4450);
nand_5 g02102(new_n4450, new_n4448, new_n4451_1);
not_8  g02103(n8920, new_n4452);
xnor_4 g02104(n12121, new_n4452, new_n4453);
not_8  g02105(new_n4453, new_n4454);
xnor_4 g02106(n26979, new_n2805, new_n4455);
not_8  g02107(new_n4455, new_n4456);
nor_5  g02108(new_n4456, new_n4454, new_n4457);
xnor_4 g02109(new_n4449, new_n4448, new_n4458);
nand_5 g02110(new_n4458, new_n4457, new_n4459);
nand_5 g02111(new_n4459, new_n4451_1, new_n4460);
nand_5 g02112(new_n4460, new_n4447, new_n4461);
xnor_4 g02113(new_n4404, new_n4396, new_n4462);
not_8  g02114(new_n4462, new_n4463);
xnor_4 g02115(new_n4460, new_n4446, new_n4464);
nand_5 g02116(new_n4464, new_n4463, new_n4465);
nand_5 g02117(new_n4465, new_n4461, new_n4466);
nand_5 g02118(new_n4466, new_n4445, new_n4467);
nand_5 g02119(new_n4467, new_n4444, new_n4468);
xnor_4 g02120(new_n4468, new_n4439, new_n4469);
xnor_4 g02121(new_n4469, new_n4383, new_n4470);
xnor_4 g02122(new_n4380, new_n4362, new_n4471);
not_8  g02123(new_n4471, new_n4472);
xnor_4 g02124(new_n4466, new_n4445, new_n4473);
nor_5  g02125(new_n4473, new_n4472, new_n4474);
xnor_4 g02126(new_n4473, new_n4472, new_n4475);
xnor_4 g02127(new_n4464, new_n4462, new_n4476_1);
not_8  g02128(new_n4476_1, new_n4477);
xnor_4 g02129(new_n4377, new_n4367, new_n4478_1);
nor_5  g02130(new_n4478_1, new_n4477, new_n4479);
xnor_4 g02131(new_n4478_1, new_n4477, new_n4480);
xnor_4 g02132(new_n4458, new_n4457, new_n4481);
not_8  g02133(new_n4481, new_n4482);
nor_5  g02134(new_n4482, new_n4374_1, new_n4483);
not_8  g02135(new_n4483, new_n4484);
xnor_4 g02136(new_n4374_1, new_n4373, new_n4485);
not_8  g02137(new_n4485, new_n4486);
nand_5 g02138(new_n4486, new_n4482, new_n4487);
not_8  g02139(n24732, new_n4488);
xnor_4 g02140(n25435, new_n4488, new_n4489);
not_8  g02141(new_n4489, new_n4490);
xnor_4 g02142(new_n4455, new_n4453, new_n4491);
nor_5  g02143(new_n4491, new_n4490, new_n4492);
not_8  g02144(new_n4492, new_n4493);
nand_5 g02145(new_n4493, new_n4487, new_n4494);
nand_5 g02146(new_n4494, new_n4484, new_n4495);
nor_5  g02147(new_n4495, new_n4480, new_n4496);
nor_5  g02148(new_n4496, new_n4479, new_n4497);
nor_5  g02149(new_n4497, new_n4475, new_n4498);
nor_5  g02150(new_n4498, new_n4474, new_n4499);
xnor_4 g02151(new_n4499, new_n4470, n266);
not_8  g02152(n21839, new_n4501);
or_5   g02153(n22270, new_n4501, new_n4502);
xnor_4 g02154(n22270, n21839, new_n4503);
not_8  g02155(n27089, new_n4504);
or_5   g02156(new_n4504, n8806, new_n4505);
xnor_4 g02157(n27089, n8806, new_n4506);
or_5   g02158(new_n2990, n2479, new_n4507);
xnor_4 g02159(n11841, n2479, new_n4508);
or_5   g02160(new_n2994, n9372, new_n4509);
xnor_4 g02161(n10710, n9372, new_n4510);
or_5   g02162(new_n2998, n6596, new_n4511);
xnor_4 g02163(n20929, n6596, new_n4512);
nor_5  g02164(n15289, new_n3002, new_n4513);
xnor_4 g02165(n15289, n8006, new_n4514_1);
not_8  g02166(new_n4514_1, new_n4515);
not_8  g02167(n25074, new_n4516);
nor_5  g02168(new_n4516, n6556, new_n4517);
xnor_4 g02169(n25074, n6556, new_n4518);
not_8  g02170(n22871, new_n4519);
nor_5  g02171(new_n4519, n16396, new_n4520);
not_8  g02172(n16396, new_n4521);
nor_5  g02173(n22871, new_n4521, new_n4522);
not_8  g02174(n14275, new_n4523);
nor_5  g02175(new_n4523, n9399, new_n4524);
not_8  g02176(n9399, new_n4525);
nor_5  g02177(n14275, new_n4525, new_n4526);
nand_5 g02178(n25023, new_n3078, new_n4527);
nor_5  g02179(new_n4527, new_n4526, new_n4528);
nor_5  g02180(new_n4528, new_n4524, new_n4529_1);
nor_5  g02181(new_n4529_1, new_n4522, new_n4530);
nor_5  g02182(new_n4530, new_n4520, new_n4531);
nand_5 g02183(new_n4531, new_n4518, new_n4532);
not_8  g02184(new_n4532, new_n4533);
nor_5  g02185(new_n4533, new_n4517, new_n4534);
nor_5  g02186(new_n4534, new_n4515, new_n4535);
nor_5  g02187(new_n4535, new_n4513, new_n4536);
not_8  g02188(new_n4536, new_n4537);
nand_5 g02189(new_n4537, new_n4512, new_n4538);
nand_5 g02190(new_n4538, new_n4511, new_n4539);
nand_5 g02191(new_n4539, new_n4510, new_n4540);
nand_5 g02192(new_n4540, new_n4509, new_n4541);
nand_5 g02193(new_n4541, new_n4508, new_n4542);
nand_5 g02194(new_n4542, new_n4507, new_n4543);
nand_5 g02195(new_n4543, new_n4506, new_n4544);
nand_5 g02196(new_n4544, new_n4505, new_n4545);
nand_5 g02197(new_n4545, new_n4503, new_n4546);
nand_5 g02198(new_n4546, new_n4502, new_n4547);
not_8  g02199(n23272, new_n4548);
xnor_4 g02200(new_n4545, new_n4503, new_n4549);
nand_5 g02201(new_n4549, new_n4548, new_n4550);
xnor_4 g02202(new_n4549, n23272, new_n4551);
not_8  g02203(n11481, new_n4552_1);
xnor_4 g02204(new_n4543, new_n4506, new_n4553);
nand_5 g02205(new_n4553, new_n4552_1, new_n4554);
xnor_4 g02206(new_n4553, n11481, new_n4555);
not_8  g02207(n16439, new_n4556);
xnor_4 g02208(new_n4541, new_n4508, new_n4557);
nand_5 g02209(new_n4557, new_n4556, new_n4558);
xnor_4 g02210(new_n4557, n16439, new_n4559);
not_8  g02211(n15241, new_n4560);
xnor_4 g02212(new_n4539, new_n4510, new_n4561);
nand_5 g02213(new_n4561, new_n4560, new_n4562);
xnor_4 g02214(new_n4561, n15241, new_n4563);
not_8  g02215(n7678, new_n4564);
xnor_4 g02216(new_n4537, new_n4512, new_n4565);
nand_5 g02217(new_n4565, new_n4564, new_n4566);
xnor_4 g02218(new_n4565, n7678, new_n4567);
not_8  g02219(n3785, new_n4568);
xnor_4 g02220(new_n4534, new_n4514_1, new_n4569);
not_8  g02221(new_n4569, new_n4570);
nand_5 g02222(new_n4570, new_n4568, new_n4571);
xnor_4 g02223(new_n4569, new_n4568, new_n4572);
not_8  g02224(n20250, new_n4573);
xnor_4 g02225(new_n4531, new_n4518, new_n4574);
nand_5 g02226(new_n4574, new_n4573, new_n4575);
xnor_4 g02227(new_n4574, n20250, new_n4576);
not_8  g02228(n5822, new_n4577);
xnor_4 g02229(n22871, n16396, new_n4578);
xnor_4 g02230(new_n4578, new_n4529_1, new_n4579);
nor_5  g02231(new_n4579, new_n4577, new_n4580);
not_8  g02232(new_n4579, new_n4581);
nor_5  g02233(new_n4581, n5822, new_n4582);
xnor_4 g02234(n14275, n9399, new_n4583);
xnor_4 g02235(new_n4583, new_n4527, new_n4584);
not_8  g02236(new_n4584, new_n4585);
nor_5  g02237(new_n4585, n26443, new_n4586);
xnor_4 g02238(n25023, n2088, new_n4587);
nor_5  g02239(new_n4587, new_n2568, new_n4588_1);
xnor_4 g02240(new_n4584, n26443, new_n4589);
not_8  g02241(new_n4589, new_n4590_1);
nor_5  g02242(new_n4590_1, new_n4588_1, new_n4591);
nor_5  g02243(new_n4591, new_n4586, new_n4592);
not_8  g02244(new_n4592, new_n4593);
nor_5  g02245(new_n4593, new_n4582, new_n4594);
nor_5  g02246(new_n4594, new_n4580, new_n4595_1);
nand_5 g02247(new_n4595_1, new_n4576, new_n4596);
nand_5 g02248(new_n4596, new_n4575, new_n4597);
nand_5 g02249(new_n4597, new_n4572, new_n4598);
nand_5 g02250(new_n4598, new_n4571, new_n4599);
nand_5 g02251(new_n4599, new_n4567, new_n4600);
nand_5 g02252(new_n4600, new_n4566, new_n4601);
nand_5 g02253(new_n4601, new_n4563, new_n4602);
nand_5 g02254(new_n4602, new_n4562, new_n4603);
nand_5 g02255(new_n4603, new_n4559, new_n4604);
nand_5 g02256(new_n4604, new_n4558, new_n4605);
nand_5 g02257(new_n4605, new_n4555, new_n4606);
nand_5 g02258(new_n4606, new_n4554, new_n4607);
nand_5 g02259(new_n4607, new_n4551, new_n4608);
nand_5 g02260(new_n4608, new_n4550, new_n4609);
nor_5  g02261(new_n4609, new_n4547, new_n4610);
nor_5  g02262(new_n4101, n19477, new_n4611);
nand_5 g02263(new_n4611, new_n2595, new_n4612);
nor_5  g02264(new_n4612, n25168, new_n4613);
nand_5 g02265(new_n4613, new_n2588, new_n4614);
or_5   g02266(new_n4614, n9396, new_n4615);
xnor_4 g02267(new_n4614, new_n2584, new_n4616);
or_5   g02268(new_n4616, n18880, new_n4617);
not_8  g02269(n25475, new_n4618);
xnor_4 g02270(new_n4613, n1999, new_n4619);
not_8  g02271(new_n4619, new_n4620);
nand_5 g02272(new_n4620, new_n4618, new_n4621);
xnor_4 g02273(new_n4619, new_n4618, new_n4622);
not_8  g02274(n23849, new_n4623);
xnor_4 g02275(new_n4612, n25168, new_n4624_1);
nand_5 g02276(new_n4624_1, new_n4623, new_n4625);
xnor_4 g02277(new_n4624_1, n23849, new_n4626);
not_8  g02278(n12446, new_n4627);
xnor_4 g02279(new_n4611, n9318, new_n4628);
not_8  g02280(new_n4628, new_n4629);
nand_5 g02281(new_n4629, new_n4627, new_n4630);
not_8  g02282(n11011, new_n4631);
nand_5 g02283(new_n4102, new_n4631, new_n4632);
nand_5 g02284(new_n4132, new_n4103_1, new_n4633);
nand_5 g02285(new_n4633, new_n4632, new_n4634);
xnor_4 g02286(new_n4628, new_n4627, new_n4635);
nand_5 g02287(new_n4635, new_n4634, new_n4636);
nand_5 g02288(new_n4636, new_n4630, new_n4637);
nand_5 g02289(new_n4637, new_n4626, new_n4638);
nand_5 g02290(new_n4638, new_n4625, new_n4639);
nand_5 g02291(new_n4639, new_n4622, new_n4640);
nand_5 g02292(new_n4640, new_n4621, new_n4641);
nand_5 g02293(new_n4616, n18880, new_n4642);
nand_5 g02294(new_n4642, new_n4641, new_n4643);
nand_5 g02295(new_n4643, new_n4617, new_n4644);
nand_5 g02296(new_n4644, new_n4615, new_n4645);
not_8  g02297(new_n4645, new_n4646_1);
not_8  g02298(n24196, new_n4647);
not_8  g02299(n25381, new_n4648);
not_8  g02300(n268, new_n4649);
not_8  g02301(n6785, new_n4650);
nor_5  g02302(n24032, n22843, new_n4651);
nand_5 g02303(new_n4651, new_n4650, new_n4652);
nor_5  g02304(new_n4652, n24879, new_n4653);
nand_5 g02305(new_n4653, new_n4649, new_n4654);
nor_5  g02306(new_n4654, n12587, new_n4655);
nand_5 g02307(new_n4655, new_n4648, new_n4656);
nor_5  g02308(new_n4656, n16376, new_n4657);
and_5  g02309(new_n4657, new_n4647, new_n4658);
xnor_4 g02310(new_n4658, n18105, new_n4659);
not_8  g02311(new_n4659, new_n4660);
not_8  g02312(n18880, new_n4661);
xnor_4 g02313(new_n4616, new_n4661, new_n4662);
xnor_4 g02314(new_n4662, new_n4641, new_n4663);
not_8  g02315(new_n4663, new_n4664);
nor_5  g02316(new_n4664, new_n4660, new_n4665_1);
not_8  g02317(new_n4665_1, new_n4666);
not_8  g02318(n18105, new_n4667);
and_5  g02319(new_n4658, new_n4667, new_n4668);
xnor_4 g02320(new_n4663, new_n4659, new_n4669);
xnor_4 g02321(new_n4657, new_n4647, new_n4670);
xnor_4 g02322(new_n4639, new_n4622, new_n4671);
not_8  g02323(new_n4671, new_n4672);
nand_5 g02324(new_n4672, new_n4670, new_n4673);
xnor_4 g02325(new_n4671, new_n4670, new_n4674_1);
xnor_4 g02326(new_n4656, n16376, new_n4675);
xnor_4 g02327(new_n4637, new_n4626, new_n4676);
not_8  g02328(new_n4676, new_n4677);
nand_5 g02329(new_n4677, new_n4675, new_n4678);
xnor_4 g02330(new_n4676, new_n4675, new_n4679);
xnor_4 g02331(new_n4655, n25381, new_n4680);
not_8  g02332(new_n4680, new_n4681);
xnor_4 g02333(new_n4635, new_n4634, new_n4682);
not_8  g02334(new_n4682, new_n4683);
nand_5 g02335(new_n4683, new_n4681, new_n4684);
xnor_4 g02336(new_n4682, new_n4681, new_n4685);
not_8  g02337(new_n4133, new_n4686);
not_8  g02338(n12587, new_n4687);
xnor_4 g02339(new_n4654, new_n4687, new_n4688);
not_8  g02340(new_n4688, new_n4689);
nand_5 g02341(new_n4689, new_n4686, new_n4690);
xnor_4 g02342(new_n4689, new_n4133, new_n4691);
not_8  g02343(new_n4135, new_n4692);
xnor_4 g02344(new_n4653, n268, new_n4693_1);
not_8  g02345(new_n4693_1, new_n4694);
nand_5 g02346(new_n4694, new_n4692, new_n4695);
not_8  g02347(n24879, new_n4696);
xnor_4 g02348(new_n4652, new_n4696, new_n4697);
not_8  g02349(new_n4697, new_n4698);
nand_5 g02350(new_n4698, new_n4140, new_n4699);
xnor_4 g02351(new_n4698, new_n4139, new_n4700);
xnor_4 g02352(new_n4651, new_n4650, new_n4701);
nor_5  g02353(new_n4701, new_n4146_1, new_n4702);
xnor_4 g02354(new_n4701, new_n4146_1, new_n4703);
not_8  g02355(n22843, new_n4704);
xnor_4 g02356(n24032, new_n4704, new_n4705);
nor_5  g02357(new_n4705, new_n4151_1, new_n4706);
not_8  g02358(new_n4706, new_n4707);
nor_5  g02359(new_n4154, new_n4704, new_n4708);
not_8  g02360(new_n4708, new_n4709);
xnor_4 g02361(new_n4705, new_n4152_1, new_n4710);
nand_5 g02362(new_n4710, new_n4709, new_n4711);
nand_5 g02363(new_n4711, new_n4707, new_n4712);
nor_5  g02364(new_n4712, new_n4703, new_n4713);
nor_5  g02365(new_n4713, new_n4702, new_n4714);
nand_5 g02366(new_n4714, new_n4700, new_n4715);
nand_5 g02367(new_n4715, new_n4699, new_n4716);
xnor_4 g02368(new_n4694, new_n4135, new_n4717);
nand_5 g02369(new_n4717, new_n4716, new_n4718);
nand_5 g02370(new_n4718, new_n4695, new_n4719);
nand_5 g02371(new_n4719, new_n4691, new_n4720);
nand_5 g02372(new_n4720, new_n4690, new_n4721);
nand_5 g02373(new_n4721, new_n4685, new_n4722_1);
nand_5 g02374(new_n4722_1, new_n4684, new_n4723);
nand_5 g02375(new_n4723, new_n4679, new_n4724);
nand_5 g02376(new_n4724, new_n4678, new_n4725);
nand_5 g02377(new_n4725, new_n4674_1, new_n4726);
nand_5 g02378(new_n4726, new_n4673, new_n4727);
nor_5  g02379(new_n4727, new_n4669, new_n4728);
nor_5  g02380(new_n4728, new_n4668, new_n4729);
nand_5 g02381(new_n4729, new_n4666, new_n4730);
nor_5  g02382(new_n4730, new_n4646_1, new_n4731_1);
not_8  g02383(new_n4731_1, new_n4732);
xnor_4 g02384(new_n4732, new_n4610, new_n4733);
not_8  g02385(new_n4547, new_n4734);
xnor_4 g02386(new_n4609, new_n4734, new_n4735);
xnor_4 g02387(new_n4730, new_n4646_1, new_n4736);
nor_5  g02388(new_n4736, new_n4735, new_n4737);
not_8  g02389(new_n4737, new_n4738);
not_8  g02390(new_n4735, new_n4739);
xnor_4 g02391(new_n4736, new_n4739, new_n4740);
not_8  g02392(new_n4669, new_n4741);
xnor_4 g02393(new_n4727, new_n4741, new_n4742);
not_8  g02394(new_n4742, new_n4743);
xnor_4 g02395(new_n4607, new_n4551, new_n4744);
not_8  g02396(new_n4744, new_n4745_1);
nand_5 g02397(new_n4745_1, new_n4743, new_n4746);
xnor_4 g02398(new_n4744, new_n4743, new_n4747_1);
xnor_4 g02399(new_n4725, new_n4674_1, new_n4748);
not_8  g02400(new_n4748, new_n4749);
not_8  g02401(new_n4555, new_n4750);
xnor_4 g02402(new_n4605, new_n4750, new_n4751);
nand_5 g02403(new_n4751, new_n4749, new_n4752);
xnor_4 g02404(new_n4751, new_n4748, new_n4753);
xnor_4 g02405(new_n4723, new_n4679, new_n4754);
not_8  g02406(new_n4754, new_n4755);
not_8  g02407(new_n4559, new_n4756);
xnor_4 g02408(new_n4603, new_n4756, new_n4757);
nand_5 g02409(new_n4757, new_n4755, new_n4758);
xnor_4 g02410(new_n4757, new_n4754, new_n4759);
xnor_4 g02411(new_n4721, new_n4685, new_n4760);
not_8  g02412(new_n4760, new_n4761);
not_8  g02413(new_n4563, new_n4762);
xnor_4 g02414(new_n4601, new_n4762, new_n4763);
nand_5 g02415(new_n4763, new_n4761, new_n4764);
xnor_4 g02416(new_n4763, new_n4760, new_n4765);
xnor_4 g02417(new_n4719, new_n4691, new_n4766_1);
not_8  g02418(new_n4766_1, new_n4767);
xnor_4 g02419(new_n4599, new_n4567, new_n4768);
not_8  g02420(new_n4768, new_n4769);
nand_5 g02421(new_n4769, new_n4767, new_n4770_1);
xnor_4 g02422(new_n4769, new_n4766_1, new_n4771);
xnor_4 g02423(new_n4597, new_n4572, new_n4772);
not_8  g02424(new_n4772, new_n4773);
not_8  g02425(new_n4717, new_n4774);
xnor_4 g02426(new_n4774, new_n4716, new_n4775);
nand_5 g02427(new_n4775, new_n4773, new_n4776);
xnor_4 g02428(new_n4775, new_n4772, new_n4777_1);
xnor_4 g02429(new_n4714, new_n4700, new_n4778);
not_8  g02430(new_n4778, new_n4779);
xnor_4 g02431(new_n4595_1, new_n4576, new_n4780);
not_8  g02432(new_n4780, new_n4781);
nand_5 g02433(new_n4781, new_n4779, new_n4782);
xnor_4 g02434(new_n4781, new_n4778, new_n4783);
xnor_4 g02435(new_n4712, new_n4703, new_n4784);
xnor_4 g02436(new_n4579, n5822, new_n4785_1);
xnor_4 g02437(new_n4785_1, new_n4593, new_n4786);
not_8  g02438(new_n4786, new_n4787);
nor_5  g02439(new_n4787, new_n4784, new_n4788);
xnor_4 g02440(new_n4589, new_n4588_1, new_n4789);
not_8  g02441(new_n4789, new_n4790);
xnor_4 g02442(new_n4710, new_n4709, new_n4791);
nor_5  g02443(new_n4791, new_n4790, new_n4792);
not_8  g02444(new_n4792, new_n4793);
xnor_4 g02445(new_n2581, new_n4704, new_n4794);
xnor_4 g02446(new_n4587, n1681, new_n4795);
and_5  g02447(new_n4795, new_n4794, new_n4796);
not_8  g02448(new_n4796, new_n4797);
xnor_4 g02449(new_n4791, new_n4789, new_n4798);
nand_5 g02450(new_n4798, new_n4797, new_n4799);
nand_5 g02451(new_n4799, new_n4793, new_n4800);
xnor_4 g02452(new_n4787, new_n4784, new_n4801);
nor_5  g02453(new_n4801, new_n4800, new_n4802);
nor_5  g02454(new_n4802, new_n4788, new_n4803);
nand_5 g02455(new_n4803, new_n4783, new_n4804_1);
nand_5 g02456(new_n4804_1, new_n4782, new_n4805);
nand_5 g02457(new_n4805, new_n4777_1, new_n4806);
nand_5 g02458(new_n4806, new_n4776, new_n4807);
nand_5 g02459(new_n4807, new_n4771, new_n4808);
nand_5 g02460(new_n4808, new_n4770_1, new_n4809);
nand_5 g02461(new_n4809, new_n4765, new_n4810_1);
nand_5 g02462(new_n4810_1, new_n4764, new_n4811);
nand_5 g02463(new_n4811, new_n4759, new_n4812_1);
nand_5 g02464(new_n4812_1, new_n4758, new_n4813);
nand_5 g02465(new_n4813, new_n4753, new_n4814_1);
nand_5 g02466(new_n4814_1, new_n4752, new_n4815);
nand_5 g02467(new_n4815, new_n4747_1, new_n4816);
nand_5 g02468(new_n4816, new_n4746, new_n4817);
nand_5 g02469(new_n4817, new_n4740, new_n4818);
nand_5 g02470(new_n4818, new_n4738, new_n4819);
xnor_4 g02471(new_n4819, new_n4733, n298);
xnor_4 g02472(n21735, n20604, new_n4821);
not_8  g02473(n24085, new_n4822);
nor_5  g02474(new_n4822, n16158, new_n4823);
not_8  g02475(new_n4823, new_n4824);
xnor_4 g02476(n24085, n16158, new_n4825);
not_8  g02477(n14071, new_n4826);
nor_5  g02478(new_n4826, n5752, new_n4827);
xnor_4 g02479(n14071, n5752, new_n4828);
not_8  g02480(n18171, new_n4829);
nor_5  g02481(new_n4829, n1738, new_n4830);
not_8  g02482(n1738, new_n4831);
nor_5  g02483(n18171, new_n4831, new_n4832);
not_8  g02484(n25073, new_n4833);
nor_5  g02485(new_n4833, n12152, new_n4834);
not_8  g02486(n12152, new_n4835);
nor_5  g02487(n25073, new_n4835, new_n4836);
not_8  g02488(n19107, new_n4837);
nand_5 g02489(n22309, new_n4837, new_n4838);
nor_5  g02490(new_n4838, new_n4836, new_n4839);
nor_5  g02491(new_n4839, new_n4834, new_n4840);
nor_5  g02492(new_n4840, new_n4832, new_n4841);
nor_5  g02493(new_n4841, new_n4830, new_n4842);
and_5  g02494(new_n4842, new_n4828, new_n4843);
nor_5  g02495(new_n4843, new_n4827, new_n4844);
not_8  g02496(new_n4844, new_n4845);
nand_5 g02497(new_n4845, new_n4825, new_n4846);
nand_5 g02498(new_n4846, new_n4824, new_n4847);
xnor_4 g02499(new_n4847, new_n4821, new_n4848);
xnor_4 g02500(n4119, n1525, new_n4849);
not_8  g02501(n16988, new_n4850_1);
nor_5  g02502(new_n4850_1, n14510, new_n4851);
xnor_4 g02503(n16988, n14510, new_n4852);
not_8  g02504(new_n4852, new_n4853);
not_8  g02505(n21779, new_n4854);
nor_5  g02506(new_n4854, n13263, new_n4855);
xnor_4 g02507(n21779, n13263, new_n4856);
nor_5  g02508(new_n3580, n5376, new_n4857);
not_8  g02509(n5376, new_n4858_1);
nor_5  g02510(n20455, new_n4858_1, new_n4859);
nor_5  g02511(n5128, new_n3585, new_n4860);
not_8  g02512(n5128, new_n4861);
nor_5  g02513(new_n4861, n1639, new_n4862);
not_8  g02514(n16968, new_n4863);
nor_5  g02515(n23120, new_n4863, new_n4864);
not_8  g02516(new_n4864, new_n4865);
nor_5  g02517(new_n4865, new_n4862, new_n4866);
nor_5  g02518(new_n4866, new_n4860, new_n4867);
nor_5  g02519(new_n4867, new_n4859, new_n4868);
nor_5  g02520(new_n4868, new_n4857, new_n4869);
nand_5 g02521(new_n4869, new_n4856, new_n4870);
not_8  g02522(new_n4870, new_n4871);
nor_5  g02523(new_n4871, new_n4855, new_n4872);
nor_5  g02524(new_n4872, new_n4853, new_n4873);
nor_5  g02525(new_n4873, new_n4851, new_n4874);
xnor_4 g02526(new_n4874, new_n4849, new_n4875);
xnor_4 g02527(n12626, n4272, new_n4876);
not_8  g02528(n24319, new_n4877);
nor_5  g02529(new_n4877, n6971, new_n4878);
xnor_4 g02530(n24319, n6971, new_n4879);
not_8  g02531(new_n4879, new_n4880);
not_8  g02532(n7460, new_n4881);
nor_5  g02533(n22068, new_n4881, new_n4882);
xnor_4 g02534(n22068, n7460, new_n4883);
not_8  g02535(n9460, new_n4884);
nor_5  g02536(new_n4884, n196, new_n4885);
not_8  g02537(n196, new_n4886);
nor_5  g02538(n9460, new_n4886, new_n4887);
not_8  g02539(n14954, new_n4888);
nor_5  g02540(new_n4888, n11749, new_n4889);
not_8  g02541(n11749, new_n4890);
nor_5  g02542(n14954, new_n4890, new_n4891_1);
not_8  g02543(n13424, new_n4892);
nand_5 g02544(n23831, new_n4892, new_n4893);
nor_5  g02545(new_n4893, new_n4891_1, new_n4894);
nor_5  g02546(new_n4894, new_n4889, new_n4895);
nor_5  g02547(new_n4895, new_n4887, new_n4896);
nor_5  g02548(new_n4896, new_n4885, new_n4897);
nand_5 g02549(new_n4897, new_n4883, new_n4898);
not_8  g02550(new_n4898, new_n4899);
nor_5  g02551(new_n4899, new_n4882, new_n4900);
nor_5  g02552(new_n4900, new_n4880, new_n4901);
nor_5  g02553(new_n4901, new_n4878, new_n4902);
xnor_4 g02554(new_n4902, new_n4876, new_n4903);
not_8  g02555(new_n4903, new_n4904);
xnor_4 g02556(new_n4904, new_n4875, new_n4905);
xnor_4 g02557(new_n4872, new_n4852, new_n4906);
not_8  g02558(new_n4906, new_n4907);
xnor_4 g02559(new_n4900, new_n4879, new_n4908);
not_8  g02560(new_n4908, new_n4909);
nor_5  g02561(new_n4909, new_n4907, new_n4910);
not_8  g02562(new_n4910, new_n4911);
xnor_4 g02563(new_n4909, new_n4906, new_n4912);
xnor_4 g02564(new_n4869, new_n4856, new_n4913_1);
not_8  g02565(new_n4913_1, new_n4914);
xnor_4 g02566(new_n4897, new_n4883, new_n4915);
not_8  g02567(new_n4915, new_n4916);
nor_5  g02568(new_n4916, new_n4914, new_n4917);
not_8  g02569(new_n4917, new_n4918);
xnor_4 g02570(new_n4916, new_n4913_1, new_n4919);
xnor_4 g02571(n20455, n5376, new_n4920);
xnor_4 g02572(new_n4920, new_n4867, new_n4921);
not_8  g02573(new_n4921, new_n4922);
xnor_4 g02574(n9460, n196, new_n4923);
xnor_4 g02575(new_n4923, new_n4895, new_n4924);
not_8  g02576(new_n4924, new_n4925_1);
nor_5  g02577(new_n4925_1, new_n4922, new_n4926);
not_8  g02578(new_n4926, new_n4927);
xnor_4 g02579(new_n4925_1, new_n4921, new_n4928);
xnor_4 g02580(n5128, n1639, new_n4929);
xnor_4 g02581(new_n4929, new_n4865, new_n4930);
xnor_4 g02582(n14954, n11749, new_n4931);
xnor_4 g02583(new_n4931, new_n4893, new_n4932);
nor_5  g02584(new_n4932, new_n4930, new_n4933);
xnor_4 g02585(n23120, n16968, new_n4934);
xnor_4 g02586(n23831, n13424, new_n4935);
nor_5  g02587(new_n4935, new_n4934, new_n4936);
not_8  g02588(new_n4932, new_n4937);
xnor_4 g02589(new_n4937, new_n4930, new_n4938);
nand_5 g02590(new_n4938, new_n4936, new_n4939_1);
not_8  g02591(new_n4939_1, new_n4940);
nor_5  g02592(new_n4940, new_n4933, new_n4941);
nand_5 g02593(new_n4941, new_n4928, new_n4942);
nand_5 g02594(new_n4942, new_n4927, new_n4943);
nand_5 g02595(new_n4943, new_n4919, new_n4944);
nand_5 g02596(new_n4944, new_n4918, new_n4945);
not_8  g02597(new_n4945, new_n4946);
nand_5 g02598(new_n4946, new_n4912, new_n4947_1);
nand_5 g02599(new_n4947_1, new_n4911, new_n4948);
xnor_4 g02600(new_n4948, new_n4905, new_n4949);
xnor_4 g02601(new_n4949, new_n4848, new_n4950);
xnor_4 g02602(new_n4844, new_n4825, new_n4951);
xnor_4 g02603(new_n4945, new_n4912, new_n4952_1);
nor_5  g02604(new_n4952_1, new_n4951, new_n4953);
not_8  g02605(new_n4953, new_n4954);
not_8  g02606(new_n4952_1, new_n4955);
xnor_4 g02607(new_n4955, new_n4951, new_n4956);
xnor_4 g02608(new_n4943, new_n4919, new_n4957_1);
xnor_4 g02609(new_n4842, new_n4828, new_n4958);
not_8  g02610(new_n4958, new_n4959);
nor_5  g02611(new_n4959, new_n4957_1, new_n4960);
not_8  g02612(new_n4960, new_n4961);
xnor_4 g02613(new_n4941, new_n4928, new_n4962);
xnor_4 g02614(n18171, n1738, new_n4963);
xnor_4 g02615(new_n4963, new_n4840, new_n4964_1);
not_8  g02616(new_n4964_1, new_n4965);
nor_5  g02617(new_n4965, new_n4962, new_n4966_1);
not_8  g02618(new_n4966_1, new_n4967_1);
xnor_4 g02619(new_n4964_1, new_n4962, new_n4968);
xnor_4 g02620(n22309, n19107, new_n4969);
not_8  g02621(new_n4934, new_n4970);
xnor_4 g02622(new_n4935, new_n4970, new_n4971);
not_8  g02623(new_n4971, new_n4972_1);
nor_5  g02624(new_n4972_1, new_n4969, new_n4973);
xnor_4 g02625(n25073, n12152, new_n4974);
xnor_4 g02626(new_n4974, new_n4838, new_n4975);
not_8  g02627(new_n4975, new_n4976);
nor_5  g02628(new_n4976, new_n4973, new_n4977);
xnor_4 g02629(new_n4938, new_n4936, new_n4978);
xnor_4 g02630(new_n4975, new_n4973, new_n4979);
and_5  g02631(new_n4979, new_n4978, new_n4980);
nor_5  g02632(new_n4980, new_n4977, new_n4981);
not_8  g02633(new_n4981, new_n4982);
nand_5 g02634(new_n4982, new_n4968, new_n4983);
nand_5 g02635(new_n4983, new_n4967_1, new_n4984);
xnor_4 g02636(new_n4958, new_n4957_1, new_n4985);
nand_5 g02637(new_n4985, new_n4984, new_n4986);
nand_5 g02638(new_n4986, new_n4961, new_n4987);
nand_5 g02639(new_n4987, new_n4956, new_n4988);
nand_5 g02640(new_n4988, new_n4954, new_n4989);
xor_4  g02641(new_n4989, new_n4950, n317);
or_5   g02642(n9934, n3506, new_n4991);
not_8  g02643(n3506, new_n4992);
xnor_4 g02644(n9934, new_n4992, new_n4993);
or_5   g02645(n18496, n14899, new_n4994);
not_8  g02646(n14899, new_n4995);
xnor_4 g02647(n18496, new_n4995, new_n4996);
or_5   g02648(n26224, n18444, new_n4997);
not_8  g02649(n18444, new_n4998);
xnor_4 g02650(n26224, new_n4998, new_n4999);
nor_5  g02651(n24638, n19327, new_n5000);
xnor_4 g02652(n24638, new_n3878, new_n5001);
not_8  g02653(new_n5001, new_n5002);
nor_5  g02654(n22597, n21674, new_n5003);
not_8  g02655(n21674, new_n5004);
xnor_4 g02656(n22597, new_n5004, new_n5005);
not_8  g02657(new_n5005, new_n5006);
nor_5  g02658(n26107, n17251, new_n5007);
not_8  g02659(n17251, new_n5008);
xnor_4 g02660(n26107, new_n5008, new_n5009);
not_8  g02661(new_n5009, new_n5010);
nor_5  g02662(n14790, n342, new_n5011_1);
xnor_4 g02663(n14790, new_n3899, new_n5012);
not_8  g02664(new_n5012, new_n5013);
nor_5  g02665(n26553, n10096, new_n5014);
xnor_4 g02666(n26553, new_n3694, new_n5015);
not_8  g02667(new_n5015, new_n5016);
nor_5  g02668(n16994, n4964, new_n5017);
nand_5 g02669(n9246, n7876, new_n5018);
not_8  g02670(new_n5018, new_n5019);
xnor_4 g02671(n16994, new_n3909_1, new_n5020_1);
not_8  g02672(new_n5020_1, new_n5021);
nor_5  g02673(new_n5021, new_n5019, new_n5022);
nor_5  g02674(new_n5022, new_n5017, new_n5023);
nor_5  g02675(new_n5023, new_n5016, new_n5024_1);
nor_5  g02676(new_n5024_1, new_n5014, new_n5025_1);
nor_5  g02677(new_n5025_1, new_n5013, new_n5026_1);
nor_5  g02678(new_n5026_1, new_n5011_1, new_n5027);
nor_5  g02679(new_n5027, new_n5010, new_n5028);
nor_5  g02680(new_n5028, new_n5007, new_n5029);
nor_5  g02681(new_n5029, new_n5006, new_n5030);
nor_5  g02682(new_n5030, new_n5003, new_n5031_1);
nor_5  g02683(new_n5031_1, new_n5002, new_n5032);
nor_5  g02684(new_n5032, new_n5000, new_n5033);
not_8  g02685(new_n5033, new_n5034);
nand_5 g02686(new_n5034, new_n4999, new_n5035);
nand_5 g02687(new_n5035, new_n4997, new_n5036);
nand_5 g02688(new_n5036, new_n4996, new_n5037);
nand_5 g02689(new_n5037, new_n4994, new_n5038);
nand_5 g02690(new_n5038, new_n4993, new_n5039);
nand_5 g02691(new_n5039, new_n4991, new_n5040);
not_8  g02692(new_n5040, new_n5041);
not_8  g02693(n2979, new_n5042);
xnor_4 g02694(n9554, new_n5042, new_n5043);
not_8  g02695(new_n5043, new_n5044);
or_5   g02696(n26408, n647, new_n5045);
not_8  g02697(n647, new_n5046_1);
xnor_4 g02698(n26408, new_n5046_1, new_n5047);
or_5   g02699(n20409, n18227, new_n5048);
not_8  g02700(n18227, new_n5049);
xnor_4 g02701(n20409, new_n5049, new_n5050);
nor_5  g02702(n25749, n7377, new_n5051);
not_8  g02703(new_n5051, new_n5052);
not_8  g02704(n7377, new_n5053);
xnor_4 g02705(n25749, new_n5053, new_n5054);
nor_5  g02706(n11630, n3161, new_n5055);
not_8  g02707(new_n5055, new_n5056);
xnor_4 g02708(n11630, new_n3929, new_n5057);
nor_5  g02709(n13453, n9003, new_n5058);
not_8  g02710(new_n5058, new_n5059);
xnor_4 g02711(n13453, new_n3933, new_n5060_1);
nor_5  g02712(n7421, n4957, new_n5061);
xnor_4 g02713(n7421, new_n3937, new_n5062_1);
not_8  g02714(new_n5062_1, new_n5063);
nor_5  g02715(n19680, n7524, new_n5064_1);
xnor_4 g02716(n19680, new_n3941, new_n5065);
not_8  g02717(new_n5065, new_n5066);
nor_5  g02718(n15743, n2809, new_n5067);
nand_5 g02719(n20658, n15508, new_n5068);
not_8  g02720(new_n5068, new_n5069);
xnor_4 g02721(n15743, n2809, new_n5070);
nor_5  g02722(new_n5070, new_n5069, new_n5071);
nor_5  g02723(new_n5071, new_n5067, new_n5072);
nor_5  g02724(new_n5072, new_n5066, new_n5073);
nor_5  g02725(new_n5073, new_n5064_1, new_n5074);
nor_5  g02726(new_n5074, new_n5063, new_n5075);
nor_5  g02727(new_n5075, new_n5061, new_n5076);
not_8  g02728(new_n5076, new_n5077_1);
nand_5 g02729(new_n5077_1, new_n5060_1, new_n5078);
nand_5 g02730(new_n5078, new_n5059, new_n5079);
nand_5 g02731(new_n5079, new_n5057, new_n5080);
nand_5 g02732(new_n5080, new_n5056, new_n5081);
nand_5 g02733(new_n5081, new_n5054, new_n5082_1);
nand_5 g02734(new_n5082_1, new_n5052, new_n5083);
nand_5 g02735(new_n5083, new_n5050, new_n5084);
nand_5 g02736(new_n5084, new_n5048, new_n5085);
nand_5 g02737(new_n5085, new_n5047, new_n5086);
nand_5 g02738(new_n5086, new_n5045, new_n5087);
xnor_4 g02739(new_n5087, new_n5044, new_n5088);
not_8  g02740(new_n5088, new_n5089);
nand_5 g02741(new_n5089, n9259, new_n5090);
xnor_4 g02742(new_n5088, n9259, new_n5091);
not_8  g02743(new_n5047, new_n5092);
xnor_4 g02744(new_n5085, new_n5092, new_n5093);
not_8  g02745(new_n5093, new_n5094);
nand_5 g02746(new_n5094, n21489, new_n5095);
xnor_4 g02747(new_n5093, n21489, new_n5096);
xnor_4 g02748(new_n5083, new_n5050, new_n5097);
nand_5 g02749(new_n5097, n20213, new_n5098_1);
xnor_4 g02750(new_n5097, new_n3746, new_n5099);
not_8  g02751(new_n5054, new_n5100);
xnor_4 g02752(new_n5081, new_n5100, new_n5101_1);
not_8  g02753(new_n5101_1, new_n5102);
nand_5 g02754(new_n5102, n13912, new_n5103);
xnor_4 g02755(new_n5101_1, n13912, new_n5104);
not_8  g02756(new_n5057, new_n5105);
xnor_4 g02757(new_n5079, new_n5105, new_n5106);
not_8  g02758(new_n5106, new_n5107);
nand_5 g02759(new_n5107, n7670, new_n5108);
xnor_4 g02760(new_n5106, n7670, new_n5109);
not_8  g02761(new_n5060_1, new_n5110);
xnor_4 g02762(new_n5076, new_n5110, new_n5111);
nand_5 g02763(new_n5111, n9598, new_n5112);
xnor_4 g02764(new_n5111, new_n3726, new_n5113);
xnor_4 g02765(new_n5074, new_n5062_1, new_n5114);
nor_5  g02766(new_n5114, new_n3768, new_n5115_1);
not_8  g02767(new_n5115_1, new_n5116);
xnor_4 g02768(new_n5114, n22290, new_n5117);
xnor_4 g02769(new_n5072, new_n5065, new_n5118);
nor_5  g02770(new_n5118, new_n3727, new_n5119);
not_8  g02771(new_n5119, new_n5120_1);
not_8  g02772(n25565, new_n5121);
xnor_4 g02773(new_n5070, new_n5068, new_n5122);
nand_5 g02774(new_n5122, new_n5121, new_n5123);
not_8  g02775(new_n5123, new_n5124);
not_8  g02776(n15508, new_n5125);
xnor_4 g02777(n20658, new_n5125, new_n5126);
nand_5 g02778(new_n5126, n21993, new_n5127);
not_8  g02779(new_n5127, new_n5128_1);
xnor_4 g02780(new_n5122, new_n5121, new_n5129);
nor_5  g02781(new_n5129, new_n5128_1, new_n5130);
nor_5  g02782(new_n5130, new_n5124, new_n5131_1);
xnor_4 g02783(new_n5118, n11273, new_n5132);
nand_5 g02784(new_n5132, new_n5131_1, new_n5133);
nand_5 g02785(new_n5133, new_n5120_1, new_n5134);
nand_5 g02786(new_n5134, new_n5117, new_n5135);
nand_5 g02787(new_n5135, new_n5116, new_n5136);
nand_5 g02788(new_n5136, new_n5113, new_n5137);
nand_5 g02789(new_n5137, new_n5112, new_n5138);
nand_5 g02790(new_n5138, new_n5109, new_n5139);
nand_5 g02791(new_n5139, new_n5108, new_n5140_1);
nand_5 g02792(new_n5140_1, new_n5104, new_n5141);
nand_5 g02793(new_n5141, new_n5103, new_n5142);
nand_5 g02794(new_n5142, new_n5099, new_n5143);
nand_5 g02795(new_n5143, new_n5098_1, new_n5144);
nand_5 g02796(new_n5144, new_n5096, new_n5145);
nand_5 g02797(new_n5145, new_n5095, new_n5146);
nand_5 g02798(new_n5146, new_n5091, new_n5147);
nand_5 g02799(new_n5147, new_n5090, new_n5148);
or_5   g02800(n9554, n2979, new_n5149);
nand_5 g02801(new_n5087, new_n5043, new_n5150);
nand_5 g02802(new_n5150, new_n5149, new_n5151);
xnor_4 g02803(new_n5151, new_n5148, new_n5152);
xnor_4 g02804(new_n5146, new_n5091, new_n5153);
nor_5  g02805(new_n5153, n3740, new_n5154);
xnor_4 g02806(new_n5153, n3740, new_n5155);
xnor_4 g02807(new_n5144, new_n5096, new_n5156);
nand_5 g02808(new_n5156, n2858, new_n5157);
not_8  g02809(n2858, new_n5158_1);
xnor_4 g02810(new_n5156, new_n5158_1, new_n5159);
xnor_4 g02811(new_n5142, new_n5099, new_n5160);
nand_5 g02812(new_n5160, n2659, new_n5161);
not_8  g02813(n2659, new_n5162);
xnor_4 g02814(new_n5160, new_n5162, new_n5163);
xnor_4 g02815(new_n5140_1, new_n5104, new_n5164);
nand_5 g02816(new_n5164, n24327, new_n5165);
not_8  g02817(n24327, new_n5166);
xnor_4 g02818(new_n5164, new_n5166, new_n5167);
xnor_4 g02819(new_n5138, new_n5109, new_n5168_1);
nand_5 g02820(new_n5168_1, n22198, new_n5169);
not_8  g02821(n22198, new_n5170);
xnor_4 g02822(new_n5168_1, new_n5170, new_n5171);
xnor_4 g02823(new_n5136, new_n5113, new_n5172);
nand_5 g02824(new_n5172, n20826, new_n5173);
not_8  g02825(n20826, new_n5174);
xnor_4 g02826(new_n5172, new_n5174, new_n5175);
not_8  g02827(n7305, new_n5176);
xnor_4 g02828(new_n5134, new_n5117, new_n5177);
not_8  g02829(new_n5177, new_n5178);
nor_5  g02830(new_n5178, new_n5176, new_n5179);
not_8  g02831(new_n5179, new_n5180);
not_8  g02832(n25872, new_n5181);
not_8  g02833(new_n5132, new_n5182);
xnor_4 g02834(new_n5182, new_n5131_1, new_n5183);
nand_5 g02835(new_n5183, new_n5181, new_n5184_1);
not_8  g02836(new_n5184_1, new_n5185);
xnor_4 g02837(new_n5183, new_n5181, new_n5186);
not_8  g02838(n20259, new_n5187);
xnor_4 g02839(new_n5129, new_n5128_1, new_n5188);
nor_5  g02840(new_n5188, new_n5187, new_n5189);
not_8  g02841(new_n5189, new_n5190);
xnor_4 g02842(new_n5126, new_n3779, new_n5191);
not_8  g02843(new_n5191, new_n5192);
nor_5  g02844(new_n5192, n3925, new_n5193);
not_8  g02845(new_n5193, new_n5194);
xnor_4 g02846(new_n5188, n20259, new_n5195);
nand_5 g02847(new_n5195, new_n5194, new_n5196);
nand_5 g02848(new_n5196, new_n5190, new_n5197);
nor_5  g02849(new_n5197, new_n5186, new_n5198);
nor_5  g02850(new_n5198, new_n5185, new_n5199);
xnor_4 g02851(new_n5177, new_n5176, new_n5200);
nand_5 g02852(new_n5200, new_n5199, new_n5201);
nand_5 g02853(new_n5201, new_n5180, new_n5202);
nand_5 g02854(new_n5202, new_n5175, new_n5203);
nand_5 g02855(new_n5203, new_n5173, new_n5204);
nand_5 g02856(new_n5204, new_n5171, new_n5205);
nand_5 g02857(new_n5205, new_n5169, new_n5206);
nand_5 g02858(new_n5206, new_n5167, new_n5207);
nand_5 g02859(new_n5207, new_n5165, new_n5208);
nand_5 g02860(new_n5208, new_n5163, new_n5209);
nand_5 g02861(new_n5209, new_n5161, new_n5210);
nand_5 g02862(new_n5210, new_n5159, new_n5211_1);
nand_5 g02863(new_n5211_1, new_n5157, new_n5212);
nor_5  g02864(new_n5212, new_n5155, new_n5213_1);
nor_5  g02865(new_n5213_1, new_n5154, new_n5214);
xnor_4 g02866(new_n5214, new_n5152, new_n5215);
xnor_4 g02867(new_n5215, new_n5041, new_n5216);
not_8  g02868(new_n5216, new_n5217);
xnor_4 g02869(new_n5038, new_n4993, new_n5218);
not_8  g02870(new_n5218, new_n5219);
not_8  g02871(n3740, new_n5220);
xnor_4 g02872(new_n5153, new_n5220, new_n5221);
xnor_4 g02873(new_n5212, new_n5221, new_n5222);
nand_5 g02874(new_n5222, new_n5219, new_n5223);
xnor_4 g02875(new_n5222, new_n5218, new_n5224);
xnor_4 g02876(new_n5036, new_n4996, new_n5225);
not_8  g02877(new_n5225, new_n5226_1);
xnor_4 g02878(new_n5210, new_n5159, new_n5227);
nand_5 g02879(new_n5227, new_n5226_1, new_n5228_1);
xnor_4 g02880(new_n5227, new_n5225, new_n5229);
xnor_4 g02881(new_n5033, new_n4999, new_n5230);
xnor_4 g02882(new_n5208, new_n5163, new_n5231);
nand_5 g02883(new_n5231, new_n5230, new_n5232);
not_8  g02884(new_n5230, new_n5233);
xnor_4 g02885(new_n5231, new_n5233, new_n5234);
xnor_4 g02886(new_n5031_1, new_n5001, new_n5235);
xnor_4 g02887(new_n5164, n24327, new_n5236);
xnor_4 g02888(new_n5206, new_n5236, new_n5237);
not_8  g02889(new_n5237, new_n5238);
nand_5 g02890(new_n5238, new_n5235, new_n5239);
xnor_4 g02891(new_n5237, new_n5235, new_n5240);
xnor_4 g02892(new_n5029, new_n5005, new_n5241);
xnor_4 g02893(new_n5168_1, n22198, new_n5242);
xnor_4 g02894(new_n5204, new_n5242, new_n5243);
not_8  g02895(new_n5243, new_n5244);
nand_5 g02896(new_n5244, new_n5241, new_n5245);
xnor_4 g02897(new_n5243, new_n5241, new_n5246);
xnor_4 g02898(new_n5027, new_n5009, new_n5247);
xnor_4 g02899(new_n5202, new_n5175, new_n5248);
nand_5 g02900(new_n5248, new_n5247, new_n5249);
not_8  g02901(new_n5247, new_n5250);
xnor_4 g02902(new_n5248, new_n5250, new_n5251);
xnor_4 g02903(new_n5025_1, new_n5012, new_n5252);
not_8  g02904(new_n5252, new_n5253);
not_8  g02905(new_n5200, new_n5254);
xnor_4 g02906(new_n5254, new_n5199, new_n5255_1);
nor_5  g02907(new_n5255_1, new_n5253, new_n5256_1);
not_8  g02908(new_n5256_1, new_n5257);
xnor_4 g02909(new_n5255_1, new_n5252, new_n5258);
not_8  g02910(new_n5186, new_n5259);
xnor_4 g02911(new_n5197, new_n5259, new_n5260);
xnor_4 g02912(new_n5023, new_n5015, new_n5261);
nand_5 g02913(new_n5261, new_n5260, new_n5262);
not_8  g02914(new_n5261, new_n5263);
xnor_4 g02915(new_n5263, new_n5260, new_n5264);
xnor_4 g02916(new_n5191, n3925, new_n5265_1);
xnor_4 g02917(n9246, new_n3946, new_n5266);
not_8  g02918(new_n5266, new_n5267);
nor_5  g02919(new_n5267, new_n5265_1, new_n5268);
not_8  g02920(new_n5268, new_n5269);
nor_5  g02921(new_n5269, new_n5021, new_n5270);
xnor_4 g02922(new_n5195, new_n5194, new_n5271);
xnor_4 g02923(new_n5020_1, new_n5019, new_n5272);
not_8  g02924(new_n5272, new_n5273_1);
nor_5  g02925(new_n5273_1, new_n5268, new_n5274_1);
nor_5  g02926(new_n5274_1, new_n5270, new_n5275);
not_8  g02927(new_n5275, new_n5276);
nor_5  g02928(new_n5276, new_n5271, new_n5277);
nor_5  g02929(new_n5277, new_n5270, new_n5278);
nand_5 g02930(new_n5278, new_n5264, new_n5279);
nand_5 g02931(new_n5279, new_n5262, new_n5280);
nand_5 g02932(new_n5280, new_n5258, new_n5281);
nand_5 g02933(new_n5281, new_n5257, new_n5282);
nand_5 g02934(new_n5282, new_n5251, new_n5283);
nand_5 g02935(new_n5283, new_n5249, new_n5284);
nand_5 g02936(new_n5284, new_n5246, new_n5285);
nand_5 g02937(new_n5285, new_n5245, new_n5286);
nand_5 g02938(new_n5286, new_n5240, new_n5287);
nand_5 g02939(new_n5287, new_n5239, new_n5288);
nand_5 g02940(new_n5288, new_n5234, new_n5289);
nand_5 g02941(new_n5289, new_n5232, new_n5290);
nand_5 g02942(new_n5290, new_n5229, new_n5291);
nand_5 g02943(new_n5291, new_n5228_1, new_n5292);
nand_5 g02944(new_n5292, new_n5224, new_n5293);
nand_5 g02945(new_n5293, new_n5223, new_n5294);
xnor_4 g02946(new_n5294, new_n5217, n332);
not_8  g02947(n8381, new_n5296);
xnor_4 g02948(n18295, n16223, new_n5297);
not_8  g02949(new_n5297, new_n5298);
nor_5  g02950(n19494, n6502, new_n5299);
nand_5 g02951(n15780, n2387, new_n5300_1);
not_8  g02952(new_n5300_1, new_n5301);
xnor_4 g02953(n19494, n6502, new_n5302_1);
nor_5  g02954(new_n5302_1, new_n5301, new_n5303);
nor_5  g02955(new_n5303, new_n5299, new_n5304);
xnor_4 g02956(new_n5304, new_n5298, new_n5305);
xnor_4 g02957(new_n5305, new_n5296, new_n5306);
not_8  g02958(n20235, new_n5307);
xnor_4 g02959(n15780, new_n2368, new_n5308);
not_8  g02960(new_n5308, new_n5309);
nor_5  g02961(new_n5309, n12495, new_n5310);
nand_5 g02962(new_n5310, new_n5307, new_n5311);
not_8  g02963(new_n5311, new_n5312);
xnor_4 g02964(new_n5310, new_n5307, new_n5313);
xnor_4 g02965(new_n5302_1, new_n5300_1, new_n5314);
nor_5  g02966(new_n5314, new_n5313, new_n5315);
nor_5  g02967(new_n5315, new_n5312, new_n5316);
xnor_4 g02968(new_n5316, new_n5306, new_n5317);
not_8  g02969(n23146, new_n5318);
nor_5  g02970(n21654, new_n3486, new_n5319);
xnor_4 g02971(n25471, n23842, new_n5320);
xnor_4 g02972(new_n5320, new_n5319, new_n5321);
not_8  g02973(new_n5321, new_n5322);
nor_5  g02974(new_n5322, new_n5318, new_n5323);
not_8  g02975(new_n5323, new_n5324);
not_8  g02976(n17968, new_n5325_1);
xnor_4 g02977(n21654, n16502, new_n5326);
nor_5  g02978(new_n5326, new_n5325_1, new_n5327);
xnor_4 g02979(new_n5321, new_n5318, new_n5328);
nand_5 g02980(new_n5328, new_n5327, new_n5329);
nand_5 g02981(new_n5329, new_n5324, new_n5330_1);
xnor_4 g02982(n15053, n3828, new_n5331);
not_8  g02983(n23842, new_n5332);
nand_5 g02984(n25471, new_n5332, new_n5333);
nand_5 g02985(new_n5320, new_n5319, new_n5334);
nand_5 g02986(new_n5334, new_n5333, new_n5335);
xnor_4 g02987(new_n5335, new_n5331, new_n5336);
xnor_4 g02988(new_n5336, n11184, new_n5337_1);
xnor_4 g02989(new_n5337_1, new_n5330_1, new_n5338);
xnor_4 g02990(new_n5338, new_n5317, new_n5339);
xnor_4 g02991(new_n5321, n23146, new_n5340);
xnor_4 g02992(new_n5340, new_n5327, new_n5341);
not_8  g02993(new_n5314, new_n5342);
xnor_4 g02994(new_n5342, new_n5313, new_n5343);
not_8  g02995(new_n5343, new_n5344);
nor_5  g02996(new_n5344, new_n5341, new_n5345);
not_8  g02997(new_n5345, new_n5346);
xnor_4 g02998(new_n5308, n12495, new_n5347);
xnor_4 g02999(new_n5326, n17968, new_n5348);
not_8  g03000(new_n5348, new_n5349);
nor_5  g03001(new_n5349, new_n5347, new_n5350);
not_8  g03002(new_n5350, new_n5351_1);
xnor_4 g03003(new_n5343, new_n5341, new_n5352);
nand_5 g03004(new_n5352, new_n5351_1, new_n5353_1);
nand_5 g03005(new_n5353_1, new_n5346, new_n5354);
xnor_4 g03006(new_n5354, new_n5339, n357);
xnor_4 g03007(n22309, new_n3650, new_n5356);
nand_5 g03008(n22309, n9251, new_n5357);
not_8  g03009(new_n5357, new_n5358);
xnor_4 g03010(n25073, n20138, new_n5359);
xnor_4 g03011(new_n5359, new_n5358, new_n5360);
nor_5  g03012(new_n5360, new_n5356, new_n5361);
not_8  g03013(new_n5361, new_n5362);
xnor_4 g03014(n18171, new_n2360, new_n5363);
nor_5  g03015(n25073, n20138, new_n5364);
nor_5  g03016(new_n5359, new_n5358, new_n5365);
nor_5  g03017(new_n5365, new_n5364, new_n5366);
xnor_4 g03018(new_n5366, new_n5363, new_n5367);
not_8  g03019(new_n5367, new_n5368);
nor_5  g03020(new_n5368, new_n5362, new_n5369);
xnor_4 g03021(n5752, new_n3576, new_n5370);
nor_5  g03022(n18171, n6385, new_n5371);
not_8  g03023(new_n5363, new_n5372);
nor_5  g03024(new_n5366, new_n5372, new_n5373);
nor_5  g03025(new_n5373, new_n5371, new_n5374);
xnor_4 g03026(new_n5374, new_n5370, new_n5375);
nand_5 g03027(new_n5375, new_n5369, new_n5376_1);
xnor_4 g03028(n16158, new_n3536, new_n5377);
not_8  g03029(new_n5377, new_n5378);
nor_5  g03030(n5752, n3136, new_n5379);
not_8  g03031(new_n5370, new_n5380);
nor_5  g03032(new_n5374, new_n5380, new_n5381);
nor_5  g03033(new_n5381, new_n5379, new_n5382);
xnor_4 g03034(new_n5382, new_n5378, new_n5383);
nor_5  g03035(new_n5383, new_n5376_1, new_n5384);
not_8  g03036(n20604, new_n5385);
xnor_4 g03037(n25643, new_n5385, new_n5386_1);
nor_5  g03038(n16158, n9557, new_n5387);
nor_5  g03039(new_n5382, new_n5378, new_n5388);
nor_5  g03040(new_n5388, new_n5387, new_n5389);
xnor_4 g03041(new_n5389, new_n5386_1, new_n5390);
xnor_4 g03042(new_n5390, new_n5384, new_n5391);
xnor_4 g03043(new_n5391, new_n3238, new_n5392);
not_8  g03044(new_n5392, new_n5393);
not_8  g03045(new_n3250, new_n5394);
not_8  g03046(new_n5383, new_n5395);
xnor_4 g03047(new_n5395, new_n5376_1, new_n5396);
not_8  g03048(new_n5396, new_n5397);
nand_5 g03049(new_n5397, new_n5394, new_n5398);
xnor_4 g03050(new_n5396, new_n5394, new_n5399_1);
xnor_4 g03051(new_n5375, new_n5369, new_n5400_1);
nand_5 g03052(new_n5400_1, new_n3254, new_n5401);
xnor_4 g03053(new_n5400_1, new_n3255, new_n5402);
xnor_4 g03054(new_n5367, new_n5361, new_n5403_1);
nor_5  g03055(new_n5403_1, new_n3259, new_n5404);
not_8  g03056(new_n5356, new_n5405);
nor_5  g03057(new_n5405, new_n3264, new_n5406);
nor_5  g03058(new_n5406, new_n3269, new_n5407);
nor_5  g03059(n22309, n9251, new_n5408);
not_8  g03060(new_n5365, new_n5409);
nor_5  g03061(new_n5409, new_n5408, new_n5410);
nor_5  g03062(new_n5410, new_n5361, new_n5411);
not_8  g03063(new_n5406, new_n5412);
nor_5  g03064(new_n5412, new_n3197, new_n5413);
nor_5  g03065(new_n5413, new_n5407, new_n5414);
not_8  g03066(new_n5414, new_n5415);
nor_5  g03067(new_n5415, new_n5411, new_n5416);
nor_5  g03068(new_n5416, new_n5407, new_n5417);
not_8  g03069(new_n5417, new_n5418);
xnor_4 g03070(new_n5403_1, new_n3259, new_n5419);
nor_5  g03071(new_n5419, new_n5418, new_n5420);
nor_5  g03072(new_n5420, new_n5404, new_n5421);
nand_5 g03073(new_n5421, new_n5402, new_n5422);
nand_5 g03074(new_n5422, new_n5401, new_n5423);
nand_5 g03075(new_n5423, new_n5399_1, new_n5424);
nand_5 g03076(new_n5424, new_n5398, new_n5425);
xnor_4 g03077(new_n5425, new_n5393, new_n5426);
xnor_4 g03078(n5255, n4119, new_n5427);
not_8  g03079(n21649, new_n5428);
nor_5  g03080(new_n5428, n14510, new_n5429);
not_8  g03081(new_n5429, new_n5430_1);
xnor_4 g03082(n21649, n14510, new_n5431);
not_8  g03083(n18274, new_n5432);
nor_5  g03084(new_n5432, n13263, new_n5433);
xnor_4 g03085(n18274, n13263, new_n5434);
nor_5  g03086(new_n3580, n3828, new_n5435);
not_8  g03087(n3828, new_n5436);
nor_5  g03088(n20455, new_n5436, new_n5437);
nor_5  g03089(n23842, new_n3585, new_n5438_1);
nor_5  g03090(new_n5332, n1639, new_n5439_1);
nor_5  g03091(n21654, new_n4863, new_n5440);
not_8  g03092(new_n5440, new_n5441);
nor_5  g03093(new_n5441, new_n5439_1, new_n5442);
nor_5  g03094(new_n5442, new_n5438_1, new_n5443_1);
nor_5  g03095(new_n5443_1, new_n5437, new_n5444);
nor_5  g03096(new_n5444, new_n5435, new_n5445);
and_5  g03097(new_n5445, new_n5434, new_n5446);
nor_5  g03098(new_n5446, new_n5433, new_n5447);
not_8  g03099(new_n5447, new_n5448);
nand_5 g03100(new_n5448, new_n5431, new_n5449);
nand_5 g03101(new_n5449, new_n5430_1, new_n5450);
xnor_4 g03102(new_n5450, new_n5427, new_n5451_1);
xnor_4 g03103(new_n5451_1, new_n5426, new_n5452);
xnor_4 g03104(new_n5447, new_n5431, new_n5453);
xnor_4 g03105(new_n5423, new_n5399_1, new_n5454);
nor_5  g03106(new_n5454, new_n5453, new_n5455);
xnor_4 g03107(new_n5454, new_n5453, new_n5456);
xnor_4 g03108(new_n5421, new_n5402, new_n5457);
xnor_4 g03109(new_n5445, new_n5434, new_n5458);
not_8  g03110(new_n5458, new_n5459);
nor_5  g03111(new_n5459, new_n5457, new_n5460);
xnor_4 g03112(new_n5459, new_n5457, new_n5461);
xnor_4 g03113(new_n5419, new_n5418, new_n5462);
xnor_4 g03114(n20455, n3828, new_n5463);
xnor_4 g03115(new_n5463, new_n5443_1, new_n5464);
nand_5 g03116(new_n5464, new_n5462, new_n5465);
not_8  g03117(new_n5465, new_n5466);
xnor_4 g03118(new_n5464, new_n5462, new_n5467);
xnor_4 g03119(n21654, n16968, new_n5468);
xnor_4 g03120(new_n5405, new_n3264, new_n5469);
nor_5  g03121(new_n5469, new_n5468, new_n5470);
xnor_4 g03122(n23842, new_n3585, new_n5471);
xnor_4 g03123(new_n5471, new_n5440, new_n5472_1);
not_8  g03124(new_n5472_1, new_n5473);
nor_5  g03125(new_n5473, new_n5470, new_n5474);
xnor_4 g03126(new_n5414, new_n5411, new_n5475);
xnor_4 g03127(new_n5472_1, new_n5470, new_n5476);
nand_5 g03128(new_n5476, new_n5475, new_n5477);
not_8  g03129(new_n5477, new_n5478);
nor_5  g03130(new_n5478, new_n5474, new_n5479);
nor_5  g03131(new_n5479, new_n5467, new_n5480);
nor_5  g03132(new_n5480, new_n5466, new_n5481);
nor_5  g03133(new_n5481, new_n5461, new_n5482);
nor_5  g03134(new_n5482, new_n5460, new_n5483);
nor_5  g03135(new_n5483, new_n5456, new_n5484);
nor_5  g03136(new_n5484, new_n5455, new_n5485_1);
xnor_4 g03137(new_n5485_1, new_n5452, n422);
not_8  g03138(n21471, new_n5487);
nor_5  g03139(n23333, n20794, new_n5488);
nand_5 g03140(new_n5488, new_n3409, new_n5489);
nor_5  g03141(new_n5489, n18737, new_n5490);
nand_5 g03142(new_n5490, new_n5487, new_n5491);
nor_5  g03143(new_n5491, n25738, new_n5492);
nand_5 g03144(new_n5492, new_n3393, new_n5493);
nor_5  g03145(new_n5493, n3228, new_n5494);
xnor_4 g03146(new_n5494, n337, new_n5495);
xnor_4 g03147(new_n5495, new_n3219_1, new_n5496);
not_8  g03148(new_n5496, new_n5497);
xnor_4 g03149(new_n5493, new_n3390_1, new_n5498);
or_5   g03150(new_n5498, n26036, new_n5499);
xnor_4 g03151(new_n5498, new_n3225, new_n5500);
xnor_4 g03152(new_n5492, n5302, new_n5501);
or_5   g03153(new_n5501, n19770, new_n5502);
xnor_4 g03154(new_n5501, new_n3231, new_n5503);
not_8  g03155(n25738, new_n5504);
xnor_4 g03156(new_n5491, new_n5504, new_n5505);
or_5   g03157(new_n5505, n8782, new_n5506);
xnor_4 g03158(new_n5505, new_n3237, new_n5507);
xnor_4 g03159(new_n5490, n21471, new_n5508);
not_8  g03160(new_n5508, new_n5509);
nand_5 g03161(new_n5509, new_n3241, new_n5510);
xnor_4 g03162(new_n5508, new_n3241, new_n5511);
not_8  g03163(n18737, new_n5512);
xnor_4 g03164(new_n5489, new_n5512, new_n5513);
not_8  g03165(new_n5513, new_n5514);
nand_5 g03166(new_n5514, new_n3253_1, new_n5515);
xnor_4 g03167(new_n5488, n14603, new_n5516);
not_8  g03168(new_n5516, new_n5517_1);
nand_5 g03169(new_n5517_1, new_n3258, new_n5518);
xnor_4 g03170(new_n5516, new_n3258, new_n5519);
xnor_4 g03171(n23333, n20794, new_n5520);
nand_5 g03172(new_n5520, new_n3263_1, new_n5521_1);
nand_5 g03173(n23333, n11424, new_n5522);
not_8  g03174(new_n5522, new_n5523);
xnor_4 g03175(new_n5520, n25336, new_n5524_1);
not_8  g03176(new_n5524_1, new_n5525);
nor_5  g03177(new_n5525, new_n5523, new_n5526);
not_8  g03178(new_n5526, new_n5527);
nand_5 g03179(new_n5527, new_n5521_1, new_n5528);
nand_5 g03180(new_n5528, new_n5519, new_n5529);
nand_5 g03181(new_n5529, new_n5518, new_n5530);
xnor_4 g03182(new_n5513, new_n3253_1, new_n5531);
nand_5 g03183(new_n5531, new_n5530, new_n5532_1);
nand_5 g03184(new_n5532_1, new_n5515, new_n5533);
nand_5 g03185(new_n5533, new_n5511, new_n5534);
nand_5 g03186(new_n5534, new_n5510, new_n5535);
nand_5 g03187(new_n5535, new_n5507, new_n5536);
nand_5 g03188(new_n5536, new_n5506, new_n5537);
nand_5 g03189(new_n5537, new_n5503, new_n5538);
nand_5 g03190(new_n5538, new_n5502, new_n5539);
nand_5 g03191(new_n5539, new_n5500, new_n5540);
nand_5 g03192(new_n5540, new_n5499, new_n5541);
xnor_4 g03193(new_n5541, new_n5497, new_n5542);
xnor_4 g03194(n22379, new_n3295, new_n5543);
or_5   g03195(n20946, n1662, new_n5544);
xnor_4 g03196(n20946, new_n2900, new_n5545);
nor_5  g03197(n12875, n7751, new_n5546);
xnor_4 g03198(n12875, new_n2430, new_n5547);
not_8  g03199(new_n5547, new_n5548);
nor_5  g03200(n26823, n2035, new_n5549);
xnor_4 g03201(n26823, new_n2906, new_n5550);
not_8  g03202(new_n5550, new_n5551);
nor_5  g03203(n5213, n4812, new_n5552);
xnor_4 g03204(n5213, new_n2438, new_n5553);
not_8  g03205(new_n5553, new_n5554);
nor_5  g03206(n24278, n4665, new_n5555);
xnor_4 g03207(n24278, new_n2912, new_n5556);
not_8  g03208(new_n5556, new_n5557);
nor_5  g03209(n24618, n19005, new_n5558);
xnor_4 g03210(n24618, new_n2917, new_n5559);
not_8  g03211(new_n5559, new_n5560);
nor_5  g03212(n4326, n3952, new_n5561);
nand_5 g03213(n12315, n5438, new_n5562);
not_8  g03214(new_n5562, new_n5563);
xnor_4 g03215(n4326, n3952, new_n5564_1);
nor_5  g03216(new_n5564_1, new_n5563, new_n5565);
nor_5  g03217(new_n5565, new_n5561, new_n5566);
nor_5  g03218(new_n5566, new_n5560, new_n5567);
nor_5  g03219(new_n5567, new_n5558, new_n5568);
nor_5  g03220(new_n5568, new_n5557, new_n5569);
nor_5  g03221(new_n5569, new_n5555, new_n5570);
nor_5  g03222(new_n5570, new_n5554, new_n5571);
nor_5  g03223(new_n5571, new_n5552, new_n5572);
nor_5  g03224(new_n5572, new_n5551, new_n5573);
nor_5  g03225(new_n5573, new_n5549, new_n5574);
nor_5  g03226(new_n5574, new_n5548, new_n5575);
nor_5  g03227(new_n5575, new_n5546, new_n5576);
not_8  g03228(new_n5576, new_n5577);
nand_5 g03229(new_n5577, new_n5545, new_n5578);
nand_5 g03230(new_n5578, new_n5544, new_n5579_1);
xnor_4 g03231(new_n5579_1, new_n5543, new_n5580);
xnor_4 g03232(n10763, new_n3168, new_n5581);
or_5   g03233(n13367, n7437, new_n5582);
xnor_4 g03234(n13367, new_n2944_1, new_n5583);
nor_5  g03235(n20700, n932, new_n5584);
xnor_4 g03236(n20700, new_n3175, new_n5585);
not_8  g03237(new_n5585, new_n5586);
nor_5  g03238(n7099, n6691, new_n5587);
xnor_4 g03239(n7099, new_n3179, new_n5588);
not_8  g03240(new_n5588, new_n5589);
nor_5  g03241(n12811, n3260, new_n5590);
xnor_4 g03242(n12811, new_n3183, new_n5591);
not_8  g03243(new_n5591, new_n5592);
nor_5  g03244(n20489, n1118, new_n5593_1);
xnor_4 g03245(n20489, new_n2959, new_n5594);
not_8  g03246(new_n5594, new_n5595);
nor_5  g03247(n25974, n2355, new_n5596);
xnor_4 g03248(n25974, n2355, new_n5597);
nor_5  g03249(n11121, n1630, new_n5598);
nand_5 g03250(n16217, n1451, new_n5599);
not_8  g03251(new_n5599, new_n5600);
xnor_4 g03252(n11121, n1630, new_n5601);
nor_5  g03253(new_n5601, new_n5600, new_n5602);
nor_5  g03254(new_n5602, new_n5598, new_n5603_1);
nor_5  g03255(new_n5603_1, new_n5597, new_n5604);
nor_5  g03256(new_n5604, new_n5596, new_n5605_1);
nor_5  g03257(new_n5605_1, new_n5595, new_n5606);
nor_5  g03258(new_n5606, new_n5593_1, new_n5607);
nor_5  g03259(new_n5607, new_n5592, new_n5608);
nor_5  g03260(new_n5608, new_n5590, new_n5609_1);
nor_5  g03261(new_n5609_1, new_n5589, new_n5610);
nor_5  g03262(new_n5610, new_n5587, new_n5611);
nor_5  g03263(new_n5611, new_n5586, new_n5612);
nor_5  g03264(new_n5612, new_n5584, new_n5613);
not_8  g03265(new_n5613, new_n5614);
nand_5 g03266(new_n5614, new_n5583, new_n5615);
nand_5 g03267(new_n5615, new_n5582, new_n5616);
xnor_4 g03268(new_n5616, new_n5581, new_n5617);
xnor_4 g03269(new_n5617, new_n5580, new_n5618);
xnor_4 g03270(new_n5613, new_n5583, new_n5619);
xnor_4 g03271(new_n5576, new_n5545, new_n5620);
not_8  g03272(new_n5620, new_n5621);
nor_5  g03273(new_n5621, new_n5619, new_n5622);
not_8  g03274(new_n5622, new_n5623);
xnor_4 g03275(new_n5620, new_n5619, new_n5624);
xnor_4 g03276(new_n5611, new_n5585, new_n5625);
not_8  g03277(new_n5625, new_n5626);
xnor_4 g03278(new_n5574, new_n5547, new_n5627);
nor_5  g03279(new_n5627, new_n5626, new_n5628);
xnor_4 g03280(new_n5627, new_n5625, new_n5629);
not_8  g03281(new_n5629, new_n5630);
xnor_4 g03282(new_n5609_1, new_n5588, new_n5631);
not_8  g03283(new_n5631, new_n5632);
xnor_4 g03284(new_n5572, new_n5550, new_n5633);
nor_5  g03285(new_n5633, new_n5632, new_n5634_1);
xnor_4 g03286(new_n5605_1, new_n5595, new_n5635);
xnor_4 g03287(new_n5568, new_n5556, new_n5636);
nor_5  g03288(new_n5636, new_n5635, new_n5637);
xnor_4 g03289(new_n5636, new_n5635, new_n5638);
xnor_4 g03290(new_n5603_1, new_n5597, new_n5639);
xnor_4 g03291(new_n5566, new_n5559, new_n5640);
nor_5  g03292(new_n5640, new_n5639, new_n5641);
xnor_4 g03293(new_n5564_1, new_n5562, new_n5642);
xnor_4 g03294(new_n5601, new_n5600, new_n5643_1);
nor_5  g03295(new_n5643_1, new_n5642, new_n5644);
xnor_4 g03296(n12315, n5438, new_n5645);
not_8  g03297(new_n5645, new_n5646);
xnor_4 g03298(n16217, n1451, new_n5647);
nand_5 g03299(new_n5647, new_n5646, new_n5648);
xnor_4 g03300(new_n5643_1, new_n5642, new_n5649);
nor_5  g03301(new_n5649, new_n5648, new_n5650);
nor_5  g03302(new_n5650, new_n5644, new_n5651);
xnor_4 g03303(new_n5640, new_n5639, new_n5652);
nor_5  g03304(new_n5652, new_n5651, new_n5653);
nor_5  g03305(new_n5653, new_n5641, new_n5654);
nor_5  g03306(new_n5654, new_n5638, new_n5655);
nor_5  g03307(new_n5655, new_n5637, new_n5656);
xnor_4 g03308(new_n5607, new_n5592, new_n5657);
nand_5 g03309(new_n5657, new_n5656, new_n5658);
xnor_4 g03310(new_n5657, new_n5656, new_n5659);
not_8  g03311(new_n5659, new_n5660);
xnor_4 g03312(new_n5570, new_n5553, new_n5661);
nand_5 g03313(new_n5661, new_n5660, new_n5662);
nand_5 g03314(new_n5662, new_n5658, new_n5663);
xnor_4 g03315(new_n5633, new_n5631, new_n5664);
not_8  g03316(new_n5664, new_n5665);
nor_5  g03317(new_n5665, new_n5663, new_n5666);
nor_5  g03318(new_n5666, new_n5634_1, new_n5667);
nor_5  g03319(new_n5667, new_n5630, new_n5668);
nor_5  g03320(new_n5668, new_n5628, new_n5669);
nand_5 g03321(new_n5669, new_n5624, new_n5670);
nand_5 g03322(new_n5670, new_n5623, new_n5671);
nand_5 g03323(new_n5671, new_n5618, new_n5672);
not_8  g03324(new_n5672, new_n5673);
nor_5  g03325(new_n5671, new_n5618, new_n5674);
nor_5  g03326(new_n5674, new_n5673, new_n5675);
xnor_4 g03327(new_n5675, new_n5542, new_n5676);
xnor_4 g03328(new_n5539, new_n5500, new_n5677);
xnor_4 g03329(new_n5669, new_n5624, new_n5678);
not_8  g03330(new_n5678, new_n5679);
nor_5  g03331(new_n5679, new_n5677, new_n5680_1);
xnor_4 g03332(new_n5679, new_n5677, new_n5681);
xnor_4 g03333(new_n5537, new_n5503, new_n5682);
xnor_4 g03334(new_n5667, new_n5630, new_n5683);
nor_5  g03335(new_n5683, new_n5682, new_n5684);
xnor_4 g03336(new_n5683, new_n5682, new_n5685);
xnor_4 g03337(new_n5535, new_n5507, new_n5686);
xnor_4 g03338(new_n5665, new_n5663, new_n5687_1);
nor_5  g03339(new_n5687_1, new_n5686, new_n5688);
xnor_4 g03340(new_n5687_1, new_n5686, new_n5689);
xnor_4 g03341(new_n5533, new_n5511, new_n5690);
not_8  g03342(new_n5661, new_n5691);
xnor_4 g03343(new_n5691, new_n5659, new_n5692);
not_8  g03344(new_n5692, new_n5693);
nor_5  g03345(new_n5693, new_n5690, new_n5694);
xnor_4 g03346(new_n5693, new_n5690, new_n5695);
not_8  g03347(new_n5638, new_n5696_1);
xnor_4 g03348(new_n5654, new_n5696_1, new_n5697);
not_8  g03349(new_n5697, new_n5698);
xnor_4 g03350(new_n5531, new_n5530, new_n5699);
nor_5  g03351(new_n5699, new_n5698, new_n5700_1);
xnor_4 g03352(new_n5699, new_n5697, new_n5701);
not_8  g03353(new_n5701, new_n5702);
xnor_4 g03354(new_n5528, new_n5519, new_n5703);
not_8  g03355(new_n5703, new_n5704_1);
not_8  g03356(new_n5652, new_n5705);
xnor_4 g03357(new_n5705, new_n5651, new_n5706);
nor_5  g03358(new_n5706, new_n5704_1, new_n5707);
not_8  g03359(new_n5707, new_n5708);
xnor_4 g03360(new_n5706, new_n5703, new_n5709);
xnor_4 g03361(new_n5649, new_n5648, new_n5710);
nor_5  g03362(new_n5710, new_n5524_1, new_n5711);
not_8  g03363(new_n5710, new_n5712);
xnor_4 g03364(new_n5524_1, new_n5523, new_n5713);
nor_5  g03365(new_n5713, new_n5712, new_n5714);
xnor_4 g03366(n23333, new_n3350, new_n5715);
not_8  g03367(new_n5715, new_n5716);
xnor_4 g03368(new_n5647, new_n5645, new_n5717);
nor_5  g03369(new_n5717, new_n5716, new_n5718);
nor_5  g03370(new_n5718, new_n5714, new_n5719);
nor_5  g03371(new_n5719, new_n5711, new_n5720);
nand_5 g03372(new_n5720, new_n5709, new_n5721);
nand_5 g03373(new_n5721, new_n5708, new_n5722);
nor_5  g03374(new_n5722, new_n5702, new_n5723);
nor_5  g03375(new_n5723, new_n5700_1, new_n5724);
nor_5  g03376(new_n5724, new_n5695, new_n5725);
nor_5  g03377(new_n5725, new_n5694, new_n5726);
nor_5  g03378(new_n5726, new_n5689, new_n5727);
nor_5  g03379(new_n5727, new_n5688, new_n5728);
nor_5  g03380(new_n5728, new_n5685, new_n5729);
nor_5  g03381(new_n5729, new_n5684, new_n5730);
nor_5  g03382(new_n5730, new_n5681, new_n5731);
nor_5  g03383(new_n5731, new_n5680_1, new_n5732_1);
nand_5 g03384(new_n5732_1, new_n5676, new_n5733);
not_8  g03385(new_n5733, new_n5734);
nor_5  g03386(new_n5732_1, new_n5676, new_n5735);
nor_5  g03387(new_n5735, new_n5734, n431);
not_8  g03388(n23895, new_n5737);
or_5   g03389(new_n5737, n8614, new_n5738);
xnor_4 g03390(n23895, n8614, new_n5739);
not_8  g03391(n17351, new_n5740);
or_5   g03392(new_n5740, n15182, new_n5741);
xnor_4 g03393(n17351, n15182, new_n5742_1);
not_8  g03394(n11736, new_n5743);
or_5   g03395(n27037, new_n5743, new_n5744);
xnor_4 g03396(n27037, n11736, new_n5745);
not_8  g03397(n23200, new_n5746);
or_5   g03398(new_n5746, n8964, new_n5747);
xnor_4 g03399(n23200, n8964, new_n5748);
not_8  g03400(n17959, new_n5749);
or_5   g03401(n20151, new_n5749, new_n5750);
xnor_4 g03402(n20151, n17959, new_n5751);
not_8  g03403(n7566, new_n5752_1);
nor_5  g03404(n7693, new_n5752_1, new_n5753);
xnor_4 g03405(n7693, n7566, new_n5754);
not_8  g03406(n7731, new_n5755);
nor_5  g03407(n10405, new_n5755, new_n5756);
not_8  g03408(new_n5756, new_n5757);
xnor_4 g03409(n10405, n7731, new_n5758);
nor_5  g03410(n12341, new_n4199, new_n5759);
not_8  g03411(n12341, new_n5760);
nor_5  g03412(new_n5760, n11302, new_n5761);
nor_5  g03413(n20986, new_n4201, new_n5762);
not_8  g03414(n20986, new_n5763);
nor_5  g03415(new_n5763, n17090, new_n5764);
nor_5  g03416(n12384, new_n2575, new_n5765_1);
not_8  g03417(new_n5765_1, new_n5766);
nor_5  g03418(new_n5766, new_n5764, new_n5767);
nor_5  g03419(new_n5767, new_n5762, new_n5768);
nor_5  g03420(new_n5768, new_n5761, new_n5769);
nor_5  g03421(new_n5769, new_n5759, new_n5770);
nand_5 g03422(new_n5770, new_n5758, new_n5771);
nand_5 g03423(new_n5771, new_n5757, new_n5772);
and_5  g03424(new_n5772, new_n5754, new_n5773);
nor_5  g03425(new_n5773, new_n5753, new_n5774);
not_8  g03426(new_n5774, new_n5775);
nand_5 g03427(new_n5775, new_n5751, new_n5776_1);
nand_5 g03428(new_n5776_1, new_n5750, new_n5777);
nand_5 g03429(new_n5777, new_n5748, new_n5778);
nand_5 g03430(new_n5778, new_n5747, new_n5779);
nand_5 g03431(new_n5779, new_n5745, new_n5780);
nand_5 g03432(new_n5780, new_n5744, new_n5781);
nand_5 g03433(new_n5781, new_n5742_1, new_n5782_1);
nand_5 g03434(new_n5782_1, new_n5741, new_n5783);
nand_5 g03435(new_n5783, new_n5739, new_n5784);
nand_5 g03436(new_n5784, new_n5738, new_n5785);
not_8  g03437(new_n5785, new_n5786);
not_8  g03438(n13494, new_n5787);
or_5   g03439(n18880, new_n5787, new_n5788);
xnor_4 g03440(n18880, n13494, new_n5789);
not_8  g03441(n25345, new_n5790);
or_5   g03442(n25475, new_n5790, new_n5791);
xnor_4 g03443(n25475, n25345, new_n5792);
not_8  g03444(n9655, new_n5793);
or_5   g03445(n23849, new_n5793, new_n5794);
xnor_4 g03446(n23849, n9655, new_n5795);
not_8  g03447(n13490, new_n5796);
or_5   g03448(new_n5796, n12446, new_n5797);
xnor_4 g03449(n13490, n12446, new_n5798);
nand_5 g03450(n22660, new_n4631, new_n5799);
xnor_4 g03451(n22660, n11011, new_n5800);
nor_5  g03452(n16029, new_n2437, new_n5801);
xnor_4 g03453(n16029, n1777, new_n5802);
not_8  g03454(new_n5802, new_n5803);
nor_5  g03455(n16476, new_n2441, new_n5804);
xnor_4 g03456(n16476, n8745, new_n5805);
nor_5  g03457(n15636, new_n4115, new_n5806);
nor_5  g03458(new_n2445, n11615, new_n5807);
nor_5  g03459(new_n4120, n20077, new_n5808);
not_8  g03460(n20077, new_n5809);
nor_5  g03461(n22433, new_n5809, new_n5810);
nor_5  g03462(new_n2580, n6794, new_n5811);
not_8  g03463(new_n5811, new_n5812);
nor_5  g03464(new_n5812, new_n5810, new_n5813);
nor_5  g03465(new_n5813, new_n5808, new_n5814);
nor_5  g03466(new_n5814, new_n5807, new_n5815);
nor_5  g03467(new_n5815, new_n5806, new_n5816);
nand_5 g03468(new_n5816, new_n5805, new_n5817);
not_8  g03469(new_n5817, new_n5818);
nor_5  g03470(new_n5818, new_n5804, new_n5819);
nor_5  g03471(new_n5819, new_n5803, new_n5820);
nor_5  g03472(new_n5820, new_n5801, new_n5821);
not_8  g03473(new_n5821, new_n5822_1);
nand_5 g03474(new_n5822_1, new_n5800, new_n5823);
nand_5 g03475(new_n5823, new_n5799, new_n5824);
nand_5 g03476(new_n5824, new_n5798, new_n5825);
nand_5 g03477(new_n5825, new_n5797, new_n5826);
nand_5 g03478(new_n5826, new_n5795, new_n5827);
nand_5 g03479(new_n5827, new_n5794, new_n5828);
nand_5 g03480(new_n5828, new_n5792, new_n5829);
nand_5 g03481(new_n5829, new_n5791, new_n5830);
nand_5 g03482(new_n5830, new_n5789, new_n5831);
nand_5 g03483(new_n5831, new_n5788, new_n5832);
not_8  g03484(new_n5832, new_n5833_1);
xnor_4 g03485(new_n5830, new_n5789, new_n5834_1);
not_8  g03486(n10201, new_n5835);
not_8  g03487(n22554, new_n5836);
not_8  g03488(n3909, new_n5837);
not_8  g03489(n2146, new_n5838);
nor_5  g03490(n22173, n583, new_n5839);
nand_5 g03491(new_n5839, new_n5838, new_n5840_1);
nor_5  g03492(new_n5840_1, n23974, new_n5841_1);
nand_5 g03493(new_n5841_1, new_n5837, new_n5842_1);
nor_5  g03494(new_n5842_1, n20429, new_n5843);
nand_5 g03495(new_n5843, new_n5836, new_n5844);
nor_5  g03496(new_n5844, n23913, new_n5845);
xnor_4 g03497(new_n5845, n26797, new_n5846);
not_8  g03498(new_n5846, new_n5847);
nand_5 g03499(new_n5847, new_n5835, new_n5848);
xnor_4 g03500(new_n5846, new_n5835, new_n5849);
not_8  g03501(n10593, new_n5850_1);
not_8  g03502(n23913, new_n5851);
xnor_4 g03503(new_n5844, new_n5851, new_n5852);
not_8  g03504(new_n5852, new_n5853);
nand_5 g03505(new_n5853, new_n5850_1, new_n5854);
xnor_4 g03506(new_n5852, new_n5850_1, new_n5855);
not_8  g03507(n18290, new_n5856);
xnor_4 g03508(new_n5843, n22554, new_n5857);
not_8  g03509(new_n5857, new_n5858);
nand_5 g03510(new_n5858, new_n5856, new_n5859);
xnor_4 g03511(new_n5857, new_n5856, new_n5860);
not_8  g03512(n11580, new_n5861);
not_8  g03513(n20429, new_n5862);
xnor_4 g03514(new_n5842_1, new_n5862, new_n5863);
not_8  g03515(new_n5863, new_n5864);
nand_5 g03516(new_n5864, new_n5861, new_n5865);
xnor_4 g03517(new_n5863, new_n5861, new_n5866);
not_8  g03518(n15884, new_n5867);
xnor_4 g03519(new_n5841_1, n3909, new_n5868);
not_8  g03520(new_n5868, new_n5869);
nand_5 g03521(new_n5869, new_n5867, new_n5870);
xnor_4 g03522(new_n5868, new_n5867, new_n5871);
not_8  g03523(n6356, new_n5872);
not_8  g03524(n23974, new_n5873);
xnor_4 g03525(new_n5840_1, new_n5873, new_n5874);
not_8  g03526(new_n5874, new_n5875);
nand_5 g03527(new_n5875, new_n5872, new_n5876);
not_8  g03528(n27104, new_n5877);
xnor_4 g03529(new_n5839, n2146, new_n5878);
not_8  g03530(new_n5878, new_n5879);
nand_5 g03531(new_n5879, new_n5877, new_n5880);
xnor_4 g03532(new_n5878, new_n5877, new_n5881);
not_8  g03533(n27188, new_n5882_1);
xnor_4 g03534(n22173, n583, new_n5883);
nand_5 g03535(new_n5883, new_n5882_1, new_n5884);
nand_5 g03536(n6611, n583, new_n5885);
xnor_4 g03537(new_n5883, n27188, new_n5886);
nand_5 g03538(new_n5886, new_n5885, new_n5887);
nand_5 g03539(new_n5887, new_n5884, new_n5888);
nand_5 g03540(new_n5888, new_n5881, new_n5889);
nand_5 g03541(new_n5889, new_n5880, new_n5890);
xnor_4 g03542(new_n5874, new_n5872, new_n5891);
nand_5 g03543(new_n5891, new_n5890, new_n5892);
nand_5 g03544(new_n5892, new_n5876, new_n5893);
nand_5 g03545(new_n5893, new_n5871, new_n5894);
nand_5 g03546(new_n5894, new_n5870, new_n5895);
nand_5 g03547(new_n5895, new_n5866, new_n5896);
nand_5 g03548(new_n5896, new_n5865, new_n5897);
nand_5 g03549(new_n5897, new_n5860, new_n5898);
nand_5 g03550(new_n5898, new_n5859, new_n5899);
nand_5 g03551(new_n5899, new_n5855, new_n5900);
nand_5 g03552(new_n5900, new_n5854, new_n5901);
nand_5 g03553(new_n5901, new_n5849, new_n5902);
nand_5 g03554(new_n5902, new_n5848, new_n5903_1);
not_8  g03555(n12650, new_n5904_1);
not_8  g03556(n12702, new_n5905);
not_8  g03557(n26797, new_n5906);
nand_5 g03558(new_n5845, new_n5906, new_n5907);
xnor_4 g03559(new_n5907, new_n5905, new_n5908);
xnor_4 g03560(new_n5908, new_n5904_1, new_n5909);
xnor_4 g03561(new_n5909, new_n5903_1, new_n5910);
not_8  g03562(new_n5910, new_n5911_1);
nand_5 g03563(new_n5911_1, new_n5834_1, new_n5912);
xnor_4 g03564(new_n5910, new_n5834_1, new_n5913);
xnor_4 g03565(new_n5828, new_n5792, new_n5914);
xnor_4 g03566(new_n5901, new_n5849, new_n5915);
not_8  g03567(new_n5915, new_n5916);
nand_5 g03568(new_n5916, new_n5914, new_n5917);
xnor_4 g03569(new_n5915, new_n5914, new_n5918);
xnor_4 g03570(new_n5826, new_n5795, new_n5919);
xnor_4 g03571(new_n5899, new_n5855, new_n5920);
not_8  g03572(new_n5920, new_n5921);
nand_5 g03573(new_n5921, new_n5919, new_n5922);
xnor_4 g03574(new_n5920, new_n5919, new_n5923);
xnor_4 g03575(new_n5824, new_n5798, new_n5924);
xnor_4 g03576(new_n5897, new_n5860, new_n5925);
not_8  g03577(new_n5925, new_n5926);
nand_5 g03578(new_n5926, new_n5924, new_n5927);
xnor_4 g03579(new_n5925, new_n5924, new_n5928);
xnor_4 g03580(new_n5821, new_n5800, new_n5929);
not_8  g03581(new_n5929, new_n5930);
not_8  g03582(new_n5866, new_n5931);
xnor_4 g03583(new_n5895, new_n5931, new_n5932);
nand_5 g03584(new_n5932, new_n5930, new_n5933);
xnor_4 g03585(new_n5932, new_n5929, new_n5934);
xnor_4 g03586(new_n5819, new_n5803, new_n5935);
xnor_4 g03587(new_n5893, new_n5871, new_n5936_1);
not_8  g03588(new_n5936_1, new_n5937);
nand_5 g03589(new_n5937, new_n5935, new_n5938);
xnor_4 g03590(new_n5936_1, new_n5935, new_n5939);
not_8  g03591(new_n5816, new_n5940);
xnor_4 g03592(new_n5940, new_n5805, new_n5941);
xnor_4 g03593(new_n5891, new_n5890, new_n5942);
nor_5  g03594(new_n5942, new_n5941, new_n5943_1);
not_8  g03595(new_n5943_1, new_n5944);
not_8  g03596(new_n5941, new_n5945);
xnor_4 g03597(new_n5942, new_n5945, new_n5946);
xnor_4 g03598(new_n5888, new_n5881, new_n5947);
xnor_4 g03599(n15636, n11615, new_n5948);
xnor_4 g03600(new_n5948, new_n5814, new_n5949);
not_8  g03601(new_n5949, new_n5950);
nand_5 g03602(new_n5950, new_n5947, new_n5951);
not_8  g03603(new_n5951, new_n5952);
xnor_4 g03604(new_n5949, new_n5947, new_n5953);
not_8  g03605(new_n5953, new_n5954);
xnor_4 g03606(new_n5886, new_n5885, new_n5955);
xnor_4 g03607(n22433, n20077, new_n5956);
xnor_4 g03608(new_n5956, new_n5811, new_n5957);
nand_5 g03609(new_n5957, new_n5955, new_n5958);
not_8  g03610(new_n5958, new_n5959);
xnor_4 g03611(n14090, n6794, new_n5960);
not_8  g03612(n583, new_n5961);
xnor_4 g03613(n6611, new_n5961, new_n5962);
not_8  g03614(new_n5962, new_n5963);
nor_5  g03615(new_n5963, new_n5960, new_n5964_1);
not_8  g03616(new_n5964_1, new_n5965);
xnor_4 g03617(new_n5957, new_n5955, new_n5966);
nor_5  g03618(new_n5966, new_n5965, new_n5967);
nor_5  g03619(new_n5967, new_n5959, new_n5968);
nor_5  g03620(new_n5968, new_n5954, new_n5969);
nor_5  g03621(new_n5969, new_n5952, new_n5970);
nand_5 g03622(new_n5970, new_n5946, new_n5971);
nand_5 g03623(new_n5971, new_n5944, new_n5972);
nand_5 g03624(new_n5972, new_n5939, new_n5973);
nand_5 g03625(new_n5973, new_n5938, new_n5974);
nand_5 g03626(new_n5974, new_n5934, new_n5975);
nand_5 g03627(new_n5975, new_n5933, new_n5976);
nand_5 g03628(new_n5976, new_n5928, new_n5977);
nand_5 g03629(new_n5977, new_n5927, new_n5978);
nand_5 g03630(new_n5978, new_n5923, new_n5979);
nand_5 g03631(new_n5979, new_n5922, new_n5980_1);
nand_5 g03632(new_n5980_1, new_n5918, new_n5981);
nand_5 g03633(new_n5981, new_n5917, new_n5982);
nand_5 g03634(new_n5982, new_n5913, new_n5983);
nand_5 g03635(new_n5983, new_n5912, new_n5984);
nor_5  g03636(new_n5907, n12702, new_n5985);
and_5  g03637(new_n5908, n12650, new_n5986);
nor_5  g03638(new_n5908, n12650, new_n5987);
nor_5  g03639(new_n5987, new_n5903_1, new_n5988);
nor_5  g03640(new_n5988, new_n5986, new_n5989);
not_8  g03641(new_n5989, new_n5990);
nor_5  g03642(new_n5990, new_n5985, new_n5991);
nor_5  g03643(new_n5991, new_n5984, new_n5992);
nand_5 g03644(new_n5992, new_n5833_1, new_n5993);
not_8  g03645(new_n5993, new_n5994);
nand_5 g03646(new_n5991, new_n5984, new_n5995);
nor_5  g03647(new_n5995, new_n5833_1, new_n5996);
nor_5  g03648(new_n5996, new_n5994, new_n5997);
xnor_4 g03649(new_n5997, new_n5786, new_n5998);
not_8  g03650(new_n5991, new_n5999);
xnor_4 g03651(new_n5999, new_n5984, new_n6000);
xnor_4 g03652(new_n6000, new_n5833_1, new_n6001);
not_8  g03653(new_n6001, new_n6002);
nor_5  g03654(new_n6002, new_n5785, new_n6003);
nor_5  g03655(new_n6001, new_n5786, new_n6004);
xnor_4 g03656(new_n5783, new_n5739, new_n6005);
xnor_4 g03657(new_n5982, new_n5913, new_n6006);
not_8  g03658(new_n6006, new_n6007);
nand_5 g03659(new_n6007, new_n6005, new_n6008);
xnor_4 g03660(new_n6006, new_n6005, new_n6009);
xnor_4 g03661(new_n5781, new_n5742_1, new_n6010);
xnor_4 g03662(new_n5980_1, new_n5918, new_n6011);
not_8  g03663(new_n6011, new_n6012_1);
nand_5 g03664(new_n6012_1, new_n6010, new_n6013);
xnor_4 g03665(new_n6011, new_n6010, new_n6014);
xnor_4 g03666(new_n5779, new_n5745, new_n6015);
xnor_4 g03667(new_n5978, new_n5923, new_n6016);
not_8  g03668(new_n6016, new_n6017);
nand_5 g03669(new_n6017, new_n6015, new_n6018);
xnor_4 g03670(new_n6016, new_n6015, new_n6019);
xnor_4 g03671(new_n5777, new_n5748, new_n6020);
xnor_4 g03672(new_n5976, new_n5928, new_n6021);
not_8  g03673(new_n6021, new_n6022_1);
nand_5 g03674(new_n6022_1, new_n6020, new_n6023);
xnor_4 g03675(new_n6021, new_n6020, new_n6024);
xnor_4 g03676(new_n5774, new_n5751, new_n6025);
not_8  g03677(new_n6025, new_n6026);
not_8  g03678(new_n5934, new_n6027);
xnor_4 g03679(new_n5974, new_n6027, new_n6028);
nand_5 g03680(new_n6028, new_n6026, new_n6029);
xnor_4 g03681(new_n6028, new_n6025, new_n6030);
not_8  g03682(new_n5754, new_n6031_1);
xnor_4 g03683(new_n5772, new_n6031_1, new_n6032);
not_8  g03684(new_n6032, new_n6033);
not_8  g03685(new_n5939, new_n6034);
xnor_4 g03686(new_n5972, new_n6034, new_n6035);
nand_5 g03687(new_n6035, new_n6033, new_n6036);
xnor_4 g03688(new_n6035, new_n6032, new_n6037);
xnor_4 g03689(new_n5970, new_n5946, new_n6038);
not_8  g03690(new_n6038, new_n6039);
xnor_4 g03691(new_n5770, new_n5758, new_n6040);
nand_5 g03692(new_n6040, new_n6039, new_n6041);
xnor_4 g03693(new_n6040, new_n6038, new_n6042);
xnor_4 g03694(new_n5968, new_n5953, new_n6043);
not_8  g03695(new_n6043, new_n6044_1);
xnor_4 g03696(n12341, n11302, new_n6045);
xnor_4 g03697(new_n6045, new_n5768, new_n6046_1);
nand_5 g03698(new_n6046_1, new_n6044_1, new_n6047);
xnor_4 g03699(new_n6046_1, new_n6043, new_n6048);
xnor_4 g03700(new_n5962, new_n5960, new_n6049);
not_8  g03701(new_n6049, new_n6050);
xnor_4 g03702(n12384, n6773, new_n6051);
nor_5  g03703(new_n6051, new_n6050, new_n6052);
xnor_4 g03704(n20986, n17090, new_n6053);
xnor_4 g03705(new_n6053, new_n5766, new_n6054);
not_8  g03706(new_n6054, new_n6055);
nor_5  g03707(new_n6055, new_n6052, new_n6056);
not_8  g03708(new_n6056, new_n6057);
xnor_4 g03709(new_n5966, new_n5964_1, new_n6058);
not_8  g03710(new_n6058, new_n6059);
xnor_4 g03711(new_n6054, new_n6052, new_n6060);
nand_5 g03712(new_n6060, new_n6059, new_n6061);
nand_5 g03713(new_n6061, new_n6057, new_n6062);
nand_5 g03714(new_n6062, new_n6048, new_n6063);
nand_5 g03715(new_n6063, new_n6047, new_n6064);
nand_5 g03716(new_n6064, new_n6042, new_n6065);
nand_5 g03717(new_n6065, new_n6041, new_n6066);
nand_5 g03718(new_n6066, new_n6037, new_n6067);
nand_5 g03719(new_n6067, new_n6036, new_n6068);
nand_5 g03720(new_n6068, new_n6030, new_n6069);
nand_5 g03721(new_n6069, new_n6029, new_n6070);
nand_5 g03722(new_n6070, new_n6024, new_n6071);
nand_5 g03723(new_n6071, new_n6023, new_n6072);
nand_5 g03724(new_n6072, new_n6019, new_n6073);
nand_5 g03725(new_n6073, new_n6018, new_n6074);
nand_5 g03726(new_n6074, new_n6014, new_n6075);
nand_5 g03727(new_n6075, new_n6013, new_n6076);
nand_5 g03728(new_n6076, new_n6009, new_n6077);
nand_5 g03729(new_n6077, new_n6008, new_n6078);
nor_5  g03730(new_n6078, new_n6004, new_n6079);
nor_5  g03731(new_n6079, new_n6003, new_n6080);
xnor_4 g03732(new_n6080, new_n5998, n457);
not_8  g03733(new_n5957, new_n6082);
xnor_4 g03734(n24323, n1681, new_n6083);
xnor_4 g03735(n13781, n2088, new_n6084_1);
xnor_4 g03736(new_n6084_1, new_n6083, new_n6085);
nor_5  g03737(new_n6085, new_n5960, new_n6086);
xnor_4 g03738(new_n6086, new_n6082, new_n6087);
not_8  g03739(new_n6087, new_n6088);
nor_5  g03740(new_n6084_1, new_n6083, new_n6089);
nor_5  g03741(n24323, new_n2568, new_n6090);
xnor_4 g03742(n26443, n25877, new_n6091);
xnor_4 g03743(new_n6091, new_n6090, new_n6092);
not_8  g03744(new_n6092, new_n6093);
xnor_4 g03745(new_n6093, new_n6089, new_n6094);
xnor_4 g03746(n9399, new_n3078, new_n6095);
not_8  g03747(new_n6095, new_n6096);
not_8  g03748(n11486, new_n6097);
nand_5 g03749(n13781, n2088, new_n6098);
nand_5 g03750(new_n6098, new_n6097, new_n6099);
nand_5 g03751(n13781, n11486, new_n6100);
nor_5  g03752(new_n6100, new_n3078, new_n6101);
not_8  g03753(new_n6101, new_n6102);
nand_5 g03754(new_n6102, new_n6099, new_n6103);
xnor_4 g03755(new_n6103, new_n6096, new_n6104_1);
xnor_4 g03756(new_n6104_1, new_n6094, new_n6105_1);
xnor_4 g03757(new_n6105_1, new_n6088, n463);
not_8  g03758(n6775, new_n6107);
xnor_4 g03759(n12121, new_n6107, new_n6108);
xnor_4 g03760(new_n6108, new_n4452, new_n6109);
not_8  g03761(new_n6109, new_n6110);
xnor_4 g03762(new_n3076_1, n5438, new_n6111);
xnor_4 g03763(new_n6111, new_n6110, n491);
xnor_4 g03764(new_n6064, new_n6042, n496);
xnor_4 g03765(n25926, n12384, new_n6114);
xnor_4 g03766(new_n6114, n6773, new_n6115);
not_8  g03767(new_n6115, new_n6116);
xnor_4 g03768(new_n5960, n16167, new_n6117);
not_8  g03769(new_n6117, new_n6118);
nor_5  g03770(new_n6118, new_n6116, new_n6119);
not_8  g03771(n16167, new_n6120);
nor_5  g03772(new_n5960, new_n6120, new_n6121);
not_8  g03773(n18745, new_n6122);
xnor_4 g03774(new_n5957, new_n6122, new_n6123);
xnor_4 g03775(new_n6123, new_n6121, new_n6124);
nand_5 g03776(n25926, n12384, new_n6125);
xnor_4 g03777(n25926, n7657, new_n6126);
xnor_4 g03778(new_n6126, new_n5763, new_n6127);
xnor_4 g03779(new_n6127, new_n6125, new_n6128);
nor_5  g03780(new_n6114, new_n2575, new_n6129);
nand_5 g03781(new_n6129, new_n4201, new_n6130);
nor_5  g03782(n17090, n6773, new_n6131);
not_8  g03783(new_n6131, new_n6132);
nand_5 g03784(n17090, n6773, new_n6133);
not_8  g03785(new_n6133, new_n6134);
nand_5 g03786(new_n6134, new_n6114, new_n6135);
nand_5 g03787(new_n6135, new_n6132, new_n6136);
not_8  g03788(new_n6136, new_n6137);
nand_5 g03789(new_n6137, new_n6130, new_n6138);
xnor_4 g03790(new_n6138, new_n6128, new_n6139);
not_8  g03791(new_n6139, new_n6140);
xnor_4 g03792(new_n6140, new_n6124, new_n6141);
not_8  g03793(new_n6141, new_n6142);
xnor_4 g03794(new_n6142, new_n6119, n498);
not_8  g03795(new_n5118, new_n6144);
xnor_4 g03796(n25872, new_n3994, new_n6145);
nor_5  g03797(n22043, n20259, new_n6146);
nand_5 g03798(n12121, n3925, new_n6147);
not_8  g03799(new_n6147, new_n6148);
xnor_4 g03800(n22043, n20259, new_n6149);
nor_5  g03801(new_n6149, new_n6148, new_n6150);
nor_5  g03802(new_n6150, new_n6146, new_n6151);
xnor_4 g03803(new_n6151, new_n6145, new_n6152);
xnor_4 g03804(new_n6152, new_n6144, new_n6153);
not_8  g03805(new_n5122, new_n6154);
xnor_4 g03806(new_n6149, new_n6147, new_n6155);
nor_5  g03807(new_n6155, new_n6154, new_n6156);
not_8  g03808(new_n5126, new_n6157);
not_8  g03809(n3925, new_n6158);
xnor_4 g03810(n12121, new_n6158, new_n6159);
nor_5  g03811(new_n6159, new_n6157, new_n6160_1);
xnor_4 g03812(new_n6155, new_n6154, new_n6161);
nor_5  g03813(new_n6161, new_n6160_1, new_n6162);
nor_5  g03814(new_n6162, new_n6156, new_n6163);
xnor_4 g03815(new_n6163, new_n6153, new_n6164);
xnor_4 g03816(new_n6164, new_n3939, new_n6165);
xnor_4 g03817(new_n6161, new_n6160_1, new_n6166);
not_8  g03818(new_n6166, new_n6167);
nor_5  g03819(new_n6167, new_n3913, new_n6168);
not_8  g03820(new_n3943, new_n6169);
nor_5  g03821(new_n6166, new_n6169, new_n6170);
xnor_4 g03822(new_n6159, new_n5126, new_n6171_1);
nor_5  g03823(new_n6171_1, new_n3948, new_n6172);
nor_5  g03824(new_n6172, new_n6170, new_n6173);
nor_5  g03825(new_n6173, new_n6168, new_n6174);
xor_4  g03826(new_n6174, new_n6165, n521);
xnor_4 g03827(new_n6051, new_n6049, n548);
xor_4  g03828(new_n4497, new_n4475, n554);
nor_5  g03829(n20658, n15743, new_n6178);
nand_5 g03830(new_n6178, new_n3941, new_n6179);
nor_5  g03831(new_n6179, n4957, new_n6180);
nand_5 g03832(new_n6180, new_n3933, new_n6181);
nor_5  g03833(new_n6181, n3161, new_n6182);
nand_5 g03834(new_n6182, new_n3877, new_n6183_1);
nor_5  g03835(new_n6183_1, n20409, new_n6184);
nand_5 g03836(new_n6184, new_n5046_1, new_n6185);
xnor_4 g03837(new_n6185, n2979, new_n6186);
not_8  g03838(new_n6186, new_n6187);
not_8  g03839(n6456, new_n6188);
xnor_4 g03840(n9259, new_n6188, new_n6189_1);
or_5   g03841(n21489, n4085, new_n6190);
not_8  g03842(n4085, new_n6191);
xnor_4 g03843(n21489, new_n6191, new_n6192);
or_5   g03844(n26725, n20213, new_n6193);
xnor_4 g03845(n26725, new_n3746, new_n6194);
nor_5  g03846(n13912, n11980, new_n6195);
not_8  g03847(n11980, new_n6196);
xnor_4 g03848(n13912, new_n6196, new_n6197);
not_8  g03849(new_n6197, new_n6198);
nor_5  g03850(n7670, n3253, new_n6199);
not_8  g03851(n3253, new_n6200);
xnor_4 g03852(n7670, new_n6200, new_n6201);
not_8  g03853(new_n6201, new_n6202);
nor_5  g03854(n9598, n7759, new_n6203);
not_8  g03855(n7759, new_n6204_1);
xnor_4 g03856(n9598, new_n6204_1, new_n6205);
not_8  g03857(new_n6205, new_n6206);
nor_5  g03858(n22290, n12562, new_n6207);
not_8  g03859(n12562, new_n6208);
xnor_4 g03860(n22290, new_n6208, new_n6209);
not_8  g03861(new_n6209, new_n6210);
nor_5  g03862(n11273, n7949, new_n6211);
not_8  g03863(n7949, new_n6212);
xnor_4 g03864(n11273, new_n6212, new_n6213);
not_8  g03865(new_n6213, new_n6214);
nor_5  g03866(n25565, n24374, new_n6215);
nand_5 g03867(n21993, n14575, new_n6216);
not_8  g03868(new_n6216, new_n6217);
xnor_4 g03869(n25565, n24374, new_n6218_1);
nor_5  g03870(new_n6218_1, new_n6217, new_n6219);
nor_5  g03871(new_n6219, new_n6215, new_n6220);
nor_5  g03872(new_n6220, new_n6214, new_n6221);
nor_5  g03873(new_n6221, new_n6211, new_n6222);
nor_5  g03874(new_n6222, new_n6210, new_n6223_1);
nor_5  g03875(new_n6223_1, new_n6207, new_n6224);
nor_5  g03876(new_n6224, new_n6206, new_n6225);
nor_5  g03877(new_n6225, new_n6203, new_n6226);
nor_5  g03878(new_n6226, new_n6202, new_n6227);
nor_5  g03879(new_n6227, new_n6199, new_n6228);
nor_5  g03880(new_n6228, new_n6198, new_n6229);
nor_5  g03881(new_n6229, new_n6195, new_n6230);
not_8  g03882(new_n6230, new_n6231);
nand_5 g03883(new_n6231, new_n6194, new_n6232);
nand_5 g03884(new_n6232, new_n6193, new_n6233_1);
nand_5 g03885(new_n6233_1, new_n6192, new_n6234);
nand_5 g03886(new_n6234, new_n6190, new_n6235);
xnor_4 g03887(new_n6235, new_n6189_1, new_n6236);
xnor_4 g03888(new_n6236, new_n6187, new_n6237);
xnor_4 g03889(new_n6184, n647, new_n6238);
not_8  g03890(new_n6238, new_n6239);
xnor_4 g03891(new_n6233_1, new_n6192, new_n6240);
nor_5  g03892(new_n6240, new_n6239, new_n6241);
xnor_4 g03893(new_n6240, new_n6239, new_n6242);
not_8  g03894(n20409, new_n6243);
xnor_4 g03895(new_n6183_1, new_n6243, new_n6244);
not_8  g03896(new_n6244, new_n6245_1);
xnor_4 g03897(new_n6230, new_n6194, new_n6246);
not_8  g03898(new_n6246, new_n6247);
nand_5 g03899(new_n6247, new_n6245_1, new_n6248_1);
xnor_4 g03900(new_n6246, new_n6245_1, new_n6249);
xnor_4 g03901(new_n6182, n25749, new_n6250);
not_8  g03902(new_n6250, new_n6251);
xnor_4 g03903(new_n6228, new_n6197, new_n6252);
not_8  g03904(new_n6252, new_n6253);
nand_5 g03905(new_n6253, new_n6251, new_n6254);
xnor_4 g03906(new_n6252, new_n6251, new_n6255);
xnor_4 g03907(new_n6181, new_n3929, new_n6256_1);
not_8  g03908(new_n6256_1, new_n6257);
xnor_4 g03909(new_n6226, new_n6201, new_n6258);
not_8  g03910(new_n6258, new_n6259);
nand_5 g03911(new_n6259, new_n6257, new_n6260);
xnor_4 g03912(new_n6258, new_n6257, new_n6261);
xnor_4 g03913(new_n6180, n9003, new_n6262);
xnor_4 g03914(new_n6224, new_n6205, new_n6263);
nor_5  g03915(new_n6263, new_n6262, new_n6264);
not_8  g03916(new_n6264, new_n6265);
not_8  g03917(new_n6262, new_n6266);
xnor_4 g03918(new_n6263, new_n6266, new_n6267);
xnor_4 g03919(new_n6179, new_n3937, new_n6268);
xnor_4 g03920(new_n6222, new_n6209, new_n6269);
nor_5  g03921(new_n6269, new_n6268, new_n6270);
not_8  g03922(new_n6270, new_n6271_1);
not_8  g03923(new_n6268, new_n6272);
xnor_4 g03924(new_n6269, new_n6272, new_n6273);
xnor_4 g03925(new_n6178, n7524, new_n6274);
not_8  g03926(new_n6274, new_n6275);
xnor_4 g03927(new_n6220, new_n6213, new_n6276_1);
not_8  g03928(new_n6276_1, new_n6277);
nor_5  g03929(new_n6277, new_n6275, new_n6278);
xnor_4 g03930(new_n6276_1, new_n6275, new_n6279);
not_8  g03931(new_n6279, new_n6280);
not_8  g03932(n14575, new_n6281);
xnor_4 g03933(n21993, new_n6281, new_n6282);
not_8  g03934(new_n6282, new_n6283);
nor_5  g03935(new_n6283, n20658, new_n6284);
nand_5 g03936(new_n6284, new_n3950, new_n6285);
xnor_4 g03937(new_n6218_1, new_n6217, new_n6286);
not_8  g03938(new_n6285, new_n6287);
xnor_4 g03939(n20658, n15743, new_n6288);
nor_5  g03940(new_n6288, new_n6284, new_n6289);
nor_5  g03941(new_n6289, new_n6287, new_n6290);
nand_5 g03942(new_n6290, new_n6286, new_n6291);
nand_5 g03943(new_n6291, new_n6285, new_n6292);
nor_5  g03944(new_n6292, new_n6280, new_n6293);
nor_5  g03945(new_n6293, new_n6278, new_n6294);
nand_5 g03946(new_n6294, new_n6273, new_n6295);
nand_5 g03947(new_n6295, new_n6271_1, new_n6296);
nand_5 g03948(new_n6296, new_n6267, new_n6297);
nand_5 g03949(new_n6297, new_n6265, new_n6298);
nand_5 g03950(new_n6298, new_n6261, new_n6299);
nand_5 g03951(new_n6299, new_n6260, new_n6300);
nand_5 g03952(new_n6300, new_n6255, new_n6301);
nand_5 g03953(new_n6301, new_n6254, new_n6302);
nand_5 g03954(new_n6302, new_n6249, new_n6303);
nand_5 g03955(new_n6303, new_n6248_1, new_n6304);
nor_5  g03956(new_n6304, new_n6242, new_n6305);
nor_5  g03957(new_n6305, new_n6241, new_n6306);
xnor_4 g03958(new_n6306, new_n6237, new_n6307);
not_8  g03959(n8526, new_n6308_1);
not_8  g03960(n3582, new_n6309);
xnor_4 g03961(n21784, new_n6309, new_n6310);
or_5   g03962(n5521, n2145, new_n6311_1);
not_8  g03963(n2145, new_n6312);
xnor_4 g03964(n5521, new_n6312, new_n6313);
or_5   g03965(n11926, n5031, new_n6314);
not_8  g03966(n5031, new_n6315);
xnor_4 g03967(n11926, new_n6315, new_n6316);
nor_5  g03968(n11044, n4325, new_n6317);
not_8  g03969(n4325, new_n6318);
xnor_4 g03970(n11044, new_n6318, new_n6319);
not_8  g03971(new_n6319, new_n6320);
nor_5  g03972(n5337, n2421, new_n6321);
not_8  g03973(n2421, new_n6322);
xnor_4 g03974(n5337, new_n6322, new_n6323_1);
not_8  g03975(new_n6323_1, new_n6324);
nor_5  g03976(n987, n626, new_n6325);
xnor_4 g03977(n987, new_n3993, new_n6326);
not_8  g03978(new_n6326, new_n6327);
nor_5  g03979(n20478, n1204, new_n6328);
xnor_4 g03980(n20478, new_n4015, new_n6329);
not_8  g03981(new_n6329, new_n6330_1);
nor_5  g03982(n26882, n19618, new_n6331);
xnor_4 g03983(n26882, new_n3994, new_n6332);
not_8  g03984(new_n6332, new_n6333);
nor_5  g03985(n22619, n22043, new_n6334);
nand_5 g03986(n12121, n6775, new_n6335);
not_8  g03987(new_n6335, new_n6336);
xnor_4 g03988(n22619, n22043, new_n6337);
nor_5  g03989(new_n6337, new_n6336, new_n6338);
nor_5  g03990(new_n6338, new_n6334, new_n6339_1);
nor_5  g03991(new_n6339_1, new_n6333, new_n6340);
nor_5  g03992(new_n6340, new_n6331, new_n6341);
nor_5  g03993(new_n6341, new_n6330_1, new_n6342);
nor_5  g03994(new_n6342, new_n6328, new_n6343);
nor_5  g03995(new_n6343, new_n6327, new_n6344);
nor_5  g03996(new_n6344, new_n6325, new_n6345);
nor_5  g03997(new_n6345, new_n6324, new_n6346);
nor_5  g03998(new_n6346, new_n6321, new_n6347);
nor_5  g03999(new_n6347, new_n6320, new_n6348);
nor_5  g04000(new_n6348, new_n6317, new_n6349);
not_8  g04001(new_n6349, new_n6350);
nand_5 g04002(new_n6350, new_n6316, new_n6351);
nand_5 g04003(new_n6351, new_n6314, new_n6352);
nand_5 g04004(new_n6352, new_n6313, new_n6353);
nand_5 g04005(new_n6353, new_n6311_1, new_n6354_1);
xnor_4 g04006(new_n6354_1, new_n6310, new_n6355);
xnor_4 g04007(new_n6355, new_n6308_1, new_n6356_1);
xnor_4 g04008(new_n6352, new_n6313, new_n6357);
nand_5 g04009(new_n6357, n2816, new_n6358);
not_8  g04010(n2816, new_n6359);
xnor_4 g04011(new_n6357, new_n6359, new_n6360);
xnor_4 g04012(new_n6349, new_n6316, new_n6361);
not_8  g04013(new_n6361, new_n6362);
nand_5 g04014(new_n6362, n20359, new_n6363);
xnor_4 g04015(new_n6361, n20359, new_n6364);
xnor_4 g04016(new_n6347, new_n6319, new_n6365);
not_8  g04017(new_n6365, new_n6366);
nand_5 g04018(new_n6366, n4409, new_n6367);
xnor_4 g04019(new_n6365, n4409, new_n6368);
xnor_4 g04020(new_n6345, new_n6323_1, new_n6369_1);
not_8  g04021(new_n6369_1, new_n6370);
nand_5 g04022(new_n6370, n3570, new_n6371);
xnor_4 g04023(new_n6369_1, n3570, new_n6372);
not_8  g04024(n13668, new_n6373);
xnor_4 g04025(new_n6343, new_n6326, new_n6374);
nor_5  g04026(new_n6374, new_n6373, new_n6375_1);
not_8  g04027(new_n6375_1, new_n6376);
xnor_4 g04028(new_n6374, n13668, new_n6377);
xnor_4 g04029(new_n6341, new_n6329, new_n6378);
nor_5  g04030(new_n6378, new_n4417, new_n6379_1);
not_8  g04031(new_n6379_1, new_n6380);
xnor_4 g04032(new_n6378, n21276, new_n6381_1);
xnor_4 g04033(new_n6339_1, new_n6332, new_n6382);
nor_5  g04034(new_n6382, new_n4411, new_n6383_1);
xnor_4 g04035(new_n6337, new_n6335, new_n6384);
not_8  g04036(new_n6384, new_n6385_1);
nor_5  g04037(new_n6385_1, n10057, new_n6386);
not_8  g04038(new_n6108, new_n6387);
nor_5  g04039(new_n6387, new_n4452, new_n6388);
xnor_4 g04040(new_n6384, n10057, new_n6389);
not_8  g04041(new_n6389, new_n6390);
nor_5  g04042(new_n6390, new_n6388, new_n6391);
nor_5  g04043(new_n6391, new_n6386, new_n6392);
xnor_4 g04044(new_n6382, n26748, new_n6393);
nand_5 g04045(new_n6393, new_n6392, new_n6394);
not_8  g04046(new_n6394, new_n6395);
nor_5  g04047(new_n6395, new_n6383_1, new_n6396);
not_8  g04048(new_n6396, new_n6397_1);
nand_5 g04049(new_n6397_1, new_n6381_1, new_n6398);
nand_5 g04050(new_n6398, new_n6380, new_n6399);
nand_5 g04051(new_n6399, new_n6377, new_n6400);
nand_5 g04052(new_n6400, new_n6376, new_n6401);
nand_5 g04053(new_n6401, new_n6372, new_n6402);
nand_5 g04054(new_n6402, new_n6371, new_n6403);
nand_5 g04055(new_n6403, new_n6368, new_n6404);
nand_5 g04056(new_n6404, new_n6367, new_n6405);
nand_5 g04057(new_n6405, new_n6364, new_n6406);
nand_5 g04058(new_n6406, new_n6363, new_n6407_1);
nand_5 g04059(new_n6407_1, new_n6360, new_n6408);
nand_5 g04060(new_n6408, new_n6358, new_n6409);
xnor_4 g04061(new_n6409, new_n6356_1, new_n6410);
xnor_4 g04062(new_n6410, new_n6307, new_n6411);
xnor_4 g04063(new_n6407_1, new_n6360, new_n6412);
not_8  g04064(new_n6304, new_n6413);
xnor_4 g04065(new_n6413, new_n6242, new_n6414);
not_8  g04066(new_n6414, new_n6415);
nand_5 g04067(new_n6415, new_n6412, new_n6416);
xnor_4 g04068(new_n6414, new_n6412, new_n6417);
xnor_4 g04069(new_n6302, new_n6249, new_n6418);
not_8  g04070(new_n6418, new_n6419);
xnor_4 g04071(new_n6405, new_n6364, new_n6420);
nand_5 g04072(new_n6420, new_n6419, new_n6421);
xnor_4 g04073(new_n6420, new_n6418, new_n6422);
xnor_4 g04074(new_n6300, new_n6255, new_n6423);
not_8  g04075(new_n6423, new_n6424);
xnor_4 g04076(new_n6403, new_n6368, new_n6425);
nand_5 g04077(new_n6425, new_n6424, new_n6426);
xnor_4 g04078(new_n6425, new_n6423, new_n6427_1);
not_8  g04079(new_n6261, new_n6428);
xnor_4 g04080(new_n6298, new_n6428, new_n6429);
not_8  g04081(new_n6372, new_n6430);
xnor_4 g04082(new_n6401, new_n6430, new_n6431_1);
not_8  g04083(new_n6431_1, new_n6432);
nand_5 g04084(new_n6432, new_n6429, new_n6433);
xnor_4 g04085(new_n6431_1, new_n6429, new_n6434);
xnor_4 g04086(new_n6296, new_n6267, new_n6435);
not_8  g04087(new_n6435, new_n6436);
xnor_4 g04088(new_n6399, new_n6377, new_n6437_1);
nand_5 g04089(new_n6437_1, new_n6436, new_n6438);
xnor_4 g04090(new_n6437_1, new_n6435, new_n6439);
xnor_4 g04091(new_n6294, new_n6273, new_n6440);
xnor_4 g04092(new_n6396, new_n6381_1, new_n6441);
nor_5  g04093(new_n6441, new_n6440, new_n6442);
not_8  g04094(new_n6442, new_n6443);
not_8  g04095(new_n6441, new_n6444);
xnor_4 g04096(new_n6444, new_n6440, new_n6445);
xnor_4 g04097(new_n6292, new_n6279, new_n6446);
xnor_4 g04098(new_n6393, new_n6392, new_n6447);
not_8  g04099(new_n6447, new_n6448);
nor_5  g04100(new_n6448, new_n6446, new_n6449);
not_8  g04101(new_n6449, new_n6450);
xnor_4 g04102(new_n6447, new_n6446, new_n6451);
xnor_4 g04103(new_n6389, new_n6388, new_n6452);
not_8  g04104(new_n6286, new_n6453);
xnor_4 g04105(new_n6290, new_n6453, new_n6454);
nor_5  g04106(new_n6454, new_n6452, new_n6455);
xnor_4 g04107(new_n6282, n20658, new_n6456_1);
nor_5  g04108(new_n6456_1, new_n6110, new_n6457_1);
not_8  g04109(new_n6457_1, new_n6458);
xnor_4 g04110(new_n6454, new_n6452, new_n6459);
nor_5  g04111(new_n6459, new_n6458, new_n6460);
nor_5  g04112(new_n6460, new_n6455, new_n6461);
nand_5 g04113(new_n6461, new_n6451, new_n6462);
nand_5 g04114(new_n6462, new_n6450, new_n6463);
nand_5 g04115(new_n6463, new_n6445, new_n6464);
nand_5 g04116(new_n6464, new_n6443, new_n6465_1);
nand_5 g04117(new_n6465_1, new_n6439, new_n6466);
nand_5 g04118(new_n6466, new_n6438, new_n6467);
nand_5 g04119(new_n6467, new_n6434, new_n6468);
nand_5 g04120(new_n6468, new_n6433, new_n6469);
nand_5 g04121(new_n6469, new_n6427_1, new_n6470_1);
nand_5 g04122(new_n6470_1, new_n6426, new_n6471);
nand_5 g04123(new_n6471, new_n6422, new_n6472);
nand_5 g04124(new_n6472, new_n6421, new_n6473);
nand_5 g04125(new_n6473, new_n6417, new_n6474);
nand_5 g04126(new_n6474, new_n6416, new_n6475);
xnor_4 g04127(new_n6475, new_n6411, n567);
or_5   g04128(n10250, n1831, new_n6477);
not_8  g04129(n1831, new_n6478);
xnor_4 g04130(n10250, new_n6478, new_n6479);
or_5   g04131(n13137, n7674, new_n6480);
not_8  g04132(n7674, new_n6481);
xnor_4 g04133(n13137, new_n6481, new_n6482);
or_5   g04134(n18452, n6397, new_n6483);
not_8  g04135(n6397, new_n6484);
xnor_4 g04136(n18452, new_n6484, new_n6485_1);
nor_5  g04137(n21317, n19196, new_n6486);
not_8  g04138(n19196, new_n6487);
xnor_4 g04139(n21317, new_n6487, new_n6488);
not_8  g04140(new_n6488, new_n6489);
nor_5  g04141(n23586, n12398, new_n6490);
xnor_4 g04142(n23586, new_n4169, new_n6491);
not_8  g04143(new_n6491, new_n6492);
nor_5  g04144(n21226, n19789, new_n6493);
xnor_4 g04145(n21226, new_n4170, new_n6494);
not_8  g04146(new_n6494, new_n6495);
nor_5  g04147(n20169, n4426, new_n6496);
not_8  g04148(n4426, new_n6497);
xnor_4 g04149(n20169, new_n6497, new_n6498);
not_8  g04150(new_n6498, new_n6499);
nor_5  g04151(n20036, n8285, new_n6500);
xnor_4 g04152(n20036, new_n4171, new_n6501);
not_8  g04153(new_n6501, new_n6502_1);
nor_5  g04154(n11192, n6729, new_n6503);
nand_5 g04155(n21687, n9380, new_n6504);
not_8  g04156(new_n6504, new_n6505);
xnor_4 g04157(n11192, n6729, new_n6506_1);
nor_5  g04158(new_n6506_1, new_n6505, new_n6507);
nor_5  g04159(new_n6507, new_n6503, new_n6508);
nor_5  g04160(new_n6508, new_n6502_1, new_n6509);
nor_5  g04161(new_n6509, new_n6500, new_n6510);
nor_5  g04162(new_n6510, new_n6499, new_n6511);
nor_5  g04163(new_n6511, new_n6496, new_n6512);
nor_5  g04164(new_n6512, new_n6495, new_n6513_1);
nor_5  g04165(new_n6513_1, new_n6493, new_n6514_1);
nor_5  g04166(new_n6514_1, new_n6492, new_n6515);
nor_5  g04167(new_n6515, new_n6490, new_n6516);
nor_5  g04168(new_n6516, new_n6489, new_n6517);
nor_5  g04169(new_n6517, new_n6486, new_n6518);
not_8  g04170(new_n6518, new_n6519);
nand_5 g04171(new_n6519, new_n6485_1, new_n6520);
nand_5 g04172(new_n6520, new_n6483, new_n6521);
nand_5 g04173(new_n6521, new_n6482, new_n6522);
nand_5 g04174(new_n6522, new_n6480, new_n6523);
nand_5 g04175(new_n6523, new_n6479, new_n6524);
nand_5 g04176(new_n6524, new_n6477, new_n6525);
not_8  g04177(n8614, new_n6526);
not_8  g04178(n1288, new_n6527);
not_8  g04179(n13110, new_n6528);
nor_5  g04180(new_n4182, n25694, new_n6529);
nand_5 g04181(new_n6529, new_n6528, new_n6530);
nor_5  g04182(new_n6530, n1752, new_n6531);
nand_5 g04183(new_n6531, new_n6527, new_n6532);
xnor_4 g04184(new_n6532, n3320, new_n6533);
nor_5  g04185(new_n6533, new_n6526, new_n6534);
nor_5  g04186(new_n6532, n3320, new_n6535);
not_8  g04187(new_n6535, new_n6536);
not_8  g04188(new_n6533, new_n6537);
nor_5  g04189(new_n6537, n8614, new_n6538);
not_8  g04190(new_n6538, new_n6539);
xnor_4 g04191(new_n6531, n1288, new_n6540);
nor_5  g04192(new_n6540, n15182, new_n6541);
not_8  g04193(n15182, new_n6542_1);
xnor_4 g04194(new_n6540, new_n6542_1, new_n6543);
not_8  g04195(new_n6543, new_n6544);
not_8  g04196(n1752, new_n6545);
xnor_4 g04197(new_n6530, new_n6545, new_n6546);
nor_5  g04198(new_n6546, n27037, new_n6547);
not_8  g04199(new_n6546, new_n6548);
xnor_4 g04200(new_n6548, n27037, new_n6549);
not_8  g04201(new_n6549, new_n6550);
not_8  g04202(n8964, new_n6551);
xnor_4 g04203(new_n6529, n13110, new_n6552);
not_8  g04204(new_n6552, new_n6553);
nor_5  g04205(new_n6553, new_n6551, new_n6554);
not_8  g04206(new_n6554, new_n6555);
xnor_4 g04207(new_n6552, new_n6551, new_n6556_1);
not_8  g04208(n20151, new_n6557);
nor_5  g04209(new_n4183, new_n6557, new_n6558_1);
not_8  g04210(new_n6558_1, new_n6559);
nand_5 g04211(new_n4216, new_n4184, new_n6560_1);
nand_5 g04212(new_n6560_1, new_n6559, new_n6561);
nand_5 g04213(new_n6561, new_n6556_1, new_n6562);
nand_5 g04214(new_n6562, new_n6555, new_n6563);
nor_5  g04215(new_n6563, new_n6550, new_n6564);
nor_5  g04216(new_n6564, new_n6547, new_n6565);
nor_5  g04217(new_n6565, new_n6544, new_n6566);
nor_5  g04218(new_n6566, new_n6541, new_n6567_1);
nand_5 g04219(new_n6567_1, new_n6539, new_n6568);
nand_5 g04220(new_n6568, new_n6536, new_n6569);
nor_5  g04221(new_n6569, new_n6534, new_n6570);
not_8  g04222(new_n6570, new_n6571);
nand_5 g04223(new_n6571, new_n6525, new_n6572);
xnor_4 g04224(new_n6570, new_n6525, new_n6573);
xnor_4 g04225(new_n6523, new_n6479, new_n6574);
not_8  g04226(new_n6574, new_n6575);
xnor_4 g04227(new_n6533, n8614, new_n6576_1);
xnor_4 g04228(new_n6576_1, new_n6567_1, new_n6577);
nor_5  g04229(new_n6577, new_n6575, new_n6578);
xnor_4 g04230(new_n6565, new_n6544, new_n6579);
not_8  g04231(new_n6579, new_n6580);
xnor_4 g04232(new_n6521, new_n6482, new_n6581);
not_8  g04233(new_n6581, new_n6582);
nand_5 g04234(new_n6582, new_n6580, new_n6583);
xnor_4 g04235(new_n6582, new_n6579, new_n6584);
xnor_4 g04236(new_n6563, new_n6550, new_n6585);
not_8  g04237(new_n6585, new_n6586);
xnor_4 g04238(new_n6518, new_n6485_1, new_n6587_1);
nand_5 g04239(new_n6587_1, new_n6586, new_n6588);
xnor_4 g04240(new_n6587_1, new_n6585, new_n6589);
xnor_4 g04241(new_n6516, new_n6488, new_n6590_1);
xnor_4 g04242(new_n6561, new_n6556_1, new_n6591);
nor_5  g04243(new_n6591, new_n6590_1, new_n6592);
xnor_4 g04244(new_n6514_1, new_n6491, new_n6593);
nand_5 g04245(new_n6593, new_n4217, new_n6594);
not_8  g04246(new_n6593, new_n6595);
xnor_4 g04247(new_n6595, new_n4217, new_n6596_1);
xnor_4 g04248(new_n6512, new_n6494, new_n6597);
xnor_4 g04249(new_n6510, new_n6498, new_n6598);
not_8  g04250(new_n6598, new_n6599);
nor_5  g04251(new_n6599, new_n4226, new_n6600);
xnor_4 g04252(new_n6508, new_n6501, new_n6601);
nor_5  g04253(new_n6601, new_n4232, new_n6602);
not_8  g04254(new_n6602, new_n6603);
xnor_4 g04255(new_n6601, new_n4231_1, new_n6604);
xnor_4 g04256(new_n6506_1, new_n6504, new_n6605);
not_8  g04257(new_n6605, new_n6606);
nand_5 g04258(new_n6606, new_n4241, new_n6607);
xnor_4 g04259(n21687, new_n4307, new_n6608);
not_8  g04260(new_n6608, new_n6609);
nor_5  g04261(new_n6609, new_n4245, new_n6610);
xnor_4 g04262(new_n6605, new_n4241, new_n6611_1);
nand_5 g04263(new_n6611_1, new_n6610, new_n6612_1);
nand_5 g04264(new_n6612_1, new_n6607, new_n6613);
nand_5 g04265(new_n6613, new_n6604, new_n6614);
nand_5 g04266(new_n6614, new_n6603, new_n6615);
xnor_4 g04267(new_n6599, new_n4226, new_n6616);
nor_5  g04268(new_n6616, new_n6615, new_n6617);
nor_5  g04269(new_n6617, new_n6600, new_n6618);
not_8  g04270(new_n6618, new_n6619);
nand_5 g04271(new_n6619, new_n6597, new_n6620);
xnor_4 g04272(new_n6618, new_n6597, new_n6621);
nand_5 g04273(new_n6621, new_n4222, new_n6622);
nand_5 g04274(new_n6622, new_n6620, new_n6623);
nand_5 g04275(new_n6623, new_n6596_1, new_n6624);
nand_5 g04276(new_n6624, new_n6594, new_n6625);
xnor_4 g04277(new_n6591, new_n6590_1, new_n6626);
nor_5  g04278(new_n6626, new_n6625, new_n6627);
nor_5  g04279(new_n6627, new_n6592, new_n6628_1);
nand_5 g04280(new_n6628_1, new_n6589, new_n6629);
nand_5 g04281(new_n6629, new_n6588, new_n6630_1);
nand_5 g04282(new_n6630_1, new_n6584, new_n6631_1);
nand_5 g04283(new_n6631_1, new_n6583, new_n6632);
xnor_4 g04284(new_n6577, new_n6575, new_n6633);
nor_5  g04285(new_n6633, new_n6632, new_n6634_1);
nor_5  g04286(new_n6634_1, new_n6578, new_n6635);
nand_5 g04287(new_n6635, new_n6573, new_n6636);
nand_5 g04288(new_n6636, new_n6572, new_n6637);
xnor_4 g04289(new_n6635, new_n6573, new_n6638);
not_8  g04290(new_n6638, new_n6639);
or_5   g04291(n15766, n6105, new_n6640);
not_8  g04292(n6105, new_n6641);
xnor_4 g04293(n15766, new_n6641, new_n6642);
nor_5  g04294(n25629, n3795, new_n6643);
not_8  g04295(new_n6643, new_n6644);
not_8  g04296(n3795, new_n6645);
xnor_4 g04297(n25629, new_n6645, new_n6646);
nor_5  g04298(n25464, n7692, new_n6647);
not_8  g04299(n7692, new_n6648);
xnor_4 g04300(n25464, new_n6648, new_n6649);
not_8  g04301(new_n6649, new_n6650);
nor_5  g04302(n23039, n4590, new_n6651);
not_8  g04303(n4590, new_n6652_1);
xnor_4 g04304(n23039, new_n6652_1, new_n6653);
not_8  g04305(new_n6653, new_n6654);
nor_5  g04306(n26752, n13677, new_n6655_1);
xnor_4 g04307(n26752, new_n4095, new_n6656);
not_8  g04308(new_n6656, new_n6657);
nor_5  g04309(n18926, n6513, new_n6658);
not_8  g04310(n6513, new_n6659_1);
xnor_4 g04311(n18926, new_n6659_1, new_n6660);
not_8  g04312(new_n6660, new_n6661);
not_8  g04313(n3918, new_n6662);
or_5   g04314(new_n4138, new_n6662, new_n6663);
nor_5  g04315(n5451, n3918, new_n6664);
not_8  g04316(new_n6664, new_n6665);
nor_5  g04317(n5330, n919, new_n6666);
not_8  g04318(new_n4328, new_n6667);
nor_5  g04319(new_n4333, new_n6667, new_n6668);
nor_5  g04320(new_n6668, new_n6666, new_n6669_1);
nand_5 g04321(new_n6669_1, new_n6665, new_n6670);
nand_5 g04322(new_n6670, new_n6663, new_n6671_1);
nor_5  g04323(new_n6671_1, new_n6661, new_n6672);
nor_5  g04324(new_n6672, new_n6658, new_n6673_1);
nor_5  g04325(new_n6673_1, new_n6657, new_n6674_1);
nor_5  g04326(new_n6674_1, new_n6655_1, new_n6675);
nor_5  g04327(new_n6675, new_n6654, new_n6676);
nor_5  g04328(new_n6676, new_n6651, new_n6677);
nor_5  g04329(new_n6677, new_n6650, new_n6678);
nor_5  g04330(new_n6678, new_n6647, new_n6679);
not_8  g04331(new_n6679, new_n6680);
nand_5 g04332(new_n6680, new_n6646, new_n6681);
nand_5 g04333(new_n6681, new_n6644, new_n6682);
nand_5 g04334(new_n6682, new_n6642, new_n6683);
nand_5 g04335(new_n6683, new_n6640, new_n6684_1);
not_8  g04336(new_n6684_1, new_n6685);
nand_5 g04337(new_n6685, new_n6639, new_n6686);
xnor_4 g04338(new_n6685, new_n6638, new_n6687);
xnor_4 g04339(new_n6682, new_n6642, new_n6688);
not_8  g04340(new_n6633, new_n6689);
xnor_4 g04341(new_n6689, new_n6632, new_n6690);
not_8  g04342(new_n6690, new_n6691_1);
nand_5 g04343(new_n6691_1, new_n6688, new_n6692);
xnor_4 g04344(new_n6690, new_n6688, new_n6693);
xnor_4 g04345(new_n6630_1, new_n6584, new_n6694);
not_8  g04346(new_n6694, new_n6695);
xnor_4 g04347(new_n6679, new_n6646, new_n6696);
not_8  g04348(new_n6696, new_n6697);
nand_5 g04349(new_n6697, new_n6695, new_n6698);
xnor_4 g04350(new_n6696, new_n6695, new_n6699);
xnor_4 g04351(new_n6628_1, new_n6589, new_n6700);
not_8  g04352(new_n6700, new_n6701);
xnor_4 g04353(new_n6677, new_n6649, new_n6702);
not_8  g04354(new_n6702, new_n6703);
nand_5 g04355(new_n6703, new_n6701, new_n6704);
xnor_4 g04356(new_n6702, new_n6701, new_n6705);
xnor_4 g04357(new_n6675, new_n6653, new_n6706_1);
not_8  g04358(new_n6706_1, new_n6707_1);
xnor_4 g04359(new_n6626, new_n6625, new_n6708);
nand_5 g04360(new_n6708, new_n6707_1, new_n6709);
xnor_4 g04361(new_n6708, new_n6706_1, new_n6710);
not_8  g04362(new_n6596_1, new_n6711);
xnor_4 g04363(new_n6623, new_n6711, new_n6712);
xnor_4 g04364(new_n6673_1, new_n6656, new_n6713);
not_8  g04365(new_n6713, new_n6714);
nand_5 g04366(new_n6714, new_n6712, new_n6715);
xnor_4 g04367(new_n6713, new_n6712, new_n6716);
xnor_4 g04368(new_n6621, new_n4222, new_n6717);
not_8  g04369(new_n6717, new_n6718);
xnor_4 g04370(new_n6671_1, new_n6661, new_n6719);
nand_5 g04371(new_n6719, new_n6718, new_n6720);
xnor_4 g04372(new_n6719, new_n6717, new_n6721);
xnor_4 g04373(new_n6616, new_n6615, new_n6722);
xnor_4 g04374(n5451, new_n6662, new_n6723);
xnor_4 g04375(new_n6723, new_n6669_1, new_n6724);
nor_5  g04376(new_n6724, new_n6722, new_n6725);
not_8  g04377(new_n6725, new_n6726);
not_8  g04378(new_n6724, new_n6727);
xnor_4 g04379(new_n6727, new_n6722, new_n6728);
xnor_4 g04380(new_n6613, new_n6604, new_n6729_1);
not_8  g04381(new_n6729_1, new_n6730);
nor_5  g04382(new_n6730, new_n4334, new_n6731);
not_8  g04383(new_n6731, new_n6732);
xnor_4 g04384(new_n6729_1, new_n4334, new_n6733);
xnor_4 g04385(new_n6611_1, new_n6610, new_n6734);
nand_5 g04386(new_n6734, new_n4340_1, new_n6735);
xnor_4 g04387(new_n6608, new_n2576, new_n6736_1);
nand_5 g04388(new_n6736_1, new_n4343, new_n6737);
xnor_4 g04389(new_n6734, new_n4339, new_n6738);
not_8  g04390(new_n6738, new_n6739);
nor_5  g04391(new_n6739, new_n6737, new_n6740);
not_8  g04392(new_n6740, new_n6741);
nand_5 g04393(new_n6741, new_n6735, new_n6742);
nand_5 g04394(new_n6742, new_n6733, new_n6743);
nand_5 g04395(new_n6743, new_n6732, new_n6744);
nand_5 g04396(new_n6744, new_n6728, new_n6745);
nand_5 g04397(new_n6745, new_n6726, new_n6746);
nand_5 g04398(new_n6746, new_n6721, new_n6747);
nand_5 g04399(new_n6747, new_n6720, new_n6748);
nand_5 g04400(new_n6748, new_n6716, new_n6749);
nand_5 g04401(new_n6749, new_n6715, new_n6750);
nand_5 g04402(new_n6750, new_n6710, new_n6751);
nand_5 g04403(new_n6751, new_n6709, new_n6752);
nand_5 g04404(new_n6752, new_n6705, new_n6753);
nand_5 g04405(new_n6753, new_n6704, new_n6754);
nand_5 g04406(new_n6754, new_n6699, new_n6755);
nand_5 g04407(new_n6755, new_n6698, new_n6756);
nand_5 g04408(new_n6756, new_n6693, new_n6757);
nand_5 g04409(new_n6757, new_n6692, new_n6758);
nand_5 g04410(new_n6758, new_n6687, new_n6759);
nand_5 g04411(new_n6759, new_n6686, new_n6760);
nand_5 g04412(new_n6760, new_n6637, new_n6761);
not_8  g04413(new_n6761, n588);
xnor_4 g04414(n19803, n18584, new_n6763);
not_8  g04415(n12626, new_n6764);
or_5   g04416(new_n6764, n4272, new_n6765);
not_8  g04417(new_n4902, new_n6766);
nand_5 g04418(new_n6766, new_n4876, new_n6767);
nand_5 g04419(new_n6767, new_n6765, new_n6768);
xnor_4 g04420(new_n6768, new_n6763, new_n6769);
not_8  g04421(new_n6769, new_n6770);
xnor_4 g04422(n16911, n7773, new_n6771);
not_8  g04423(n7721, new_n6772);
nand_5 g04424(new_n6772, n376, new_n6773_1);
xnor_4 g04425(n7721, n376, new_n6774);
not_8  g04426(n5517, new_n6775_1);
nor_5  g04427(n21981, new_n6775_1, new_n6776);
xnor_4 g04428(n21981, n5517, new_n6777);
not_8  g04429(new_n6777, new_n6778);
not_8  g04430(n12113, new_n6779);
nor_5  g04431(n12917, new_n6779, new_n6780);
xnor_4 g04432(n12917, n12113, new_n6781);
not_8  g04433(n21898, new_n6782);
nor_5  g04434(new_n6782, n10614, new_n6783);
not_8  g04435(n10614, new_n6784);
nor_5  g04436(n21898, new_n6784, new_n6785_1);
not_8  g04437(n9926, new_n6786);
nor_5  g04438(n11266, new_n6786, new_n6787);
nand_5 g04439(n11266, new_n6786, new_n6788);
not_8  g04440(new_n6788, new_n6789);
not_8  g04441(n2646, new_n6790_1);
nand_5 g04442(n22072, new_n6790_1, new_n6791_1);
nor_5  g04443(new_n6791_1, new_n6789, new_n6792);
nor_5  g04444(new_n6792, new_n6787, new_n6793);
nor_5  g04445(new_n6793, new_n6785_1, new_n6794_1);
nor_5  g04446(new_n6794_1, new_n6783, new_n6795);
nand_5 g04447(new_n6795, new_n6781, new_n6796);
not_8  g04448(new_n6796, new_n6797);
nor_5  g04449(new_n6797, new_n6780, new_n6798);
nor_5  g04450(new_n6798, new_n6778, new_n6799);
nor_5  g04451(new_n6799, new_n6776, new_n6800);
not_8  g04452(new_n6800, new_n6801);
nand_5 g04453(new_n6801, new_n6774, new_n6802_1);
nand_5 g04454(new_n6802_1, new_n6773_1, new_n6803);
xnor_4 g04455(new_n6803, new_n6771, new_n6804);
not_8  g04456(n1742, new_n6805);
not_8  g04457(n14576, new_n6806);
not_8  g04458(n5605, new_n6807);
nor_5  g04459(n15652, n4939, new_n6808);
nand_5 g04460(new_n6808, new_n6807, new_n6809);
nor_5  g04461(new_n6809, n2985, new_n6810);
nand_5 g04462(new_n6810, new_n6806, new_n6811);
nor_5  g04463(new_n6811, n1269, new_n6812);
xnor_4 g04464(new_n6812, n16818, new_n6813);
xnor_4 g04465(new_n6813, new_n6805, new_n6814_1);
not_8  g04466(n4858, new_n6815);
not_8  g04467(n1269, new_n6816);
xnor_4 g04468(new_n6811, new_n6816, new_n6817);
not_8  g04469(new_n6817, new_n6818);
nand_5 g04470(new_n6818, new_n6815, new_n6819);
xnor_4 g04471(new_n6817, new_n6815, new_n6820);
not_8  g04472(n8244, new_n6821);
xnor_4 g04473(new_n6810, n14576, new_n6822);
not_8  g04474(new_n6822, new_n6823);
nand_5 g04475(new_n6823, new_n6821, new_n6824);
xnor_4 g04476(new_n6822, new_n6821, new_n6825);
not_8  g04477(n9493, new_n6826_1);
not_8  g04478(n2985, new_n6827);
xnor_4 g04479(new_n6809, new_n6827, new_n6828);
not_8  g04480(new_n6828, new_n6829);
nand_5 g04481(new_n6829, new_n6826_1, new_n6830);
not_8  g04482(n15167, new_n6831);
xnor_4 g04483(new_n6808, n5605, new_n6832);
not_8  g04484(new_n6832, new_n6833);
nand_5 g04485(new_n6833, new_n6831, new_n6834);
xnor_4 g04486(new_n6832, new_n6831, new_n6835_1);
not_8  g04487(n21095, new_n6836);
xnor_4 g04488(n15652, n4939, new_n6837);
nand_5 g04489(new_n6837, new_n6836, new_n6838);
nand_5 g04490(n8656, n4939, new_n6839);
xnor_4 g04491(new_n6837, n21095, new_n6840);
nand_5 g04492(new_n6840, new_n6839, new_n6841);
nand_5 g04493(new_n6841, new_n6838, new_n6842);
nand_5 g04494(new_n6842, new_n6835_1, new_n6843);
nand_5 g04495(new_n6843, new_n6834, new_n6844);
xnor_4 g04496(new_n6828, new_n6826_1, new_n6845);
nand_5 g04497(new_n6845, new_n6844, new_n6846);
nand_5 g04498(new_n6846, new_n6830, new_n6847);
nand_5 g04499(new_n6847, new_n6825, new_n6848);
nand_5 g04500(new_n6848, new_n6824, new_n6849);
nand_5 g04501(new_n6849, new_n6820, new_n6850);
nand_5 g04502(new_n6850, new_n6819, new_n6851);
xnor_4 g04503(new_n6851, new_n6814_1, new_n6852);
xnor_4 g04504(new_n6852, new_n6804, new_n6853_1);
xnor_4 g04505(new_n6800, new_n6774, new_n6854);
not_8  g04506(new_n6854, new_n6855);
not_8  g04507(new_n6820, new_n6856);
xnor_4 g04508(new_n6849, new_n6856, new_n6857);
nor_5  g04509(new_n6857, new_n6855, new_n6858);
not_8  g04510(new_n6858, new_n6859);
xnor_4 g04511(new_n6857, new_n6854, new_n6860);
xnor_4 g04512(new_n6798, new_n6777, new_n6861_1);
xnor_4 g04513(new_n6847, new_n6825, new_n6862_1);
nor_5  g04514(new_n6862_1, new_n6861_1, new_n6863_1);
xnor_4 g04515(new_n6862_1, new_n6861_1, new_n6864);
not_8  g04516(new_n6795, new_n6865);
xnor_4 g04517(new_n6865, new_n6781, new_n6866);
not_8  g04518(new_n6866, new_n6867_1);
not_8  g04519(new_n6845, new_n6868);
xnor_4 g04520(new_n6868, new_n6844, new_n6869);
nor_5  g04521(new_n6869, new_n6867_1, new_n6870);
not_8  g04522(new_n6870, new_n6871);
xnor_4 g04523(new_n6842, new_n6835_1, new_n6872);
not_8  g04524(new_n6793, new_n6873);
xnor_4 g04525(n21898, n10614, new_n6874);
xnor_4 g04526(new_n6874, new_n6873, new_n6875);
nor_5  g04527(new_n6875, new_n6872, new_n6876);
not_8  g04528(new_n6875, new_n6877);
xnor_4 g04529(new_n6877, new_n6872, new_n6878);
not_8  g04530(new_n6878, new_n6879);
not_8  g04531(n4939, new_n6880);
xnor_4 g04532(n8656, new_n6880, new_n6881);
not_8  g04533(new_n6881, new_n6882);
xnor_4 g04534(n22072, n2646, new_n6883);
nor_5  g04535(new_n6883, new_n6882, new_n6884);
xnor_4 g04536(n11266, n9926, new_n6885);
xnor_4 g04537(new_n6885, new_n6791_1, new_n6886);
not_8  g04538(new_n6886, new_n6887);
nor_5  g04539(new_n6887, new_n6884, new_n6888);
xnor_4 g04540(new_n6840, new_n6839, new_n6889);
xnor_4 g04541(new_n6887, new_n6884, new_n6890);
nor_5  g04542(new_n6890, new_n6889, new_n6891);
nor_5  g04543(new_n6891, new_n6888, new_n6892);
nor_5  g04544(new_n6892, new_n6879, new_n6893);
nor_5  g04545(new_n6893, new_n6876, new_n6894);
xnor_4 g04546(new_n6869, new_n6866, new_n6895);
nand_5 g04547(new_n6895, new_n6894, new_n6896);
nand_5 g04548(new_n6896, new_n6871, new_n6897);
nor_5  g04549(new_n6897, new_n6864, new_n6898);
nor_5  g04550(new_n6898, new_n6863_1, new_n6899);
nand_5 g04551(new_n6899, new_n6860, new_n6900);
nand_5 g04552(new_n6900, new_n6859, new_n6901);
xnor_4 g04553(new_n6901, new_n6853_1, new_n6902);
xnor_4 g04554(new_n6902, new_n6770, new_n6903);
xnor_4 g04555(new_n6899, new_n6860, new_n6904);
nand_5 g04556(new_n6904, new_n4904, new_n6905);
xnor_4 g04557(new_n6904, new_n4903, new_n6906);
xnor_4 g04558(new_n6897, new_n6864, new_n6907);
not_8  g04559(new_n6907, new_n6908);
nand_5 g04560(new_n6908, new_n4909, new_n6909);
xnor_4 g04561(new_n6907, new_n4909, new_n6910);
not_8  g04562(new_n6894, new_n6911);
xnor_4 g04563(new_n6895, new_n6911, new_n6912);
not_8  g04564(new_n6912, new_n6913);
nand_5 g04565(new_n6913, new_n4915, new_n6914);
xnor_4 g04566(new_n6912, new_n4915, new_n6915);
xnor_4 g04567(new_n6892, new_n6878, new_n6916);
not_8  g04568(new_n6916, new_n6917);
nor_5  g04569(new_n6917, new_n4925_1, new_n6918);
xnor_4 g04570(new_n6916, new_n4925_1, new_n6919);
not_8  g04571(new_n6919, new_n6920);
xnor_4 g04572(new_n6883, new_n6881, new_n6921);
not_8  g04573(new_n6921, new_n6922);
nor_5  g04574(new_n6922, new_n4935, new_n6923);
nor_5  g04575(new_n6923, new_n4937, new_n6924);
xnor_4 g04576(new_n6890, new_n6889, new_n6925);
xnor_4 g04577(new_n6923, new_n4932, new_n6926);
not_8  g04578(new_n6926, new_n6927);
nor_5  g04579(new_n6927, new_n6925, new_n6928);
nor_5  g04580(new_n6928, new_n6924, new_n6929);
nor_5  g04581(new_n6929, new_n6920, new_n6930);
nor_5  g04582(new_n6930, new_n6918, new_n6931);
not_8  g04583(new_n6931, new_n6932);
nand_5 g04584(new_n6932, new_n6915, new_n6933);
nand_5 g04585(new_n6933, new_n6914, new_n6934);
nand_5 g04586(new_n6934, new_n6910, new_n6935);
nand_5 g04587(new_n6935, new_n6909, new_n6936);
nand_5 g04588(new_n6936, new_n6906, new_n6937);
nand_5 g04589(new_n6937, new_n6905, new_n6938);
xnor_4 g04590(new_n6938, new_n6903, n597);
not_8  g04591(n14230, new_n6940);
xnor_4 g04592(n25926, n9646, new_n6941);
xnor_4 g04593(new_n6941, new_n6940, new_n6942);
xnor_4 g04594(new_n6942, new_n6117, n637);
not_8  g04595(n10611, new_n6944);
xnor_4 g04596(n25797, new_n6944, new_n6945);
nor_5  g04597(n15967, n2783, new_n6946);
not_8  g04598(n2783, new_n6947);
xnor_4 g04599(n15967, new_n6947, new_n6948);
not_8  g04600(new_n6948, new_n6949);
nor_5  g04601(n15490, n13319, new_n6950);
nand_5 g04602(n25435, n18, new_n6951);
not_8  g04603(new_n6951, new_n6952);
xnor_4 g04604(n15490, n13319, new_n6953);
nor_5  g04605(new_n6953, new_n6952, new_n6954);
nor_5  g04606(new_n6954, new_n6950, new_n6955);
nor_5  g04607(new_n6955, new_n6949, new_n6956);
nor_5  g04608(new_n6956, new_n6946, new_n6957);
xnor_4 g04609(new_n6957, new_n6945, new_n6958);
xnor_4 g04610(new_n6958, n7421, new_n6959);
not_8  g04611(n19680, new_n6960);
xnor_4 g04612(new_n6955, new_n6948, new_n6961);
nor_5  g04613(new_n6961, new_n6960, new_n6962);
xnor_4 g04614(new_n6961, n19680, new_n6963);
xnor_4 g04615(new_n6953, new_n6951, new_n6964);
not_8  g04616(new_n6964, new_n6965_1);
nor_5  g04617(new_n6965_1, n2809, new_n6966);
not_8  g04618(n18, new_n6967_1);
xnor_4 g04619(n25435, new_n6967_1, new_n6968);
not_8  g04620(new_n6968, new_n6969);
nor_5  g04621(new_n6969, new_n5125, new_n6970);
xnor_4 g04622(new_n6964, n2809, new_n6971_1);
not_8  g04623(new_n6971_1, new_n6972);
nor_5  g04624(new_n6972, new_n6970, new_n6973);
nor_5  g04625(new_n6973, new_n6966, new_n6974);
nand_5 g04626(new_n6974, new_n6963, new_n6975_1);
not_8  g04627(new_n6975_1, new_n6976);
nor_5  g04628(new_n6976, new_n6962, new_n6977);
xnor_4 g04629(new_n6977, new_n6959, new_n6978);
not_8  g04630(n11056, new_n6979);
xnor_4 g04631(n18157, new_n6979, new_n6980);
nor_5  g04632(n15271, n12161, new_n6981);
not_8  g04633(n12161, new_n6982);
xnor_4 g04634(n15271, new_n6982, new_n6983_1);
not_8  g04635(new_n6983_1, new_n6984);
nor_5  g04636(n25877, n5026, new_n6985_1);
nand_5 g04637(n24323, n8581, new_n6986);
not_8  g04638(new_n6986, new_n6987);
xnor_4 g04639(n25877, n5026, new_n6988);
nor_5  g04640(new_n6988, new_n6987, new_n6989);
nor_5  g04641(new_n6989, new_n6985_1, new_n6990);
nor_5  g04642(new_n6990, new_n6984, new_n6991);
nor_5  g04643(new_n6991, new_n6981, new_n6992);
xnor_4 g04644(new_n6992, new_n6980, new_n6993);
xnor_4 g04645(new_n6993, n20250, new_n6994);
xnor_4 g04646(new_n6990, new_n6983_1, new_n6995);
nand_5 g04647(new_n6995, new_n4577, new_n6996);
not_8  g04648(new_n6996, new_n6997);
not_8  g04649(n26443, new_n6998_1);
xnor_4 g04650(new_n6988, new_n6986, new_n6999);
nand_5 g04651(new_n6999, new_n6998_1, new_n7000);
not_8  g04652(new_n7000, new_n7001);
xnor_4 g04653(n24323, n8581, new_n7002);
nor_5  g04654(new_n7002, new_n2568, new_n7003);
xnor_4 g04655(new_n6999, new_n6998_1, new_n7004);
nor_5  g04656(new_n7004, new_n7003, new_n7005);
nor_5  g04657(new_n7005, new_n7001, new_n7006);
xnor_4 g04658(new_n6995, n5822, new_n7007);
not_8  g04659(new_n7007, new_n7008);
nor_5  g04660(new_n7008, new_n7006, new_n7009);
nor_5  g04661(new_n7009, new_n6997, new_n7010);
xnor_4 g04662(new_n7010, new_n6994, new_n7011);
not_8  g04663(new_n7011, new_n7012);
xnor_4 g04664(new_n7012, new_n6978, new_n7013);
xnor_4 g04665(new_n6974, new_n6963, new_n7014);
not_8  g04666(new_n7014, new_n7015);
xnor_4 g04667(new_n7007, new_n7006, new_n7016);
nor_5  g04668(new_n7016, new_n7015, new_n7017);
xnor_4 g04669(new_n7016, new_n7014, new_n7018);
not_8  g04670(new_n7018, new_n7019);
xnor_4 g04671(new_n6971_1, new_n6970, new_n7020);
xnor_4 g04672(new_n7004, new_n7003, new_n7021);
nor_5  g04673(new_n7021, new_n7020, new_n7022);
xnor_4 g04674(new_n6968, n15508, new_n7023);
xnor_4 g04675(new_n7002, n1681, new_n7024);
nor_5  g04676(new_n7024, new_n7023, new_n7025);
not_8  g04677(new_n7025, new_n7026_1);
not_8  g04678(new_n7020, new_n7027);
xnor_4 g04679(new_n7021, new_n7027, new_n7028);
not_8  g04680(new_n7028, new_n7029);
nor_5  g04681(new_n7029, new_n7026_1, new_n7030);
nor_5  g04682(new_n7030, new_n7022, new_n7031);
not_8  g04683(new_n7031, new_n7032_1);
nor_5  g04684(new_n7032_1, new_n7019, new_n7033);
nor_5  g04685(new_n7033, new_n7017, new_n7034);
xnor_4 g04686(new_n7034, new_n7013, n646);
nor_5  g04687(n19494, n2387, new_n7036);
nand_5 g04688(new_n7036, new_n2362, new_n7037);
nor_5  g04689(new_n7037, n26913, new_n7038_1);
xnor_4 g04690(new_n7038_1, n21832, new_n7039);
xnor_4 g04691(new_n2476, new_n5752_1, new_n7040);
nand_5 g04692(new_n2481, n7731, new_n7041);
xnor_4 g04693(new_n2481, new_n5755, new_n7042);
nand_5 g04694(new_n2485, n12341, new_n7043);
xnor_4 g04695(new_n2485, new_n5760, new_n7044);
nor_5  g04696(new_n2489, n12384, new_n7045);
not_8  g04697(new_n7045, new_n7046);
nor_5  g04698(new_n7046, n20986, new_n7047);
xnor_4 g04699(new_n7045, new_n5763, new_n7048);
nor_5  g04700(new_n7048, new_n2492, new_n7049);
nor_5  g04701(new_n7049, new_n7047, new_n7050);
nand_5 g04702(new_n7050, new_n7044, new_n7051);
nand_5 g04703(new_n7051, new_n7043, new_n7052);
nand_5 g04704(new_n7052, new_n7042, new_n7053);
nand_5 g04705(new_n7053, new_n7041, new_n7054);
xnor_4 g04706(new_n7054, new_n7040, new_n7055);
xnor_4 g04707(new_n7055, new_n7039, new_n7056);
not_8  g04708(new_n7056, new_n7057_1);
xnor_4 g04709(new_n7037, new_n2356, new_n7058);
xnor_4 g04710(new_n7052, new_n7042, new_n7059);
not_8  g04711(new_n7059, new_n7060);
nand_5 g04712(new_n7060, new_n7058, new_n7061);
xnor_4 g04713(new_n7059, new_n7058, new_n7062);
xnor_4 g04714(new_n2489, n12384, new_n7063);
nand_5 g04715(new_n7063, n2387, new_n7064);
nor_5  g04716(new_n7064, n19494, new_n7065);
not_8  g04717(new_n7065, new_n7066);
xnor_4 g04718(new_n7048, new_n2492, new_n7067);
not_8  g04719(n12384, new_n7068);
xnor_4 g04720(new_n2489, new_n7068, new_n7069);
nor_5  g04721(new_n7069, new_n2368, new_n7070);
xnor_4 g04722(n19494, new_n2368, new_n7071);
nor_5  g04723(new_n7071, new_n7070, new_n7072);
nor_5  g04724(new_n7072, new_n7065, new_n7073);
nand_5 g04725(new_n7073, new_n7067, new_n7074);
nand_5 g04726(new_n7074, new_n7066, new_n7075);
xnor_4 g04727(new_n7036, n16223, new_n7076);
nand_5 g04728(new_n7076, new_n7075, new_n7077);
not_8  g04729(new_n7044, new_n7078);
xnor_4 g04730(new_n7050, new_n7078, new_n7079_1);
not_8  g04731(new_n7076, new_n7080);
xnor_4 g04732(new_n7080, new_n7075, new_n7081);
nand_5 g04733(new_n7081, new_n7079_1, new_n7082);
nand_5 g04734(new_n7082, new_n7077, new_n7083);
nand_5 g04735(new_n7083, new_n7062, new_n7084);
nand_5 g04736(new_n7084, new_n7061, new_n7085);
xnor_4 g04737(new_n7085, new_n7057_1, new_n7086);
xnor_4 g04738(new_n7086, new_n3471, new_n7087);
not_8  g04739(new_n7062, new_n7088);
xnor_4 g04740(new_n7083, new_n7088, new_n7089);
not_8  g04741(new_n7089, new_n7090);
nand_5 g04742(new_n7090, new_n3478, new_n7091);
xnor_4 g04743(new_n7081, new_n7079_1, new_n7092);
nor_5  g04744(new_n7092, new_n3482, new_n7093);
xnor_4 g04745(new_n7092, new_n3482, new_n7094);
xnor_4 g04746(new_n7069, n2387, new_n7095);
not_8  g04747(new_n7095, new_n7096);
nor_5  g04748(new_n7096, new_n3488, new_n7097);
nor_5  g04749(new_n7097, new_n3493, new_n7098);
not_8  g04750(new_n7067, new_n7099_1);
xnor_4 g04751(new_n7073, new_n7099_1, new_n7100);
not_8  g04752(new_n7097, new_n7101);
nor_5  g04753(new_n7101, new_n3417, new_n7102);
nor_5  g04754(new_n7102, new_n7098, new_n7103);
not_8  g04755(new_n7103, new_n7104);
nor_5  g04756(new_n7104, new_n7100, new_n7105);
nor_5  g04757(new_n7105, new_n7098, new_n7106);
not_8  g04758(new_n7106, new_n7107);
nor_5  g04759(new_n7107, new_n7094, new_n7108);
nor_5  g04760(new_n7108, new_n7093, new_n7109);
xnor_4 g04761(new_n7089, new_n3478, new_n7110);
nand_5 g04762(new_n7110, new_n7109, new_n7111);
nand_5 g04763(new_n7111, new_n7091, new_n7112);
xnor_4 g04764(new_n7112, new_n7087, n696);
not_8  g04765(n23697, new_n7114);
xnor_4 g04766(n25475, new_n7114, new_n7115);
not_8  g04767(new_n7115, new_n7116);
or_5   g04768(n23849, n2289, new_n7117);
not_8  g04769(n2289, new_n7118);
xnor_4 g04770(n23849, new_n7118, new_n7119);
nor_5  g04771(n12446, n1112, new_n7120);
not_8  g04772(new_n7120, new_n7121);
not_8  g04773(n1112, new_n7122);
xnor_4 g04774(n12446, new_n7122, new_n7123);
nor_5  g04775(n20179, n11011, new_n7124);
not_8  g04776(new_n7124, new_n7125);
xnor_4 g04777(n20179, new_n4631, new_n7126);
nor_5  g04778(n19228, n16029, new_n7127);
not_8  g04779(new_n7127, new_n7128);
xnor_4 g04780(n19228, new_n4104, new_n7129);
nor_5  g04781(n16476, n15539, new_n7130);
not_8  g04782(new_n7130, new_n7131);
not_8  g04783(n15539, new_n7132);
xnor_4 g04784(n16476, new_n7132, new_n7133);
nor_5  g04785(n11615, n8052, new_n7134);
not_8  g04786(new_n7134, new_n7135);
not_8  g04787(n8052, new_n7136);
xnor_4 g04788(n11615, new_n7136, new_n7137);
nor_5  g04789(n22433, n10158, new_n7138);
not_8  g04790(new_n7138, new_n7139_1);
nand_5 g04791(n18962, n14090, new_n7140);
xnor_4 g04792(n22433, n10158, new_n7141);
not_8  g04793(new_n7141, new_n7142);
nand_5 g04794(new_n7142, new_n7140, new_n7143);
nand_5 g04795(new_n7143, new_n7139_1, new_n7144);
nand_5 g04796(new_n7144, new_n7137, new_n7145);
nand_5 g04797(new_n7145, new_n7135, new_n7146);
nand_5 g04798(new_n7146, new_n7133, new_n7147);
nand_5 g04799(new_n7147, new_n7131, new_n7148);
nand_5 g04800(new_n7148, new_n7129, new_n7149_1);
nand_5 g04801(new_n7149_1, new_n7128, new_n7150);
nand_5 g04802(new_n7150, new_n7126, new_n7151);
nand_5 g04803(new_n7151, new_n7125, new_n7152);
nand_5 g04804(new_n7152, new_n7123, new_n7153);
nand_5 g04805(new_n7153, new_n7121, new_n7154);
nand_5 g04806(new_n7154, new_n7119, new_n7155);
nand_5 g04807(new_n7155, new_n7117, new_n7156);
xnor_4 g04808(new_n7156, new_n7116, new_n7157);
xnor_4 g04809(new_n7157, n25345, new_n7158);
not_8  g04810(new_n7158, new_n7159);
xnor_4 g04811(new_n7154, new_n7119, new_n7160);
nand_5 g04812(new_n7160, n9655, new_n7161);
xnor_4 g04813(new_n7160, new_n5793, new_n7162);
not_8  g04814(new_n7123, new_n7163);
xnor_4 g04815(new_n7152, new_n7163, new_n7164);
not_8  g04816(new_n7164, new_n7165);
nand_5 g04817(new_n7165, n13490, new_n7166);
xnor_4 g04818(new_n7164, n13490, new_n7167);
not_8  g04819(new_n7126, new_n7168);
xnor_4 g04820(new_n7150, new_n7168, new_n7169);
nor_5  g04821(new_n7169, new_n2433, new_n7170);
xnor_4 g04822(new_n7148, new_n7129, new_n7171);
nor_5  g04823(new_n7171, n1777, new_n7172);
not_8  g04824(new_n7172, new_n7173);
xnor_4 g04825(new_n7171, new_n2437, new_n7174);
not_8  g04826(new_n7137, new_n7175);
not_8  g04827(new_n7140, new_n7176);
nor_5  g04828(new_n7141, new_n7176, new_n7177);
nor_5  g04829(new_n7177, new_n7138, new_n7178);
nor_5  g04830(new_n7178, new_n7175, new_n7179);
nor_5  g04831(new_n7179, new_n7134, new_n7180);
xnor_4 g04832(new_n7180, new_n7133, new_n7181);
not_8  g04833(new_n7181, new_n7182);
nor_5  g04834(new_n7182, n8745, new_n7183);
not_8  g04835(new_n7183, new_n7184);
xnor_4 g04836(new_n7181, n8745, new_n7185);
xnor_4 g04837(new_n7178, new_n7137, new_n7186);
nor_5  g04838(new_n7186, new_n2445, new_n7187);
not_8  g04839(new_n7187, new_n7188);
xnor_4 g04840(new_n7186, n15636, new_n7189);
not_8  g04841(n6794, new_n7190_1);
xnor_4 g04842(n18962, n14090, new_n7191);
nor_5  g04843(new_n7191, new_n7190_1, new_n7192);
nor_5  g04844(new_n7192, n20077, new_n7193);
xnor_4 g04845(new_n7141, new_n7176, new_n7194);
xnor_4 g04846(new_n7192, new_n5809, new_n7195);
not_8  g04847(new_n7195, new_n7196);
nor_5  g04848(new_n7196, new_n7194, new_n7197);
nor_5  g04849(new_n7197, new_n7193, new_n7198);
nand_5 g04850(new_n7198, new_n7189, new_n7199);
nand_5 g04851(new_n7199, new_n7188, new_n7200);
not_8  g04852(new_n7200, new_n7201);
nand_5 g04853(new_n7201, new_n7185, new_n7202);
nand_5 g04854(new_n7202, new_n7184, new_n7203);
nand_5 g04855(new_n7203, new_n7174, new_n7204);
nand_5 g04856(new_n7204, new_n7173, new_n7205);
xnor_4 g04857(new_n7169, n22660, new_n7206);
not_8  g04858(new_n7206, new_n7207);
nor_5  g04859(new_n7207, new_n7205, new_n7208);
nor_5  g04860(new_n7208, new_n7170, new_n7209);
not_8  g04861(new_n7209, new_n7210);
nand_5 g04862(new_n7210, new_n7167, new_n7211);
nand_5 g04863(new_n7211, new_n7166, new_n7212);
nand_5 g04864(new_n7212, new_n7162, new_n7213);
nand_5 g04865(new_n7213, new_n7161, new_n7214);
xnor_4 g04866(new_n7214, new_n7159, new_n7215);
not_8  g04867(new_n7215, new_n7216);
xnor_4 g04868(n21915, new_n6542_1, new_n7217);
nor_5  g04869(n27037, n13775, new_n7218);
not_8  g04870(n13775, new_n7219);
xnor_4 g04871(n27037, new_n7219, new_n7220);
not_8  g04872(new_n7220, new_n7221);
nor_5  g04873(n8964, n1293, new_n7222);
not_8  g04874(n1293, new_n7223);
xnor_4 g04875(n8964, new_n7223, new_n7224);
not_8  g04876(new_n7224, new_n7225);
nor_5  g04877(n20151, n19042, new_n7226);
not_8  g04878(n19042, new_n7227);
xnor_4 g04879(n20151, new_n7227, new_n7228);
not_8  g04880(new_n7228, new_n7229_1);
nor_5  g04881(n19472, n7693, new_n7230_1);
xnor_4 g04882(n19472, new_n4185, new_n7231);
not_8  g04883(new_n7231, new_n7232);
nand_5 g04884(n25370, n10405, new_n7233_1);
nor_5  g04885(n25370, n10405, new_n7234);
not_8  g04886(new_n7234, new_n7235);
nor_5  g04887(n24786, n11302, new_n7236_1);
not_8  g04888(new_n4293, new_n7237);
nor_5  g04889(new_n4299, new_n7237, new_n7238);
nor_5  g04890(new_n7238, new_n7236_1, new_n7239);
nand_5 g04891(new_n7239, new_n7235, new_n7240);
nand_5 g04892(new_n7240, new_n7233_1, new_n7241);
nor_5  g04893(new_n7241, new_n7232, new_n7242);
nor_5  g04894(new_n7242, new_n7230_1, new_n7243);
nor_5  g04895(new_n7243, new_n7229_1, new_n7244);
nor_5  g04896(new_n7244, new_n7226, new_n7245);
nor_5  g04897(new_n7245, new_n7225, new_n7246);
nor_5  g04898(new_n7246, new_n7222, new_n7247);
nor_5  g04899(new_n7247, new_n7221, new_n7248);
nor_5  g04900(new_n7248, new_n7218, new_n7249);
xnor_4 g04901(new_n7249, new_n7217, new_n7250);
xnor_4 g04902(new_n7250, n17351, new_n7251);
xnor_4 g04903(new_n7247, new_n7220, new_n7252);
not_8  g04904(new_n7252, new_n7253_1);
nand_5 g04905(new_n7253_1, n11736, new_n7254);
xnor_4 g04906(new_n7252, n11736, new_n7255);
xnor_4 g04907(new_n7245, new_n7224, new_n7256_1);
nor_5  g04908(new_n7256_1, new_n5746, new_n7257);
not_8  g04909(new_n7257, new_n7258);
xnor_4 g04910(new_n7256_1, n23200, new_n7259);
xnor_4 g04911(new_n7243, new_n7228, new_n7260);
nor_5  g04912(new_n7260, new_n5749, new_n7261);
not_8  g04913(new_n7261, new_n7262);
xnor_4 g04914(new_n7260, n17959, new_n7263);
xnor_4 g04915(new_n7241, new_n7231, new_n7264);
not_8  g04916(new_n7264, new_n7265);
nand_5 g04917(new_n7265, n7566, new_n7266);
xnor_4 g04918(new_n7264, n7566, new_n7267);
xnor_4 g04919(n25370, new_n4189, new_n7268_1);
not_8  g04920(new_n7268_1, new_n7269);
xnor_4 g04921(new_n7269, new_n7239, new_n7270);
nand_5 g04922(new_n7270, n7731, new_n7271);
xnor_4 g04923(new_n7270, new_n5755, new_n7272);
nor_5  g04924(new_n4300, new_n5760, new_n7273);
not_8  g04925(new_n7273, new_n7274);
not_8  g04926(new_n4313, new_n7275);
nor_5  g04927(new_n7275, n20986, new_n7276);
nor_5  g04928(new_n4317, new_n7068, new_n7277_1);
xnor_4 g04929(new_n4313, new_n5763, new_n7278);
nor_5  g04930(new_n7278, new_n7277_1, new_n7279);
nor_5  g04931(new_n7279, new_n7276, new_n7280_1);
xnor_4 g04932(new_n4300, n12341, new_n7281);
nand_5 g04933(new_n7281, new_n7280_1, new_n7282);
nand_5 g04934(new_n7282, new_n7274, new_n7283);
nand_5 g04935(new_n7283, new_n7272, new_n7284);
nand_5 g04936(new_n7284, new_n7271, new_n7285);
nand_5 g04937(new_n7285, new_n7267, new_n7286);
nand_5 g04938(new_n7286, new_n7266, new_n7287);
nand_5 g04939(new_n7287, new_n7263, new_n7288);
nand_5 g04940(new_n7288, new_n7262, new_n7289);
nand_5 g04941(new_n7289, new_n7259, new_n7290);
nand_5 g04942(new_n7290, new_n7258, new_n7291);
nand_5 g04943(new_n7291, new_n7255, new_n7292);
nand_5 g04944(new_n7292, new_n7254, new_n7293);
xnor_4 g04945(new_n7293, new_n7251, new_n7294);
xnor_4 g04946(new_n7294, new_n7216, new_n7295);
xnor_4 g04947(new_n7291, new_n7255, new_n7296);
not_8  g04948(new_n7162, new_n7297);
xnor_4 g04949(new_n7212, new_n7297, new_n7298_1);
nand_5 g04950(new_n7298_1, new_n7296, new_n7299);
not_8  g04951(new_n7298_1, new_n7300);
xnor_4 g04952(new_n7300, new_n7296, new_n7301);
xnor_4 g04953(new_n7289, new_n7259, new_n7302);
xnor_4 g04954(new_n7209, new_n7167, new_n7303);
nand_5 g04955(new_n7303, new_n7302, new_n7304);
not_8  g04956(new_n7303, new_n7305_1);
xnor_4 g04957(new_n7305_1, new_n7302, new_n7306);
xnor_4 g04958(new_n7287, new_n7263, new_n7307);
xnor_4 g04959(new_n7206, new_n7205, new_n7308_1);
nand_5 g04960(new_n7308_1, new_n7307, new_n7309);
not_8  g04961(new_n7308_1, new_n7310);
xnor_4 g04962(new_n7310, new_n7307, new_n7311);
xnor_4 g04963(new_n7203, new_n7174, new_n7312);
not_8  g04964(new_n7312, new_n7313_1);
xnor_4 g04965(new_n7285, new_n7267, new_n7314);
not_8  g04966(new_n7314, new_n7315);
nor_5  g04967(new_n7315, new_n7313_1, new_n7316);
xnor_4 g04968(new_n7315, new_n7312, new_n7317);
not_8  g04969(new_n7317, new_n7318);
xnor_4 g04970(new_n7200, new_n7185, new_n7319);
not_8  g04971(new_n7319, new_n7320);
xnor_4 g04972(new_n7283, new_n7272, new_n7321);
and_5  g04973(new_n7321, new_n7320, new_n7322);
xnor_4 g04974(new_n7321, new_n7319, new_n7323);
not_8  g04975(new_n7323, new_n7324);
xnor_4 g04976(new_n7281, new_n7280_1, new_n7325);
xnor_4 g04977(new_n7198, new_n7189, new_n7326);
not_8  g04978(new_n7326, new_n7327);
and_5  g04979(new_n7327, new_n7325, new_n7328);
xnor_4 g04980(new_n7326, new_n7325, new_n7329);
not_8  g04981(new_n7329, new_n7330_1);
xnor_4 g04982(new_n7278, new_n7277_1, new_n7331);
xnor_4 g04983(new_n7195, new_n7194, new_n7332);
nor_5  g04984(new_n7332, new_n7331, new_n7333);
xnor_4 g04985(new_n7191, n6794, new_n7334);
not_8  g04986(new_n7334, new_n7335_1);
xnor_4 g04987(new_n4317, n12384, new_n7336);
nor_5  g04988(new_n7336, new_n7335_1, new_n7337);
not_8  g04989(new_n7337, new_n7338);
not_8  g04990(new_n7332, new_n7339_1);
xnor_4 g04991(new_n7339_1, new_n7331, new_n7340);
not_8  g04992(new_n7340, new_n7341);
nor_5  g04993(new_n7341, new_n7338, new_n7342);
nor_5  g04994(new_n7342, new_n7333, new_n7343);
nor_5  g04995(new_n7343, new_n7330_1, new_n7344);
nor_5  g04996(new_n7344, new_n7328, new_n7345);
nor_5  g04997(new_n7345, new_n7324, new_n7346_1);
nor_5  g04998(new_n7346_1, new_n7322, new_n7347);
nor_5  g04999(new_n7347, new_n7318, new_n7348);
nor_5  g05000(new_n7348, new_n7316, new_n7349_1);
not_8  g05001(new_n7349_1, new_n7350);
nand_5 g05002(new_n7350, new_n7311, new_n7351);
nand_5 g05003(new_n7351, new_n7309, new_n7352);
nand_5 g05004(new_n7352, new_n7306, new_n7353);
nand_5 g05005(new_n7353, new_n7304, new_n7354);
nand_5 g05006(new_n7354, new_n7301, new_n7355);
nand_5 g05007(new_n7355, new_n7299, new_n7356);
xnor_4 g05008(new_n7356, new_n7295, n723);
xnor_4 g05009(n26986, n2272, new_n7358);
not_8  g05010(n25331, new_n7359);
or_5   g05011(new_n7359, n21287, new_n7360);
xnor_4 g05012(n25331, n21287, new_n7361);
not_8  g05013(n18483, new_n7362);
or_5   g05014(new_n7362, n4256, new_n7363_1);
xnor_4 g05015(n18483, n4256, new_n7364);
not_8  g05016(n21934, new_n7365);
or_5   g05017(n22332, new_n7365, new_n7366);
xnor_4 g05018(n22332, n21934, new_n7367);
not_8  g05019(n18901, new_n7368);
or_5   g05020(n18907, new_n7368, new_n7369);
xnor_4 g05021(n18907, n18901, new_n7370);
not_8  g05022(n4376, new_n7371);
nor_5  g05023(new_n7371, n2731, new_n7372);
xnor_4 g05024(n4376, n2731, new_n7373);
not_8  g05025(new_n7373, new_n7374);
not_8  g05026(n14570, new_n7375);
nor_5  g05027(n19911, new_n7375, new_n7376);
xnor_4 g05028(n19911, n14570, new_n7377_1);
nor_5  g05029(n23775, new_n2390, new_n7378);
not_8  g05030(n23775, new_n7379);
nor_5  g05031(new_n7379, n13708, new_n7380);
nor_5  g05032(new_n3977, n8259, new_n7381);
not_8  g05033(n8259, new_n7382);
nor_5  g05034(n18409, new_n7382, new_n7383);
not_8  g05035(n11479, new_n7384);
nand_5 g05036(new_n7384, n5704, new_n7385);
nor_5  g05037(new_n7385, new_n7383, new_n7386);
nor_5  g05038(new_n7386, new_n7381, new_n7387);
nor_5  g05039(new_n7387, new_n7380, new_n7388);
nor_5  g05040(new_n7388, new_n7378, new_n7389);
and_5  g05041(new_n7389, new_n7377_1, new_n7390_1);
nor_5  g05042(new_n7390_1, new_n7376, new_n7391);
nor_5  g05043(new_n7391, new_n7374, new_n7392);
nor_5  g05044(new_n7392, new_n7372, new_n7393);
not_8  g05045(new_n7393, new_n7394);
nand_5 g05046(new_n7394, new_n7370, new_n7395);
nand_5 g05047(new_n7395, new_n7369, new_n7396);
nand_5 g05048(new_n7396, new_n7367, new_n7397);
nand_5 g05049(new_n7397, new_n7366, new_n7398);
nand_5 g05050(new_n7398, new_n7364, new_n7399);
nand_5 g05051(new_n7399, new_n7363_1, new_n7400);
nand_5 g05052(new_n7400, new_n7361, new_n7401);
nand_5 g05053(new_n7401, new_n7360, new_n7402);
xnor_4 g05054(new_n7402, new_n7358, new_n7403_1);
not_8  g05055(n468, new_n7404);
xnor_4 g05056(n1255, new_n7404, new_n7405);
not_8  g05057(new_n7405, new_n7406);
or_5   g05058(n9512, n5400, new_n7407);
not_8  g05059(n5400, new_n7408_1);
xnor_4 g05060(n9512, new_n7408_1, new_n7409);
nor_5  g05061(n23923, n16608, new_n7410);
not_8  g05062(new_n7410, new_n7411);
not_8  g05063(n16608, new_n7412);
xnor_4 g05064(n23923, new_n7412, new_n7413);
nor_5  g05065(n21735, n329, new_n7414);
not_8  g05066(n329, new_n7415);
xnor_4 g05067(n21735, new_n7415, new_n7416);
not_8  g05068(new_n7416, new_n7417);
nor_5  g05069(n24170, n24085, new_n7418);
xnor_4 g05070(n24170, new_n4822, new_n7419);
not_8  g05071(new_n7419, new_n7420);
nor_5  g05072(n14071, n2409, new_n7421_1);
not_8  g05073(n2409, new_n7422);
xnor_4 g05074(n14071, new_n7422, new_n7423);
not_8  g05075(new_n7423, new_n7424);
nor_5  g05076(n8869, n1738, new_n7425);
xnor_4 g05077(n8869, new_n4831, new_n7426);
not_8  g05078(new_n7426, new_n7427);
nor_5  g05079(n12152, n10372, new_n7428_1);
nand_5 g05080(n19107, n7428, new_n7429);
not_8  g05081(new_n7429, new_n7430);
not_8  g05082(n10372, new_n7431);
xnor_4 g05083(n12152, new_n7431, new_n7432_1);
not_8  g05084(new_n7432_1, new_n7433);
nor_5  g05085(new_n7433, new_n7430, new_n7434);
nor_5  g05086(new_n7434, new_n7428_1, new_n7435);
nor_5  g05087(new_n7435, new_n7427, new_n7436);
nor_5  g05088(new_n7436, new_n7425, new_n7437_1);
nor_5  g05089(new_n7437_1, new_n7424, new_n7438);
nor_5  g05090(new_n7438, new_n7421_1, new_n7439);
nor_5  g05091(new_n7439, new_n7420, new_n7440);
nor_5  g05092(new_n7440, new_n7418, new_n7441);
nor_5  g05093(new_n7441, new_n7417, new_n7442);
nor_5  g05094(new_n7442, new_n7414, new_n7443);
not_8  g05095(new_n7443, new_n7444);
nand_5 g05096(new_n7444, new_n7413, new_n7445);
nand_5 g05097(new_n7445, new_n7411, new_n7446);
nand_5 g05098(new_n7446, new_n7409, new_n7447);
nand_5 g05099(new_n7447, new_n7407, new_n7448);
xnor_4 g05100(new_n7448, new_n7406, new_n7449);
not_8  g05101(n12861, new_n7450);
xnor_4 g05102(n14130, new_n7450, new_n7451);
not_8  g05103(new_n7451, new_n7452);
or_5   g05104(n16482, n13333, new_n7453);
not_8  g05105(n13333, new_n7454);
xnor_4 g05106(n16482, new_n7454, new_n7455);
nor_5  g05107(n9942, n2210, new_n7456);
not_8  g05108(n2210, new_n7457);
xnor_4 g05109(n9942, new_n7457, new_n7458);
not_8  g05110(new_n7458, new_n7459);
nor_5  g05111(n25643, n20604, new_n7460_1);
not_8  g05112(new_n5386_1, new_n7461);
nor_5  g05113(new_n5389, new_n7461, new_n7462);
nor_5  g05114(new_n7462, new_n7460_1, new_n7463);
nor_5  g05115(new_n7463, new_n7459, new_n7464);
nor_5  g05116(new_n7464, new_n7456, new_n7465);
not_8  g05117(new_n7465, new_n7466);
nand_5 g05118(new_n7466, new_n7455, new_n7467);
nand_5 g05119(new_n7467, new_n7453, new_n7468);
xnor_4 g05120(new_n7468, new_n7452, new_n7469);
not_8  g05121(new_n7469, new_n7470);
nand_5 g05122(new_n7470, new_n7449, new_n7471);
xnor_4 g05123(new_n7469, new_n7449, new_n7472);
not_8  g05124(new_n7409, new_n7473);
xnor_4 g05125(new_n7446, new_n7473, new_n7474);
xnor_4 g05126(new_n7465, new_n7455, new_n7475_1);
not_8  g05127(new_n7475_1, new_n7476);
nand_5 g05128(new_n7476, new_n7474, new_n7477_1);
xnor_4 g05129(new_n7475_1, new_n7474, new_n7478);
xnor_4 g05130(new_n7463, new_n7458, new_n7479);
not_8  g05131(new_n7479, new_n7480);
xnor_4 g05132(new_n7443, new_n7413, new_n7481);
nand_5 g05133(new_n7481, new_n7480, new_n7482);
xnor_4 g05134(new_n7481, new_n7479, new_n7483);
not_8  g05135(new_n5390, new_n7484);
xnor_4 g05136(new_n7441, new_n7416, new_n7485);
nand_5 g05137(new_n7485, new_n7484, new_n7486);
xnor_4 g05138(new_n7485, new_n5390, new_n7487);
xnor_4 g05139(new_n7439, new_n7419, new_n7488);
nand_5 g05140(new_n7488, new_n5383, new_n7489);
xnor_4 g05141(new_n7488, new_n5395, new_n7490);
not_8  g05142(new_n5375, new_n7491);
xnor_4 g05143(new_n7437_1, new_n7423, new_n7492);
nand_5 g05144(new_n7492, new_n7491, new_n7493);
xnor_4 g05145(new_n7492, new_n5375, new_n7494);
xnor_4 g05146(new_n7435, new_n7426, new_n7495);
nand_5 g05147(new_n7495, new_n5368, new_n7496);
not_8  g05148(new_n7496, new_n7497);
xnor_4 g05149(new_n7495, new_n5367, new_n7498);
not_8  g05150(new_n7498, new_n7499);
not_8  g05151(new_n5360, new_n7500);
xnor_4 g05152(new_n7432_1, new_n7430, new_n7501);
not_8  g05153(new_n7501, new_n7502);
nor_5  g05154(new_n7502, new_n7500, new_n7503);
not_8  g05155(n7428, new_n7504);
xnor_4 g05156(n19107, new_n7504, new_n7505);
nor_5  g05157(new_n7505, new_n5405, new_n7506);
xnor_4 g05158(new_n7501, new_n7500, new_n7507_1);
nand_5 g05159(new_n7507_1, new_n7506, new_n7508);
not_8  g05160(new_n7508, new_n7509);
nor_5  g05161(new_n7509, new_n7503, new_n7510);
nor_5  g05162(new_n7510, new_n7499, new_n7511);
nor_5  g05163(new_n7511, new_n7497, new_n7512);
not_8  g05164(new_n7512, new_n7513);
nand_5 g05165(new_n7513, new_n7494, new_n7514_1);
nand_5 g05166(new_n7514_1, new_n7493, new_n7515);
nand_5 g05167(new_n7515, new_n7490, new_n7516);
nand_5 g05168(new_n7516, new_n7489, new_n7517);
nand_5 g05169(new_n7517, new_n7487, new_n7518);
nand_5 g05170(new_n7518, new_n7486, new_n7519);
nand_5 g05171(new_n7519, new_n7483, new_n7520);
nand_5 g05172(new_n7520, new_n7482, new_n7521);
nand_5 g05173(new_n7521, new_n7478, new_n7522);
nand_5 g05174(new_n7522, new_n7477_1, new_n7523);
nand_5 g05175(new_n7523, new_n7472, new_n7524_1);
nand_5 g05176(new_n7524_1, new_n7471, new_n7525);
not_8  g05177(n22253, new_n7526);
xnor_4 g05178(n22442, new_n7526, new_n7527);
not_8  g05179(new_n7527, new_n7528);
or_5   g05180(n1255, n468, new_n7529);
nand_5 g05181(new_n7448, new_n7405, new_n7530);
nand_5 g05182(new_n7530, new_n7529, new_n7531);
xnor_4 g05183(new_n7531, new_n7528, new_n7532);
not_8  g05184(n8305, new_n7533);
xnor_4 g05185(n8856, new_n7533, new_n7534);
not_8  g05186(new_n7534, new_n7535);
or_5   g05187(n14130, n12861, new_n7536);
nand_5 g05188(new_n7468, new_n7451, new_n7537);
nand_5 g05189(new_n7537, new_n7536, new_n7538);
xnor_4 g05190(new_n7538, new_n7535, new_n7539);
xnor_4 g05191(new_n7539, new_n7532, new_n7540);
xnor_4 g05192(new_n7540, new_n7525, new_n7541);
not_8  g05193(new_n7541, new_n7542);
nand_5 g05194(new_n7542, new_n7403_1, new_n7543);
xnor_4 g05195(new_n7541, new_n7403_1, new_n7544);
xnor_4 g05196(new_n7400, new_n7361, new_n7545);
xnor_4 g05197(new_n7523, new_n7472, new_n7546);
not_8  g05198(new_n7546, new_n7547);
nand_5 g05199(new_n7547, new_n7545, new_n7548);
xnor_4 g05200(new_n7546, new_n7545, new_n7549);
xnor_4 g05201(new_n7398, new_n7364, new_n7550);
xnor_4 g05202(new_n7521, new_n7478, new_n7551);
not_8  g05203(new_n7551, new_n7552);
nand_5 g05204(new_n7552, new_n7550, new_n7553);
xnor_4 g05205(new_n7551, new_n7550, new_n7554);
xnor_4 g05206(new_n7396, new_n7367, new_n7555);
xnor_4 g05207(new_n7519, new_n7483, new_n7556);
not_8  g05208(new_n7556, new_n7557);
nand_5 g05209(new_n7557, new_n7555, new_n7558_1);
xnor_4 g05210(new_n7556, new_n7555, new_n7559);
xnor_4 g05211(new_n7393, new_n7370, new_n7560);
not_8  g05212(new_n7560, new_n7561);
not_8  g05213(new_n7487, new_n7562);
xnor_4 g05214(new_n7517, new_n7562, new_n7563);
nand_5 g05215(new_n7563, new_n7561, new_n7564);
xnor_4 g05216(new_n7563, new_n7560, new_n7565);
xnor_4 g05217(new_n7391, new_n7374, new_n7566_1);
xnor_4 g05218(new_n7515, new_n7490, new_n7567);
not_8  g05219(new_n7567, new_n7568);
nand_5 g05220(new_n7568, new_n7566_1, new_n7569_1);
xnor_4 g05221(new_n7567, new_n7566_1, new_n7570);
xnor_4 g05222(new_n7512, new_n7494, new_n7571);
not_8  g05223(new_n7571, new_n7572_1);
xnor_4 g05224(new_n7389, new_n7377_1, new_n7573);
not_8  g05225(new_n7573, new_n7574);
nor_5  g05226(new_n7574, new_n7572_1, new_n7575_1);
not_8  g05227(new_n7575_1, new_n7576);
xnor_4 g05228(new_n7510, new_n7498, new_n7577);
not_8  g05229(new_n7577, new_n7578);
xnor_4 g05230(n23775, n13708, new_n7579);
xnor_4 g05231(new_n7579, new_n7387, new_n7580);
not_8  g05232(new_n7580, new_n7581);
nor_5  g05233(new_n7581, new_n7578, new_n7582);
not_8  g05234(new_n7582, new_n7583);
xnor_4 g05235(new_n7581, new_n7577, new_n7584);
xnor_4 g05236(new_n7505, new_n5356, new_n7585_1);
xnor_4 g05237(n11479, n5704, new_n7586);
nor_5  g05238(new_n7586, new_n7585_1, new_n7587);
xnor_4 g05239(n18409, n8259, new_n7588_1);
xnor_4 g05240(new_n7588_1, new_n7385, new_n7589);
not_8  g05241(new_n7589, new_n7590);
and_5  g05242(new_n7590, new_n7587, new_n7591);
xnor_4 g05243(new_n7507_1, new_n7506, new_n7592);
xnor_4 g05244(new_n7589, new_n7587, new_n7593_1);
and_5  g05245(new_n7593_1, new_n7592, new_n7594);
nor_5  g05246(new_n7594, new_n7591, new_n7595);
nand_5 g05247(new_n7595, new_n7584, new_n7596);
nand_5 g05248(new_n7596, new_n7583, new_n7597);
xnor_4 g05249(new_n7574, new_n7571, new_n7598_1);
nand_5 g05250(new_n7598_1, new_n7597, new_n7599);
nand_5 g05251(new_n7599, new_n7576, new_n7600);
nand_5 g05252(new_n7600, new_n7570, new_n7601);
nand_5 g05253(new_n7601, new_n7569_1, new_n7602);
nand_5 g05254(new_n7602, new_n7565, new_n7603);
nand_5 g05255(new_n7603, new_n7564, new_n7604);
nand_5 g05256(new_n7604, new_n7559, new_n7605);
nand_5 g05257(new_n7605, new_n7558_1, new_n7606);
nand_5 g05258(new_n7606, new_n7554, new_n7607_1);
nand_5 g05259(new_n7607_1, new_n7553, new_n7608);
nand_5 g05260(new_n7608, new_n7549, new_n7609);
nand_5 g05261(new_n7609, new_n7548, new_n7610_1);
nand_5 g05262(new_n7610_1, new_n7544, new_n7611);
nand_5 g05263(new_n7611, new_n7543, new_n7612);
not_8  g05264(n2272, new_n7613);
or_5   g05265(n26986, new_n7613, new_n7614);
nand_5 g05266(new_n7402, new_n7358, new_n7615);
nand_5 g05267(new_n7615, new_n7614, new_n7616_1);
not_8  g05268(new_n7616_1, new_n7617);
or_5   g05269(n22442, n22253, new_n7618);
nand_5 g05270(new_n7531, new_n7527, new_n7619);
nand_5 g05271(new_n7619, new_n7618, new_n7620);
nor_5  g05272(n8856, n8305, new_n7621);
not_8  g05273(new_n7621, new_n7622);
nand_5 g05274(new_n7538, new_n7534, new_n7623);
nand_5 g05275(new_n7623, new_n7622, new_n7624);
xnor_4 g05276(new_n7624, new_n7620, new_n7625);
not_8  g05277(new_n7625, new_n7626);
not_8  g05278(new_n7539, new_n7627);
nand_5 g05279(new_n7627, new_n7532, new_n7628);
nand_5 g05280(new_n7540, new_n7525, new_n7629);
nand_5 g05281(new_n7629, new_n7628, new_n7630_1);
xnor_4 g05282(new_n7630_1, new_n7626, new_n7631);
xnor_4 g05283(new_n7631, new_n7617, new_n7632);
xnor_4 g05284(new_n7632, new_n7612, n735);
xnor_4 g05285(n21138, new_n6940, new_n7634);
not_8  g05286(new_n7634, new_n7635);
not_8  g05287(n19234, new_n7636);
xnor_4 g05288(new_n7191, new_n7636, new_n7637);
xnor_4 g05289(new_n7637, n26167, new_n7638);
xnor_4 g05290(new_n7638, new_n7635, n779);
or_5   g05291(n17458, new_n6308_1, new_n7640);
xnor_4 g05292(n17458, n8526, new_n7641);
or_5   g05293(new_n6359, n1222, new_n7642);
xnor_4 g05294(n2816, n1222, new_n7643_1);
not_8  g05295(n20359, new_n7644);
or_5   g05296(n25240, new_n7644, new_n7645);
xnor_4 g05297(n25240, n20359, new_n7646);
not_8  g05298(n10125, new_n7647_1);
nand_5 g05299(new_n7647_1, n4409, new_n7648);
xnor_4 g05300(n10125, n4409, new_n7649);
not_8  g05301(n8067, new_n7650);
nand_5 g05302(new_n7650, n3570, new_n7651);
xnor_4 g05303(n8067, n3570, new_n7652);
nor_5  g05304(n20923, new_n6373, new_n7653);
not_8  g05305(new_n7653, new_n7654);
xnor_4 g05306(n20923, n13668, new_n7655);
nor_5  g05307(new_n4417, n18157, new_n7656);
not_8  g05308(new_n7656, new_n7657_1);
xnor_4 g05309(n21276, n18157, new_n7658);
nor_5  g05310(n26748, new_n6982, new_n7659);
nor_5  g05311(new_n4411, n12161, new_n7660);
not_8  g05312(n5026, new_n7661);
nor_5  g05313(n10057, new_n7661, new_n7662);
nand_5 g05314(n10057, new_n7661, new_n7663);
not_8  g05315(n8581, new_n7664);
nor_5  g05316(n8920, new_n7664, new_n7665);
nand_5 g05317(new_n7665, new_n7663, new_n7666);
not_8  g05318(new_n7666, new_n7667);
nor_5  g05319(new_n7667, new_n7662, new_n7668);
nor_5  g05320(new_n7668, new_n7660, new_n7669);
nor_5  g05321(new_n7669, new_n7659, new_n7670_1);
nand_5 g05322(new_n7670_1, new_n7658, new_n7671);
nand_5 g05323(new_n7671, new_n7657_1, new_n7672);
nand_5 g05324(new_n7672, new_n7655, new_n7673);
nand_5 g05325(new_n7673, new_n7654, new_n7674_1);
nand_5 g05326(new_n7674_1, new_n7652, new_n7675);
nand_5 g05327(new_n7675, new_n7651, new_n7676);
nand_5 g05328(new_n7676, new_n7649, new_n7677);
nand_5 g05329(new_n7677, new_n7648, new_n7678_1);
nand_5 g05330(new_n7678_1, new_n7646, new_n7679_1);
nand_5 g05331(new_n7679_1, new_n7645, new_n7680);
nand_5 g05332(new_n7680, new_n7643_1, new_n7681);
nand_5 g05333(new_n7681, new_n7642, new_n7682);
nand_5 g05334(new_n7682, new_n7641, new_n7683);
nand_5 g05335(new_n7683, new_n7640, new_n7684);
not_8  g05336(new_n7684, new_n7685);
not_8  g05337(n26986, new_n7686_1);
or_5   g05338(new_n7686_1, n19282, new_n7687);
xnor_4 g05339(n26986, n19282, new_n7688);
not_8  g05340(n21287, new_n7689);
or_5   g05341(new_n7689, n12657, new_n7690);
xnor_4 g05342(n21287, n12657, new_n7691);
not_8  g05343(n4256, new_n7692_1);
or_5   g05344(n17077, new_n7692_1, new_n7693_1);
xnor_4 g05345(n17077, n4256, new_n7694);
not_8  g05346(n22332, new_n7695);
or_5   g05347(n26510, new_n7695, new_n7696);
nand_5 g05348(new_n3991, new_n3963, new_n7697);
nand_5 g05349(new_n7697, new_n7696, new_n7698_1);
nand_5 g05350(new_n7698_1, new_n7694, new_n7699);
nand_5 g05351(new_n7699, new_n7693_1, new_n7700);
nand_5 g05352(new_n7700, new_n7691, new_n7701);
nand_5 g05353(new_n7701, new_n7690, new_n7702);
nand_5 g05354(new_n7702, new_n7688, new_n7703);
nand_5 g05355(new_n7703, new_n7687, new_n7704);
xnor_4 g05356(new_n7704, new_n7685, new_n7705);
xnor_4 g05357(new_n7682, new_n7641, new_n7706);
xnor_4 g05358(new_n7702, new_n7688, new_n7707);
nor_5  g05359(new_n7707, new_n7706, new_n7708_1);
xnor_4 g05360(new_n7707, new_n7706, new_n7709);
xnor_4 g05361(new_n7680, new_n7643_1, new_n7710);
xnor_4 g05362(new_n7700, new_n7691, new_n7711);
nand_5 g05363(new_n7711, new_n7710, new_n7712);
not_8  g05364(new_n7710, new_n7713);
xnor_4 g05365(new_n7711, new_n7713, new_n7714);
not_8  g05366(new_n7646, new_n7715);
xnor_4 g05367(new_n7678_1, new_n7715, new_n7716);
not_8  g05368(new_n7716, new_n7717);
xnor_4 g05369(new_n7698_1, new_n7694, new_n7718);
nand_5 g05370(new_n7718, new_n7717, new_n7719);
xnor_4 g05371(new_n7718, new_n7716, new_n7720);
not_8  g05372(new_n7649, new_n7721_1);
xnor_4 g05373(new_n7676, new_n7721_1, new_n7722);
not_8  g05374(new_n7722, new_n7723);
nand_5 g05375(new_n7723, new_n3992, new_n7724);
xnor_4 g05376(new_n7722, new_n3992, new_n7725);
xnor_4 g05377(new_n7674_1, new_n7652, new_n7726);
nand_5 g05378(new_n7726, new_n4002, new_n7727);
not_8  g05379(new_n7726, new_n7728);
xnor_4 g05380(new_n7728, new_n4002, new_n7729);
xnor_4 g05381(new_n7672, new_n7655, new_n7730);
nand_5 g05382(new_n7730, new_n4010_1, new_n7731_1);
xnor_4 g05383(new_n7730, new_n4009, new_n7732);
xnor_4 g05384(new_n7670_1, new_n7658, new_n7733);
nand_5 g05385(new_n7733, new_n4020, new_n7734);
xnor_4 g05386(new_n7733, new_n4019, new_n7735);
xnor_4 g05387(n26748, n12161, new_n7736);
xnor_4 g05388(new_n7736, new_n7668, new_n7737);
nand_5 g05389(new_n7737, new_n4028, new_n7738);
xnor_4 g05390(new_n7737, new_n4027, new_n7739);
xnor_4 g05391(n10057, n5026, new_n7740);
xnor_4 g05392(new_n7740, new_n7665, new_n7741);
not_8  g05393(new_n7741, new_n7742);
nor_5  g05394(new_n7742, new_n4036, new_n7743);
xnor_4 g05395(n8920, n8581, new_n7744);
nor_5  g05396(new_n7744, new_n4038, new_n7745);
not_8  g05397(new_n7745, new_n7746);
xnor_4 g05398(new_n7741, new_n4035, new_n7747);
nor_5  g05399(new_n7747, new_n7746, new_n7748);
nor_5  g05400(new_n7748, new_n7743, new_n7749);
nand_5 g05401(new_n7749, new_n7739, new_n7750);
nand_5 g05402(new_n7750, new_n7738, new_n7751_1);
nand_5 g05403(new_n7751_1, new_n7735, new_n7752);
nand_5 g05404(new_n7752, new_n7734, new_n7753);
nand_5 g05405(new_n7753, new_n7732, new_n7754);
nand_5 g05406(new_n7754, new_n7731_1, new_n7755);
nand_5 g05407(new_n7755, new_n7729, new_n7756);
nand_5 g05408(new_n7756, new_n7727, new_n7757);
nand_5 g05409(new_n7757, new_n7725, new_n7758);
nand_5 g05410(new_n7758, new_n7724, new_n7759_1);
nand_5 g05411(new_n7759_1, new_n7720, new_n7760);
nand_5 g05412(new_n7760, new_n7719, new_n7761);
nand_5 g05413(new_n7761, new_n7714, new_n7762);
nand_5 g05414(new_n7762, new_n7712, new_n7763);
nor_5  g05415(new_n7763, new_n7709, new_n7764);
nor_5  g05416(new_n7764, new_n7708_1, new_n7765);
xnor_4 g05417(new_n7765, new_n7705, new_n7766);
or_5   g05418(n11898, new_n5042, new_n7767);
xnor_4 g05419(n11898, n2979, new_n7768);
or_5   g05420(n19941, new_n5046_1, new_n7769_1);
xnor_4 g05421(n19941, n647, new_n7770);
or_5   g05422(new_n6243, n1099, new_n7771);
xnor_4 g05423(n20409, n1099, new_n7772);
or_5   g05424(new_n3877, n2113, new_n7773_1);
xnor_4 g05425(n25749, n2113, new_n7774);
or_5   g05426(n21134, new_n3929, new_n7775);
xnor_4 g05427(n21134, n3161, new_n7776);
nor_5  g05428(new_n3933, n6369, new_n7777);
xnor_4 g05429(n9003, n6369, new_n7778);
not_8  g05430(new_n7778, new_n7779);
nor_5  g05431(n25797, new_n3937, new_n7780_1);
not_8  g05432(new_n7780_1, new_n7781);
xnor_4 g05433(n25797, n4957, new_n7782);
nor_5  g05434(new_n3880, n7524, new_n7783);
nor_5  g05435(n15967, new_n3941, new_n7784);
nor_5  g05436(n15743, new_n4368, new_n7785);
nor_5  g05437(new_n3950, n13319, new_n7786);
and_5  g05438(n25435, new_n3945_1, new_n7787);
not_8  g05439(new_n7787, new_n7788_1);
nor_5  g05440(new_n7788_1, new_n7786, new_n7789);
nor_5  g05441(new_n7789, new_n7785, new_n7790);
nor_5  g05442(new_n7790, new_n7784, new_n7791);
nor_5  g05443(new_n7791, new_n7783, new_n7792);
nand_5 g05444(new_n7792, new_n7782, new_n7793);
nand_5 g05445(new_n7793, new_n7781, new_n7794_1);
not_8  g05446(new_n7794_1, new_n7795);
nor_5  g05447(new_n7795, new_n7779, new_n7796);
nor_5  g05448(new_n7796, new_n7777, new_n7797);
not_8  g05449(new_n7797, new_n7798);
nand_5 g05450(new_n7798, new_n7776, new_n7799);
nand_5 g05451(new_n7799, new_n7775, new_n7800);
nand_5 g05452(new_n7800, new_n7774, new_n7801);
nand_5 g05453(new_n7801, new_n7773_1, new_n7802);
nand_5 g05454(new_n7802, new_n7772, new_n7803);
nand_5 g05455(new_n7803, new_n7771, new_n7804);
nand_5 g05456(new_n7804, new_n7770, new_n7805);
nand_5 g05457(new_n7805, new_n7769_1, new_n7806);
nand_5 g05458(new_n7806, new_n7768, new_n7807);
nand_5 g05459(new_n7807, new_n7767, new_n7808);
xnor_4 g05460(new_n7808, new_n7766, new_n7809);
xnor_4 g05461(new_n7806, new_n7768, new_n7810);
xnor_4 g05462(new_n7763, new_n7709, new_n7811_1);
nand_5 g05463(new_n7811_1, new_n7810, new_n7812);
not_8  g05464(new_n7811_1, new_n7813);
xnor_4 g05465(new_n7813, new_n7810, new_n7814);
xnor_4 g05466(new_n7804, new_n7770, new_n7815);
xnor_4 g05467(new_n7761, new_n7714, new_n7816);
not_8  g05468(new_n7816, new_n7817);
nand_5 g05469(new_n7817, new_n7815, new_n7818);
xnor_4 g05470(new_n7816, new_n7815, new_n7819);
xnor_4 g05471(new_n7802, new_n7772, new_n7820);
xnor_4 g05472(new_n7759_1, new_n7720, new_n7821);
not_8  g05473(new_n7821, new_n7822);
nand_5 g05474(new_n7822, new_n7820, new_n7823);
xnor_4 g05475(new_n7821, new_n7820, new_n7824);
xnor_4 g05476(new_n7800, new_n7774, new_n7825);
xnor_4 g05477(new_n7757, new_n7725, new_n7826);
not_8  g05478(new_n7826, new_n7827);
nand_5 g05479(new_n7827, new_n7825, new_n7828);
xnor_4 g05480(new_n7826, new_n7825, new_n7829);
xnor_4 g05481(new_n7797, new_n7776, new_n7830_1);
not_8  g05482(new_n7830_1, new_n7831);
not_8  g05483(new_n7729, new_n7832);
xnor_4 g05484(new_n7755, new_n7832, new_n7833);
nand_5 g05485(new_n7833, new_n7831, new_n7834_1);
xnor_4 g05486(new_n7833, new_n7830_1, new_n7835);
xnor_4 g05487(new_n7794_1, new_n7779, new_n7836);
not_8  g05488(new_n7836, new_n7837);
not_8  g05489(new_n7732, new_n7838);
xnor_4 g05490(new_n7753, new_n7838, new_n7839);
nand_5 g05491(new_n7839, new_n7837, new_n7840);
xnor_4 g05492(new_n7839, new_n7836, new_n7841_1);
xnor_4 g05493(new_n7751_1, new_n7735, new_n7842);
not_8  g05494(new_n7842, new_n7843);
xnor_4 g05495(new_n7792, new_n7782, new_n7844);
nand_5 g05496(new_n7844, new_n7843, new_n7845);
xnor_4 g05497(new_n7749, new_n7739, new_n7846);
xnor_4 g05498(n15967, n7524, new_n7847);
xnor_4 g05499(new_n7847, new_n7790, new_n7848);
not_8  g05500(new_n7848, new_n7849);
nor_5  g05501(new_n7849, new_n7846, new_n7850);
xnor_4 g05502(new_n7848, new_n7846, new_n7851);
not_8  g05503(new_n7851, new_n7852);
xnor_4 g05504(n25435, n20658, new_n7853);
not_8  g05505(new_n7744, new_n7854);
xnor_4 g05506(new_n7854, new_n4038, new_n7855);
not_8  g05507(new_n7855, new_n7856);
nor_5  g05508(new_n7856, new_n7853, new_n7857);
xnor_4 g05509(n15743, n13319, new_n7858);
xnor_4 g05510(new_n7858, new_n7788_1, new_n7859);
not_8  g05511(new_n7859, new_n7860);
nor_5  g05512(new_n7860, new_n7857, new_n7861);
xnor_4 g05513(new_n7747, new_n7745, new_n7862);
xnor_4 g05514(new_n7859, new_n7857, new_n7863);
not_8  g05515(new_n7863, new_n7864);
nor_5  g05516(new_n7864, new_n7862, new_n7865);
nor_5  g05517(new_n7865, new_n7861, new_n7866);
nor_5  g05518(new_n7866, new_n7852, new_n7867);
nor_5  g05519(new_n7867, new_n7850, new_n7868);
not_8  g05520(new_n7868, new_n7869);
xnor_4 g05521(new_n7844, new_n7842, new_n7870);
nand_5 g05522(new_n7870, new_n7869, new_n7871);
nand_5 g05523(new_n7871, new_n7845, new_n7872);
nand_5 g05524(new_n7872, new_n7841_1, new_n7873);
nand_5 g05525(new_n7873, new_n7840, new_n7874);
nand_5 g05526(new_n7874, new_n7835, new_n7875);
nand_5 g05527(new_n7875, new_n7834_1, new_n7876_1);
nand_5 g05528(new_n7876_1, new_n7829, new_n7877);
nand_5 g05529(new_n7877, new_n7828, new_n7878);
nand_5 g05530(new_n7878, new_n7824, new_n7879);
nand_5 g05531(new_n7879, new_n7823, new_n7880);
nand_5 g05532(new_n7880, new_n7819, new_n7881);
nand_5 g05533(new_n7881, new_n7818, new_n7882);
nand_5 g05534(new_n7882, new_n7814, new_n7883);
nand_5 g05535(new_n7883, new_n7812, new_n7884_1);
xnor_4 g05536(new_n7884_1, new_n7809, n809);
not_8  g05537(n2978, new_n7886);
or_5   g05538(n19282, new_n7886, new_n7887);
xnor_4 g05539(n19282, n2978, new_n7888);
or_5   g05540(new_n7114, n12657, new_n7889);
xnor_4 g05541(n23697, n12657, new_n7890);
or_5   g05542(n17077, new_n7118, new_n7891);
xnor_4 g05543(n17077, n2289, new_n7892);
or_5   g05544(n26510, new_n7122, new_n7893);
xnor_4 g05545(n26510, n1112, new_n7894);
not_8  g05546(n20179, new_n7895);
or_5   g05547(n23068, new_n7895, new_n7896);
xnor_4 g05548(n23068, n20179, new_n7897);
not_8  g05549(n19228, new_n7898);
nor_5  g05550(n19514, new_n7898, new_n7899);
xnor_4 g05551(n19514, n19228, new_n7900);
nor_5  g05552(new_n7132, n10053, new_n7901);
not_8  g05553(new_n7901, new_n7902);
xnor_4 g05554(n15539, n10053, new_n7903);
nor_5  g05555(new_n3009, n8052, new_n7904);
nor_5  g05556(n8399, new_n7136, new_n7905);
nor_5  g05557(n10158, new_n3975, new_n7906);
not_8  g05558(n10158, new_n7907);
nor_5  g05559(new_n7907, n9507, new_n7908);
nor_5  g05560(new_n3979, n18962, new_n7909);
not_8  g05561(new_n7909, new_n7910);
nor_5  g05562(new_n7910, new_n7908, new_n7911);
nor_5  g05563(new_n7911, new_n7906, new_n7912);
nor_5  g05564(new_n7912, new_n7905, new_n7913);
nor_5  g05565(new_n7913, new_n7904, new_n7914);
nand_5 g05566(new_n7914, new_n7903, new_n7915);
nand_5 g05567(new_n7915, new_n7902, new_n7916);
and_5  g05568(new_n7916, new_n7900, new_n7917_1);
nor_5  g05569(new_n7917_1, new_n7899, new_n7918);
not_8  g05570(new_n7918, new_n7919);
nand_5 g05571(new_n7919, new_n7897, new_n7920);
nand_5 g05572(new_n7920, new_n7896, new_n7921);
nand_5 g05573(new_n7921, new_n7894, new_n7922);
nand_5 g05574(new_n7922, new_n7893, new_n7923);
nand_5 g05575(new_n7923, new_n7892, new_n7924);
nand_5 g05576(new_n7924, new_n7891, new_n7925);
nand_5 g05577(new_n7925, new_n7890, new_n7926);
nand_5 g05578(new_n7926, new_n7889, new_n7927);
nand_5 g05579(new_n7927, new_n7888, new_n7928);
nand_5 g05580(new_n7928, new_n7887, new_n7929);
not_8  g05581(new_n7929, new_n7930);
nor_5  g05582(n26986, n22626, new_n7931);
not_8  g05583(new_n7931, new_n7932);
not_8  g05584(new_n2428, new_n7933);
nor_5  g05585(new_n7933, new_n2421_1, new_n7934);
not_8  g05586(n1654, new_n7935);
xnor_4 g05587(n4256, new_n7935, new_n7936);
not_8  g05588(new_n7936, new_n7937_1);
nor_5  g05589(n22332, n13783, new_n7938);
not_8  g05590(new_n7938, new_n7939);
not_8  g05591(new_n2427, new_n7940);
nand_5 g05592(new_n7940, new_n2423, new_n7941);
nand_5 g05593(new_n7941, new_n7939, new_n7942);
xnor_4 g05594(new_n7942, new_n7937_1, new_n7943_1);
nand_5 g05595(new_n7943_1, new_n7934, new_n7944);
not_8  g05596(new_n7944, new_n7945);
not_8  g05597(n14440, new_n7946);
xnor_4 g05598(n21287, new_n7946, new_n7947);
not_8  g05599(new_n7947, new_n7948);
or_5   g05600(n4256, n1654, new_n7949_1);
nand_5 g05601(new_n7942, new_n7936, new_n7950_1);
nand_5 g05602(new_n7950_1, new_n7949_1, new_n7951);
xnor_4 g05603(new_n7951, new_n7948, new_n7952);
nand_5 g05604(new_n7952, new_n7945, new_n7953);
not_8  g05605(new_n7953, new_n7954);
not_8  g05606(n22626, new_n7955);
xnor_4 g05607(n26986, new_n7955, new_n7956);
or_5   g05608(n21287, n14440, new_n7957);
nand_5 g05609(new_n7951, new_n7947, new_n7958);
nand_5 g05610(new_n7958, new_n7957, new_n7959_1);
xnor_4 g05611(new_n7959_1, new_n7956, new_n7960);
not_8  g05612(new_n7960, new_n7961);
nand_5 g05613(new_n7961, new_n7954, new_n7962);
nor_5  g05614(new_n7962, new_n7932, new_n7963_1);
nand_5 g05615(new_n7959_1, new_n7956, new_n7964);
nand_5 g05616(new_n7964, new_n7932, new_n7965);
not_8  g05617(new_n7965, new_n7966);
nand_5 g05618(new_n7966, new_n7962, new_n7967);
not_8  g05619(new_n7967, new_n7968_1);
nor_5  g05620(new_n7968_1, new_n7963_1, new_n7969);
not_8  g05621(new_n7969, new_n7970);
or_5   g05622(n13494, n3425, new_n7971);
xnor_4 g05623(n13494, new_n3294, new_n7972);
or_5   g05624(n25345, n9967, new_n7973);
xnor_4 g05625(n25345, new_n3295, new_n7974);
nand_5 g05626(n20946, n9655, new_n7975);
not_8  g05627(new_n7975, new_n7976);
nor_5  g05628(n20946, n9655, new_n7977);
nand_5 g05629(new_n5796, new_n2430, new_n7978);
nand_5 g05630(new_n2463, new_n2431, new_n7979);
nand_5 g05631(new_n7979, new_n7978, new_n7980);
nor_5  g05632(new_n7980, new_n7977, new_n7981);
nor_5  g05633(new_n7981, new_n7976, new_n7982);
nand_5 g05634(new_n7982, new_n7974, new_n7983);
nand_5 g05635(new_n7983, new_n7973, new_n7984);
nand_5 g05636(new_n7984, new_n7972, new_n7985);
nand_5 g05637(new_n7985, new_n7971, new_n7986);
nor_5  g05638(new_n7986, new_n7970, new_n7987);
not_8  g05639(new_n7987, new_n7988);
not_8  g05640(new_n7986, new_n7989);
nor_5  g05641(new_n7989, new_n7969, new_n7990);
xnor_4 g05642(new_n7960, new_n7954, new_n7991);
not_8  g05643(new_n7991, new_n7992_1);
not_8  g05644(new_n7972, new_n7993);
xnor_4 g05645(new_n7984, new_n7993, new_n7994);
nand_5 g05646(new_n7994, new_n7992_1, new_n7995);
xnor_4 g05647(new_n7994, new_n7991, new_n7996);
xnor_4 g05648(new_n7952, new_n7945, new_n7997);
xnor_4 g05649(new_n7982, new_n7974, new_n7998);
not_8  g05650(new_n7998, new_n7999_1);
nand_5 g05651(new_n7999_1, new_n7997, new_n8000);
xnor_4 g05652(new_n7998, new_n7997, new_n8001);
xnor_4 g05653(new_n7943_1, new_n7934, new_n8002);
xnor_4 g05654(n20946, new_n5793, new_n8003);
xnor_4 g05655(new_n8003, new_n7980, new_n8004);
not_8  g05656(new_n8004, new_n8005);
nand_5 g05657(new_n8005, new_n8002, new_n8006_1);
xnor_4 g05658(new_n8004, new_n8002, new_n8007);
not_8  g05659(new_n2429, new_n8008);
nand_5 g05660(new_n2464, new_n8008, new_n8009);
nand_5 g05661(new_n2516, new_n2465, new_n8010);
nand_5 g05662(new_n8010, new_n8009, new_n8011);
nand_5 g05663(new_n8011, new_n8007, new_n8012);
nand_5 g05664(new_n8012, new_n8006_1, new_n8013);
nand_5 g05665(new_n8013, new_n8001, new_n8014);
nand_5 g05666(new_n8014, new_n8000, new_n8015);
nand_5 g05667(new_n8015, new_n7996, new_n8016);
nand_5 g05668(new_n8016, new_n7995, new_n8017);
nor_5  g05669(new_n8017, new_n7990, new_n8018);
nor_5  g05670(new_n8018, new_n7963_1, new_n8019);
nand_5 g05671(new_n8019, new_n7988, new_n8020);
xnor_4 g05672(new_n8020, new_n7930, new_n8021);
xnor_4 g05673(new_n7989, new_n7969, new_n8022);
xnor_4 g05674(new_n8022, new_n8017, new_n8023);
nand_5 g05675(new_n8023, new_n7929, new_n8024);
xnor_4 g05676(new_n8023, new_n7930, new_n8025);
xnor_4 g05677(new_n7927, new_n7888, new_n8026);
xnor_4 g05678(new_n8015, new_n7996, new_n8027_1);
not_8  g05679(new_n8027_1, new_n8028);
nand_5 g05680(new_n8028, new_n8026, new_n8029);
xnor_4 g05681(new_n8027_1, new_n8026, new_n8030);
xnor_4 g05682(new_n7925, new_n7890, new_n8031_1);
xnor_4 g05683(new_n8013, new_n8001, new_n8032);
not_8  g05684(new_n8032, new_n8033);
nand_5 g05685(new_n8033, new_n8031_1, new_n8034);
xnor_4 g05686(new_n8032, new_n8031_1, new_n8035);
xnor_4 g05687(new_n7923, new_n7892, new_n8036);
xnor_4 g05688(new_n8011, new_n8007, new_n8037);
not_8  g05689(new_n8037, new_n8038);
nand_5 g05690(new_n8038, new_n8036, new_n8039);
xnor_4 g05691(new_n8037, new_n8036, new_n8040);
xnor_4 g05692(new_n7921, new_n7894, new_n8041);
nand_5 g05693(new_n8041, new_n2518, new_n8042_1);
xnor_4 g05694(new_n8041, new_n2517, new_n8043);
xnor_4 g05695(new_n7918, new_n7897, new_n8044);
not_8  g05696(new_n8044, new_n8045);
nand_5 g05697(new_n8045, new_n2523, new_n8046);
xnor_4 g05698(new_n8044, new_n2523, new_n8047);
not_8  g05699(new_n7900, new_n8048);
xnor_4 g05700(new_n7916, new_n8048, new_n8049);
not_8  g05701(new_n8049, new_n8050);
nand_5 g05702(new_n8050, new_n2529, new_n8051);
xnor_4 g05703(new_n8049, new_n2529, new_n8052_1);
xnor_4 g05704(new_n7914, new_n7903, new_n8053);
not_8  g05705(new_n8053, new_n8054);
nor_5  g05706(new_n8054, new_n2534, new_n8055);
not_8  g05707(new_n8055, new_n8056);
xnor_4 g05708(new_n8053, new_n2534, new_n8057);
xnor_4 g05709(n8399, n8052, new_n8058);
xnor_4 g05710(new_n8058, new_n7912, new_n8059);
not_8  g05711(new_n8059, new_n8060);
nor_5  g05712(new_n8060, new_n2538, new_n8061);
not_8  g05713(new_n8061, new_n8062);
xnor_4 g05714(new_n8059, new_n2538, new_n8063);
xnor_4 g05715(n26979, n18962, new_n8064);
nor_5  g05716(new_n8064, new_n2548, new_n8065);
xnor_4 g05717(n10158, n9507, new_n8066);
xnor_4 g05718(new_n8066, new_n7910, new_n8067_1);
not_8  g05719(new_n8067_1, new_n8068);
nor_5  g05720(new_n8068, new_n8065, new_n8069);
not_8  g05721(new_n8069, new_n8070);
xnor_4 g05722(new_n8067_1, new_n8065, new_n8071);
nand_5 g05723(new_n8071, new_n2555_1, new_n8072);
nand_5 g05724(new_n8072, new_n8070, new_n8073);
nand_5 g05725(new_n8073, new_n8063, new_n8074);
nand_5 g05726(new_n8074, new_n8062, new_n8075);
nand_5 g05727(new_n8075, new_n8057, new_n8076);
nand_5 g05728(new_n8076, new_n8056, new_n8077);
nand_5 g05729(new_n8077, new_n8052_1, new_n8078);
nand_5 g05730(new_n8078, new_n8051, new_n8079);
nand_5 g05731(new_n8079, new_n8047, new_n8080);
nand_5 g05732(new_n8080, new_n8046, new_n8081);
nand_5 g05733(new_n8081, new_n8043, new_n8082);
nand_5 g05734(new_n8082, new_n8042_1, new_n8083);
nand_5 g05735(new_n8083, new_n8040, new_n8084);
nand_5 g05736(new_n8084, new_n8039, new_n8085);
nand_5 g05737(new_n8085, new_n8035, new_n8086);
nand_5 g05738(new_n8086, new_n8034, new_n8087);
nand_5 g05739(new_n8087, new_n8030, new_n8088);
nand_5 g05740(new_n8088, new_n8029, new_n8089);
nand_5 g05741(new_n8089, new_n8025, new_n8090);
nand_5 g05742(new_n8090, new_n8024, new_n8091);
xnor_4 g05743(new_n8091, new_n8021, n819);
or_5   g05744(n22626, new_n3533, new_n8093);
xnor_4 g05745(n22626, n8856, new_n8094);
or_5   g05746(n14440, new_n3534, new_n8095_1);
xnor_4 g05747(n14440, n14130, new_n8096);
or_5   g05748(new_n3554, n1654, new_n8097);
xnor_4 g05749(n16482, n1654, new_n8098);
or_5   g05750(n13783, new_n3535, new_n8099);
xnor_4 g05751(n13783, n9942, new_n8100);
not_8  g05752(n26660, new_n8101);
nand_5 g05753(new_n8101, n25643, new_n8102);
xnor_4 g05754(n26660, n25643, new_n8103_1);
nor_5  g05755(new_n3536, n3018, new_n8104);
xnor_4 g05756(n9557, n3018, new_n8105);
not_8  g05757(new_n8105, new_n8106);
nor_5  g05758(n3480, new_n3576, new_n8107);
xnor_4 g05759(n3480, n3136, new_n8108);
not_8  g05760(new_n8108, new_n8109_1);
not_8  g05761(n16722, new_n8110);
nor_5  g05762(new_n8110, n6385, new_n8111);
not_8  g05763(new_n8111, new_n8112);
nor_5  g05764(n16722, new_n2360, new_n8113);
not_8  g05765(new_n8113, new_n8114);
nor_5  g05766(n20138, new_n6097, new_n8115);
not_8  g05767(new_n8115, new_n8116);
nor_5  g05768(new_n2364, n11486, new_n8117);
not_8  g05769(new_n8117, new_n8118);
not_8  g05770(n13781, new_n8119);
nor_5  g05771(new_n8119, n9251, new_n8120);
nand_5 g05772(new_n8120, new_n8118, new_n8121);
nand_5 g05773(new_n8121, new_n8116, new_n8122);
nand_5 g05774(new_n8122, new_n8114, new_n8123);
nand_5 g05775(new_n8123, new_n8112, new_n8124);
nor_5  g05776(new_n8124, new_n8109_1, new_n8125);
nor_5  g05777(new_n8125, new_n8107, new_n8126);
nor_5  g05778(new_n8126, new_n8106, new_n8127_1);
nor_5  g05779(new_n8127_1, new_n8104, new_n8128);
not_8  g05780(new_n8128, new_n8129);
nand_5 g05781(new_n8129, new_n8103_1, new_n8130_1);
nand_5 g05782(new_n8130_1, new_n8102, new_n8131);
nand_5 g05783(new_n8131, new_n8100, new_n8132);
nand_5 g05784(new_n8132, new_n8099, new_n8133);
nand_5 g05785(new_n8133, new_n8098, new_n8134);
nand_5 g05786(new_n8134, new_n8097, new_n8135_1);
nand_5 g05787(new_n8135_1, new_n8096, new_n8136);
nand_5 g05788(new_n8136, new_n8095_1, new_n8137);
nand_5 g05789(new_n8137, new_n8094, new_n8138);
nand_5 g05790(new_n8138, new_n8093, new_n8139_1);
not_8  g05791(new_n8139_1, new_n8140);
or_5   g05792(n25120, new_n6309, new_n8141);
xnor_4 g05793(n25120, n3582, new_n8142);
or_5   g05794(n8363, new_n6312, new_n8143);
xnor_4 g05795(n8363, n2145, new_n8144);
or_5   g05796(n14680, new_n6315, new_n8145);
xnor_4 g05797(n14680, n5031, new_n8146);
not_8  g05798(n11044, new_n8147);
or_5   g05799(n17250, new_n8147, new_n8148_1);
xnor_4 g05800(n17250, n11044, new_n8149_1);
or_5   g05801(n23160, new_n6322, new_n8150);
xnor_4 g05802(n23160, n2421, new_n8151);
not_8  g05803(n987, new_n8152);
nor_5  g05804(n16524, new_n8152, new_n8153);
xnor_4 g05805(n16524, n987, new_n8154);
not_8  g05806(new_n8154, new_n8155);
not_8  g05807(n20478, new_n8156);
nor_5  g05808(new_n8156, n11056, new_n8157);
xnor_4 g05809(n20478, n11056, new_n8158);
not_8  g05810(n15271, new_n8159_1);
nor_5  g05811(n26882, new_n8159_1, new_n8160);
not_8  g05812(n26882, new_n8161);
nor_5  g05813(new_n8161, n15271, new_n8162);
not_8  g05814(n25877, new_n8163);
nor_5  g05815(new_n8163, n22619, new_n8164);
not_8  g05816(n22619, new_n8165);
nor_5  g05817(n25877, new_n8165, new_n8166);
nand_5 g05818(n24323, new_n6107, new_n8167);
nor_5  g05819(new_n8167, new_n8166, new_n8168);
nor_5  g05820(new_n8168, new_n8164, new_n8169);
nor_5  g05821(new_n8169, new_n8162, new_n8170);
nor_5  g05822(new_n8170, new_n8160, new_n8171);
nand_5 g05823(new_n8171, new_n8158, new_n8172);
not_8  g05824(new_n8172, new_n8173);
nor_5  g05825(new_n8173, new_n8157, new_n8174);
nor_5  g05826(new_n8174, new_n8155, new_n8175);
nor_5  g05827(new_n8175, new_n8153, new_n8176);
not_8  g05828(new_n8176, new_n8177);
nand_5 g05829(new_n8177, new_n8151, new_n8178);
nand_5 g05830(new_n8178, new_n8150, new_n8179_1);
nand_5 g05831(new_n8179_1, new_n8149_1, new_n8180);
nand_5 g05832(new_n8180, new_n8148_1, new_n8181);
nand_5 g05833(new_n8181, new_n8146, new_n8182);
nand_5 g05834(new_n8182, new_n8145, new_n8183);
nand_5 g05835(new_n8183, new_n8144, new_n8184);
nand_5 g05836(new_n8184, new_n8143, new_n8185);
nand_5 g05837(new_n8185, new_n8142, new_n8186);
nand_5 g05838(new_n8186, new_n8141, new_n8187);
xnor_4 g05839(new_n8187, new_n8140, new_n8188);
not_8  g05840(new_n8188, new_n8189);
xnor_4 g05841(new_n8185, new_n8142, new_n8190);
xnor_4 g05842(new_n8137, new_n8094, new_n8191);
nand_5 g05843(new_n8191, new_n8190, new_n8192);
not_8  g05844(new_n8190, new_n8193);
xnor_4 g05845(new_n8191, new_n8193, new_n8194_1);
not_8  g05846(new_n8144, new_n8195);
xnor_4 g05847(new_n8183, new_n8195, new_n8196);
not_8  g05848(new_n8196, new_n8197);
xnor_4 g05849(new_n8135_1, new_n8096, new_n8198);
nand_5 g05850(new_n8198, new_n8197, new_n8199);
xnor_4 g05851(new_n8198, new_n8196, new_n8200);
xnor_4 g05852(new_n8181, new_n8146, new_n8201);
xnor_4 g05853(new_n8133, new_n8098, new_n8202);
nand_5 g05854(new_n8202, new_n8201, new_n8203);
xnor_4 g05855(new_n8202, new_n8201, new_n8204);
not_8  g05856(new_n8204, new_n8205);
xnor_4 g05857(new_n8179_1, new_n8149_1, new_n8206);
xnor_4 g05858(new_n8131, new_n8100, new_n8207);
nand_5 g05859(new_n8207, new_n8206, new_n8208);
not_8  g05860(new_n8206, new_n8209);
xnor_4 g05861(new_n8207, new_n8209, new_n8210);
xnor_4 g05862(new_n8176, new_n8151, new_n8211);
not_8  g05863(new_n8211, new_n8212);
xnor_4 g05864(new_n8128, new_n8103_1, new_n8213);
not_8  g05865(new_n8213, new_n8214);
nand_5 g05866(new_n8214, new_n8212, new_n8215_1);
xnor_4 g05867(new_n8214, new_n8211, new_n8216);
xnor_4 g05868(new_n8174, new_n8154, new_n8217);
not_8  g05869(new_n8217, new_n8218);
xnor_4 g05870(new_n8126, new_n8105, new_n8219);
not_8  g05871(new_n8219, new_n8220);
nand_5 g05872(new_n8220, new_n8218, new_n8221);
xnor_4 g05873(new_n8220, new_n8217, new_n8222);
xnor_4 g05874(new_n8171, new_n8158, new_n8223);
xnor_4 g05875(new_n8124, new_n8108, new_n8224);
not_8  g05876(new_n8224, new_n8225);
nand_5 g05877(new_n8225, new_n8223, new_n8226);
xnor_4 g05878(new_n8224, new_n8223, new_n8227);
xnor_4 g05879(n26882, n15271, new_n8228);
xnor_4 g05880(new_n8228, new_n8169, new_n8229);
xnor_4 g05881(n16722, n6385, new_n8230);
not_8  g05882(new_n8230, new_n8231);
xnor_4 g05883(new_n8231, new_n8122, new_n8232);
nand_5 g05884(new_n8232, new_n8229, new_n8233);
not_8  g05885(new_n8229, new_n8234);
xnor_4 g05886(new_n8232, new_n8234, new_n8235);
xnor_4 g05887(n25877, n22619, new_n8236);
xnor_4 g05888(new_n8236, new_n8167, new_n8237);
not_8  g05889(new_n8237, new_n8238);
xnor_4 g05890(n20138, n11486, new_n8239);
xnor_4 g05891(new_n8239, new_n8120, new_n8240);
nor_5  g05892(new_n8240, new_n8238, new_n8241);
xnor_4 g05893(n24323, n6775, new_n8242);
xnor_4 g05894(n13781, n9251, new_n8243);
nor_5  g05895(new_n8243, new_n8242, new_n8244_1);
xnor_4 g05896(new_n8240, new_n8237, new_n8245);
not_8  g05897(new_n8245, new_n8246);
nor_5  g05898(new_n8246, new_n8244_1, new_n8247);
nor_5  g05899(new_n8247, new_n8241, new_n8248);
not_8  g05900(new_n8248, new_n8249);
nand_5 g05901(new_n8249, new_n8235, new_n8250);
nand_5 g05902(new_n8250, new_n8233, new_n8251);
nand_5 g05903(new_n8251, new_n8227, new_n8252);
nand_5 g05904(new_n8252, new_n8226, new_n8253);
nand_5 g05905(new_n8253, new_n8222, new_n8254);
nand_5 g05906(new_n8254, new_n8221, new_n8255_1);
nand_5 g05907(new_n8255_1, new_n8216, new_n8256_1);
nand_5 g05908(new_n8256_1, new_n8215_1, new_n8257);
nand_5 g05909(new_n8257, new_n8210, new_n8258);
nand_5 g05910(new_n8258, new_n8208, new_n8259_1);
nand_5 g05911(new_n8259_1, new_n8205, new_n8260);
nand_5 g05912(new_n8260, new_n8203, new_n8261);
nand_5 g05913(new_n8261, new_n8200, new_n8262);
nand_5 g05914(new_n8262, new_n8199, new_n8263);
nand_5 g05915(new_n8263, new_n8194_1, new_n8264);
nand_5 g05916(new_n8264, new_n8192, new_n8265);
xnor_4 g05917(new_n8265, new_n8189, new_n8266);
not_8  g05918(n26408, new_n8267_1);
not_8  g05919(n13453, new_n8268);
nor_5  g05920(n15508, n2809, new_n8269);
nand_5 g05921(new_n8269, new_n6960, new_n8270);
nor_5  g05922(new_n8270, n7421, new_n8271);
nand_5 g05923(new_n8271, new_n8268, new_n8272);
nor_5  g05924(new_n8272, n11630, new_n8273);
nand_5 g05925(new_n8273, new_n5053, new_n8274);
nor_5  g05926(new_n8274, n18227, new_n8275);
nand_5 g05927(new_n8275, new_n8267_1, new_n8276_1);
or_5   g05928(new_n8276_1, n9554, new_n8277);
not_8  g05929(n9554, new_n8278);
xnor_4 g05930(new_n8276_1, new_n8278, new_n8279);
or_5   g05931(new_n8279, n9259, new_n8280);
xnor_4 g05932(new_n8275, n26408, new_n8281);
or_5   g05933(new_n8281, n21489, new_n8282);
xnor_4 g05934(new_n8281, new_n3724, new_n8283);
xnor_4 g05935(new_n8274, new_n5049, new_n8284);
or_5   g05936(new_n8284, n20213, new_n8285_1);
xnor_4 g05937(new_n8284, new_n3746, new_n8286);
xnor_4 g05938(new_n8273, n7377, new_n8287);
or_5   g05939(new_n8287, n13912, new_n8288_1);
xnor_4 g05940(new_n8287, new_n3725_1, new_n8289);
not_8  g05941(n11630, new_n8290);
xnor_4 g05942(new_n8272, new_n8290, new_n8291);
not_8  g05943(new_n8291, new_n8292);
nand_5 g05944(new_n8292, new_n3757, new_n8293);
xnor_4 g05945(new_n8291, new_n3757, new_n8294);
xnor_4 g05946(new_n8271, n13453, new_n8295);
not_8  g05947(new_n8295, new_n8296);
nand_5 g05948(new_n8296, new_n3726, new_n8297);
xnor_4 g05949(new_n8295, new_n3726, new_n8298);
not_8  g05950(n7421, new_n8299);
xnor_4 g05951(new_n8270, new_n8299, new_n8300);
not_8  g05952(new_n8300, new_n8301);
nand_5 g05953(new_n8301, new_n3768, new_n8302);
xnor_4 g05954(new_n8269, n19680, new_n8303);
not_8  g05955(new_n8303, new_n8304);
nand_5 g05956(new_n8304, new_n3727, new_n8305_1);
xnor_4 g05957(new_n8303, new_n3727, new_n8306_1);
xnor_4 g05958(n15508, n2809, new_n8307);
nand_5 g05959(new_n8307, new_n5121, new_n8308);
nand_5 g05960(n21993, n15508, new_n8309_1);
xnor_4 g05961(new_n8307, n25565, new_n8310);
nand_5 g05962(new_n8310, new_n8309_1, new_n8311);
nand_5 g05963(new_n8311, new_n8308, new_n8312);
nand_5 g05964(new_n8312, new_n8306_1, new_n8313);
nand_5 g05965(new_n8313, new_n8305_1, new_n8314);
xnor_4 g05966(new_n8300, new_n3768, new_n8315);
nand_5 g05967(new_n8315, new_n8314, new_n8316);
nand_5 g05968(new_n8316, new_n8302, new_n8317);
nand_5 g05969(new_n8317, new_n8298, new_n8318);
nand_5 g05970(new_n8318, new_n8297, new_n8319);
nand_5 g05971(new_n8319, new_n8294, new_n8320_1);
nand_5 g05972(new_n8320_1, new_n8293, new_n8321_1);
nand_5 g05973(new_n8321_1, new_n8289, new_n8322);
nand_5 g05974(new_n8322, new_n8288_1, new_n8323);
nand_5 g05975(new_n8323, new_n8286, new_n8324_1);
nand_5 g05976(new_n8324_1, new_n8285_1, new_n8325);
nand_5 g05977(new_n8325, new_n8283, new_n8326);
nand_5 g05978(new_n8326, new_n8282, new_n8327);
nand_5 g05979(new_n8279, n9259, new_n8328);
nand_5 g05980(new_n8328, new_n8327, new_n8329);
nand_5 g05981(new_n8329, new_n8280, new_n8330);
nand_5 g05982(new_n8330, new_n8277, new_n8331);
xnor_4 g05983(new_n8331, new_n8266, new_n8332);
not_8  g05984(new_n8332, new_n8333);
xnor_4 g05985(new_n8263, new_n8194_1, new_n8334);
not_8  g05986(new_n8334, new_n8335);
xnor_4 g05987(new_n8279, new_n3723, new_n8336);
not_8  g05988(new_n8336, new_n8337);
xnor_4 g05989(new_n8337, new_n8327, new_n8338);
nand_5 g05990(new_n8338, new_n8335, new_n8339_1);
xnor_4 g05991(new_n8338, new_n8334, new_n8340);
xnor_4 g05992(new_n8261, new_n8200, new_n8341);
not_8  g05993(new_n8341, new_n8342);
not_8  g05994(new_n8283, new_n8343);
xnor_4 g05995(new_n8325, new_n8343, new_n8344);
nor_5  g05996(new_n8344, new_n8342, new_n8345);
xnor_4 g05997(new_n8344, new_n8342, new_n8346);
xnor_4 g05998(new_n8259_1, new_n8204, new_n8347);
not_8  g05999(new_n8286, new_n8348);
xnor_4 g06000(new_n8323, new_n8348, new_n8349);
nor_5  g06001(new_n8349, new_n8347, new_n8350);
xnor_4 g06002(new_n8349, new_n8347, new_n8351);
xnor_4 g06003(new_n8257, new_n8210, new_n8352);
not_8  g06004(new_n8352, new_n8353);
xnor_4 g06005(new_n8321_1, new_n8289, new_n8354);
not_8  g06006(new_n8354, new_n8355);
nand_5 g06007(new_n8355, new_n8353, new_n8356);
nand_5 g06008(new_n8354, new_n8352, new_n8357);
not_8  g06009(new_n8255_1, new_n8358);
xnor_4 g06010(new_n8358, new_n8216, new_n8359);
xnor_4 g06011(new_n8319, new_n8294, new_n8360);
not_8  g06012(new_n8360, new_n8361);
nand_5 g06013(new_n8361, new_n8359, new_n8362);
xnor_4 g06014(new_n8360, new_n8359, new_n8363_1);
xnor_4 g06015(new_n8317, new_n8298, new_n8364);
not_8  g06016(new_n8364, new_n8365);
not_8  g06017(new_n8222, new_n8366);
xnor_4 g06018(new_n8253, new_n8366, new_n8367);
nand_5 g06019(new_n8367, new_n8365, new_n8368);
xnor_4 g06020(new_n8367, new_n8364, new_n8369);
xnor_4 g06021(new_n8251, new_n8227, new_n8370);
xnor_4 g06022(new_n8315, new_n8314, new_n8371);
nor_5  g06023(new_n8371, new_n8370, new_n8372);
not_8  g06024(new_n8372, new_n8373);
not_8  g06025(new_n8370, new_n8374);
not_8  g06026(new_n8371, new_n8375);
nor_5  g06027(new_n8375, new_n8374, new_n8376_1);
not_8  g06028(new_n8376_1, new_n8377);
xnor_4 g06029(new_n8248, new_n8235, new_n8378);
xnor_4 g06030(new_n8245, new_n8244_1, new_n8379);
not_8  g06031(new_n8379, new_n8380);
xnor_4 g06032(new_n8310, new_n8309_1, new_n8381_1);
nor_5  g06033(new_n8381_1, new_n8380, new_n8382);
xnor_4 g06034(n21993, new_n5125, new_n8383);
not_8  g06035(new_n8383, new_n8384);
not_8  g06036(new_n8242, new_n8385);
xnor_4 g06037(new_n8243, new_n8385, new_n8386);
not_8  g06038(new_n8386, new_n8387);
nor_5  g06039(new_n8387, new_n8384, new_n8388);
xnor_4 g06040(new_n8381_1, new_n8379, new_n8389);
not_8  g06041(new_n8389, new_n8390);
nor_5  g06042(new_n8390, new_n8388, new_n8391);
nor_5  g06043(new_n8391, new_n8382, new_n8392);
not_8  g06044(new_n8392, new_n8393);
nor_5  g06045(new_n8393, new_n8378, new_n8394);
xnor_4 g06046(new_n8312, new_n8306_1, new_n8395);
not_8  g06047(new_n8395, new_n8396);
not_8  g06048(new_n8378, new_n8397);
xnor_4 g06049(new_n8392, new_n8397, new_n8398);
nor_5  g06050(new_n8398, new_n8396, new_n8399_1);
nor_5  g06051(new_n8399_1, new_n8394, new_n8400);
nand_5 g06052(new_n8400, new_n8377, new_n8401);
nand_5 g06053(new_n8401, new_n8373, new_n8402);
nand_5 g06054(new_n8402, new_n8369, new_n8403);
nand_5 g06055(new_n8403, new_n8368, new_n8404);
nand_5 g06056(new_n8404, new_n8363_1, new_n8405_1);
nand_5 g06057(new_n8405_1, new_n8362, new_n8406);
nand_5 g06058(new_n8406, new_n8357, new_n8407);
nand_5 g06059(new_n8407, new_n8356, new_n8408_1);
nor_5  g06060(new_n8408_1, new_n8351, new_n8409);
nor_5  g06061(new_n8409, new_n8350, new_n8410);
nor_5  g06062(new_n8410, new_n8346, new_n8411);
nor_5  g06063(new_n8411, new_n8345, new_n8412);
nand_5 g06064(new_n8412, new_n8340, new_n8413);
nand_5 g06065(new_n8413, new_n8339_1, new_n8414);
xnor_4 g06066(new_n8414, new_n8333, n829);
not_8  g06067(n22764, new_n8416);
not_8  g06068(n14826, new_n8417_1);
xnor_4 g06069(n23272, new_n8417_1, new_n8418);
or_5   g06070(n23493, n11481, new_n8419);
xnor_4 g06071(n23493, new_n4552_1, new_n8420);
or_5   g06072(n16439, n10275, new_n8421);
not_8  g06073(n10275, new_n8422);
xnor_4 g06074(n16439, new_n8422, new_n8423);
nor_5  g06075(n15241, n15146, new_n8424);
not_8  g06076(n15146, new_n8425);
xnor_4 g06077(n15241, new_n8425, new_n8426);
not_8  g06078(new_n8426, new_n8427);
nor_5  g06079(n11579, n7678, new_n8428);
xnor_4 g06080(n11579, new_n4564, new_n8429);
not_8  g06081(new_n8429, new_n8430);
nor_5  g06082(n3785, n21, new_n8431);
not_8  g06083(n21, new_n8432_1);
xnor_4 g06084(n3785, new_n8432_1, new_n8433);
not_8  g06085(new_n8433, new_n8434);
nor_5  g06086(n20250, n1682, new_n8435);
not_8  g06087(n1682, new_n8436);
xnor_4 g06088(n20250, new_n8436, new_n8437);
not_8  g06089(new_n8437, new_n8438);
nor_5  g06090(n7963, n5822, new_n8439_1);
xnor_4 g06091(n7963, new_n4577, new_n8440);
not_8  g06092(new_n8440, new_n8441);
nor_5  g06093(n26443, n10017, new_n8442);
nand_5 g06094(n3618, n1681, new_n8443);
not_8  g06095(new_n8443, new_n8444);
xnor_4 g06096(n26443, n10017, new_n8445);
nor_5  g06097(new_n8445, new_n8444, new_n8446);
nor_5  g06098(new_n8446, new_n8442, new_n8447);
nor_5  g06099(new_n8447, new_n8441, new_n8448);
nor_5  g06100(new_n8448, new_n8439_1, new_n8449);
nor_5  g06101(new_n8449, new_n8438, new_n8450);
nor_5  g06102(new_n8450, new_n8435, new_n8451);
nor_5  g06103(new_n8451, new_n8434, new_n8452);
nor_5  g06104(new_n8452, new_n8431, new_n8453_1);
nor_5  g06105(new_n8453_1, new_n8430, new_n8454);
nor_5  g06106(new_n8454, new_n8428, new_n8455);
nor_5  g06107(new_n8455, new_n8427, new_n8456);
nor_5  g06108(new_n8456, new_n8424, new_n8457);
not_8  g06109(new_n8457, new_n8458);
nand_5 g06110(new_n8458, new_n8423, new_n8459);
nand_5 g06111(new_n8459, new_n8421, new_n8460);
nand_5 g06112(new_n8460, new_n8420, new_n8461);
nand_5 g06113(new_n8461, new_n8419, new_n8462);
xnor_4 g06114(new_n8462, new_n8418, new_n8463);
nand_5 g06115(new_n8463, new_n8416, new_n8464);
xnor_4 g06116(new_n8463, n22764, new_n8465);
not_8  g06117(n26264, new_n8466);
xnor_4 g06118(new_n8460, new_n8420, new_n8467);
nand_5 g06119(new_n8467, new_n8466, new_n8468);
xnor_4 g06120(new_n8467, n26264, new_n8469);
not_8  g06121(n7841, new_n8470);
xnor_4 g06122(new_n8457, new_n8423, new_n8471);
not_8  g06123(new_n8471, new_n8472);
nand_5 g06124(new_n8472, new_n8470, new_n8473);
xnor_4 g06125(new_n8471, new_n8470, new_n8474);
not_8  g06126(n16812, new_n8475);
xnor_4 g06127(new_n8455, new_n8426, new_n8476);
not_8  g06128(new_n8476, new_n8477);
nand_5 g06129(new_n8477, new_n8475, new_n8478);
xnor_4 g06130(new_n8476, new_n8475, new_n8479);
not_8  g06131(n25068, new_n8480_1);
xnor_4 g06132(new_n8453_1, new_n8429, new_n8481);
not_8  g06133(new_n8481, new_n8482);
nand_5 g06134(new_n8482, new_n8480_1, new_n8483);
xnor_4 g06135(new_n8481, new_n8480_1, new_n8484);
xnor_4 g06136(new_n8451, new_n8433, new_n8485);
nor_5  g06137(new_n8485, n2331, new_n8486);
not_8  g06138(new_n8486, new_n8487);
not_8  g06139(n2331, new_n8488);
xnor_4 g06140(new_n8485, new_n8488, new_n8489_1);
xnor_4 g06141(new_n8449, new_n8437, new_n8490);
nor_5  g06142(new_n8490, n22631, new_n8491);
not_8  g06143(new_n8491, new_n8492);
not_8  g06144(n22631, new_n8493);
xnor_4 g06145(new_n8490, new_n8493, new_n8494);
not_8  g06146(n16743, new_n8495);
xnor_4 g06147(new_n8447, new_n8440, new_n8496);
not_8  g06148(new_n8496, new_n8497);
nor_5  g06149(new_n8497, new_n8495, new_n8498);
xnor_4 g06150(new_n8496, new_n8495, new_n8499);
not_8  g06151(new_n8499, new_n8500);
not_8  g06152(n15258, new_n8501);
not_8  g06153(new_n2569, new_n8502);
nor_5  g06154(new_n8502, n4588, new_n8503);
nand_5 g06155(new_n8503, new_n8501, new_n8504);
xnor_4 g06156(new_n8445, new_n8443, new_n8505_1);
not_8  g06157(new_n8505_1, new_n8506);
xnor_4 g06158(new_n8503, n15258, new_n8507);
nand_5 g06159(new_n8507, new_n8506, new_n8508);
nand_5 g06160(new_n8508, new_n8504, new_n8509);
nor_5  g06161(new_n8509, new_n8500, new_n8510_1);
nor_5  g06162(new_n8510_1, new_n8498, new_n8511);
nand_5 g06163(new_n8511, new_n8494, new_n8512);
nand_5 g06164(new_n8512, new_n8492, new_n8513);
nand_5 g06165(new_n8513, new_n8489_1, new_n8514);
nand_5 g06166(new_n8514, new_n8487, new_n8515);
nand_5 g06167(new_n8515, new_n8484, new_n8516);
nand_5 g06168(new_n8516, new_n8483, new_n8517);
nand_5 g06169(new_n8517, new_n8479, new_n8518);
nand_5 g06170(new_n8518, new_n8478, new_n8519_1);
nand_5 g06171(new_n8519_1, new_n8474, new_n8520);
nand_5 g06172(new_n8520, new_n8473, new_n8521);
nand_5 g06173(new_n8521, new_n8469, new_n8522);
nand_5 g06174(new_n8522, new_n8468, new_n8523);
nand_5 g06175(new_n8523, new_n8465, new_n8524);
nand_5 g06176(new_n8524, new_n8464, new_n8525);
or_5   g06177(n23272, n14826, new_n8526_1);
nand_5 g06178(new_n8462, new_n8418, new_n8527);
nand_5 g06179(new_n8527, new_n8526_1, new_n8528);
not_8  g06180(new_n8528, new_n8529);
nor_5  g06181(new_n8529, new_n8525, new_n8530);
or_5   g06182(n18105, new_n5905, new_n8531);
xnor_4 g06183(n18105, n12702, new_n8532);
or_5   g06184(new_n5906, n24196, new_n8533);
xnor_4 g06185(n26797, n24196, new_n8534);
or_5   g06186(new_n5851, n16376, new_n8535_1);
xnor_4 g06187(n23913, n16376, new_n8536);
or_5   g06188(n25381, new_n5836, new_n8537);
xnor_4 g06189(n25381, n22554, new_n8538);
or_5   g06190(new_n5862, n12587, new_n8539);
xnor_4 g06191(n20429, n12587, new_n8540);
nor_5  g06192(new_n5837, n268, new_n8541);
not_8  g06193(new_n8541, new_n8542);
xnor_4 g06194(n3909, n268, new_n8543);
nor_5  g06195(n24879, new_n5873, new_n8544);
not_8  g06196(new_n8544, new_n8545);
xnor_4 g06197(n24879, n23974, new_n8546);
nor_5  g06198(new_n4650, n2146, new_n8547);
nor_5  g06199(n6785, new_n5838, new_n8548);
not_8  g06200(n24032, new_n8549);
nor_5  g06201(new_n8549, n22173, new_n8550_1);
nor_5  g06202(new_n4704, n583, new_n8551);
not_8  g06203(new_n8551, new_n8552);
not_8  g06204(n22173, new_n8553);
nor_5  g06205(n24032, new_n8553, new_n8554);
nor_5  g06206(new_n8554, new_n8552, new_n8555);
nor_5  g06207(new_n8555, new_n8550_1, new_n8556);
nor_5  g06208(new_n8556, new_n8548, new_n8557);
nor_5  g06209(new_n8557, new_n8547, new_n8558);
nand_5 g06210(new_n8558, new_n8546, new_n8559);
nand_5 g06211(new_n8559, new_n8545, new_n8560);
nand_5 g06212(new_n8560, new_n8543, new_n8561);
nand_5 g06213(new_n8561, new_n8542, new_n8562);
nand_5 g06214(new_n8562, new_n8540, new_n8563_1);
nand_5 g06215(new_n8563_1, new_n8539, new_n8564);
nand_5 g06216(new_n8564, new_n8538, new_n8565);
nand_5 g06217(new_n8565, new_n8537, new_n8566);
nand_5 g06218(new_n8566, new_n8536, new_n8567);
nand_5 g06219(new_n8567, new_n8535_1, new_n8568);
nand_5 g06220(new_n8568, new_n8534, new_n8569);
nand_5 g06221(new_n8569, new_n8533, new_n8570);
nand_5 g06222(new_n8570, new_n8532, new_n8571);
nand_5 g06223(new_n8571, new_n8531, new_n8572);
not_8  g06224(n1536, new_n8573);
xnor_4 g06225(new_n8570, new_n8532, new_n8574);
nand_5 g06226(new_n8574, new_n8573, new_n8575);
xnor_4 g06227(new_n8574, n1536, new_n8576);
not_8  g06228(n19454, new_n8577);
xnor_4 g06229(new_n8568, new_n8534, new_n8578);
nand_5 g06230(new_n8578, new_n8577, new_n8579);
xnor_4 g06231(new_n8578, n19454, new_n8580);
not_8  g06232(n9445, new_n8581_1);
xnor_4 g06233(new_n8566, new_n8536, new_n8582);
nand_5 g06234(new_n8582, new_n8581_1, new_n8583);
xnor_4 g06235(new_n8582, n9445, new_n8584);
not_8  g06236(n1279, new_n8585);
xnor_4 g06237(new_n8564, new_n8538, new_n8586);
nand_5 g06238(new_n8586, new_n8585, new_n8587);
xnor_4 g06239(new_n8586, n1279, new_n8588);
not_8  g06240(n8324, new_n8589);
xnor_4 g06241(new_n8562, new_n8540, new_n8590);
nand_5 g06242(new_n8590, new_n8589, new_n8591);
xnor_4 g06243(new_n8590, n8324, new_n8592);
not_8  g06244(n12546, new_n8593);
xnor_4 g06245(new_n8560, new_n8543, new_n8594_1);
nand_5 g06246(new_n8594_1, new_n8593, new_n8595);
xnor_4 g06247(new_n8594_1, n12546, new_n8596);
not_8  g06248(n21078, new_n8597);
xnor_4 g06249(new_n8558, new_n8546, new_n8598);
nand_5 g06250(new_n8598, new_n8597, new_n8599);
xnor_4 g06251(new_n8598, n21078, new_n8600);
not_8  g06252(n24485, new_n8601);
xnor_4 g06253(n6785, n2146, new_n8602);
xnor_4 g06254(new_n8602, new_n8556, new_n8603);
nor_5  g06255(new_n8603, new_n8601, new_n8604);
not_8  g06256(new_n8603, new_n8605);
nor_5  g06257(new_n8605, n24485, new_n8606);
xnor_4 g06258(n24032, n22173, new_n8607);
xnor_4 g06259(new_n8607, new_n8552, new_n8608_1);
not_8  g06260(new_n8608_1, new_n8609);
nor_5  g06261(new_n8609, n2420, new_n8610);
not_8  g06262(new_n8610, new_n8611);
not_8  g06263(n22201, new_n8612);
nor_5  g06264(new_n2571, new_n8612, new_n8613);
not_8  g06265(new_n8613, new_n8614_1);
xnor_4 g06266(new_n8608_1, n2420, new_n8615);
nand_5 g06267(new_n8615, new_n8614_1, new_n8616);
nand_5 g06268(new_n8616, new_n8611, new_n8617);
nor_5  g06269(new_n8617, new_n8606, new_n8618);
nor_5  g06270(new_n8618, new_n8604, new_n8619);
nand_5 g06271(new_n8619, new_n8600, new_n8620_1);
nand_5 g06272(new_n8620_1, new_n8599, new_n8621);
nand_5 g06273(new_n8621, new_n8596, new_n8622);
nand_5 g06274(new_n8622, new_n8595, new_n8623);
nand_5 g06275(new_n8623, new_n8592, new_n8624);
nand_5 g06276(new_n8624, new_n8591, new_n8625);
nand_5 g06277(new_n8625, new_n8588, new_n8626);
nand_5 g06278(new_n8626, new_n8587, new_n8627);
nand_5 g06279(new_n8627, new_n8584, new_n8628);
nand_5 g06280(new_n8628, new_n8583, new_n8629);
nand_5 g06281(new_n8629, new_n8580, new_n8630);
nand_5 g06282(new_n8630, new_n8579, new_n8631);
nand_5 g06283(new_n8631, new_n8576, new_n8632);
nand_5 g06284(new_n8632, new_n8575, new_n8633);
nor_5  g06285(new_n8633, new_n8572, new_n8634);
xnor_4 g06286(new_n8529, new_n8525, new_n8635);
not_8  g06287(new_n8572, new_n8636);
xnor_4 g06288(new_n8633, new_n8636, new_n8637_1);
not_8  g06289(new_n8637_1, new_n8638_1);
nand_5 g06290(new_n8638_1, new_n8635, new_n8639);
xnor_4 g06291(new_n8637_1, new_n8635, new_n8640);
xnor_4 g06292(new_n8523, new_n8465, new_n8641);
not_8  g06293(new_n8641, new_n8642);
xnor_4 g06294(new_n8574, new_n8573, new_n8643);
xnor_4 g06295(new_n8631, new_n8643, new_n8644);
nand_5 g06296(new_n8644, new_n8642, new_n8645);
xnor_4 g06297(new_n8644, new_n8641, new_n8646);
xnor_4 g06298(new_n8521, new_n8469, new_n8647);
not_8  g06299(new_n8647, new_n8648);
xnor_4 g06300(new_n8578, new_n8577, new_n8649);
xnor_4 g06301(new_n8629, new_n8649, new_n8650);
nand_5 g06302(new_n8650, new_n8648, new_n8651);
xnor_4 g06303(new_n8650, new_n8647, new_n8652);
not_8  g06304(new_n8474, new_n8653);
xnor_4 g06305(new_n8519_1, new_n8653, new_n8654);
xnor_4 g06306(new_n8627, new_n8584, new_n8655);
not_8  g06307(new_n8655, new_n8656_1);
nand_5 g06308(new_n8656_1, new_n8654, new_n8657);
xnor_4 g06309(new_n8655, new_n8654, new_n8658);
xnor_4 g06310(new_n8517, new_n8479, new_n8659);
not_8  g06311(new_n8659, new_n8660);
xnor_4 g06312(new_n8586, new_n8585, new_n8661);
xnor_4 g06313(new_n8625, new_n8661, new_n8662_1);
nand_5 g06314(new_n8662_1, new_n8660, new_n8663);
xnor_4 g06315(new_n8662_1, new_n8659, new_n8664);
xnor_4 g06316(new_n8515, new_n8484, new_n8665);
not_8  g06317(new_n8665, new_n8666);
xnor_4 g06318(new_n8623, new_n8592, new_n8667);
not_8  g06319(new_n8667, new_n8668);
nand_5 g06320(new_n8668, new_n8666, new_n8669);
xnor_4 g06321(new_n8668, new_n8665, new_n8670);
xnor_4 g06322(new_n8513, new_n8489_1, new_n8671);
not_8  g06323(new_n8671, new_n8672);
not_8  g06324(new_n8596, new_n8673);
xnor_4 g06325(new_n8621, new_n8673, new_n8674);
nand_5 g06326(new_n8674, new_n8672, new_n8675);
xnor_4 g06327(new_n8674, new_n8671, new_n8676);
xnor_4 g06328(new_n8511, new_n8494, new_n8677);
xnor_4 g06329(new_n8619, new_n8600, new_n8678_1);
nor_5  g06330(new_n8678_1, new_n8677, new_n8679);
not_8  g06331(new_n8679, new_n8680);
not_8  g06332(new_n8677, new_n8681);
xnor_4 g06333(new_n8678_1, new_n8681, new_n8682);
xnor_4 g06334(new_n8509, new_n8499, new_n8683);
xnor_4 g06335(new_n8603, n24485, new_n8684);
xnor_4 g06336(new_n8684, new_n8617, new_n8685);
nor_5  g06337(new_n8685, new_n8683, new_n8686);
not_8  g06338(new_n8686, new_n8687_1);
not_8  g06339(new_n8683, new_n8688);
xnor_4 g06340(new_n8685, new_n8688, new_n8689);
xnor_4 g06341(new_n8615, new_n8613, new_n8690);
xnor_4 g06342(new_n8507, new_n8505_1, new_n8691);
nor_5  g06343(new_n8691, new_n8690, new_n8692);
not_8  g06344(new_n2570_1, new_n8693);
nand_5 g06345(new_n2572, new_n8693, new_n8694_1);
xnor_4 g06346(new_n8691, new_n8690, new_n8695);
nor_5  g06347(new_n8695, new_n8694_1, new_n8696);
nor_5  g06348(new_n8696, new_n8692, new_n8697);
nand_5 g06349(new_n8697, new_n8689, new_n8698);
nand_5 g06350(new_n8698, new_n8687_1, new_n8699);
nand_5 g06351(new_n8699, new_n8682, new_n8700);
nand_5 g06352(new_n8700, new_n8680, new_n8701);
nand_5 g06353(new_n8701, new_n8676, new_n8702);
nand_5 g06354(new_n8702, new_n8675, new_n8703);
nand_5 g06355(new_n8703, new_n8670, new_n8704);
nand_5 g06356(new_n8704, new_n8669, new_n8705);
nand_5 g06357(new_n8705, new_n8664, new_n8706);
nand_5 g06358(new_n8706, new_n8663, new_n8707);
nand_5 g06359(new_n8707, new_n8658, new_n8708);
nand_5 g06360(new_n8708, new_n8657, new_n8709);
nand_5 g06361(new_n8709, new_n8652, new_n8710);
nand_5 g06362(new_n8710, new_n8651, new_n8711);
nand_5 g06363(new_n8711, new_n8646, new_n8712);
nand_5 g06364(new_n8712, new_n8645, new_n8713);
nand_5 g06365(new_n8713, new_n8640, new_n8714);
nand_5 g06366(new_n8714, new_n8639, new_n8715);
xnor_4 g06367(new_n8715, new_n8634, new_n8716_1);
xnor_4 g06368(new_n8716_1, new_n8530, n849);
xnor_4 g06369(new_n2556, new_n2555_1, n858);
not_8  g06370(n22442, new_n8719);
not_8  g06371(n1314, new_n8720);
not_8  g06372(n24638, new_n8721_1);
nor_5  g06373(n16994, n9246, new_n8722);
nand_5 g06374(new_n8722, new_n3694, new_n8723);
nor_5  g06375(new_n8723, n14790, new_n8724);
nand_5 g06376(new_n8724, new_n5008, new_n8725);
nor_5  g06377(new_n8725, n21674, new_n8726);
nand_5 g06378(new_n8726, new_n8721_1, new_n8727);
nor_5  g06379(new_n8727, n18444, new_n8728);
nand_5 g06380(new_n8728, new_n4995, new_n8729);
xnor_4 g06381(new_n8729, new_n4992, new_n8730);
xnor_4 g06382(new_n8730, new_n8720, new_n8731);
xnor_4 g06383(new_n8728, n14899, new_n8732);
and_5  g06384(new_n8732, n3306, new_n8733);
nor_5  g06385(new_n8732, n3306, new_n8734);
not_8  g06386(n22335, new_n8735);
xnor_4 g06387(new_n8727, new_n4998, new_n8736);
not_8  g06388(new_n8736, new_n8737);
nand_5 g06389(new_n8737, new_n8735, new_n8738);
xnor_4 g06390(new_n8736, new_n8735, new_n8739);
not_8  g06391(n24048, new_n8740);
xnor_4 g06392(new_n8726, n24638, new_n8741);
not_8  g06393(new_n8741, new_n8742);
nand_5 g06394(new_n8742, new_n8740, new_n8743);
xnor_4 g06395(new_n8741, new_n8740, new_n8744_1);
not_8  g06396(n1525, new_n8745_1);
xnor_4 g06397(new_n8725, new_n5004, new_n8746);
not_8  g06398(new_n8746, new_n8747);
nand_5 g06399(new_n8747, new_n8745_1, new_n8748);
xnor_4 g06400(new_n8746, new_n8745_1, new_n8749);
xnor_4 g06401(new_n8724, n17251, new_n8750);
not_8  g06402(new_n8750, new_n8751);
nand_5 g06403(new_n8751, new_n4850_1, new_n8752);
xnor_4 g06404(new_n8750, new_n4850_1, new_n8753);
not_8  g06405(n14790, new_n8754);
xnor_4 g06406(new_n8723, new_n8754, new_n8755);
not_8  g06407(new_n8755, new_n8756);
nand_5 g06408(new_n8756, new_n4854, new_n8757);
xnor_4 g06409(new_n8722, n10096, new_n8758);
not_8  g06410(new_n8758, new_n8759);
nand_5 g06411(new_n8759, new_n4858_1, new_n8760);
xnor_4 g06412(new_n8758, new_n4858_1, new_n8761);
xnor_4 g06413(n16994, n9246, new_n8762);
nand_5 g06414(new_n8762, new_n4861, new_n8763);
nand_5 g06415(n23120, n9246, new_n8764);
xnor_4 g06416(new_n8762, n5128, new_n8765);
nand_5 g06417(new_n8765, new_n8764, new_n8766);
nand_5 g06418(new_n8766, new_n8763, new_n8767);
nand_5 g06419(new_n8767, new_n8761, new_n8768);
nand_5 g06420(new_n8768, new_n8760, new_n8769);
xnor_4 g06421(new_n8755, new_n4854, new_n8770);
nand_5 g06422(new_n8770, new_n8769, new_n8771);
nand_5 g06423(new_n8771, new_n8757, new_n8772);
nand_5 g06424(new_n8772, new_n8753, new_n8773);
nand_5 g06425(new_n8773, new_n8752, new_n8774);
nand_5 g06426(new_n8774, new_n8749, new_n8775);
nand_5 g06427(new_n8775, new_n8748, new_n8776);
nand_5 g06428(new_n8776, new_n8744_1, new_n8777);
nand_5 g06429(new_n8777, new_n8743, new_n8778);
nand_5 g06430(new_n8778, new_n8739, new_n8779);
nand_5 g06431(new_n8779, new_n8738, new_n8780);
nor_5  g06432(new_n8780, new_n8734, new_n8781);
nor_5  g06433(new_n8781, new_n8733, new_n8782_1);
xnor_4 g06434(new_n8782_1, new_n8731, new_n8783);
nand_5 g06435(new_n8783, new_n8719, new_n8784);
xnor_4 g06436(new_n8783, n22442, new_n8785);
not_8  g06437(n3306, new_n8786);
xnor_4 g06438(new_n8732, new_n8786, new_n8787);
xnor_4 g06439(new_n8787, new_n8780, new_n8788);
nor_5  g06440(new_n8788, new_n7404, new_n8789);
xnor_4 g06441(new_n8788, n468, new_n8790);
not_8  g06442(new_n8790, new_n8791);
xnor_4 g06443(new_n8778, new_n8739, new_n8792);
nand_5 g06444(new_n8792, new_n7408_1, new_n8793);
xnor_4 g06445(new_n8792, n5400, new_n8794);
not_8  g06446(n23923, new_n8795);
xnor_4 g06447(new_n8776, new_n8744_1, new_n8796);
nand_5 g06448(new_n8796, new_n8795, new_n8797);
xnor_4 g06449(new_n8796, n23923, new_n8798);
xnor_4 g06450(new_n8774, new_n8749, new_n8799);
nor_5  g06451(new_n8799, new_n7415, new_n8800);
not_8  g06452(new_n8799, new_n8801);
nor_5  g06453(new_n8801, n329, new_n8802);
not_8  g06454(n24170, new_n8803_1);
xnor_4 g06455(new_n8770, new_n8769, new_n8804);
nand_5 g06456(new_n8804, new_n7422, new_n8805);
xnor_4 g06457(new_n8804, n2409, new_n8806_1);
not_8  g06458(n8869, new_n8807);
xnor_4 g06459(new_n8767, new_n8761, new_n8808);
nand_5 g06460(new_n8808, new_n8807, new_n8809_1);
xnor_4 g06461(new_n8765, new_n8764, new_n8810);
nand_5 g06462(new_n8810, new_n7431, new_n8811);
xnor_4 g06463(n23120, n9246, new_n8812);
nand_5 g06464(new_n8812, n7428, new_n8813);
xnor_4 g06465(new_n8810, n10372, new_n8814);
nand_5 g06466(new_n8814, new_n8813, new_n8815);
nand_5 g06467(new_n8815, new_n8811, new_n8816);
xnor_4 g06468(new_n8808, n8869, new_n8817);
nand_5 g06469(new_n8817, new_n8816, new_n8818);
nand_5 g06470(new_n8818, new_n8809_1, new_n8819);
nand_5 g06471(new_n8819, new_n8806_1, new_n8820);
nand_5 g06472(new_n8820, new_n8805, new_n8821_1);
nand_5 g06473(new_n8821_1, new_n8803_1, new_n8822);
xnor_4 g06474(new_n8772, new_n8753, new_n8823);
xnor_4 g06475(new_n8821_1, n24170, new_n8824_1);
nand_5 g06476(new_n8824_1, new_n8823, new_n8825);
nand_5 g06477(new_n8825, new_n8822, new_n8826);
nor_5  g06478(new_n8826, new_n8802, new_n8827_1);
nor_5  g06479(new_n8827_1, new_n8800, new_n8828);
nand_5 g06480(new_n8828, new_n8798, new_n8829);
nand_5 g06481(new_n8829, new_n8797, new_n8830);
nand_5 g06482(new_n8830, new_n8794, new_n8831);
nand_5 g06483(new_n8831, new_n8793, new_n8832);
nor_5  g06484(new_n8832, new_n8791, new_n8833);
nor_5  g06485(new_n8833, new_n8789, new_n8834);
nand_5 g06486(new_n8834, new_n8785, new_n8835);
nand_5 g06487(new_n8835, new_n8784, new_n8836);
nor_5  g06488(new_n8730, n1314, new_n8837);
nor_5  g06489(new_n8782_1, new_n8837, new_n8838);
nor_5  g06490(new_n8729, n3506, new_n8839);
and_5  g06491(new_n8730, n1314, new_n8840);
nor_5  g06492(new_n8840, new_n8839, new_n8841);
not_8  g06493(new_n8841, new_n8842);
nor_5  g06494(new_n8842, new_n8838, new_n8843);
xnor_4 g06495(new_n8843, new_n8836, new_n8844);
not_8  g06496(new_n3607, new_n8845);
nand_5 g06497(new_n8845, new_n3532, new_n8846);
nand_5 g06498(new_n3671, new_n3608, new_n8847);
nand_5 g06499(new_n8847, new_n8846, new_n8848);
or_5   g06500(new_n3544, n8856, new_n8849_1);
or_5   g06501(new_n3545, n25494, new_n8850);
nand_5 g06502(new_n3545, n25494, new_n8851);
nand_5 g06503(new_n3606, new_n8851, new_n8852);
nand_5 g06504(new_n8852, new_n8850, new_n8853);
nand_5 g06505(new_n8853, new_n8849_1, new_n8854);
not_8  g06506(new_n8854, new_n8855);
xnor_4 g06507(new_n8855, new_n8848, new_n8856_1);
not_8  g06508(new_n8856_1, new_n8857);
xnor_4 g06509(new_n8857, new_n8844, new_n8858);
xnor_4 g06510(new_n8834, new_n8785, new_n8859);
nand_5 g06511(new_n8859, new_n3673, new_n8860);
xnor_4 g06512(new_n8859, new_n3672, new_n8861_1);
xnor_4 g06513(new_n8832, new_n8790, new_n8862_1);
nand_5 g06514(new_n8862_1, new_n3810, new_n8863);
xnor_4 g06515(new_n8862_1, new_n3809, new_n8864);
xnor_4 g06516(new_n8830, new_n8794, new_n8865);
nand_5 g06517(new_n8865, new_n3817, new_n8866);
xnor_4 g06518(new_n8865, new_n3816, new_n8867);
xnor_4 g06519(new_n8828, new_n8798, new_n8868);
nand_5 g06520(new_n8868, new_n3823, new_n8869_1);
xnor_4 g06521(new_n8799, n329, new_n8870);
xnor_4 g06522(new_n8870, new_n8826, new_n8871);
nand_5 g06523(new_n8871, new_n3829, new_n8872);
xnor_4 g06524(new_n8871, new_n3828_1, new_n8873);
xnor_4 g06525(new_n8824_1, new_n8823, new_n8874);
nand_5 g06526(new_n8874, new_n3835, new_n8875);
not_8  g06527(new_n3841, new_n8876);
not_8  g06528(new_n8806_1, new_n8877);
xnor_4 g06529(new_n8819, new_n8877, new_n8878);
nor_5  g06530(new_n8878, new_n8876, new_n8879);
not_8  g06531(new_n8879, new_n8880);
xnor_4 g06532(new_n8878, new_n3841, new_n8881);
xnor_4 g06533(new_n8817, new_n8816, new_n8882);
not_8  g06534(new_n8882, new_n8883);
nor_5  g06535(new_n8883, new_n3846, new_n8884_1);
not_8  g06536(new_n8884_1, new_n8885);
not_8  g06537(new_n8813, new_n8886);
xnor_4 g06538(new_n8814, new_n8886, new_n8887);
nor_5  g06539(new_n8887, new_n3858, new_n8888);
not_8  g06540(new_n8888, new_n8889);
not_8  g06541(new_n3854, new_n8890);
xnor_4 g06542(new_n8812, new_n7504, new_n8891);
nor_5  g06543(new_n8891, new_n8890, new_n8892);
not_8  g06544(new_n8892, new_n8893);
xnor_4 g06545(new_n8887, new_n3852, new_n8894);
nand_5 g06546(new_n8894, new_n8893, new_n8895);
nand_5 g06547(new_n8895, new_n8889, new_n8896);
xnor_4 g06548(new_n8882, new_n3846, new_n8897);
nand_5 g06549(new_n8897, new_n8896, new_n8898);
nand_5 g06550(new_n8898, new_n8885, new_n8899);
nand_5 g06551(new_n8899, new_n8881, new_n8900);
nand_5 g06552(new_n8900, new_n8880, new_n8901);
xnor_4 g06553(new_n8874, new_n3834, new_n8902);
nand_5 g06554(new_n8902, new_n8901, new_n8903);
nand_5 g06555(new_n8903, new_n8875, new_n8904);
nand_5 g06556(new_n8904, new_n8873, new_n8905);
nand_5 g06557(new_n8905, new_n8872, new_n8906);
xnor_4 g06558(new_n8868, new_n3822, new_n8907);
nand_5 g06559(new_n8907, new_n8906, new_n8908);
nand_5 g06560(new_n8908, new_n8869_1, new_n8909_1);
nand_5 g06561(new_n8909_1, new_n8867, new_n8910);
nand_5 g06562(new_n8910, new_n8866, new_n8911_1);
nand_5 g06563(new_n8911_1, new_n8864, new_n8912);
nand_5 g06564(new_n8912, new_n8863, new_n8913);
nand_5 g06565(new_n8913, new_n8861_1, new_n8914);
nand_5 g06566(new_n8914, new_n8860, new_n8915);
xnor_4 g06567(new_n8915, new_n8858, n873);
not_8  g06568(new_n5454, new_n8917);
xnor_4 g06569(n4812, n2731, new_n8918);
not_8  g06570(new_n8918, new_n8919);
nor_5  g06571(new_n2442, n19911, new_n8920_1);
xnor_4 g06572(n24278, n19911, new_n8921);
nor_5  g06573(n24618, new_n2390, new_n8922);
nor_5  g06574(new_n2446, n13708, new_n8923);
nor_5  g06575(new_n3977, n3952, new_n8924);
nor_5  g06576(n18409, new_n3348, new_n8925);
nand_5 g06577(new_n3349_1, n5704, new_n8926);
nor_5  g06578(new_n8926, new_n8925, new_n8927);
nor_5  g06579(new_n8927, new_n8924, new_n8928);
nor_5  g06580(new_n8928, new_n8923, new_n8929);
nor_5  g06581(new_n8929, new_n8922, new_n8930);
and_5  g06582(new_n8930, new_n8921, new_n8931);
nor_5  g06583(new_n8931, new_n8920_1, new_n8932);
xnor_4 g06584(new_n8932, new_n8919, new_n8933);
xnor_4 g06585(new_n8933, new_n8917, new_n8934);
xnor_4 g06586(new_n8930, new_n8921, new_n8935);
not_8  g06587(new_n8935, new_n8936);
nor_5  g06588(new_n8936, new_n5457, new_n8937);
not_8  g06589(new_n8937, new_n8938);
xnor_4 g06590(n24618, n13708, new_n8939);
xnor_4 g06591(new_n8939, new_n8928, new_n8940);
nor_5  g06592(new_n8940, new_n5462, new_n8941);
xnor_4 g06593(new_n8940, new_n5462, new_n8942);
xnor_4 g06594(n12315, n5704, new_n8943_1);
nor_5  g06595(new_n8943_1, new_n5469, new_n8944);
not_8  g06596(new_n8944, new_n8945);
nor_5  g06597(new_n8945, new_n5475, new_n8946);
xnor_4 g06598(new_n8945, new_n5475, new_n8947);
xnor_4 g06599(n18409, n3952, new_n8948);
xnor_4 g06600(new_n8948, new_n8926, new_n8949);
nor_5  g06601(new_n8949, new_n8947, new_n8950);
nor_5  g06602(new_n8950, new_n8946, new_n8951);
nor_5  g06603(new_n8951, new_n8942, new_n8952);
nor_5  g06604(new_n8952, new_n8941, new_n8953);
xnor_4 g06605(new_n8935, new_n5457, new_n8954);
nand_5 g06606(new_n8954, new_n8953, new_n8955);
nand_5 g06607(new_n8955, new_n8938, new_n8956);
xor_4  g06608(new_n8956, new_n8934, n879);
xnor_4 g06609(new_n8490, n18157, new_n8958);
nor_5  g06610(new_n8497, n12161, new_n8959);
nor_5  g06611(new_n8505_1, new_n7661, new_n8960);
nor_5  g06612(new_n8502, new_n7664, new_n8961);
not_8  g06613(new_n8961, new_n8962);
xnor_4 g06614(new_n8505_1, new_n7661, new_n8963);
nor_5  g06615(new_n8963, new_n8962, new_n8964_1);
nor_5  g06616(new_n8964_1, new_n8960, new_n8965);
not_8  g06617(new_n8965, new_n8966);
xnor_4 g06618(new_n8496, new_n6982, new_n8967);
nor_5  g06619(new_n8967, new_n8966, new_n8968);
nor_5  g06620(new_n8968, new_n8959, new_n8969);
xnor_4 g06621(new_n8969, new_n8958, new_n8970);
xnor_4 g06622(new_n8967, new_n8965, new_n8971_1);
xnor_4 g06623(new_n6961, n14684, new_n8972);
nor_5  g06624(new_n6965_1, n6631, new_n8973);
nor_5  g06625(new_n6969, new_n4488, new_n8974);
not_8  g06626(n6631, new_n8975);
xnor_4 g06627(new_n6964, new_n8975, new_n8976);
nor_5  g06628(new_n8976, new_n8974, new_n8977);
nor_5  g06629(new_n8977, new_n8973, new_n8978);
xnor_4 g06630(new_n8978, new_n8972, new_n8979);
not_8  g06631(new_n8979, new_n8980);
nand_5 g06632(new_n8980, new_n8971_1, new_n8981);
xnor_4 g06633(new_n8979, new_n8971_1, new_n8982_1);
xnor_4 g06634(new_n8976, new_n8974, new_n8983);
not_8  g06635(new_n8983, new_n8984);
xnor_4 g06636(new_n8963, new_n8961, new_n8985);
nor_5  g06637(new_n8985, new_n8984, new_n8986);
not_8  g06638(new_n8986, new_n8987);
xnor_4 g06639(new_n6968, new_n4488, new_n8988);
not_8  g06640(new_n8988, new_n8989);
xnor_4 g06641(new_n2569, new_n7664, new_n8990);
nor_5  g06642(new_n8990, new_n8989, new_n8991);
xnor_4 g06643(new_n8985, new_n8983, new_n8992);
nand_5 g06644(new_n8992, new_n8991, new_n8993_1);
nand_5 g06645(new_n8993_1, new_n8987, new_n8994);
nand_5 g06646(new_n8994, new_n8982_1, new_n8995);
nand_5 g06647(new_n8995, new_n8981, new_n8996);
xnor_4 g06648(new_n8996, new_n8970, new_n8997);
xnor_4 g06649(new_n6958, n17035, new_n8998);
nand_5 g06650(new_n6961, new_n4353, new_n8999);
not_8  g06651(new_n8999, new_n9000);
not_8  g06652(new_n8972, new_n9001);
nor_5  g06653(new_n8978, new_n9001, new_n9002);
nor_5  g06654(new_n9002, new_n9000, new_n9003_1);
xnor_4 g06655(new_n9003_1, new_n8998, new_n9004);
xnor_4 g06656(new_n9004, new_n8997, n887);
xnor_4 g06657(new_n6365, n24327, new_n9006);
nand_5 g06658(new_n6370, n22198, new_n9007);
xnor_4 g06659(new_n6369_1, n22198, new_n9008);
nor_5  g06660(new_n6374, new_n5174, new_n9009);
not_8  g06661(new_n9009, new_n9010);
xnor_4 g06662(new_n6374, n20826, new_n9011);
nor_5  g06663(new_n6378, new_n5176, new_n9012_1);
not_8  g06664(new_n9012_1, new_n9013);
xnor_4 g06665(new_n6378, n7305, new_n9014);
nor_5  g06666(new_n6382, new_n5181, new_n9015);
not_8  g06667(new_n9015, new_n9016);
nor_5  g06668(new_n6385_1, n20259, new_n9017);
nor_5  g06669(new_n6387, new_n6158, new_n9018);
xnor_4 g06670(new_n6384, n20259, new_n9019);
not_8  g06671(new_n9019, new_n9020);
nor_5  g06672(new_n9020, new_n9018, new_n9021);
nor_5  g06673(new_n9021, new_n9017, new_n9022);
xnor_4 g06674(new_n6382, n25872, new_n9023);
nand_5 g06675(new_n9023, new_n9022, new_n9024);
nand_5 g06676(new_n9024, new_n9016, new_n9025);
nand_5 g06677(new_n9025, new_n9014, new_n9026);
nand_5 g06678(new_n9026, new_n9013, new_n9027);
nand_5 g06679(new_n9027, new_n9011, new_n9028);
nand_5 g06680(new_n9028, new_n9010, new_n9029);
nand_5 g06681(new_n9029, new_n9008, new_n9030);
nand_5 g06682(new_n9030, new_n9007, new_n9031);
xnor_4 g06683(new_n9031, new_n9006, new_n9032_1);
xnor_4 g06684(new_n3040, n25119, new_n9033);
not_8  g06685(new_n9033, new_n9034);
not_8  g06686(n1163, new_n9035);
nor_5  g06687(new_n3047, new_n9035, new_n9036);
nor_5  g06688(new_n3055, n18537, new_n9037);
xnor_4 g06689(new_n3054, n18537, new_n9038);
not_8  g06690(new_n9038, new_n9039);
nor_5  g06691(new_n3062, n7057, new_n9040);
xnor_4 g06692(new_n3061, n7057, new_n9041);
nor_5  g06693(new_n3067_1, new_n5296, new_n9042_1);
xnor_4 g06694(new_n3067_1, new_n5296, new_n9043);
not_8  g06695(n12495, new_n9044);
nor_5  g06696(new_n3076_1, new_n9044, new_n9045);
nor_5  g06697(new_n9045, n20235, new_n9046_1);
xnor_4 g06698(new_n9045, n20235, new_n9047_1);
nor_5  g06699(new_n9047_1, new_n3073, new_n9048);
nor_5  g06700(new_n9048, new_n9046_1, new_n9049);
not_8  g06701(new_n9049, new_n9050);
nor_5  g06702(new_n9050, new_n9043, new_n9051);
nor_5  g06703(new_n9051, new_n9042_1, new_n9052);
nand_5 g06704(new_n9052, new_n9041, new_n9053);
not_8  g06705(new_n9053, new_n9054);
nor_5  g06706(new_n9054, new_n9040, new_n9055);
nor_5  g06707(new_n9055, new_n9039, new_n9056);
nor_5  g06708(new_n9056, new_n9037, new_n9057);
xnor_4 g06709(new_n3047, n1163, new_n9058);
nand_5 g06710(new_n9058, new_n9057, new_n9059);
not_8  g06711(new_n9059, new_n9060);
nor_5  g06712(new_n9060, new_n9036, new_n9061);
xnor_4 g06713(new_n9061, new_n9034, new_n9062);
xnor_4 g06714(new_n9062, new_n9032_1, new_n9063);
xnor_4 g06715(new_n9029, new_n9008, new_n9064);
not_8  g06716(new_n9064, new_n9065);
xnor_4 g06717(new_n9058, new_n9057, new_n9066);
nand_5 g06718(new_n9066, new_n9065, new_n9067);
xnor_4 g06719(new_n9066, new_n9064, new_n9068);
xnor_4 g06720(new_n9055, new_n9038, new_n9069);
not_8  g06721(new_n9069, new_n9070);
xnor_4 g06722(new_n9027, new_n9011, new_n9071);
nor_5  g06723(new_n9071, new_n9070, new_n9072);
xnor_4 g06724(new_n9071, new_n9069, new_n9073);
not_8  g06725(new_n9073, new_n9074);
xnor_4 g06726(new_n9052, new_n9041, new_n9075);
xnor_4 g06727(new_n9025, new_n9014, new_n9076);
nor_5  g06728(new_n9076, new_n9075, new_n9077);
not_8  g06729(new_n9076, new_n9078);
xnor_4 g06730(new_n9078, new_n9075, new_n9079);
not_8  g06731(new_n9079, new_n9080);
xnor_4 g06732(new_n9049, new_n9043, new_n9081);
xnor_4 g06733(new_n9023, new_n9022, new_n9082);
nor_5  g06734(new_n9082, new_n9081, new_n9083);
not_8  g06735(new_n9082, new_n9084);
xnor_4 g06736(new_n9084, new_n9081, new_n9085);
not_8  g06737(new_n9085, new_n9086);
xnor_4 g06738(new_n9019, new_n9018, new_n9087);
not_8  g06739(new_n9087, new_n9088);
xnor_4 g06740(new_n9047_1, new_n3082, new_n9089);
and_5  g06741(new_n9089, new_n9088, new_n9090_1);
xnor_4 g06742(new_n6108, new_n6158, new_n9091);
not_8  g06743(new_n9091, new_n9092);
xnor_4 g06744(new_n3076_1, n12495, new_n9093);
nor_5  g06745(new_n9093, new_n9092, new_n9094);
not_8  g06746(new_n9094, new_n9095);
xnor_4 g06747(new_n9089, new_n9087, new_n9096);
not_8  g06748(new_n9096, new_n9097);
nor_5  g06749(new_n9097, new_n9095, new_n9098);
nor_5  g06750(new_n9098, new_n9090_1, new_n9099);
nor_5  g06751(new_n9099, new_n9086, new_n9100);
nor_5  g06752(new_n9100, new_n9083, new_n9101);
nor_5  g06753(new_n9101, new_n9080, new_n9102);
nor_5  g06754(new_n9102, new_n9077, new_n9103);
nor_5  g06755(new_n9103, new_n9074, new_n9104_1);
nor_5  g06756(new_n9104_1, new_n9072, new_n9105);
not_8  g06757(new_n9105, new_n9106);
nand_5 g06758(new_n9106, new_n9068, new_n9107);
nand_5 g06759(new_n9107, new_n9067, new_n9108);
xnor_4 g06760(new_n9108, new_n9063, n904);
not_8  g06761(new_n7055, new_n9110);
not_8  g06762(n19472, new_n9111);
nor_5  g06763(n18962, n10158, new_n9112);
nand_5 g06764(new_n9112, new_n7136, new_n9113);
nor_5  g06765(new_n9113, n15539, new_n9114);
xnor_4 g06766(new_n9114, n19228, new_n9115);
xnor_4 g06767(new_n9115, new_n5487, new_n9116);
xnor_4 g06768(new_n9113, new_n7132, new_n9117);
not_8  g06769(new_n9117, new_n9118);
nor_5  g06770(new_n9118, new_n5512, new_n9119);
xnor_4 g06771(new_n9117, new_n5512, new_n9120);
not_8  g06772(new_n9120, new_n9121);
xnor_4 g06773(new_n9112, new_n7136, new_n9122);
nor_5  g06774(new_n9122, new_n3409, new_n9123);
xnor_4 g06775(new_n9122, n14603, new_n9124);
not_8  g06776(new_n9124, new_n9125);
xnor_4 g06777(n18962, n10158, new_n9126);
nand_5 g06778(new_n9126, new_n3415, new_n9127);
nand_5 g06779(n23333, n18962, new_n9128);
xnor_4 g06780(new_n9126, n20794, new_n9129_1);
nand_5 g06781(new_n9129_1, new_n9128, new_n9130);
nand_5 g06782(new_n9130, new_n9127, new_n9131);
nor_5  g06783(new_n9131, new_n9125, new_n9132);
nor_5  g06784(new_n9132, new_n9123, new_n9133);
nor_5  g06785(new_n9133, new_n9121, new_n9134);
nor_5  g06786(new_n9134, new_n9119, new_n9135);
xnor_4 g06787(new_n9135, new_n9116, new_n9136);
xnor_4 g06788(new_n9136, new_n9111, new_n9137);
not_8  g06789(new_n9137, new_n9138);
xnor_4 g06790(new_n9133, new_n9120, new_n9139);
nor_5  g06791(new_n9139, n25370, new_n9140);
not_8  g06792(new_n9140, new_n9141);
xnor_4 g06793(new_n9131, new_n9124, new_n9142);
nand_5 g06794(new_n9142, n24786, new_n9143);
not_8  g06795(new_n9143, new_n9144);
not_8  g06796(n24786, new_n9145);
xnor_4 g06797(new_n9142, new_n9145, new_n9146_1);
not_8  g06798(new_n9146_1, new_n9147);
not_8  g06799(n23065, new_n9148);
not_8  g06800(n18962, new_n9149);
xnor_4 g06801(n23333, new_n9149, new_n9150);
not_8  g06802(new_n9150, new_n9151);
nor_5  g06803(new_n9151, new_n9148, new_n9152);
nand_5 g06804(new_n9152, new_n9129_1, new_n9153);
not_8  g06805(new_n9153, new_n9154);
not_8  g06806(n27120, new_n9155);
not_8  g06807(new_n9152, new_n9156);
not_8  g06808(new_n9128, new_n9157);
xnor_4 g06809(new_n9129_1, new_n9157, new_n9158);
nand_5 g06810(new_n9158, new_n9156, new_n9159);
nand_5 g06811(new_n9159, new_n9153, new_n9160);
nor_5  g06812(new_n9160, new_n9155, new_n9161);
nor_5  g06813(new_n9161, new_n9154, new_n9162);
nor_5  g06814(new_n9162, new_n9147, new_n9163);
nor_5  g06815(new_n9163, new_n9144, new_n9164_1);
not_8  g06816(n25370, new_n9165);
xnor_4 g06817(new_n9139, new_n9165, new_n9166_1);
nand_5 g06818(new_n9166_1, new_n9164_1, new_n9167);
nand_5 g06819(new_n9167, new_n9141, new_n9168);
xnor_4 g06820(new_n9168, new_n9138, new_n9169);
xnor_4 g06821(new_n9169, new_n9110, new_n9170);
xnor_4 g06822(new_n9166_1, new_n9164_1, new_n9171);
not_8  g06823(new_n9171, new_n9172_1);
nand_5 g06824(new_n9172_1, new_n7059, new_n9173);
xnor_4 g06825(new_n9171, new_n7059, new_n9174);
not_8  g06826(new_n7079_1, new_n9175);
xnor_4 g06827(new_n9160, n27120, new_n9176);
not_8  g06828(new_n9176, new_n9177);
nand_5 g06829(new_n9177, new_n7099_1, new_n9178);
xnor_4 g06830(new_n9150, new_n9148, new_n9179);
not_8  g06831(new_n9179, new_n9180);
nor_5  g06832(new_n9180, new_n7069, new_n9181);
not_8  g06833(new_n9181, new_n9182_1);
xnor_4 g06834(new_n9176, new_n7099_1, new_n9183);
nand_5 g06835(new_n9183, new_n9182_1, new_n9184);
nand_5 g06836(new_n9184, new_n9178, new_n9185);
nand_5 g06837(new_n9185, new_n9175, new_n9186);
xnor_4 g06838(new_n9162, new_n9146_1, new_n9187);
not_8  g06839(new_n9187, new_n9188);
xnor_4 g06840(new_n9185, new_n7079_1, new_n9189);
nand_5 g06841(new_n9189, new_n9188, new_n9190);
nand_5 g06842(new_n9190, new_n9186, new_n9191_1);
nand_5 g06843(new_n9191_1, new_n9174, new_n9192);
nand_5 g06844(new_n9192, new_n9173, new_n9193);
xnor_4 g06845(new_n9193, new_n9170, n948);
xnor_4 g06846(n25972, n10250, new_n9195);
not_8  g06847(n21915, new_n9196);
or_5   g06848(new_n9196, n7674, new_n9197);
xnor_4 g06849(n21915, n7674, new_n9198);
or_5   g06850(new_n7219, n6397, new_n9199);
xnor_4 g06851(n13775, n6397, new_n9200);
or_5   g06852(n19196, new_n7223, new_n9201);
xnor_4 g06853(n19196, n1293, new_n9202);
or_5   g06854(n23586, new_n7227, new_n9203);
xnor_4 g06855(n23586, n19042, new_n9204);
nor_5  g06856(n21226, new_n9111, new_n9205);
xnor_4 g06857(n21226, n19472, new_n9206);
nor_5  g06858(new_n9165, n4426, new_n9207);
not_8  g06859(new_n9207, new_n9208);
xnor_4 g06860(n25370, n4426, new_n9209);
not_8  g06861(n20036, new_n9210);
nor_5  g06862(n24786, new_n9210, new_n9211);
nor_5  g06863(new_n9145, n20036, new_n9212);
nor_5  g06864(n27120, new_n4305, new_n9213);
nor_5  g06865(new_n9155, n11192, new_n9214);
nor_5  g06866(n23065, new_n4307, new_n9215);
not_8  g06867(new_n9215, new_n9216);
nor_5  g06868(new_n9216, new_n9214, new_n9217_1);
nor_5  g06869(new_n9217_1, new_n9213, new_n9218);
nor_5  g06870(new_n9218, new_n9212, new_n9219);
nor_5  g06871(new_n9219, new_n9211, new_n9220_1);
nand_5 g06872(new_n9220_1, new_n9209, new_n9221);
nand_5 g06873(new_n9221, new_n9208, new_n9222);
and_5  g06874(new_n9222, new_n9206, new_n9223);
nor_5  g06875(new_n9223, new_n9205, new_n9224);
not_8  g06876(new_n9224, new_n9225);
nand_5 g06877(new_n9225, new_n9204, new_n9226);
nand_5 g06878(new_n9226, new_n9203, new_n9227);
nand_5 g06879(new_n9227, new_n9202, new_n9228);
nand_5 g06880(new_n9228, new_n9201, new_n9229);
nand_5 g06881(new_n9229, new_n9200, new_n9230);
nand_5 g06882(new_n9230, new_n9199, new_n9231);
nand_5 g06883(new_n9231, new_n9198, new_n9232);
nand_5 g06884(new_n9232, new_n9197, new_n9233);
xnor_4 g06885(new_n9233, new_n9195, new_n9234);
xnor_4 g06886(n20040, n2978, new_n9235);
or_5   g06887(new_n7114, n19531, new_n9236);
xnor_4 g06888(n23697, n19531, new_n9237);
or_5   g06889(n18345, new_n7118, new_n9238);
xnor_4 g06890(n18345, n2289, new_n9239);
or_5   g06891(n13190, new_n7122, new_n9240);
xnor_4 g06892(n13190, n1112, new_n9241);
or_5   g06893(new_n7895, n3460, new_n9242);
xnor_4 g06894(n20179, n3460, new_n9243);
nor_5  g06895(new_n7898, n5226, new_n9244);
not_8  g06896(new_n9244, new_n9245);
xnor_4 g06897(n19228, n5226, new_n9246_1);
nor_5  g06898(n17664, new_n7132, new_n9247);
not_8  g06899(new_n9247, new_n9248);
xnor_4 g06900(n17664, n15539, new_n9249);
nor_5  g06901(new_n2610, n8052, new_n9250);
nor_5  g06902(n23369, new_n7136, new_n9251_1);
not_8  g06903(n1136, new_n9252);
nor_5  g06904(n10158, new_n9252, new_n9253);
nor_5  g06905(new_n7907, n1136, new_n9254);
nor_5  g06906(new_n7636, n18962, new_n9255);
not_8  g06907(new_n9255, new_n9256);
nor_5  g06908(new_n9256, new_n9254, new_n9257);
nor_5  g06909(new_n9257, new_n9253, new_n9258);
nor_5  g06910(new_n9258, new_n9251_1, new_n9259_1);
nor_5  g06911(new_n9259_1, new_n9250, new_n9260);
nand_5 g06912(new_n9260, new_n9249, new_n9261_1);
nand_5 g06913(new_n9261_1, new_n9248, new_n9262);
nand_5 g06914(new_n9262, new_n9246_1, new_n9263);
nand_5 g06915(new_n9263, new_n9245, new_n9264);
nand_5 g06916(new_n9264, new_n9243, new_n9265);
nand_5 g06917(new_n9265, new_n9242, new_n9266);
nand_5 g06918(new_n9266, new_n9241, new_n9267);
nand_5 g06919(new_n9267, new_n9240, new_n9268);
nand_5 g06920(new_n9268, new_n9239, new_n9269);
nand_5 g06921(new_n9269, new_n9238, new_n9270);
nand_5 g06922(new_n9270, new_n9237, new_n9271);
nand_5 g06923(new_n9271, new_n9236, new_n9272);
xnor_4 g06924(new_n9272, new_n9235, new_n9273);
not_8  g06925(n12507, new_n9274);
nor_5  g06926(n15258, n4588, new_n9275);
nand_5 g06927(new_n9275, new_n8495, new_n9276);
nor_5  g06928(new_n9276, n22631, new_n9277);
nand_5 g06929(new_n9277, new_n8488, new_n9278);
nor_5  g06930(new_n9278, n25068, new_n9279);
nand_5 g06931(new_n9279, new_n8475, new_n9280);
nor_5  g06932(new_n9280, n7841, new_n9281);
nand_5 g06933(new_n9281, new_n8466, new_n9282);
xnor_4 g06934(new_n9282, new_n8416, new_n9283);
xnor_4 g06935(new_n9283, new_n9274, new_n9284);
xnor_4 g06936(new_n9281, n26264, new_n9285);
and_5  g06937(new_n9285, n15077, new_n9286);
nor_5  g06938(new_n9285, n15077, new_n9287_1);
xnor_4 g06939(new_n9280, new_n8470, new_n9288);
and_5  g06940(new_n9288, n3710, new_n9289);
nor_5  g06941(new_n9288, n3710, new_n9290);
not_8  g06942(n26318, new_n9291);
xnor_4 g06943(new_n9279, n16812, new_n9292);
not_8  g06944(new_n9292, new_n9293);
nand_5 g06945(new_n9293, new_n9291, new_n9294);
xnor_4 g06946(new_n9292, new_n9291, new_n9295);
not_8  g06947(n26054, new_n9296);
xnor_4 g06948(new_n9278, new_n8480_1, new_n9297);
not_8  g06949(new_n9297, new_n9298);
nand_5 g06950(new_n9298, new_n9296, new_n9299);
xnor_4 g06951(new_n9297, new_n9296, new_n9300);
not_8  g06952(n19081, new_n9301);
xnor_4 g06953(new_n9277, n2331, new_n9302);
not_8  g06954(new_n9302, new_n9303);
nand_5 g06955(new_n9303, new_n9301, new_n9304);
xnor_4 g06956(new_n9302, new_n9301, new_n9305);
not_8  g06957(n8309, new_n9306);
xnor_4 g06958(new_n9276, new_n8493, new_n9307);
not_8  g06959(new_n9307, new_n9308_1);
nand_5 g06960(new_n9308_1, new_n9306, new_n9309);
not_8  g06961(n19144, new_n9310);
xnor_4 g06962(new_n9275, n16743, new_n9311);
not_8  g06963(new_n9311, new_n9312);
nand_5 g06964(new_n9312, new_n9310, new_n9313);
xnor_4 g06965(new_n9311, new_n9310, new_n9314);
not_8  g06966(n12593, new_n9315);
xnor_4 g06967(n15258, n4588, new_n9316);
nand_5 g06968(new_n9316, new_n9315, new_n9317);
nand_5 g06969(n13714, n4588, new_n9318_1);
xnor_4 g06970(new_n9316, n12593, new_n9319);
nand_5 g06971(new_n9319, new_n9318_1, new_n9320);
nand_5 g06972(new_n9320, new_n9317, new_n9321);
nand_5 g06973(new_n9321, new_n9314, new_n9322);
nand_5 g06974(new_n9322, new_n9313, new_n9323_1);
xnor_4 g06975(new_n9307, new_n9306, new_n9324);
nand_5 g06976(new_n9324, new_n9323_1, new_n9325);
nand_5 g06977(new_n9325, new_n9309, new_n9326);
nand_5 g06978(new_n9326, new_n9305, new_n9327);
nand_5 g06979(new_n9327, new_n9304, new_n9328);
nand_5 g06980(new_n9328, new_n9300, new_n9329);
nand_5 g06981(new_n9329, new_n9299, new_n9330);
nand_5 g06982(new_n9330, new_n9295, new_n9331);
nand_5 g06983(new_n9331, new_n9294, new_n9332);
nor_5  g06984(new_n9332, new_n9290, new_n9333);
nor_5  g06985(new_n9333, new_n9289, new_n9334);
nor_5  g06986(new_n9334, new_n9287_1, new_n9335);
nor_5  g06987(new_n9335, new_n9286, new_n9336);
xnor_4 g06988(new_n9336, new_n9284, new_n9337);
xnor_4 g06989(new_n9337, new_n9273, new_n9338);
not_8  g06990(new_n9338, new_n9339);
xnor_4 g06991(new_n9270, new_n9237, new_n9340);
not_8  g06992(n15077, new_n9341);
xnor_4 g06993(new_n9285, new_n9341, new_n9342);
xnor_4 g06994(new_n9342, new_n9334, new_n9343);
not_8  g06995(new_n9343, new_n9344_1);
nor_5  g06996(new_n9344_1, new_n9340, new_n9345);
xnor_4 g06997(new_n9343, new_n9340, new_n9346);
not_8  g06998(new_n9346, new_n9347);
xnor_4 g06999(new_n9268, new_n9239, new_n9348);
not_8  g07000(n3710, new_n9349);
xnor_4 g07001(new_n9288, new_n9349, new_n9350);
xnor_4 g07002(new_n9350, new_n9332, new_n9351);
not_8  g07003(new_n9351, new_n9352);
nand_5 g07004(new_n9352, new_n9348, new_n9353);
xnor_4 g07005(new_n9351, new_n9348, new_n9354);
xnor_4 g07006(new_n9266, new_n9241, new_n9355);
xnor_4 g07007(new_n9330, new_n9295, new_n9356);
not_8  g07008(new_n9356, new_n9357);
nand_5 g07009(new_n9357, new_n9355, new_n9358);
xnor_4 g07010(new_n9356, new_n9355, new_n9359);
xnor_4 g07011(new_n9264, new_n9243, new_n9360);
not_8  g07012(new_n9300, new_n9361);
xnor_4 g07013(new_n9328, new_n9361, new_n9362);
nand_5 g07014(new_n9362, new_n9360, new_n9363);
not_8  g07015(new_n9360, new_n9364_1);
xnor_4 g07016(new_n9362, new_n9364_1, new_n9365);
xnor_4 g07017(new_n9262, new_n9246_1, new_n9366);
xnor_4 g07018(new_n9326, new_n9305, new_n9367);
not_8  g07019(new_n9367, new_n9368);
nand_5 g07020(new_n9368, new_n9366, new_n9369);
xnor_4 g07021(new_n9367, new_n9366, new_n9370);
xnor_4 g07022(new_n9260, new_n9249, new_n9371_1);
not_8  g07023(new_n9371_1, new_n9372_1);
xnor_4 g07024(new_n9324, new_n9323_1, new_n9373);
nor_5  g07025(new_n9373, new_n9372_1, new_n9374);
not_8  g07026(new_n9374, new_n9375);
xnor_4 g07027(new_n9373, new_n9371_1, new_n9376);
xnor_4 g07028(new_n9321, new_n9314, new_n9377);
xnor_4 g07029(n23369, n8052, new_n9378);
xnor_4 g07030(new_n9378, new_n9258, new_n9379);
not_8  g07031(new_n9379, new_n9380_1);
nand_5 g07032(new_n9380_1, new_n9377, new_n9381);
xnor_4 g07033(new_n9379, new_n9377, new_n9382_1);
xnor_4 g07034(new_n9319, new_n9318_1, new_n9383);
xnor_4 g07035(n10158, n1136, new_n9384);
xnor_4 g07036(new_n9384, new_n9256, new_n9385);
not_8  g07037(new_n9385, new_n9386);
nand_5 g07038(new_n9386, new_n9383, new_n9387);
xnor_4 g07039(n19234, n18962, new_n9388);
not_8  g07040(n4588, new_n9389);
xnor_4 g07041(n13714, new_n9389, new_n9390);
not_8  g07042(new_n9390, new_n9391);
nor_5  g07043(new_n9391, new_n9388, new_n9392);
xnor_4 g07044(new_n9385, new_n9383, new_n9393);
nand_5 g07045(new_n9393, new_n9392, new_n9394);
nand_5 g07046(new_n9394, new_n9387, new_n9395);
nand_5 g07047(new_n9395, new_n9382_1, new_n9396_1);
nand_5 g07048(new_n9396_1, new_n9381, new_n9397);
not_8  g07049(new_n9397, new_n9398);
nand_5 g07050(new_n9398, new_n9376, new_n9399_1);
nand_5 g07051(new_n9399_1, new_n9375, new_n9400);
nand_5 g07052(new_n9400, new_n9370, new_n9401);
nand_5 g07053(new_n9401, new_n9369, new_n9402);
nand_5 g07054(new_n9402, new_n9365, new_n9403_1);
nand_5 g07055(new_n9403_1, new_n9363, new_n9404);
nand_5 g07056(new_n9404, new_n9359, new_n9405);
nand_5 g07057(new_n9405, new_n9358, new_n9406);
nand_5 g07058(new_n9406, new_n9354, new_n9407);
nand_5 g07059(new_n9407, new_n9353, new_n9408);
nor_5  g07060(new_n9408, new_n9347, new_n9409);
nor_5  g07061(new_n9409, new_n9345, new_n9410);
xnor_4 g07062(new_n9410, new_n9339, new_n9411);
xnor_4 g07063(new_n9411, new_n9234, new_n9412);
xnor_4 g07064(new_n9231, new_n9198, new_n9413);
xnor_4 g07065(new_n9408, new_n9346, new_n9414);
not_8  g07066(new_n9414, new_n9415);
nand_5 g07067(new_n9415, new_n9413, new_n9416);
xnor_4 g07068(new_n9414, new_n9413, new_n9417);
xnor_4 g07069(new_n9229, new_n9200, new_n9418);
xnor_4 g07070(new_n9406, new_n9354, new_n9419_1);
not_8  g07071(new_n9419_1, new_n9420);
nand_5 g07072(new_n9420, new_n9418, new_n9421);
xnor_4 g07073(new_n9419_1, new_n9418, new_n9422);
xnor_4 g07074(new_n9227, new_n9202, new_n9423_1);
xnor_4 g07075(new_n9404, new_n9359, new_n9424);
not_8  g07076(new_n9424, new_n9425);
nand_5 g07077(new_n9425, new_n9423_1, new_n9426);
xnor_4 g07078(new_n9424, new_n9423_1, new_n9427);
xnor_4 g07079(new_n9224, new_n9204, new_n9428);
not_8  g07080(new_n9428, new_n9429);
not_8  g07081(new_n9365, new_n9430_1);
xnor_4 g07082(new_n9402, new_n9430_1, new_n9431);
nand_5 g07083(new_n9431, new_n9429, new_n9432);
xnor_4 g07084(new_n9431, new_n9428, new_n9433);
not_8  g07085(new_n9206, new_n9434);
xnor_4 g07086(new_n9222, new_n9434, new_n9435_1);
not_8  g07087(new_n9435_1, new_n9436);
not_8  g07088(new_n9370, new_n9437);
xnor_4 g07089(new_n9400, new_n9437, new_n9438);
nand_5 g07090(new_n9438, new_n9436, new_n9439);
xnor_4 g07091(new_n9438, new_n9435_1, new_n9440);
xnor_4 g07092(new_n9397, new_n9376, new_n9441);
xnor_4 g07093(new_n9220_1, new_n9209, new_n9442);
nand_5 g07094(new_n9442, new_n9441, new_n9443);
not_8  g07095(new_n9442, new_n9444);
xnor_4 g07096(new_n9444, new_n9441, new_n9445_1);
xnor_4 g07097(new_n9395, new_n9382_1, new_n9446);
xnor_4 g07098(n24786, n20036, new_n9447);
xnor_4 g07099(new_n9447, new_n9218, new_n9448);
nand_5 g07100(new_n9448, new_n9446, new_n9449);
not_8  g07101(new_n9446, new_n9450);
xnor_4 g07102(new_n9448, new_n9450, new_n9451_1);
xnor_4 g07103(n23065, n9380, new_n9452);
xnor_4 g07104(new_n9390, new_n9388, new_n9453);
not_8  g07105(new_n9453, new_n9454);
nor_5  g07106(new_n9454, new_n9452, new_n9455);
xnor_4 g07107(n27120, n11192, new_n9456);
xnor_4 g07108(new_n9456, new_n9216, new_n9457);
not_8  g07109(new_n9457, new_n9458_1);
nor_5  g07110(new_n9458_1, new_n9455, new_n9459_1);
not_8  g07111(new_n9459_1, new_n9460_1);
xnor_4 g07112(new_n9393, new_n9392, new_n9461);
xnor_4 g07113(new_n9457, new_n9455, new_n9462);
nand_5 g07114(new_n9462, new_n9461, new_n9463);
nand_5 g07115(new_n9463, new_n9460_1, new_n9464);
nand_5 g07116(new_n9464, new_n9451_1, new_n9465);
nand_5 g07117(new_n9465, new_n9449, new_n9466);
nand_5 g07118(new_n9466, new_n9445_1, new_n9467);
nand_5 g07119(new_n9467, new_n9443, new_n9468);
nand_5 g07120(new_n9468, new_n9440, new_n9469);
nand_5 g07121(new_n9469, new_n9439, new_n9470);
nand_5 g07122(new_n9470, new_n9433, new_n9471);
nand_5 g07123(new_n9471, new_n9432, new_n9472);
nand_5 g07124(new_n9472, new_n9427, new_n9473);
nand_5 g07125(new_n9473, new_n9426, new_n9474);
nand_5 g07126(new_n9474, new_n9422, new_n9475);
nand_5 g07127(new_n9475, new_n9421, new_n9476);
nand_5 g07128(new_n9476, new_n9417, new_n9477);
nand_5 g07129(new_n9477, new_n9416, new_n9478);
not_8  g07130(new_n9478, new_n9479);
xnor_4 g07131(new_n9479, new_n9412, n957);
xnor_4 g07132(new_n9388, n20385, new_n9481);
not_8  g07133(n21138, new_n9482);
xnor_4 g07134(n26167, n24129, new_n9483);
xnor_4 g07135(new_n9483, new_n9482, new_n9484);
xnor_4 g07136(new_n9484, new_n9481, n980);
nor_5  g07137(new_n8190, new_n4549, new_n9486);
xnor_4 g07138(new_n8190, new_n4549, new_n9487);
nand_5 g07139(new_n8197, new_n4553, new_n9488);
xnor_4 g07140(new_n8196, new_n4553, new_n9489);
nand_5 g07141(new_n8201, new_n4557, new_n9490);
xnor_4 g07142(new_n8201, new_n4557, new_n9491);
not_8  g07143(new_n9491, new_n9492);
nand_5 g07144(new_n8206, new_n4561, new_n9493_1);
xnor_4 g07145(new_n8206, new_n4561, new_n9494);
not_8  g07146(new_n9494, new_n9495);
nand_5 g07147(new_n8212, new_n4565, new_n9496);
xnor_4 g07148(new_n8211, new_n4565, new_n9497);
nand_5 g07149(new_n8218, new_n4570, new_n9498);
xnor_4 g07150(new_n8218, new_n4569, new_n9499);
nand_5 g07151(new_n8223, new_n4574, new_n9500);
not_8  g07152(new_n8223, new_n9501);
xnor_4 g07153(new_n9501, new_n4574, new_n9502);
nand_5 g07154(new_n8229, new_n4579, new_n9503);
xnor_4 g07155(new_n8229, new_n4581, new_n9504);
nor_5  g07156(new_n8237, new_n4584, new_n9505);
nor_5  g07157(new_n8242, new_n4587, new_n9506);
not_8  g07158(new_n9506, new_n9507_1);
xnor_4 g07159(new_n8237, new_n4585, new_n9508_1);
not_8  g07160(new_n9508_1, new_n9509);
nor_5  g07161(new_n9509, new_n9507_1, new_n9510);
nor_5  g07162(new_n9510, new_n9505, new_n9511);
nand_5 g07163(new_n9511, new_n9504, new_n9512_1);
nand_5 g07164(new_n9512_1, new_n9503, new_n9513);
nand_5 g07165(new_n9513, new_n9502, new_n9514);
nand_5 g07166(new_n9514, new_n9500, new_n9515);
nand_5 g07167(new_n9515, new_n9499, new_n9516);
nand_5 g07168(new_n9516, new_n9498, new_n9517);
nand_5 g07169(new_n9517, new_n9497, new_n9518);
nand_5 g07170(new_n9518, new_n9496, new_n9519);
nand_5 g07171(new_n9519, new_n9495, new_n9520);
nand_5 g07172(new_n9520, new_n9493_1, new_n9521);
nand_5 g07173(new_n9521, new_n9492, new_n9522);
nand_5 g07174(new_n9522, new_n9490, new_n9523);
nand_5 g07175(new_n9523, new_n9489, new_n9524);
nand_5 g07176(new_n9524, new_n9488, new_n9525);
nor_5  g07177(new_n9525, new_n9487, new_n9526);
nor_5  g07178(new_n9526, new_n9486, new_n9527);
xnor_4 g07179(new_n8187, new_n4547, new_n9528);
xnor_4 g07180(new_n9528, new_n9527, new_n9529);
not_8  g07181(n16544, new_n9530);
or_5   g07182(new_n9530, n12650, new_n9531);
xnor_4 g07183(n16544, n12650, new_n9532);
or_5   g07184(n10201, new_n2941, new_n9533);
xnor_4 g07185(n10201, n6814, new_n9534);
not_8  g07186(n19701, new_n9535);
or_5   g07187(new_n9535, n10593, new_n9536);
xnor_4 g07188(n19701, n10593, new_n9537);
not_8  g07189(n23529, new_n9538);
or_5   g07190(new_n9538, n18290, new_n9539);
xnor_4 g07191(n23529, n18290, new_n9540);
not_8  g07192(n24620, new_n9541);
or_5   g07193(new_n9541, n11580, new_n9542);
xnor_4 g07194(n24620, n11580, new_n9543);
nor_5  g07195(n15884, new_n2955, new_n9544);
xnor_4 g07196(n15884, n5211, new_n9545);
not_8  g07197(n12956, new_n9546);
nor_5  g07198(new_n9546, n6356, new_n9547);
not_8  g07199(new_n9547, new_n9548);
xnor_4 g07200(n12956, n6356, new_n9549);
nor_5  g07201(new_n5877, n18295, new_n9550);
nor_5  g07202(n27104, new_n2963, new_n9551);
nor_5  g07203(new_n5882_1, n6502, new_n9552_1);
not_8  g07204(n6502, new_n9553);
nor_5  g07205(n27188, new_n9553, new_n9554_1);
not_8  g07206(n6611, new_n9555);
nor_5  g07207(n15780, new_n9555, new_n9556_1);
not_8  g07208(new_n9556_1, new_n9557_1);
nor_5  g07209(new_n9557_1, new_n9554_1, new_n9558_1);
nor_5  g07210(new_n9558_1, new_n9552_1, new_n9559);
nor_5  g07211(new_n9559, new_n9551, new_n9560);
nor_5  g07212(new_n9560, new_n9550, new_n9561);
nand_5 g07213(new_n9561, new_n9549, new_n9562);
nand_5 g07214(new_n9562, new_n9548, new_n9563);
and_5  g07215(new_n9563, new_n9545, new_n9564);
nor_5  g07216(new_n9564, new_n9544, new_n9565);
not_8  g07217(new_n9565, new_n9566);
nand_5 g07218(new_n9566, new_n9543, new_n9567);
nand_5 g07219(new_n9567, new_n9542, new_n9568);
nand_5 g07220(new_n9568, new_n9540, new_n9569);
nand_5 g07221(new_n9569, new_n9539, new_n9570);
nand_5 g07222(new_n9570, new_n9537, new_n9571);
nand_5 g07223(new_n9571, new_n9536, new_n9572);
nand_5 g07224(new_n9572, new_n9534, new_n9573);
nand_5 g07225(new_n9573, new_n9533, new_n9574);
nand_5 g07226(new_n9574, new_n9532, new_n9575);
nand_5 g07227(new_n9575, new_n9531, new_n9576);
not_8  g07228(new_n9576, new_n9577);
xnor_4 g07229(new_n9577, new_n9529, new_n9578);
xnor_4 g07230(new_n9574, new_n9532, new_n9579);
not_8  g07231(new_n9487, new_n9580);
xnor_4 g07232(new_n9525, new_n9580, new_n9581);
not_8  g07233(new_n9581, new_n9582);
nand_5 g07234(new_n9582, new_n9579, new_n9583);
xnor_4 g07235(new_n9581, new_n9579, new_n9584);
xnor_4 g07236(new_n9572, new_n9534, new_n9585);
xnor_4 g07237(new_n9523, new_n9489, new_n9586);
not_8  g07238(new_n9586, new_n9587);
nand_5 g07239(new_n9587, new_n9585, new_n9588);
xnor_4 g07240(new_n9586, new_n9585, new_n9589);
xnor_4 g07241(new_n9570, new_n9537, new_n9590);
xnor_4 g07242(new_n9521, new_n9491, new_n9591);
nand_5 g07243(new_n9591, new_n9590, new_n9592);
not_8  g07244(new_n9591, new_n9593);
xnor_4 g07245(new_n9593, new_n9590, new_n9594);
xnor_4 g07246(new_n9568, new_n9540, new_n9595);
xnor_4 g07247(new_n9519, new_n9494, new_n9596);
nand_5 g07248(new_n9596, new_n9595, new_n9597);
not_8  g07249(new_n9596, new_n9598_1);
xnor_4 g07250(new_n9598_1, new_n9595, new_n9599);
xnor_4 g07251(new_n9565, new_n9543, new_n9600);
not_8  g07252(new_n9600, new_n9601);
xnor_4 g07253(new_n9517, new_n9497, new_n9602);
not_8  g07254(new_n9602, new_n9603);
nand_5 g07255(new_n9603, new_n9601, new_n9604);
xnor_4 g07256(new_n9603, new_n9600, new_n9605);
nor_5  g07257(new_n9563, new_n9545, new_n9606);
nor_5  g07258(new_n9606, new_n9564, new_n9607);
not_8  g07259(new_n9607, new_n9608);
xnor_4 g07260(new_n9515, new_n9499, new_n9609);
not_8  g07261(new_n9609, new_n9610);
nand_5 g07262(new_n9610, new_n9608, new_n9611);
xnor_4 g07263(new_n9610, new_n9607, new_n9612);
xnor_4 g07264(new_n9513, new_n9502, new_n9613);
not_8  g07265(new_n9613, new_n9614);
xnor_4 g07266(new_n9561, new_n9549, new_n9615);
nand_5 g07267(new_n9615, new_n9614, new_n9616_1);
xnor_4 g07268(new_n9511, new_n9504, new_n9617);
xnor_4 g07269(n27104, n18295, new_n9618);
xnor_4 g07270(new_n9618, new_n9559, new_n9619);
not_8  g07271(new_n9619, new_n9620);
nor_5  g07272(new_n9620, new_n9617, new_n9621);
xnor_4 g07273(new_n9619, new_n9617, new_n9622_1);
not_8  g07274(new_n9622_1, new_n9623);
xnor_4 g07275(n15780, n6611, new_n9624);
xnor_4 g07276(new_n8385, new_n4587, new_n9625);
not_8  g07277(new_n9625, new_n9626_1);
nor_5  g07278(new_n9626_1, new_n9624, new_n9627);
xnor_4 g07279(n27188, n6502, new_n9628);
xnor_4 g07280(new_n9628, new_n9557_1, new_n9629);
not_8  g07281(new_n9629, new_n9630);
nor_5  g07282(new_n9630, new_n9627, new_n9631);
xnor_4 g07283(new_n9508_1, new_n9507_1, new_n9632);
xnor_4 g07284(new_n9629, new_n9627, new_n9633_1);
not_8  g07285(new_n9633_1, new_n9634);
nor_5  g07286(new_n9634, new_n9632, new_n9635_1);
nor_5  g07287(new_n9635_1, new_n9631, new_n9636);
nor_5  g07288(new_n9636, new_n9623, new_n9637);
nor_5  g07289(new_n9637, new_n9621, new_n9638);
not_8  g07290(new_n9638, new_n9639);
xnor_4 g07291(new_n9615, new_n9613, new_n9640);
nand_5 g07292(new_n9640, new_n9639, new_n9641);
nand_5 g07293(new_n9641, new_n9616_1, new_n9642);
nand_5 g07294(new_n9642, new_n9612, new_n9643);
nand_5 g07295(new_n9643, new_n9611, new_n9644);
nand_5 g07296(new_n9644, new_n9605, new_n9645);
nand_5 g07297(new_n9645, new_n9604, new_n9646_1);
nand_5 g07298(new_n9646_1, new_n9599, new_n9647);
nand_5 g07299(new_n9647, new_n9597, new_n9648_1);
nand_5 g07300(new_n9648_1, new_n9594, new_n9649);
nand_5 g07301(new_n9649, new_n9592, new_n9650);
nand_5 g07302(new_n9650, new_n9589, new_n9651);
nand_5 g07303(new_n9651, new_n9588, new_n9652);
nand_5 g07304(new_n9652, new_n9584, new_n9653);
nand_5 g07305(new_n9653, new_n9583, new_n9654);
xnor_4 g07306(new_n9654, new_n9578, n982);
not_8  g07307(n4306, new_n9656);
not_8  g07308(n3279, new_n9657);
not_8  g07309(n14702, new_n9658);
not_8  g07310(n2547, new_n9659);
not_8  g07311(n1667, new_n9660);
nor_5  g07312(n26808, n7339, new_n9661);
nand_5 g07313(new_n9661, new_n9660, new_n9662);
nor_5  g07314(new_n9662, n2680, new_n9663);
nand_5 g07315(new_n9663, new_n9659, new_n9664);
nor_5  g07316(new_n9664, n2999, new_n9665);
nand_5 g07317(new_n9665, new_n9658, new_n9666);
nor_5  g07318(new_n9666, n13914, new_n9667);
nand_5 g07319(new_n9667, new_n9657, new_n9668);
xnor_4 g07320(new_n9668, new_n9656, new_n9669);
not_8  g07321(new_n9669, new_n9670);
xnor_4 g07322(n23166, n18105, new_n9671);
not_8  g07323(n10577, new_n9672);
or_5   g07324(n24196, new_n9672, new_n9673);
xnor_4 g07325(n24196, n10577, new_n9674);
not_8  g07326(n6381, new_n9675);
or_5   g07327(n16376, new_n9675, new_n9676);
xnor_4 g07328(n16376, n6381, new_n9677);
not_8  g07329(n14345, new_n9678);
or_5   g07330(n25381, new_n9678, new_n9679);
xnor_4 g07331(n25381, n14345, new_n9680);
nand_5 g07332(new_n4687, n11356, new_n9681);
xnor_4 g07333(n12587, n11356, new_n9682);
not_8  g07334(n3164, new_n9683);
nor_5  g07335(new_n9683, n268, new_n9684);
xnor_4 g07336(n3164, n268, new_n9685);
not_8  g07337(new_n9685, new_n9686);
nor_5  g07338(n24879, new_n6944, new_n9687);
xnor_4 g07339(n24879, n10611, new_n9688);
not_8  g07340(new_n9688, new_n9689_1);
nor_5  g07341(new_n4650, n2783, new_n9690);
not_8  g07342(new_n9690, new_n9691);
nand_5 g07343(new_n4650, n2783, new_n9692);
not_8  g07344(n15490, new_n9693);
nand_5 g07345(n24032, new_n9693, new_n9694);
nand_5 g07346(new_n8549, n15490, new_n9695_1);
nor_5  g07347(new_n4704, n18, new_n9696);
nand_5 g07348(new_n9696, new_n9695_1, new_n9697);
nand_5 g07349(new_n9697, new_n9694, new_n9698);
nand_5 g07350(new_n9698, new_n9692, new_n9699_1);
nand_5 g07351(new_n9699_1, new_n9691, new_n9700);
nor_5  g07352(new_n9700, new_n9689_1, new_n9701);
nor_5  g07353(new_n9701, new_n9687, new_n9702);
nor_5  g07354(new_n9702, new_n9686, new_n9703);
nor_5  g07355(new_n9703, new_n9684, new_n9704);
not_8  g07356(new_n9704, new_n9705);
nand_5 g07357(new_n9705, new_n9682, new_n9706);
nand_5 g07358(new_n9706, new_n9681, new_n9707);
nand_5 g07359(new_n9707, new_n9680, new_n9708);
nand_5 g07360(new_n9708, new_n9679, new_n9709);
nand_5 g07361(new_n9709, new_n9677, new_n9710);
nand_5 g07362(new_n9710, new_n9676, new_n9711);
nand_5 g07363(new_n9711, new_n9674, new_n9712);
nand_5 g07364(new_n9712, new_n9673, new_n9713);
xnor_4 g07365(new_n9713, new_n9671, new_n9714);
xnor_4 g07366(new_n9714, new_n9670, new_n9715);
not_8  g07367(new_n9715, new_n9716);
xnor_4 g07368(new_n9667, n3279, new_n9717);
not_8  g07369(new_n9717, new_n9718);
xnor_4 g07370(new_n9711, new_n9674, new_n9719);
nor_5  g07371(new_n9719, new_n9718, new_n9720);
xnor_4 g07372(new_n9719, new_n9717, new_n9721);
not_8  g07373(new_n9721, new_n9722);
xnor_4 g07374(new_n9666, n13914, new_n9723);
xnor_4 g07375(new_n9709, new_n9677, new_n9724);
nand_5 g07376(new_n9724, new_n9723, new_n9725);
not_8  g07377(new_n9724, new_n9726_1);
xnor_4 g07378(new_n9726_1, new_n9723, new_n9727);
xnor_4 g07379(new_n9665, n14702, new_n9728);
not_8  g07380(new_n9728, new_n9729);
xnor_4 g07381(new_n9707, new_n9680, new_n9730);
nand_5 g07382(new_n9730, new_n9729, new_n9731);
xnor_4 g07383(new_n9730, new_n9728, new_n9732);
not_8  g07384(n2999, new_n9733);
xnor_4 g07385(new_n9664, new_n9733, new_n9734);
xnor_4 g07386(new_n9704, new_n9682, new_n9735);
nor_5  g07387(new_n9735, new_n9734, new_n9736);
not_8  g07388(new_n9736, new_n9737);
xnor_4 g07389(new_n9663, n2547, new_n9738);
xnor_4 g07390(new_n9702, new_n9685, new_n9739);
nor_5  g07391(new_n9739, new_n9738, new_n9740);
not_8  g07392(new_n9740, new_n9741);
not_8  g07393(new_n9739, new_n9742);
xnor_4 g07394(new_n9742, new_n9738, new_n9743);
xnor_4 g07395(new_n9662, n2680, new_n9744);
xnor_4 g07396(new_n9700, new_n9688, new_n9745);
not_8  g07397(new_n9745, new_n9746);
nand_5 g07398(new_n9746, new_n9744, new_n9747);
xnor_4 g07399(new_n9661, new_n9660, new_n9748);
xnor_4 g07400(n6785, new_n6947, new_n9749);
not_8  g07401(new_n9749, new_n9750);
xnor_4 g07402(new_n9750, new_n9698, new_n9751);
not_8  g07403(new_n9751, new_n9752);
nand_5 g07404(new_n9752, new_n9748, new_n9753_1);
xnor_4 g07405(new_n9751, new_n9748, new_n9754);
not_8  g07406(n7339, new_n9755);
xnor_4 g07407(n26808, new_n9755, new_n9756);
not_8  g07408(new_n9756, new_n9757);
xnor_4 g07409(n24032, n15490, new_n9758);
xnor_4 g07410(new_n9758, new_n9696, new_n9759);
not_8  g07411(new_n9759, new_n9760);
nor_5  g07412(new_n9760, new_n9757, new_n9761_1);
not_8  g07413(n26808, new_n9762);
xnor_4 g07414(n22843, n18, new_n9763_1);
nor_5  g07415(new_n9763_1, new_n9762, new_n9764);
not_8  g07416(new_n9764, new_n9765);
xnor_4 g07417(new_n9759, new_n9756, new_n9766);
nor_5  g07418(new_n9766, new_n9765, new_n9767_1);
nor_5  g07419(new_n9767_1, new_n9761_1, new_n9768);
nand_5 g07420(new_n9768, new_n9754, new_n9769);
nand_5 g07421(new_n9769, new_n9753_1, new_n9770);
xnor_4 g07422(new_n9745, new_n9744, new_n9771_1);
nand_5 g07423(new_n9771_1, new_n9770, new_n9772);
nand_5 g07424(new_n9772, new_n9747, new_n9773);
nand_5 g07425(new_n9773, new_n9743, new_n9774);
nand_5 g07426(new_n9774, new_n9741, new_n9775);
xnor_4 g07427(new_n9735, new_n9734, new_n9776);
not_8  g07428(new_n9776, new_n9777);
nand_5 g07429(new_n9777, new_n9775, new_n9778_1);
nand_5 g07430(new_n9778_1, new_n9737, new_n9779);
nand_5 g07431(new_n9779, new_n9732, new_n9780);
nand_5 g07432(new_n9780, new_n9731, new_n9781);
nand_5 g07433(new_n9781, new_n9727, new_n9782);
nand_5 g07434(new_n9782, new_n9725, new_n9783_1);
nor_5  g07435(new_n9783_1, new_n9722, new_n9784);
nor_5  g07436(new_n9784, new_n9720, new_n9785);
xnor_4 g07437(new_n9785, new_n9716, new_n9786);
xnor_4 g07438(new_n9786, new_n4745_1, new_n9787);
xnor_4 g07439(new_n9783_1, new_n9721, new_n9788);
not_8  g07440(new_n9788, new_n9789);
nand_5 g07441(new_n9789, new_n4751, new_n9790);
xnor_4 g07442(new_n9788, new_n4751, new_n9791);
xnor_4 g07443(new_n9781, new_n9727, new_n9792);
not_8  g07444(new_n9792, new_n9793);
nand_5 g07445(new_n9793, new_n4757, new_n9794);
xnor_4 g07446(new_n9792, new_n4757, new_n9795);
xnor_4 g07447(new_n9779, new_n9732, new_n9796);
not_8  g07448(new_n9796, new_n9797);
nand_5 g07449(new_n9797, new_n4763, new_n9798);
xnor_4 g07450(new_n9796, new_n4763, new_n9799);
xnor_4 g07451(new_n9776, new_n9775, new_n9800);
nand_5 g07452(new_n9800, new_n4769, new_n9801);
xnor_4 g07453(new_n9800, new_n4768, new_n9802);
xnor_4 g07454(new_n9773, new_n9743, new_n9803_1);
not_8  g07455(new_n9803_1, new_n9804);
nand_5 g07456(new_n9804, new_n4773, new_n9805);
xnor_4 g07457(new_n9804, new_n4772, new_n9806);
xnor_4 g07458(new_n9771_1, new_n9770, new_n9807);
nor_5  g07459(new_n9807, new_n4780, new_n9808);
not_8  g07460(new_n9808, new_n9809);
xnor_4 g07461(new_n9807, new_n4781, new_n9810);
not_8  g07462(new_n9754, new_n9811);
xnor_4 g07463(new_n9768, new_n9811, new_n9812);
nor_5  g07464(new_n9812, new_n4787, new_n9813);
xnor_4 g07465(new_n9812, new_n4787, new_n9814);
xnor_4 g07466(new_n9766, new_n9764, new_n9815);
and_5  g07467(new_n9815, new_n4790, new_n9816);
xnor_4 g07468(new_n9763_1, n26808, new_n9817);
and_5  g07469(new_n9817, new_n4795, new_n9818);
not_8  g07470(new_n9818, new_n9819);
xnor_4 g07471(new_n9815, new_n4790, new_n9820);
nor_5  g07472(new_n9820, new_n9819, new_n9821);
nor_5  g07473(new_n9821, new_n9816, new_n9822);
nor_5  g07474(new_n9822, new_n9814, new_n9823);
nor_5  g07475(new_n9823, new_n9813, new_n9824);
nand_5 g07476(new_n9824, new_n9810, new_n9825);
nand_5 g07477(new_n9825, new_n9809, new_n9826);
nand_5 g07478(new_n9826, new_n9806, new_n9827);
nand_5 g07479(new_n9827, new_n9805, new_n9828);
nand_5 g07480(new_n9828, new_n9802, new_n9829);
nand_5 g07481(new_n9829, new_n9801, new_n9830);
nand_5 g07482(new_n9830, new_n9799, new_n9831);
nand_5 g07483(new_n9831, new_n9798, new_n9832_1);
nand_5 g07484(new_n9832_1, new_n9795, new_n9833_1);
nand_5 g07485(new_n9833_1, new_n9794, new_n9834);
nand_5 g07486(new_n9834, new_n9791, new_n9835);
nand_5 g07487(new_n9835, new_n9790, new_n9836);
xnor_4 g07488(new_n9836, new_n9787, n984);
xnor_4 g07489(new_n9830, new_n9799, n1005);
xnor_4 g07490(new_n3513, new_n3458, n1016);
xnor_4 g07491(new_n4287, new_n4268, n1020);
xnor_4 g07492(n18290, new_n2903, new_n9841);
nor_5  g07493(n11580, n2035, new_n9842);
xnor_4 g07494(n11580, new_n2906, new_n9843);
not_8  g07495(new_n9843, new_n9844);
nor_5  g07496(n15884, n5213, new_n9845);
xnor_4 g07497(n15884, new_n2909, new_n9846);
not_8  g07498(new_n9846, new_n9847);
nor_5  g07499(n6356, n4665, new_n9848);
xnor_4 g07500(n6356, new_n2912, new_n9849);
not_8  g07501(new_n9849, new_n9850);
nor_5  g07502(n27104, n19005, new_n9851);
xnor_4 g07503(n27104, new_n2917, new_n9852);
not_8  g07504(new_n9852, new_n9853);
nor_5  g07505(n27188, n4326, new_n9854);
nand_5 g07506(n6611, n5438, new_n9855);
not_8  g07507(new_n9855, new_n9856);
xnor_4 g07508(n27188, n4326, new_n9857);
nor_5  g07509(new_n9857, new_n9856, new_n9858);
nor_5  g07510(new_n9858, new_n9854, new_n9859);
nor_5  g07511(new_n9859, new_n9853, new_n9860);
nor_5  g07512(new_n9860, new_n9851, new_n9861);
nor_5  g07513(new_n9861, new_n9850, new_n9862);
nor_5  g07514(new_n9862, new_n9848, new_n9863);
nor_5  g07515(new_n9863, new_n9847, new_n9864);
nor_5  g07516(new_n9864, new_n9845, new_n9865);
nor_5  g07517(new_n9865, new_n9844, new_n9866);
nor_5  g07518(new_n9866, new_n9842, new_n9867_1);
xnor_4 g07519(new_n9867_1, new_n9841, new_n9868);
xnor_4 g07520(new_n9868, n23529, new_n9869);
not_8  g07521(new_n9869, new_n9870);
xnor_4 g07522(new_n9865, new_n9843, new_n9871);
nand_5 g07523(new_n9871, new_n9541, new_n9872_1);
xnor_4 g07524(new_n9871, n24620, new_n9873);
xnor_4 g07525(new_n9863, new_n9846, new_n9874);
nand_5 g07526(new_n9874, new_n2955, new_n9875);
xnor_4 g07527(new_n9874, n5211, new_n9876);
xnor_4 g07528(new_n9861, new_n9849, new_n9877);
not_8  g07529(new_n9877, new_n9878);
nor_5  g07530(new_n9878, n12956, new_n9879);
xnor_4 g07531(new_n9877, n12956, new_n9880);
not_8  g07532(new_n9880, new_n9881);
xnor_4 g07533(new_n9859, new_n9852, new_n9882);
not_8  g07534(new_n9882, new_n9883);
nor_5  g07535(new_n9883, n18295, new_n9884);
not_8  g07536(new_n9884, new_n9885);
xnor_4 g07537(new_n9857, new_n9855, new_n9886);
nor_5  g07538(new_n9886, new_n9553, new_n9887);
not_8  g07539(n15780, new_n9888);
not_8  g07540(n5438, new_n9889);
xnor_4 g07541(n6611, new_n9889, new_n9890_1);
not_8  g07542(new_n9890_1, new_n9891);
nor_5  g07543(new_n9891, new_n9888, new_n9892);
not_8  g07544(new_n9892, new_n9893);
xnor_4 g07545(new_n9886, new_n9553, new_n9894);
nor_5  g07546(new_n9894, new_n9893, new_n9895);
nor_5  g07547(new_n9895, new_n9887, new_n9896);
xnor_4 g07548(new_n9882, n18295, new_n9897);
nand_5 g07549(new_n9897, new_n9896, new_n9898);
nand_5 g07550(new_n9898, new_n9885, new_n9899);
not_8  g07551(new_n9899, new_n9900);
nor_5  g07552(new_n9900, new_n9881, new_n9901);
nor_5  g07553(new_n9901, new_n9879, new_n9902);
not_8  g07554(new_n9902, new_n9903);
nand_5 g07555(new_n9903, new_n9876, new_n9904);
nand_5 g07556(new_n9904, new_n9875, new_n9905);
nand_5 g07557(new_n9905, new_n9873, new_n9906);
nand_5 g07558(new_n9906, new_n9872_1, new_n9907);
xnor_4 g07559(new_n9907, new_n9870, new_n9908);
not_8  g07560(n4409, new_n9909);
xnor_4 g07561(n17250, new_n9909, new_n9910);
nor_5  g07562(n23160, n3570, new_n9911);
not_8  g07563(n3570, new_n9912);
xnor_4 g07564(n23160, new_n9912, new_n9913);
not_8  g07565(new_n9913, new_n9914);
nor_5  g07566(n16524, n13668, new_n9915);
xnor_4 g07567(n16524, new_n6373, new_n9916);
not_8  g07568(new_n9916, new_n9917_1);
nor_5  g07569(n21276, n11056, new_n9918);
xnor_4 g07570(n21276, new_n6979, new_n9919_1);
not_8  g07571(new_n9919_1, new_n9920);
nor_5  g07572(n26748, n15271, new_n9921);
xnor_4 g07573(n26748, new_n8159_1, new_n9922);
not_8  g07574(new_n9922, new_n9923);
nor_5  g07575(n25877, n10057, new_n9924);
nand_5 g07576(n24323, n8920, new_n9925);
not_8  g07577(new_n9925, new_n9926_1);
xnor_4 g07578(n25877, n10057, new_n9927);
nor_5  g07579(new_n9927, new_n9926_1, new_n9928);
nor_5  g07580(new_n9928, new_n9924, new_n9929);
nor_5  g07581(new_n9929, new_n9923, new_n9930);
nor_5  g07582(new_n9930, new_n9921, new_n9931);
nor_5  g07583(new_n9931, new_n9920, new_n9932);
nor_5  g07584(new_n9932, new_n9918, new_n9933);
nor_5  g07585(new_n9933, new_n9917_1, new_n9934_1);
nor_5  g07586(new_n9934_1, new_n9915, new_n9935);
nor_5  g07587(new_n9935, new_n9914, new_n9936);
nor_5  g07588(new_n9936, new_n9911, new_n9937);
xnor_4 g07589(new_n9937, new_n9910, new_n9938_1);
xnor_4 g07590(new_n9938_1, n11044, new_n9939);
not_8  g07591(new_n9939, new_n9940);
xnor_4 g07592(new_n9935, new_n9913, new_n9941);
nor_5  g07593(new_n9941, new_n6322, new_n9942_1);
xnor_4 g07594(new_n9941, n2421, new_n9943);
not_8  g07595(new_n9943, new_n9944);
xnor_4 g07596(new_n9933, new_n9917_1, new_n9945);
not_8  g07597(new_n9945, new_n9946_1);
nor_5  g07598(new_n9946_1, new_n8152, new_n9947);
xnor_4 g07599(new_n9945, new_n8152, new_n9948);
not_8  g07600(new_n9948, new_n9949);
xnor_4 g07601(new_n9931, new_n9919_1, new_n9950);
nor_5  g07602(new_n9950, new_n8156, new_n9951);
xnor_4 g07603(new_n9950, n20478, new_n9952);
not_8  g07604(new_n9952, new_n9953);
xnor_4 g07605(new_n9929, new_n9922, new_n9954);
nor_5  g07606(new_n9954, new_n8161, new_n9955);
xnor_4 g07607(new_n9927, new_n9925, new_n9956);
not_8  g07608(new_n9956, new_n9957);
nor_5  g07609(new_n9957, n22619, new_n9958);
not_8  g07610(new_n9958, new_n9959);
xnor_4 g07611(n24323, new_n4452, new_n9960);
not_8  g07612(new_n9960, new_n9961);
nor_5  g07613(new_n9961, new_n6107, new_n9962);
not_8  g07614(new_n9962, new_n9963);
xnor_4 g07615(new_n9956, n22619, new_n9964);
nand_5 g07616(new_n9964, new_n9963, new_n9965);
nand_5 g07617(new_n9965, new_n9959, new_n9966);
xnor_4 g07618(new_n9954, new_n8161, new_n9967_1);
nor_5  g07619(new_n9967_1, new_n9966, new_n9968_1);
nor_5  g07620(new_n9968_1, new_n9955, new_n9969);
nor_5  g07621(new_n9969, new_n9953, new_n9970);
nor_5  g07622(new_n9970, new_n9951, new_n9971);
nor_5  g07623(new_n9971, new_n9949, new_n9972);
nor_5  g07624(new_n9972, new_n9947, new_n9973);
nor_5  g07625(new_n9973, new_n9944, new_n9974);
nor_5  g07626(new_n9974, new_n9942_1, new_n9975);
xnor_4 g07627(new_n9975, new_n9940, new_n9976);
xnor_4 g07628(new_n9976, new_n9908, new_n9977);
not_8  g07629(new_n9873, new_n9978);
xnor_4 g07630(new_n9905, new_n9978, new_n9979);
xnor_4 g07631(new_n9973, new_n9943, new_n9980);
nand_5 g07632(new_n9980, new_n9979, new_n9981);
not_8  g07633(new_n9980, new_n9982);
xnor_4 g07634(new_n9982, new_n9979, new_n9983);
xnor_4 g07635(new_n9902, new_n9876, new_n9984);
xnor_4 g07636(new_n9971, new_n9948, new_n9985);
and_5  g07637(new_n9985, new_n9984, new_n9986);
not_8  g07638(new_n9985, new_n9987);
xnor_4 g07639(new_n9987, new_n9984, new_n9988);
not_8  g07640(new_n9988, new_n9989);
xnor_4 g07641(new_n9900, new_n9880, new_n9990);
xnor_4 g07642(new_n9969, new_n9952, new_n9991);
and_5  g07643(new_n9991, new_n9990, new_n9992);
not_8  g07644(new_n9991, new_n9993);
xnor_4 g07645(new_n9993, new_n9990, new_n9994);
not_8  g07646(new_n9994, new_n9995);
xnor_4 g07647(new_n9897, new_n9896, new_n9996);
xnor_4 g07648(new_n9967_1, new_n9966, new_n9997);
nor_5  g07649(new_n9997, new_n9996, new_n9998);
not_8  g07650(new_n9997, new_n9999);
xnor_4 g07651(new_n9999, new_n9996, new_n10000);
not_8  g07652(new_n10000, new_n10001);
xnor_4 g07653(new_n9964, new_n9962, new_n10002);
xnor_4 g07654(new_n9894, new_n9892, new_n10003);
nor_5  g07655(new_n10003, new_n10002, new_n10004);
xnor_4 g07656(new_n9960, new_n6107, new_n10005);
not_8  g07657(new_n10005, new_n10006);
xnor_4 g07658(new_n9890_1, new_n9888, new_n10007);
nor_5  g07659(new_n10007, new_n10006, new_n10008);
not_8  g07660(new_n10008, new_n10009_1);
not_8  g07661(new_n10002, new_n10010_1);
xnor_4 g07662(new_n10003, new_n10010_1, new_n10011);
not_8  g07663(new_n10011, new_n10012);
nor_5  g07664(new_n10012, new_n10009_1, new_n10013);
nor_5  g07665(new_n10013, new_n10004, new_n10014);
nor_5  g07666(new_n10014, new_n10001, new_n10015);
nor_5  g07667(new_n10015, new_n9998, new_n10016);
nor_5  g07668(new_n10016, new_n9995, new_n10017_1);
nor_5  g07669(new_n10017_1, new_n9992, new_n10018_1);
nor_5  g07670(new_n10018_1, new_n9989, new_n10019_1);
nor_5  g07671(new_n10019_1, new_n9986, new_n10020);
not_8  g07672(new_n10020, new_n10021_1);
nand_5 g07673(new_n10021_1, new_n9983, new_n10022);
nand_5 g07674(new_n10022, new_n9981, new_n10023);
xnor_4 g07675(new_n10023, new_n9977, n1044);
nor_5  g07676(n22619, n6775, new_n10025);
nand_5 g07677(new_n10025, new_n8161, new_n10026);
xnor_4 g07678(new_n10026, new_n8156, new_n10027);
xnor_4 g07679(new_n10027, new_n5176, new_n10028);
xnor_4 g07680(new_n10025, n26882, new_n10029);
nand_5 g07681(new_n10029, n25872, new_n10030);
xnor_4 g07682(new_n10029, new_n5181, new_n10031);
xnor_4 g07683(n22619, n6775, new_n10032);
nor_5  g07684(new_n10032, new_n5187, new_n10033);
not_8  g07685(new_n10033, new_n10034);
nand_5 g07686(n6775, n3925, new_n10035);
not_8  g07687(new_n10035, new_n10036);
xnor_4 g07688(new_n10032, n20259, new_n10037);
nand_5 g07689(new_n10037, new_n10036, new_n10038);
nand_5 g07690(new_n10038, new_n10034, new_n10039);
nand_5 g07691(new_n10039, new_n10031, new_n10040);
nand_5 g07692(new_n10040, new_n10030, new_n10041);
xnor_4 g07693(new_n10041, new_n10028, new_n10042);
nor_5  g07694(n9399, n2088, new_n10043);
nand_5 g07695(new_n10043, new_n4521, new_n10044);
xnor_4 g07696(new_n10044, new_n4516, new_n10045);
xnor_4 g07697(new_n10045, new_n2398, new_n10046);
xnor_4 g07698(new_n10043, n16396, new_n10047);
not_8  g07699(new_n10047, new_n10048);
nor_5  g07700(new_n10048, new_n8110, new_n10049);
xnor_4 g07701(new_n10047, new_n8110, new_n10050);
not_8  g07702(new_n10050, new_n10051);
not_8  g07703(new_n6099, new_n10052);
nor_5  g07704(new_n6101, new_n10052, new_n10053_1);
nand_5 g07705(new_n10053_1, new_n6096, new_n10054);
nand_5 g07706(new_n10054, new_n6099, new_n10055_1);
nor_5  g07707(new_n10055_1, new_n10051, new_n10056);
nor_5  g07708(new_n10056, new_n10049, new_n10057_1);
xnor_4 g07709(new_n10057_1, new_n10046, new_n10058);
xnor_4 g07710(new_n10058, new_n10042, new_n10059);
xnor_4 g07711(new_n10055_1, new_n10051, new_n10060);
not_8  g07712(new_n10060, new_n10061);
xnor_4 g07713(new_n10039, new_n10031, new_n10062);
not_8  g07714(new_n10062, new_n10063);
nand_5 g07715(new_n10063, new_n10061, new_n10064);
xnor_4 g07716(new_n10062, new_n10061, new_n10065);
not_8  g07717(new_n6104_1, new_n10066);
xnor_4 g07718(new_n10037, new_n10036, new_n10067);
not_8  g07719(new_n10067, new_n10068);
nand_5 g07720(new_n10068, new_n10066, new_n10069);
xnor_4 g07721(n6775, new_n6158, new_n10070);
not_8  g07722(new_n10070, new_n10071);
nor_5  g07723(new_n10071, new_n6084_1, new_n10072);
xnor_4 g07724(new_n10067, new_n10066, new_n10073);
nand_5 g07725(new_n10073, new_n10072, new_n10074);
nand_5 g07726(new_n10074, new_n10069, new_n10075);
nand_5 g07727(new_n10075, new_n10065, new_n10076);
nand_5 g07728(new_n10076, new_n10064, new_n10077);
xnor_4 g07729(new_n10077, new_n10059, new_n10078);
not_8  g07730(new_n10078, new_n10079);
xnor_4 g07731(n12956, n7057, new_n10080);
nor_5  g07732(new_n2963, n8381, new_n10081);
nor_5  g07733(n18295, new_n5296, new_n10082);
nor_5  g07734(n20235, new_n9553, new_n10083);
not_8  g07735(new_n10083, new_n10084);
nor_5  g07736(new_n5307, n6502, new_n10085);
not_8  g07737(new_n10085, new_n10086);
nor_5  g07738(new_n9888, n12495, new_n10087);
nand_5 g07739(new_n10087, new_n10086, new_n10088);
nand_5 g07740(new_n10088, new_n10084, new_n10089);
not_8  g07741(new_n10089, new_n10090);
nor_5  g07742(new_n10090, new_n10082, new_n10091);
nor_5  g07743(new_n10091, new_n10081, new_n10092);
xnor_4 g07744(new_n10092, new_n10080, new_n10093);
xnor_4 g07745(new_n10093, new_n10079, new_n10094);
xnor_4 g07746(new_n10075, new_n10065, new_n10095);
not_8  g07747(new_n10095, new_n10096_1);
xnor_4 g07748(n18295, n8381, new_n10097);
xnor_4 g07749(new_n10097, new_n10090, new_n10098);
not_8  g07750(new_n10098, new_n10099);
nor_5  g07751(new_n10099, new_n10096_1, new_n10100);
not_8  g07752(new_n10100, new_n10101_1);
xnor_4 g07753(new_n10099, new_n10095, new_n10102);
xnor_4 g07754(n15780, n12495, new_n10103);
xnor_4 g07755(new_n10070, new_n6084_1, new_n10104);
not_8  g07756(new_n10104, new_n10105);
nor_5  g07757(new_n10105, new_n10103, new_n10106);
xnor_4 g07758(n20235, n6502, new_n10107);
xnor_4 g07759(new_n10107, new_n10087, new_n10108);
nor_5  g07760(new_n10108, new_n10106, new_n10109);
xnor_4 g07761(new_n10073, new_n10072, new_n10110);
xnor_4 g07762(new_n10108, new_n10106, new_n10111_1);
not_8  g07763(new_n10111_1, new_n10112);
nand_5 g07764(new_n10112, new_n10110, new_n10113);
not_8  g07765(new_n10113, new_n10114);
nor_5  g07766(new_n10114, new_n10109, new_n10115);
not_8  g07767(new_n10115, new_n10116);
nand_5 g07768(new_n10116, new_n10102, new_n10117_1);
nand_5 g07769(new_n10117_1, new_n10101_1, new_n10118);
xnor_4 g07770(new_n10118, new_n10094, n1060);
xnor_4 g07771(new_n3511, new_n3463, n1069);
not_8  g07772(n3959, new_n10121);
xnor_4 g07773(n9832, new_n10121, new_n10122);
nor_5  g07774(n11566, n1558, new_n10123);
not_8  g07775(n1558, new_n10124);
xnor_4 g07776(n11566, new_n10124, new_n10125_1);
not_8  g07777(new_n10125_1, new_n10126);
nor_5  g07778(n26744, n21749, new_n10127);
not_8  g07779(n21749, new_n10128);
xnor_4 g07780(n26744, new_n10128, new_n10129);
not_8  g07781(new_n10129, new_n10130);
nor_5  g07782(n26625, n7769, new_n10131);
nand_5 g07783(n21138, n14230, new_n10132);
not_8  g07784(n7769, new_n10133);
xnor_4 g07785(n26625, new_n10133, new_n10134);
and_5  g07786(new_n10134, new_n10132, new_n10135);
nor_5  g07787(new_n10135, new_n10131, new_n10136);
nor_5  g07788(new_n10136, new_n10130, new_n10137);
nor_5  g07789(new_n10137, new_n10127, new_n10138);
nor_5  g07790(new_n10138, new_n10126, new_n10139);
nor_5  g07791(new_n10139, new_n10123, new_n10140);
xnor_4 g07792(new_n10140, new_n10122, new_n10141);
not_8  g07793(n17095, new_n10142);
nor_5  g07794(n26167, n22591, new_n10143);
nand_5 g07795(new_n10143, new_n10142, new_n10144);
nor_5  g07796(new_n10144, n15378, new_n10145);
xnor_4 g07797(new_n10145, n19575, new_n10146);
xnor_4 g07798(new_n7171, new_n2603, new_n10147);
not_8  g07799(n17664, new_n10148);
nor_5  g07800(new_n7181, new_n10148, new_n10149);
not_8  g07801(new_n10149, new_n10150);
xnor_4 g07802(new_n7181, n17664, new_n10151);
nor_5  g07803(new_n7186, new_n2610, new_n10152);
not_8  g07804(new_n10152, new_n10153);
xnor_4 g07805(new_n7186, n23369, new_n10154);
not_8  g07806(new_n7194, new_n10155);
nand_5 g07807(new_n10155, new_n9252, new_n10156);
not_8  g07808(new_n10156, new_n10157);
nor_5  g07809(new_n7191, new_n7636, new_n10158_1);
xnor_4 g07810(new_n7194, n1136, new_n10159);
nor_5  g07811(new_n10159, new_n10158_1, new_n10160);
nor_5  g07812(new_n10160, new_n10157, new_n10161);
nand_5 g07813(new_n10161, new_n10154, new_n10162);
nand_5 g07814(new_n10162, new_n10153, new_n10163);
nand_5 g07815(new_n10163, new_n10151, new_n10164);
nand_5 g07816(new_n10164, new_n10150, new_n10165_1);
not_8  g07817(new_n10165_1, new_n10166);
xnor_4 g07818(new_n10166, new_n10147, new_n10167);
xnor_4 g07819(new_n10167, new_n10146, new_n10168);
xnor_4 g07820(new_n7181, new_n10148, new_n10169);
xnor_4 g07821(new_n10163, new_n10169, new_n10170);
not_8  g07822(n15378, new_n10171);
xnor_4 g07823(new_n10144, new_n10171, new_n10172);
nor_5  g07824(new_n10172, new_n10170, new_n10173);
xnor_4 g07825(new_n10172, new_n10170, new_n10174);
xnor_4 g07826(new_n7186, new_n2610, new_n10175);
xnor_4 g07827(new_n10161, new_n10175, new_n10176);
xnor_4 g07828(new_n10143, n17095, new_n10177);
nor_5  g07829(new_n10177, new_n10176, new_n10178);
xnor_4 g07830(new_n10177, new_n10176, new_n10179);
not_8  g07831(new_n10159, new_n10180);
xnor_4 g07832(new_n10180, new_n10158_1, new_n10181);
not_8  g07833(new_n10181, new_n10182);
not_8  g07834(n22591, new_n10183);
not_8  g07835(n26167, new_n10184);
not_8  g07836(new_n7637, new_n10185);
nor_5  g07837(new_n10185, new_n10184, new_n10186);
xnor_4 g07838(new_n10186, new_n10183, new_n10187);
nand_5 g07839(new_n10187, new_n10182, new_n10188);
nor_5  g07840(new_n7637, new_n10184, new_n10189);
nand_5 g07841(new_n10189, new_n10183, new_n10190);
nand_5 g07842(new_n10190, new_n10188, new_n10191);
nor_5  g07843(new_n10191, new_n10179, new_n10192);
nor_5  g07844(new_n10192, new_n10178, new_n10193);
nor_5  g07845(new_n10193, new_n10174, new_n10194);
nor_5  g07846(new_n10194, new_n10173, new_n10195);
xnor_4 g07847(new_n10195, new_n10168, new_n10196);
xnor_4 g07848(new_n10196, new_n10141, new_n10197);
xnor_4 g07849(new_n10193, new_n10174, new_n10198);
xnor_4 g07850(new_n10138, new_n10125_1, new_n10199);
nor_5  g07851(new_n10199, new_n10198, new_n10200);
not_8  g07852(new_n10200, new_n10201_1);
not_8  g07853(new_n10199, new_n10202);
xnor_4 g07854(new_n10202, new_n10198, new_n10203);
not_8  g07855(new_n10191, new_n10204);
xnor_4 g07856(new_n10204, new_n10179, new_n10205);
xnor_4 g07857(new_n10136, new_n10129, new_n10206);
not_8  g07858(new_n10206, new_n10207);
nor_5  g07859(new_n10207, new_n10205, new_n10208);
xnor_4 g07860(new_n10207, new_n10205, new_n10209);
xnor_4 g07861(new_n10187, new_n10181, new_n10210);
not_8  g07862(new_n10132, new_n10211);
xnor_4 g07863(new_n10134, new_n10211, new_n10212);
nor_5  g07864(new_n10212, new_n10210, new_n10213);
not_8  g07865(new_n10213, new_n10214);
nor_5  g07866(new_n7638, new_n7635, new_n10215);
not_8  g07867(new_n10212, new_n10216);
xnor_4 g07868(new_n10216, new_n10210, new_n10217);
nand_5 g07869(new_n10217, new_n10215, new_n10218);
nand_5 g07870(new_n10218, new_n10214, new_n10219);
nor_5  g07871(new_n10219, new_n10209, new_n10220);
nor_5  g07872(new_n10220, new_n10208, new_n10221);
nand_5 g07873(new_n10221, new_n10203, new_n10222);
nand_5 g07874(new_n10222, new_n10201_1, new_n10223);
xor_4  g07875(new_n10223, new_n10197, n1111);
xnor_4 g07876(new_n2638, n25475, new_n10225);
nor_5  g07877(new_n2644, new_n4623, new_n10226);
xnor_4 g07878(new_n2644, new_n4623, new_n10227);
nor_5  g07879(new_n2649, new_n4627, new_n10228);
nand_5 g07880(new_n2654, new_n4631, new_n10229);
xnor_4 g07881(new_n2654, n11011, new_n10230);
nand_5 g07882(new_n2659_1, new_n4104, new_n10231);
xnor_4 g07883(new_n2659_1, n16029, new_n10232);
nor_5  g07884(new_n2665, new_n4109, new_n10233);
xnor_4 g07885(new_n2665, n16476, new_n10234);
not_8  g07886(new_n10234, new_n10235);
nor_5  g07887(new_n2670, new_n4115, new_n10236_1);
nand_5 g07888(new_n2672, new_n4120, new_n10237);
nor_5  g07889(new_n2677, new_n2580, new_n10238);
not_8  g07890(new_n10238, new_n10239_1);
xnor_4 g07891(new_n2672, n22433, new_n10240);
nand_5 g07892(new_n10240, new_n10239_1, new_n10241);
nand_5 g07893(new_n10241, new_n10237, new_n10242);
xnor_4 g07894(new_n2670, n11615, new_n10243);
not_8  g07895(new_n10243, new_n10244_1);
nor_5  g07896(new_n10244_1, new_n10242, new_n10245);
nor_5  g07897(new_n10245, new_n10236_1, new_n10246);
nor_5  g07898(new_n10246, new_n10235, new_n10247);
nor_5  g07899(new_n10247, new_n10233, new_n10248);
nand_5 g07900(new_n10248, new_n10232, new_n10249);
nand_5 g07901(new_n10249, new_n10231, new_n10250_1);
nand_5 g07902(new_n10250_1, new_n10230, new_n10251);
nand_5 g07903(new_n10251, new_n10229, new_n10252);
xnor_4 g07904(new_n2649, new_n4627, new_n10253);
nor_5  g07905(new_n10253, new_n10252, new_n10254);
nor_5  g07906(new_n10254, new_n10228, new_n10255);
nor_5  g07907(new_n10255, new_n10227, new_n10256);
nor_5  g07908(new_n10256, new_n10226, new_n10257);
xnor_4 g07909(new_n10257, new_n10225, new_n10258);
nor_5  g07910(new_n10044, n25074, new_n10259);
nand_5 g07911(new_n10259, new_n3002, new_n10260);
nor_5  g07912(new_n10260, n20929, new_n10261_1);
nand_5 g07913(new_n10261_1, new_n2994, new_n10262_1);
nor_5  g07914(new_n10262_1, n11841, new_n10263);
xnor_4 g07915(new_n10263, n27089, new_n10264);
xnor_4 g07916(new_n10264, new_n2771, new_n10265);
xnor_4 g07917(new_n10262_1, new_n2990, new_n10266);
not_8  g07918(new_n10266, new_n10267);
nor_5  g07919(new_n10267, new_n2776, new_n10268);
xnor_4 g07920(new_n10266, new_n2775, new_n10269);
xnor_4 g07921(new_n10261_1, n10710, new_n10270);
nor_5  g07922(new_n10270, new_n2780, new_n10271);
not_8  g07923(new_n10270, new_n10272);
xnor_4 g07924(new_n10272, new_n2780, new_n10273);
not_8  g07925(new_n10273, new_n10274);
xnor_4 g07926(new_n10260, new_n2998, new_n10275_1);
nor_5  g07927(new_n10275_1, new_n2785, new_n10276);
not_8  g07928(new_n10275_1, new_n10277);
xnor_4 g07929(new_n10277, new_n2785, new_n10278);
not_8  g07930(new_n10278, new_n10279);
xnor_4 g07931(new_n10259, n8006, new_n10280);
nor_5  g07932(new_n10280, new_n2790, new_n10281);
nor_5  g07933(new_n10045, new_n2794, new_n10282);
not_8  g07934(new_n10045, new_n10283);
xnor_4 g07935(new_n10283, new_n2794, new_n10284);
not_8  g07936(new_n10284, new_n10285);
nor_5  g07937(new_n10047, new_n2798, new_n10286);
xnor_4 g07938(new_n10048, new_n2798, new_n10287_1);
not_8  g07939(new_n10287_1, new_n10288);
nor_5  g07940(new_n6095, new_n2803, new_n10289);
nor_5  g07941(new_n2807, n2088, new_n10290);
xnor_4 g07942(new_n6096, new_n2803, new_n10291);
nand_5 g07943(new_n10291, new_n10290, new_n10292);
not_8  g07944(new_n10292, new_n10293);
nor_5  g07945(new_n10293, new_n10289, new_n10294);
nor_5  g07946(new_n10294, new_n10288, new_n10295_1);
nor_5  g07947(new_n10295_1, new_n10286, new_n10296);
nor_5  g07948(new_n10296, new_n10285, new_n10297);
nor_5  g07949(new_n10297, new_n10282, new_n10298);
not_8  g07950(new_n10280, new_n10299);
xnor_4 g07951(new_n10299, new_n2790, new_n10300);
not_8  g07952(new_n10300, new_n10301);
nor_5  g07953(new_n10301, new_n10298, new_n10302);
nor_5  g07954(new_n10302, new_n10281, new_n10303);
nor_5  g07955(new_n10303, new_n10279, new_n10304);
nor_5  g07956(new_n10304, new_n10276, new_n10305);
nor_5  g07957(new_n10305, new_n10274, new_n10306);
nor_5  g07958(new_n10306, new_n10271, new_n10307);
not_8  g07959(new_n10307, new_n10308);
nor_5  g07960(new_n10308, new_n10269, new_n10309);
nor_5  g07961(new_n10309, new_n10268, new_n10310);
xnor_4 g07962(new_n10310, new_n10265, new_n10311);
xnor_4 g07963(new_n10311, new_n10258, new_n10312);
xnor_4 g07964(new_n10255, new_n10227, new_n10313);
xnor_4 g07965(new_n10307, new_n10269, new_n10314);
not_8  g07966(new_n10314, new_n10315);
nor_5  g07967(new_n10315, new_n10313, new_n10316);
not_8  g07968(new_n10316, new_n10317);
xnor_4 g07969(new_n10314, new_n10313, new_n10318);
xnor_4 g07970(new_n10253, new_n10252, new_n10319);
not_8  g07971(new_n10319, new_n10320);
xnor_4 g07972(new_n10305, new_n10274, new_n10321_1);
nor_5  g07973(new_n10321_1, new_n10320, new_n10322);
xnor_4 g07974(new_n10321_1, new_n10320, new_n10323);
xnor_4 g07975(new_n2654, new_n4631, new_n10324);
xnor_4 g07976(new_n10250_1, new_n10324, new_n10325);
xnor_4 g07977(new_n10303, new_n10279, new_n10326_1);
not_8  g07978(new_n10326_1, new_n10327_1);
nor_5  g07979(new_n10327_1, new_n10325, new_n10328);
not_8  g07980(new_n10328, new_n10329);
xnor_4 g07981(new_n10326_1, new_n10325, new_n10330_1);
xnor_4 g07982(new_n10248, new_n10232, new_n10331);
not_8  g07983(new_n10331, new_n10332);
xnor_4 g07984(new_n10300, new_n10298, new_n10333);
nor_5  g07985(new_n10333, new_n10332, new_n10334);
not_8  g07986(new_n10334, new_n10335);
xnor_4 g07987(new_n10333, new_n10331, new_n10336);
xnor_4 g07988(new_n10296, new_n10284, new_n10337);
xnor_4 g07989(new_n10246, new_n10235, new_n10338);
nor_5  g07990(new_n10338, new_n10337, new_n10339);
not_8  g07991(new_n10339, new_n10340_1);
not_8  g07992(new_n10338, new_n10341);
xnor_4 g07993(new_n10341, new_n10337, new_n10342);
xnor_4 g07994(new_n10294, new_n10287_1, new_n10343);
xnor_4 g07995(new_n10243, new_n10242, new_n10344);
not_8  g07996(new_n10344, new_n10345_1);
nor_5  g07997(new_n10345_1, new_n10343, new_n10346);
not_8  g07998(new_n10346, new_n10347);
xnor_4 g07999(new_n10344, new_n10343, new_n10348);
xnor_4 g08000(new_n10291, new_n10290, new_n10349);
xnor_4 g08001(new_n10240, new_n10238, new_n10350);
not_8  g08002(new_n10350, new_n10351);
nor_5  g08003(new_n10351, new_n10349, new_n10352);
xnor_4 g08004(new_n2677, n14090, new_n10353);
not_8  g08005(new_n10353, new_n10354);
xnor_4 g08006(new_n2806, n2088, new_n10355);
nor_5  g08007(new_n10355, new_n10354, new_n10356_1);
xnor_4 g08008(new_n10350, new_n10349, new_n10357);
not_8  g08009(new_n10357, new_n10358);
nor_5  g08010(new_n10358, new_n10356_1, new_n10359);
nor_5  g08011(new_n10359, new_n10352, new_n10360);
nand_5 g08012(new_n10360, new_n10348, new_n10361);
nand_5 g08013(new_n10361, new_n10347, new_n10362);
nand_5 g08014(new_n10362, new_n10342, new_n10363);
nand_5 g08015(new_n10363, new_n10340_1, new_n10364);
nand_5 g08016(new_n10364, new_n10336, new_n10365);
nand_5 g08017(new_n10365, new_n10335, new_n10366);
nand_5 g08018(new_n10366, new_n10330_1, new_n10367);
nand_5 g08019(new_n10367, new_n10329, new_n10368);
nor_5  g08020(new_n10368, new_n10323, new_n10369);
nor_5  g08021(new_n10369, new_n10322, new_n10370);
nand_5 g08022(new_n10370, new_n10318, new_n10371);
nand_5 g08023(new_n10371, new_n10317, new_n10372_1);
xnor_4 g08024(new_n10372_1, new_n10312, n1119);
xnor_4 g08025(new_n8375, new_n8370, new_n10374);
xnor_4 g08026(new_n10374, new_n8400, n1120);
xnor_4 g08027(n9246, new_n6158, new_n10376);
xnor_4 g08028(new_n10376, new_n8243, new_n10377);
xnor_4 g08029(n12495, n7428, new_n10378);
xnor_4 g08030(new_n10378, new_n10377, n1196);
xnor_4 g08031(n16223, n15636, new_n10380);
nor_5  g08032(new_n5809, n19494, new_n10381);
nor_5  g08033(n20077, new_n2366, new_n10382);
nand_5 g08034(n6794, new_n2368, new_n10383);
nor_5  g08035(new_n10383, new_n10382, new_n10384);
nor_5  g08036(new_n10384, new_n10381, new_n10385_1);
xnor_4 g08037(new_n10385_1, new_n10380, new_n10386);
xnor_4 g08038(new_n10386, new_n8397, new_n10387_1);
xnor_4 g08039(n6794, n2387, new_n10388_1);
nor_5  g08040(new_n10388_1, new_n8387, new_n10389);
xnor_4 g08041(n20077, n19494, new_n10390_1);
xnor_4 g08042(new_n10390_1, new_n10383, new_n10391);
not_8  g08043(new_n10391, new_n10392);
nor_5  g08044(new_n10392, new_n10389, new_n10393);
xnor_4 g08045(new_n10391, new_n10389, new_n10394);
not_8  g08046(new_n10394, new_n10395);
nor_5  g08047(new_n10395, new_n8380, new_n10396);
nor_5  g08048(new_n10396, new_n10393, new_n10397);
not_8  g08049(new_n10397, new_n10398);
xnor_4 g08050(new_n10398, new_n10387_1, n1237);
xnor_4 g08051(new_n6001, new_n5785, new_n10400);
xnor_4 g08052(new_n10400, new_n6078, n1239);
not_8  g08053(n2416, new_n10402);
xnor_4 g08054(n22764, new_n8573, new_n10403);
not_8  g08055(new_n10403, new_n10404_1);
or_5   g08056(n26264, n19454, new_n10405_1);
xnor_4 g08057(n26264, new_n8577, new_n10406);
or_5   g08058(n9445, n7841, new_n10407);
xnor_4 g08059(n9445, new_n8470, new_n10408);
nor_5  g08060(n16812, n1279, new_n10409_1);
xnor_4 g08061(n16812, new_n8585, new_n10410);
not_8  g08062(new_n10410, new_n10411_1);
nor_5  g08063(n25068, n8324, new_n10412);
xnor_4 g08064(n25068, new_n8589, new_n10413);
not_8  g08065(new_n10413, new_n10414);
nor_5  g08066(n12546, n2331, new_n10415);
xnor_4 g08067(n12546, new_n8488, new_n10416);
not_8  g08068(new_n10416, new_n10417);
nor_5  g08069(n22631, n21078, new_n10418);
xnor_4 g08070(n22631, new_n8597, new_n10419);
not_8  g08071(new_n10419, new_n10420_1);
nor_5  g08072(n24485, n16743, new_n10421);
xnor_4 g08073(n24485, new_n8495, new_n10422);
not_8  g08074(new_n10422, new_n10423);
nor_5  g08075(n15258, n2420, new_n10424);
nand_5 g08076(n22201, n4588, new_n10425);
not_8  g08077(new_n10425, new_n10426);
xnor_4 g08078(n15258, n2420, new_n10427);
nor_5  g08079(new_n10427, new_n10426, new_n10428);
nor_5  g08080(new_n10428, new_n10424, new_n10429);
nor_5  g08081(new_n10429, new_n10423, new_n10430);
nor_5  g08082(new_n10430, new_n10421, new_n10431);
nor_5  g08083(new_n10431, new_n10420_1, new_n10432_1);
nor_5  g08084(new_n10432_1, new_n10418, new_n10433);
nor_5  g08085(new_n10433, new_n10417, new_n10434);
nor_5  g08086(new_n10434, new_n10415, new_n10435);
nor_5  g08087(new_n10435, new_n10414, new_n10436);
nor_5  g08088(new_n10436, new_n10412, new_n10437);
nor_5  g08089(new_n10437, new_n10411_1, new_n10438);
nor_5  g08090(new_n10438, new_n10409_1, new_n10439);
not_8  g08091(new_n10439, new_n10440);
nand_5 g08092(new_n10440, new_n10408, new_n10441);
nand_5 g08093(new_n10441, new_n10407, new_n10442);
nand_5 g08094(new_n10442, new_n10406, new_n10443);
nand_5 g08095(new_n10443, new_n10405_1, new_n10444);
xnor_4 g08096(new_n10444, new_n10404_1, new_n10445);
nand_5 g08097(new_n10445, new_n10402, new_n10446);
xnor_4 g08098(new_n10445, n2416, new_n10447);
not_8  g08099(n21905, new_n10448);
not_8  g08100(new_n10406, new_n10449);
xnor_4 g08101(new_n10442, new_n10449, new_n10450);
nand_5 g08102(new_n10450, new_n10448, new_n10451);
xnor_4 g08103(new_n10450, n21905, new_n10452);
not_8  g08104(n22918, new_n10453);
xnor_4 g08105(new_n10439, new_n10408, new_n10454);
nand_5 g08106(new_n10454, new_n10453, new_n10455);
xnor_4 g08107(new_n10454, n22918, new_n10456);
not_8  g08108(n25923, new_n10457);
xnor_4 g08109(new_n10437, new_n10410, new_n10458);
nand_5 g08110(new_n10458, new_n10457, new_n10459);
xnor_4 g08111(new_n10458, n25923, new_n10460);
not_8  g08112(n6790, new_n10461);
xnor_4 g08113(new_n10435, new_n10413, new_n10462);
nand_5 g08114(new_n10462, new_n10461, new_n10463);
xnor_4 g08115(new_n10462, n6790, new_n10464);
not_8  g08116(n22879, new_n10465);
xnor_4 g08117(new_n10433, new_n10416, new_n10466);
nand_5 g08118(new_n10466, new_n10465, new_n10467);
xnor_4 g08119(new_n10466, n22879, new_n10468);
not_8  g08120(n2117, new_n10469);
xnor_4 g08121(new_n10431, new_n10419, new_n10470);
nand_5 g08122(new_n10470, new_n10469, new_n10471);
not_8  g08123(new_n10471, new_n10472);
xnor_4 g08124(new_n10470, n2117, new_n10473);
not_8  g08125(new_n10473, new_n10474);
not_8  g08126(n5882, new_n10475);
xnor_4 g08127(new_n10429, new_n10422, new_n10476);
nand_5 g08128(new_n10476, new_n10475, new_n10477);
not_8  g08129(new_n10477, new_n10478);
xnor_4 g08130(new_n10427, new_n10425, new_n10479);
not_8  g08131(new_n10479, new_n10480);
nor_5  g08132(new_n10480, n11775, new_n10481);
not_8  g08133(n27134, new_n10482);
xnor_4 g08134(n22201, n4588, new_n10483);
nor_5  g08135(new_n10483, new_n10482, new_n10484_1);
not_8  g08136(n11775, new_n10485);
xnor_4 g08137(new_n10479, new_n10485, new_n10486);
nor_5  g08138(new_n10486, new_n10484_1, new_n10487);
nor_5  g08139(new_n10487, new_n10481, new_n10488);
xnor_4 g08140(new_n10476, new_n10475, new_n10489_1);
nor_5  g08141(new_n10489_1, new_n10488, new_n10490);
nor_5  g08142(new_n10490, new_n10478, new_n10491);
nor_5  g08143(new_n10491, new_n10474, new_n10492);
nor_5  g08144(new_n10492, new_n10472, new_n10493);
not_8  g08145(new_n10493, new_n10494);
nand_5 g08146(new_n10494, new_n10468, new_n10495);
nand_5 g08147(new_n10495, new_n10467, new_n10496);
nand_5 g08148(new_n10496, new_n10464, new_n10497);
nand_5 g08149(new_n10497, new_n10463, new_n10498);
nand_5 g08150(new_n10498, new_n10460, new_n10499);
nand_5 g08151(new_n10499, new_n10459, new_n10500);
nand_5 g08152(new_n10500, new_n10456, new_n10501);
nand_5 g08153(new_n10501, new_n10455, new_n10502);
nand_5 g08154(new_n10502, new_n10452, new_n10503);
nand_5 g08155(new_n10503, new_n10451, new_n10504);
nand_5 g08156(new_n10504, new_n10447, new_n10505);
nand_5 g08157(new_n10505, new_n10446, new_n10506);
or_5   g08158(n22764, n1536, new_n10507);
nand_5 g08159(new_n10444, new_n10403, new_n10508);
nand_5 g08160(new_n10508, new_n10507, new_n10509);
nor_5  g08161(new_n10509, new_n10506, new_n10510);
or_5   g08162(n23493, n8405, new_n10511);
or_5   g08163(n22359, n10275, new_n10512);
or_5   g08164(n15146, n5532, new_n10513);
or_5   g08165(n11579, n3962, new_n10514_1);
or_5   g08166(n23513, n21, new_n10515);
xnor_4 g08167(n23513, n21, new_n10516);
not_8  g08168(new_n10516, new_n10517);
not_8  g08169(n6427, new_n10518);
nand_5 g08170(new_n10518, new_n8436, new_n10519);
nand_5 g08171(n6427, n1682, new_n10520);
not_8  g08172(n6590, new_n10521);
not_8  g08173(n7963, new_n10522);
nand_5 g08174(new_n10522, new_n10521, new_n10523);
not_8  g08175(n10017, new_n10524);
not_8  g08176(n20349, new_n10525_1);
nand_5 g08177(new_n10525_1, new_n10524, new_n10526);
nand_5 g08178(n15936, n3618, new_n10527);
nand_5 g08179(n20349, n10017, new_n10528);
nand_5 g08180(new_n10528, new_n10527, new_n10529);
nand_5 g08181(new_n10529, new_n10526, new_n10530);
nand_5 g08182(n7963, n6590, new_n10531);
nand_5 g08183(new_n10531, new_n10530, new_n10532);
nand_5 g08184(new_n10532, new_n10523, new_n10533);
nand_5 g08185(new_n10533, new_n10520, new_n10534);
nand_5 g08186(new_n10534, new_n10519, new_n10535);
nand_5 g08187(new_n10535, new_n10517, new_n10536);
nand_5 g08188(new_n10536, new_n10515, new_n10537);
xnor_4 g08189(n11579, n3962, new_n10538);
not_8  g08190(new_n10538, new_n10539);
nand_5 g08191(new_n10539, new_n10537, new_n10540_1);
nand_5 g08192(new_n10540_1, new_n10514_1, new_n10541);
xnor_4 g08193(n15146, n5532, new_n10542);
not_8  g08194(new_n10542, new_n10543);
nand_5 g08195(new_n10543, new_n10541, new_n10544);
nand_5 g08196(new_n10544, new_n10513, new_n10545);
xnor_4 g08197(n22359, n10275, new_n10546);
not_8  g08198(new_n10546, new_n10547);
nand_5 g08199(new_n10547, new_n10545, new_n10548);
nand_5 g08200(new_n10548, new_n10512, new_n10549);
xnor_4 g08201(n23493, n8405, new_n10550);
not_8  g08202(new_n10550, new_n10551);
nand_5 g08203(new_n10551, new_n10549, new_n10552);
nand_5 g08204(new_n10552, new_n10511, new_n10553);
xnor_4 g08205(n14826, n13549, new_n10554);
xnor_4 g08206(new_n10554, new_n10553, new_n10555);
nand_5 g08207(new_n10555, new_n4667, new_n10556);
xnor_4 g08208(new_n10555, n18105, new_n10557);
xnor_4 g08209(new_n10550, new_n10549, new_n10558);
nand_5 g08210(new_n10558, new_n4647, new_n10559);
xnor_4 g08211(new_n10558, n24196, new_n10560);
not_8  g08212(n16376, new_n10561_1);
xnor_4 g08213(new_n10546, new_n10545, new_n10562);
nand_5 g08214(new_n10562, new_n10561_1, new_n10563);
xnor_4 g08215(new_n10562, n16376, new_n10564_1);
xnor_4 g08216(new_n10542, new_n10541, new_n10565);
nand_5 g08217(new_n10565, new_n4648, new_n10566);
xnor_4 g08218(new_n10565, n25381, new_n10567);
xnor_4 g08219(new_n10538, new_n10537, new_n10568);
nand_5 g08220(new_n10568, new_n4687, new_n10569);
xnor_4 g08221(new_n10568, n12587, new_n10570);
xnor_4 g08222(new_n10535, new_n10516, new_n10571);
nand_5 g08223(new_n10571, new_n4649, new_n10572);
xnor_4 g08224(new_n10571, n268, new_n10573);
xnor_4 g08225(n6427, new_n8436, new_n10574);
not_8  g08226(new_n10574, new_n10575);
xnor_4 g08227(new_n10575, new_n10533, new_n10576);
nand_5 g08228(new_n10576, new_n4696, new_n10577_1);
xnor_4 g08229(new_n10576, n24879, new_n10578);
xnor_4 g08230(n7963, n6590, new_n10579);
xnor_4 g08231(new_n10579, new_n10530, new_n10580);
nand_5 g08232(new_n10580, new_n4650, new_n10581);
xnor_4 g08233(n20349, n10017, new_n10582);
not_8  g08234(new_n10582, new_n10583);
xnor_4 g08235(new_n10583, new_n10527, new_n10584);
not_8  g08236(new_n10584, new_n10585);
nand_5 g08237(new_n10585, new_n8549, new_n10586);
xnor_4 g08238(n15936, n3618, new_n10587);
nor_5  g08239(new_n10587, new_n4704, new_n10588_1);
not_8  g08240(new_n10588_1, new_n10589);
xnor_4 g08241(new_n10584, new_n8549, new_n10590);
nand_5 g08242(new_n10590, new_n10589, new_n10591);
nand_5 g08243(new_n10591, new_n10586, new_n10592);
xnor_4 g08244(new_n10580, n6785, new_n10593_1);
nand_5 g08245(new_n10593_1, new_n10592, new_n10594);
nand_5 g08246(new_n10594, new_n10581, new_n10595_1);
nand_5 g08247(new_n10595_1, new_n10578, new_n10596);
nand_5 g08248(new_n10596, new_n10577_1, new_n10597);
nand_5 g08249(new_n10597, new_n10573, new_n10598);
nand_5 g08250(new_n10598, new_n10572, new_n10599);
nand_5 g08251(new_n10599, new_n10570, new_n10600);
nand_5 g08252(new_n10600, new_n10569, new_n10601);
nand_5 g08253(new_n10601, new_n10567, new_n10602);
nand_5 g08254(new_n10602, new_n10566, new_n10603);
nand_5 g08255(new_n10603, new_n10564_1, new_n10604);
nand_5 g08256(new_n10604, new_n10563, new_n10605);
nand_5 g08257(new_n10605, new_n10560, new_n10606);
nand_5 g08258(new_n10606, new_n10559, new_n10607);
nand_5 g08259(new_n10607, new_n10557, new_n10608);
nand_5 g08260(new_n10608, new_n10556, new_n10609);
not_8  g08261(new_n10554, new_n10610);
nand_5 g08262(new_n10610, new_n10553, new_n10611_1);
or_5   g08263(n14826, n13549, new_n10612);
nand_5 g08264(new_n10612, new_n10611_1, new_n10613);
nor_5  g08265(new_n10613, new_n10609, new_n10614_1);
xnor_4 g08266(new_n10614_1, new_n10510, new_n10615);
xnor_4 g08267(new_n10509, new_n10506, new_n10616);
xnor_4 g08268(new_n10613, new_n10609, new_n10617_1);
not_8  g08269(new_n10617_1, new_n10618);
nand_5 g08270(new_n10618, new_n10616, new_n10619);
xnor_4 g08271(new_n10617_1, new_n10616, new_n10620);
xnor_4 g08272(new_n10504, new_n10447, new_n10621);
not_8  g08273(new_n10621, new_n10622);
xnor_4 g08274(new_n10607, new_n10557, new_n10623);
nand_5 g08275(new_n10623, new_n10622, new_n10624);
xnor_4 g08276(new_n10623, new_n10621, new_n10625);
xnor_4 g08277(new_n10502, new_n10452, new_n10626);
not_8  g08278(new_n10626, new_n10627);
xnor_4 g08279(new_n10605, new_n10560, new_n10628_1);
nand_5 g08280(new_n10628_1, new_n10627, new_n10629);
xnor_4 g08281(new_n10628_1, new_n10626, new_n10630);
xnor_4 g08282(new_n10500, new_n10456, new_n10631);
not_8  g08283(new_n10631, new_n10632);
xnor_4 g08284(new_n10603, new_n10564_1, new_n10633);
nand_5 g08285(new_n10633, new_n10632, new_n10634);
xnor_4 g08286(new_n10633, new_n10631, new_n10635);
xnor_4 g08287(new_n10498, new_n10460, new_n10636);
not_8  g08288(new_n10636, new_n10637);
xnor_4 g08289(new_n10601, new_n10567, new_n10638);
nand_5 g08290(new_n10638, new_n10637, new_n10639);
xnor_4 g08291(new_n10638, new_n10636, new_n10640);
not_8  g08292(new_n10464, new_n10641);
xnor_4 g08293(new_n10496, new_n10641, new_n10642);
xnor_4 g08294(new_n10599, new_n10570, new_n10643);
nand_5 g08295(new_n10643, new_n10642, new_n10644);
xnor_4 g08296(new_n10496, new_n10464, new_n10645);
xnor_4 g08297(new_n10643, new_n10645, new_n10646);
xnor_4 g08298(new_n10493, new_n10468, new_n10647_1);
xnor_4 g08299(new_n10597, new_n10573, new_n10648);
nand_5 g08300(new_n10648, new_n10647_1, new_n10649);
xnor_4 g08301(new_n10648, new_n10647_1, new_n10650_1);
not_8  g08302(new_n10650_1, new_n10651);
xnor_4 g08303(new_n10491, new_n10473, new_n10652);
not_8  g08304(new_n10652, new_n10653_1);
xnor_4 g08305(new_n10595_1, new_n10578, new_n10654);
not_8  g08306(new_n10654, new_n10655);
nor_5  g08307(new_n10655, new_n10653_1, new_n10656);
xnor_4 g08308(new_n10654, new_n10653_1, new_n10657);
not_8  g08309(new_n10657, new_n10658);
xnor_4 g08310(new_n10489_1, new_n10488, new_n10659);
xnor_4 g08311(new_n10593_1, new_n10592, new_n10660);
not_8  g08312(new_n10660, new_n10661);
nor_5  g08313(new_n10661, new_n10659, new_n10662);
xnor_4 g08314(new_n10660, new_n10659, new_n10663);
not_8  g08315(new_n10663, new_n10664);
xnor_4 g08316(new_n10486, new_n10484_1, new_n10665);
xnor_4 g08317(new_n10590, new_n10588_1, new_n10666);
nor_5  g08318(new_n10666, new_n10665, new_n10667);
xnor_4 g08319(new_n10483, n27134, new_n10668);
xnor_4 g08320(new_n10587, n22843, new_n10669);
not_8  g08321(new_n10669, new_n10670);
nor_5  g08322(new_n10670, new_n10668, new_n10671);
not_8  g08323(new_n10671, new_n10672);
not_8  g08324(new_n10666, new_n10673);
xnor_4 g08325(new_n10673, new_n10665, new_n10674);
not_8  g08326(new_n10674, new_n10675);
nor_5  g08327(new_n10675, new_n10672, new_n10676);
nor_5  g08328(new_n10676, new_n10667, new_n10677);
nor_5  g08329(new_n10677, new_n10664, new_n10678);
nor_5  g08330(new_n10678, new_n10662, new_n10679);
nor_5  g08331(new_n10679, new_n10658, new_n10680);
nor_5  g08332(new_n10680, new_n10656, new_n10681);
not_8  g08333(new_n10681, new_n10682);
nand_5 g08334(new_n10682, new_n10651, new_n10683);
nand_5 g08335(new_n10683, new_n10649, new_n10684);
nand_5 g08336(new_n10684, new_n10646, new_n10685);
nand_5 g08337(new_n10685, new_n10644, new_n10686);
nand_5 g08338(new_n10686, new_n10640, new_n10687);
nand_5 g08339(new_n10687, new_n10639, new_n10688);
nand_5 g08340(new_n10688, new_n10635, new_n10689);
nand_5 g08341(new_n10689, new_n10634, new_n10690);
nand_5 g08342(new_n10690, new_n10630, new_n10691);
nand_5 g08343(new_n10691, new_n10629, new_n10692_1);
nand_5 g08344(new_n10692_1, new_n10625, new_n10693);
nand_5 g08345(new_n10693, new_n10624, new_n10694_1);
nand_5 g08346(new_n10694_1, new_n10620, new_n10695);
nand_5 g08347(new_n10695, new_n10619, new_n10696);
xnor_4 g08348(new_n10696, new_n10615, n1302);
or_5   g08349(n13951, new_n9274, new_n10698);
xnor_4 g08350(n13951, n12507, new_n10699);
or_5   g08351(n22793, new_n9341, new_n10700);
xnor_4 g08352(n22793, n15077, new_n10701_1);
or_5   g08353(n8439, new_n9349, new_n10702);
xnor_4 g08354(n8439, n3710, new_n10703);
or_5   g08355(new_n9291, n25523, new_n10704);
xnor_4 g08356(n26318, n25523, new_n10705);
or_5   g08357(new_n9296, n5579, new_n10706);
xnor_4 g08358(n26054, n5579, new_n10707);
nor_5  g08359(n23430, new_n9301, new_n10708);
xnor_4 g08360(n23430, n19081, new_n10709);
nor_5  g08361(n10411, new_n9306, new_n10710_1);
not_8  g08362(new_n10710_1, new_n10711);
xnor_4 g08363(n10411, n8309, new_n10712_1);
nor_5  g08364(n19144, new_n2705, new_n10713);
nor_5  g08365(new_n9310, n16971, new_n10714);
nor_5  g08366(n12593, new_n2801, new_n10715);
nor_5  g08367(new_n9315, n11503, new_n10716);
not_8  g08368(n18151, new_n10717);
nor_5  g08369(new_n10717, n13714, new_n10718);
not_8  g08370(new_n10718, new_n10719);
nor_5  g08371(new_n10719, new_n10716, new_n10720);
nor_5  g08372(new_n10720, new_n10715, new_n10721);
nor_5  g08373(new_n10721, new_n10714, new_n10722);
nor_5  g08374(new_n10722, new_n10713, new_n10723);
nand_5 g08375(new_n10723, new_n10712_1, new_n10724);
nand_5 g08376(new_n10724, new_n10711, new_n10725);
and_5  g08377(new_n10725, new_n10709, new_n10726);
nor_5  g08378(new_n10726, new_n10708, new_n10727);
not_8  g08379(new_n10727, new_n10728);
nand_5 g08380(new_n10728, new_n10707, new_n10729);
nand_5 g08381(new_n10729, new_n10706, new_n10730);
nand_5 g08382(new_n10730, new_n10705, new_n10731);
nand_5 g08383(new_n10731, new_n10704, new_n10732);
nand_5 g08384(new_n10732, new_n10703, new_n10733);
nand_5 g08385(new_n10733, new_n10702, new_n10734);
nand_5 g08386(new_n10734, new_n10701_1, new_n10735);
nand_5 g08387(new_n10735, new_n10700, new_n10736);
nand_5 g08388(new_n10736, new_n10699, new_n10737);
nand_5 g08389(new_n10737, new_n10698, new_n10738);
not_8  g08390(new_n10738, new_n10739_1);
or_5   g08391(n12650, n11220, new_n10740);
not_8  g08392(n11220, new_n10741);
xnor_4 g08393(n12650, new_n10741, new_n10742);
or_5   g08394(n22379, n10201, new_n10743);
xnor_4 g08395(n22379, new_n5835, new_n10744);
or_5   g08396(n10593, n1662, new_n10745);
xnor_4 g08397(n10593, new_n2900, new_n10746);
nor_5  g08398(n18290, n12875, new_n10747);
not_8  g08399(new_n9841, new_n10748);
nor_5  g08400(new_n9867_1, new_n10748, new_n10749);
nor_5  g08401(new_n10749, new_n10747, new_n10750);
not_8  g08402(new_n10750, new_n10751);
nand_5 g08403(new_n10751, new_n10746, new_n10752);
nand_5 g08404(new_n10752, new_n10745, new_n10753);
nand_5 g08405(new_n10753, new_n10744, new_n10754);
nand_5 g08406(new_n10754, new_n10743, new_n10755);
nand_5 g08407(new_n10755, new_n10742, new_n10756_1);
nand_5 g08408(new_n10756_1, new_n10740, new_n10757);
or_5   g08409(n22270, n2944, new_n10758);
nand_5 g08410(new_n2765, new_n2718, new_n10759);
nand_5 g08411(new_n10759, new_n10758, new_n10760);
xnor_4 g08412(new_n10760, new_n10757, new_n10761);
not_8  g08413(new_n10761, new_n10762);
xnor_4 g08414(new_n10755, new_n10742, new_n10763_1);
not_8  g08415(new_n10763_1, new_n10764);
nor_5  g08416(new_n10764, new_n2766, new_n10765);
not_8  g08417(new_n2771, new_n10766);
xnor_4 g08418(new_n10753, new_n10744, new_n10767);
nor_5  g08419(new_n10767, new_n10766, new_n10768);
xnor_4 g08420(new_n10767, new_n2771, new_n10769);
not_8  g08421(new_n10769, new_n10770);
xnor_4 g08422(new_n10750, new_n10746, new_n10771);
not_8  g08423(new_n10771, new_n10772);
nor_5  g08424(new_n10772, new_n2775, new_n10773);
xnor_4 g08425(new_n10771, new_n2775, new_n10774);
not_8  g08426(new_n10774, new_n10775_1);
not_8  g08427(new_n9868, new_n10776);
nor_5  g08428(new_n10776, new_n2780, new_n10777);
not_8  g08429(new_n9871, new_n10778);
nor_5  g08430(new_n10778, new_n2785, new_n10779);
xnor_4 g08431(new_n9871, new_n2785, new_n10780_1);
not_8  g08432(new_n10780_1, new_n10781);
not_8  g08433(new_n2790, new_n10782);
nor_5  g08434(new_n9874, new_n10782, new_n10783);
not_8  g08435(new_n10783, new_n10784);
nor_5  g08436(new_n9878, new_n2794, new_n10785);
xnor_4 g08437(new_n9877, new_n2794, new_n10786);
not_8  g08438(new_n10786, new_n10787);
nor_5  g08439(new_n9883, new_n2798, new_n10788);
xnor_4 g08440(new_n9882, new_n2798, new_n10789);
not_8  g08441(new_n10789, new_n10790);
not_8  g08442(new_n9886, new_n10791);
nor_5  g08443(new_n10791, new_n2803, new_n10792_1);
nor_5  g08444(new_n9890_1, new_n2807, new_n10793);
xnor_4 g08445(new_n9886, new_n2803, new_n10794);
nand_5 g08446(new_n10794, new_n10793, new_n10795);
not_8  g08447(new_n10795, new_n10796);
nor_5  g08448(new_n10796, new_n10792_1, new_n10797);
nor_5  g08449(new_n10797, new_n10790, new_n10798);
nor_5  g08450(new_n10798, new_n10788, new_n10799);
nor_5  g08451(new_n10799, new_n10787, new_n10800);
nor_5  g08452(new_n10800, new_n10785, new_n10801);
xnor_4 g08453(new_n9874, new_n2790, new_n10802);
nand_5 g08454(new_n10802, new_n10801, new_n10803);
nand_5 g08455(new_n10803, new_n10784, new_n10804);
nor_5  g08456(new_n10804, new_n10781, new_n10805);
nor_5  g08457(new_n10805, new_n10779, new_n10806);
xnor_4 g08458(new_n9868, new_n2780, new_n10807);
not_8  g08459(new_n10807, new_n10808);
nor_5  g08460(new_n10808, new_n10806, new_n10809);
nor_5  g08461(new_n10809, new_n10777, new_n10810);
nor_5  g08462(new_n10810, new_n10775_1, new_n10811);
nor_5  g08463(new_n10811, new_n10773, new_n10812);
nor_5  g08464(new_n10812, new_n10770, new_n10813);
nor_5  g08465(new_n10813, new_n10768, new_n10814);
not_8  g08466(new_n10814, new_n10815);
xnor_4 g08467(new_n10763_1, new_n2766, new_n10816);
not_8  g08468(new_n10816, new_n10817_1);
nor_5  g08469(new_n10817_1, new_n10815, new_n10818);
nor_5  g08470(new_n10818, new_n10765, new_n10819);
xnor_4 g08471(new_n10819, new_n10762, new_n10820);
xnor_4 g08472(new_n10820, new_n10739_1, new_n10821);
xnor_4 g08473(new_n10736, new_n10699, new_n10822);
xnor_4 g08474(new_n10817_1, new_n10814, new_n10823);
not_8  g08475(new_n10823, new_n10824);
nand_5 g08476(new_n10824, new_n10822, new_n10825);
xnor_4 g08477(new_n10823, new_n10822, new_n10826);
xnor_4 g08478(new_n10734, new_n10701_1, new_n10827);
xnor_4 g08479(new_n10812, new_n10769, new_n10828);
nand_5 g08480(new_n10828, new_n10827, new_n10829);
not_8  g08481(new_n10828, new_n10830);
xnor_4 g08482(new_n10830, new_n10827, new_n10831);
xnor_4 g08483(new_n10732, new_n10703, new_n10832);
xnor_4 g08484(new_n10810, new_n10774, new_n10833);
nand_5 g08485(new_n10833, new_n10832, new_n10834_1);
not_8  g08486(new_n10833, new_n10835);
xnor_4 g08487(new_n10835, new_n10832, new_n10836);
xnor_4 g08488(new_n10730, new_n10705, new_n10837);
xnor_4 g08489(new_n10807, new_n10806, new_n10838);
nand_5 g08490(new_n10838, new_n10837, new_n10839);
not_8  g08491(new_n10838, new_n10840);
xnor_4 g08492(new_n10840, new_n10837, new_n10841);
xnor_4 g08493(new_n10728, new_n10707, new_n10842);
xnor_4 g08494(new_n10804, new_n10780_1, new_n10843);
nand_5 g08495(new_n10843, new_n10842, new_n10844);
not_8  g08496(new_n10709, new_n10845);
xnor_4 g08497(new_n10725, new_n10845, new_n10846);
not_8  g08498(new_n10846, new_n10847);
xnor_4 g08499(new_n10802, new_n10801, new_n10848);
nand_5 g08500(new_n10848, new_n10847, new_n10849);
xnor_4 g08501(new_n10848, new_n10846, new_n10850);
xnor_4 g08502(new_n10799, new_n10786, new_n10851_1);
not_8  g08503(new_n10851_1, new_n10852);
xnor_4 g08504(new_n10723, new_n10712_1, new_n10853);
not_8  g08505(new_n10853, new_n10854);
nor_5  g08506(new_n10854, new_n10852, new_n10855);
not_8  g08507(new_n10855, new_n10856);
xnor_4 g08508(new_n10797, new_n10789, new_n10857);
not_8  g08509(new_n10857, new_n10858);
xnor_4 g08510(n19144, n16971, new_n10859);
xnor_4 g08511(new_n10859, new_n10721, new_n10860);
not_8  g08512(new_n10860, new_n10861);
nor_5  g08513(new_n10861, new_n10858, new_n10862);
not_8  g08514(new_n10862, new_n10863);
xnor_4 g08515(new_n10861, new_n10857, new_n10864);
xnor_4 g08516(new_n9890_1, new_n2806, new_n10865);
xnor_4 g08517(n18151, n13714, new_n10866);
nor_5  g08518(new_n10866, new_n10865, new_n10867);
xnor_4 g08519(n12593, n11503, new_n10868);
xnor_4 g08520(new_n10868, new_n10719, new_n10869);
not_8  g08521(new_n10869, new_n10870);
and_5  g08522(new_n10870, new_n10867, new_n10871);
xnor_4 g08523(new_n10794, new_n10793, new_n10872);
xnor_4 g08524(new_n10869, new_n10867, new_n10873);
and_5  g08525(new_n10873, new_n10872, new_n10874_1);
nor_5  g08526(new_n10874_1, new_n10871, new_n10875);
nand_5 g08527(new_n10875, new_n10864, new_n10876);
nand_5 g08528(new_n10876, new_n10863, new_n10877);
xnor_4 g08529(new_n10854, new_n10851_1, new_n10878);
nand_5 g08530(new_n10878, new_n10877, new_n10879);
nand_5 g08531(new_n10879, new_n10856, new_n10880);
nand_5 g08532(new_n10880, new_n10850, new_n10881);
nand_5 g08533(new_n10881, new_n10849, new_n10882);
not_8  g08534(new_n10843, new_n10883);
xnor_4 g08535(new_n10883, new_n10842, new_n10884);
nand_5 g08536(new_n10884, new_n10882, new_n10885);
nand_5 g08537(new_n10885, new_n10844, new_n10886);
nand_5 g08538(new_n10886, new_n10841, new_n10887);
nand_5 g08539(new_n10887, new_n10839, new_n10888);
nand_5 g08540(new_n10888, new_n10836, new_n10889);
nand_5 g08541(new_n10889, new_n10834_1, new_n10890);
nand_5 g08542(new_n10890, new_n10831, new_n10891);
nand_5 g08543(new_n10891, new_n10829, new_n10892);
nand_5 g08544(new_n10892, new_n10826, new_n10893);
nand_5 g08545(new_n10893, new_n10825, new_n10894);
xnor_4 g08546(new_n10894, new_n10821, n1332);
not_8  g08547(n14692, new_n10896);
nand_5 g08548(new_n5834_1, new_n10896, new_n10897);
xnor_4 g08549(new_n5834_1, n14692, new_n10898);
not_8  g08550(n4100, new_n10899);
nand_5 g08551(new_n5914, new_n10899, new_n10900);
xnor_4 g08552(new_n5914, n4100, new_n10901);
not_8  g08553(n21957, new_n10902);
nand_5 g08554(new_n5919, new_n10902, new_n10903);
xnor_4 g08555(new_n5919, n21957, new_n10904);
not_8  g08556(n15761, new_n10905);
nand_5 g08557(new_n5924, new_n10905, new_n10906);
xnor_4 g08558(new_n5924, n15761, new_n10907);
not_8  g08559(n11201, new_n10908);
nand_5 g08560(new_n5930, new_n10908, new_n10909);
xnor_4 g08561(new_n5929, new_n10908, new_n10910);
not_8  g08562(n18690, new_n10911);
nand_5 g08563(new_n5935, new_n10911, new_n10912);
xnor_4 g08564(new_n5935, n18690, new_n10913);
not_8  g08565(n12153, new_n10914);
nand_5 g08566(new_n5945, new_n10914, new_n10915);
xnor_4 g08567(new_n5941, new_n10914, new_n10916);
not_8  g08568(n13044, new_n10917);
nor_5  g08569(new_n5949, new_n10917, new_n10918);
nor_5  g08570(new_n5950, n13044, new_n10919);
nor_5  g08571(new_n5957, n18745, new_n10920);
not_8  g08572(new_n10920, new_n10921);
not_8  g08573(new_n6121, new_n10922);
nand_5 g08574(new_n6123, new_n10922, new_n10923);
nand_5 g08575(new_n10923, new_n10921, new_n10924_1);
nor_5  g08576(new_n10924_1, new_n10919, new_n10925);
nor_5  g08577(new_n10925, new_n10918, new_n10926);
nand_5 g08578(new_n10926, new_n10916, new_n10927);
nand_5 g08579(new_n10927, new_n10915, new_n10928);
nand_5 g08580(new_n10928, new_n10913, new_n10929);
nand_5 g08581(new_n10929, new_n10912, new_n10930);
nand_5 g08582(new_n10930, new_n10910, new_n10931);
nand_5 g08583(new_n10931, new_n10909, new_n10932);
nand_5 g08584(new_n10932, new_n10907, new_n10933);
nand_5 g08585(new_n10933, new_n10906, new_n10934);
nand_5 g08586(new_n10934, new_n10904, new_n10935);
nand_5 g08587(new_n10935, new_n10903, new_n10936);
nand_5 g08588(new_n10936, new_n10901, new_n10937);
nand_5 g08589(new_n10937, new_n10900, new_n10938);
nand_5 g08590(new_n10938, new_n10898, new_n10939);
nand_5 g08591(new_n10939, new_n10897, new_n10940);
nor_5  g08592(new_n10940, new_n5832, new_n10941);
nand_5 g08593(new_n6131, new_n4199, new_n10942);
nor_5  g08594(new_n10942, n10405, new_n10943_1);
nand_5 g08595(new_n10943_1, new_n4185, new_n10944);
nor_5  g08596(new_n10944, n20151, new_n10945);
nand_5 g08597(new_n10945, new_n6551, new_n10946);
nor_5  g08598(new_n10946, n27037, new_n10947);
nand_5 g08599(new_n10947, new_n6542_1, new_n10948);
or_5   g08600(new_n10948, n8614, new_n10949);
not_8  g08601(n25629, new_n10950);
not_8  g08602(n23039, new_n10951);
nor_5  g08603(n25926, n7657, new_n10952);
nand_5 g08604(new_n10952, new_n4144, new_n10953);
nor_5  g08605(new_n10953, n5451, new_n10954);
nand_5 g08606(new_n10954, new_n4164, new_n10955);
nor_5  g08607(new_n10955, n13677, new_n10956);
nand_5 g08608(new_n10956, new_n10951, new_n10957);
nor_5  g08609(new_n10957, n7692, new_n10958);
nand_5 g08610(new_n10958, new_n10950, new_n10959);
nor_5  g08611(new_n10959, n15766, new_n10960);
not_8  g08612(new_n10960, new_n10961_1);
not_8  g08613(n15766, new_n10962);
xnor_4 g08614(new_n10959, new_n10962, new_n10963);
or_5   g08615(new_n10963, n23895, new_n10964);
xnor_4 g08616(new_n10958, n25629, new_n10965);
not_8  g08617(new_n10965, new_n10966);
nand_5 g08618(new_n10966, new_n5740, new_n10967);
xnor_4 g08619(new_n10965, new_n5740, new_n10968);
xnor_4 g08620(new_n10957, new_n6648, new_n10969);
not_8  g08621(new_n10969, new_n10970);
nand_5 g08622(new_n10970, new_n5743, new_n10971);
xnor_4 g08623(new_n10969, new_n5743, new_n10972);
xnor_4 g08624(new_n10956, n23039, new_n10973);
nor_5  g08625(new_n10973, n23200, new_n10974);
not_8  g08626(new_n10974, new_n10975);
xnor_4 g08627(new_n10973, new_n5746, new_n10976);
xnor_4 g08628(new_n10955, new_n4095, new_n10977);
nor_5  g08629(new_n10977, n17959, new_n10978);
not_8  g08630(new_n10978, new_n10979);
xnor_4 g08631(new_n10954, n18926, new_n10980);
nor_5  g08632(new_n10980, n7566, new_n10981);
xnor_4 g08633(new_n10980, new_n5752_1, new_n10982);
not_8  g08634(new_n10982, new_n10983);
xnor_4 g08635(new_n10953, new_n4138, new_n10984);
not_8  g08636(new_n10984, new_n10985);
nor_5  g08637(new_n10985, new_n5755, new_n10986);
nor_5  g08638(new_n10984, n7731, new_n10987);
xnor_4 g08639(new_n10952, n5330, new_n10988);
not_8  g08640(new_n10988, new_n10989);
nor_5  g08641(new_n10989, new_n5760, new_n10990);
xnor_4 g08642(new_n10988, new_n5760, new_n10991);
not_8  g08643(new_n10991, new_n10992);
nor_5  g08644(new_n6126, new_n5763, new_n10993);
nor_5  g08645(new_n6127, new_n6125, new_n10994);
nor_5  g08646(new_n10994, new_n10993, new_n10995);
nor_5  g08647(new_n10995, new_n10992, new_n10996);
nor_5  g08648(new_n10996, new_n10990, new_n10997);
nor_5  g08649(new_n10997, new_n10987, new_n10998);
nor_5  g08650(new_n10998, new_n10986, new_n10999);
not_8  g08651(new_n10999, new_n11000);
nor_5  g08652(new_n11000, new_n10983, new_n11001);
nor_5  g08653(new_n11001, new_n10981, new_n11002);
not_8  g08654(new_n11002, new_n11003);
xnor_4 g08655(new_n10977, new_n5749, new_n11004);
nand_5 g08656(new_n11004, new_n11003, new_n11005_1);
nand_5 g08657(new_n11005_1, new_n10979, new_n11006);
nand_5 g08658(new_n11006, new_n10976, new_n11007);
nand_5 g08659(new_n11007, new_n10975, new_n11008);
nand_5 g08660(new_n11008, new_n10972, new_n11009);
nand_5 g08661(new_n11009, new_n10971, new_n11010);
nand_5 g08662(new_n11010, new_n10968, new_n11011_1);
nand_5 g08663(new_n11011_1, new_n10967, new_n11012);
nand_5 g08664(new_n10963, n23895, new_n11013);
nand_5 g08665(new_n11013, new_n11012, new_n11014);
nand_5 g08666(new_n11014, new_n10964, new_n11015);
nand_5 g08667(new_n11015, new_n10961_1, new_n11016);
nand_5 g08668(new_n11016, new_n10949, new_n11017);
xnor_4 g08669(new_n10948, new_n6526, new_n11018);
not_8  g08670(new_n11018, new_n11019);
xnor_4 g08671(new_n10963, new_n5737, new_n11020);
not_8  g08672(new_n11020, new_n11021);
xnor_4 g08673(new_n11021, new_n11012, new_n11022);
nor_5  g08674(new_n11022, new_n11019, new_n11023_1);
xnor_4 g08675(new_n10947, n15182, new_n11024);
not_8  g08676(new_n11024, new_n11025_1);
xnor_4 g08677(new_n11010, new_n10968, new_n11026);
not_8  g08678(new_n11026, new_n11027);
nand_5 g08679(new_n11027, new_n11025_1, new_n11028);
xnor_4 g08680(new_n11026, new_n11025_1, new_n11029);
xnor_4 g08681(new_n10946, n27037, new_n11030);
xnor_4 g08682(new_n11008, new_n10972, new_n11031);
not_8  g08683(new_n11031, new_n11032);
nand_5 g08684(new_n11032, new_n11030, new_n11033);
xnor_4 g08685(new_n11031, new_n11030, new_n11034);
xnor_4 g08686(new_n10945, n8964, new_n11035);
not_8  g08687(new_n11035, new_n11036);
not_8  g08688(new_n10976, new_n11037);
xnor_4 g08689(new_n11006, new_n11037, new_n11038);
nand_5 g08690(new_n11038, new_n11036, new_n11039);
xnor_4 g08691(new_n11038, new_n11035, new_n11040);
xnor_4 g08692(new_n10944, new_n6557, new_n11041);
not_8  g08693(new_n11041, new_n11042);
xnor_4 g08694(new_n11004, new_n11002, new_n11043);
nand_5 g08695(new_n11043, new_n11042, new_n11044_1);
xnor_4 g08696(new_n11043, new_n11041, new_n11045);
xnor_4 g08697(new_n10943_1, n7693, new_n11046);
not_8  g08698(new_n11046, new_n11047);
xnor_4 g08699(new_n10999, new_n10982, new_n11048);
not_8  g08700(new_n11048, new_n11049);
nand_5 g08701(new_n11049, new_n11047, new_n11050);
xnor_4 g08702(new_n11048, new_n11046, new_n11051);
not_8  g08703(new_n11051, new_n11052);
xnor_4 g08704(new_n10942, new_n4189, new_n11053);
not_8  g08705(new_n11053, new_n11054);
xnor_4 g08706(new_n10984, new_n5755, new_n11055);
xnor_4 g08707(new_n11055, new_n10997, new_n11056_1);
not_8  g08708(new_n11056_1, new_n11057);
nand_5 g08709(new_n11057, new_n11054, new_n11058);
xnor_4 g08710(new_n11056_1, new_n11054, new_n11059);
xnor_4 g08711(new_n10995, new_n10992, new_n11060);
xnor_4 g08712(new_n6131, n11302, new_n11061);
not_8  g08713(new_n11061, new_n11062);
nand_5 g08714(new_n11062, new_n11060, new_n11063_1);
xnor_4 g08715(new_n11061, new_n11060, new_n11064);
not_8  g08716(new_n6128, new_n11065);
nor_5  g08717(new_n6138, new_n11065, new_n11066);
nor_5  g08718(new_n11066, new_n6136, new_n11067);
not_8  g08719(new_n11067, new_n11068);
nand_5 g08720(new_n11068, new_n11064, new_n11069);
nand_5 g08721(new_n11069, new_n11063_1, new_n11070);
nand_5 g08722(new_n11070, new_n11059, new_n11071);
nand_5 g08723(new_n11071, new_n11058, new_n11072);
nand_5 g08724(new_n11072, new_n11052, new_n11073);
nand_5 g08725(new_n11073, new_n11050, new_n11074);
nand_5 g08726(new_n11074, new_n11045, new_n11075);
nand_5 g08727(new_n11075, new_n11044_1, new_n11076);
nand_5 g08728(new_n11076, new_n11040, new_n11077);
nand_5 g08729(new_n11077, new_n11039, new_n11078_1);
nand_5 g08730(new_n11078_1, new_n11034, new_n11079);
nand_5 g08731(new_n11079, new_n11033, new_n11080_1);
nand_5 g08732(new_n11080_1, new_n11029, new_n11081);
nand_5 g08733(new_n11081, new_n11028, new_n11082);
xnor_4 g08734(new_n11022, new_n11019, new_n11083);
nor_5  g08735(new_n11083, new_n11082, new_n11084);
nor_5  g08736(new_n11084, new_n11023_1, new_n11085);
not_8  g08737(new_n11085, new_n11086);
nor_5  g08738(new_n11086, new_n11017, new_n11087);
xnor_4 g08739(new_n11087, new_n10941, new_n11088);
xnor_4 g08740(new_n10940, new_n5833_1, new_n11089);
xnor_4 g08741(new_n11016, new_n10949, new_n11090);
xnor_4 g08742(new_n11090, new_n11085, new_n11091);
nor_5  g08743(new_n11091, new_n11089, new_n11092);
not_8  g08744(new_n11089, new_n11093);
xnor_4 g08745(new_n11091, new_n11093, new_n11094_1);
not_8  g08746(new_n11094_1, new_n11095);
xnor_4 g08747(new_n10938, new_n10898, new_n11096);
not_8  g08748(new_n11096, new_n11097);
xnor_4 g08749(new_n11083, new_n11082, new_n11098);
nor_5  g08750(new_n11098, new_n11097, new_n11099);
not_8  g08751(new_n11099, new_n11100);
xnor_4 g08752(new_n11098, new_n11096, new_n11101_1);
not_8  g08753(new_n11029, new_n11102);
xnor_4 g08754(new_n11080_1, new_n11102, new_n11103_1);
xnor_4 g08755(new_n10936, new_n10901, new_n11104);
not_8  g08756(new_n11104, new_n11105);
nor_5  g08757(new_n11105, new_n11103_1, new_n11106);
not_8  g08758(new_n11106, new_n11107);
xnor_4 g08759(new_n11078_1, new_n11034, new_n11108);
xnor_4 g08760(new_n10934, new_n10904, new_n11109);
nor_5  g08761(new_n11109, new_n11108, new_n11110);
not_8  g08762(new_n11109, new_n11111);
xnor_4 g08763(new_n11111, new_n11108, new_n11112);
not_8  g08764(new_n11112, new_n11113);
not_8  g08765(new_n11040, new_n11114);
xnor_4 g08766(new_n11076, new_n11114, new_n11115);
xnor_4 g08767(new_n10932, new_n10907, new_n11116);
not_8  g08768(new_n11116, new_n11117);
nor_5  g08769(new_n11117, new_n11115, new_n11118);
not_8  g08770(new_n11118, new_n11119);
not_8  g08771(new_n11045, new_n11120_1);
xnor_4 g08772(new_n11074, new_n11120_1, new_n11121_1);
xnor_4 g08773(new_n10930, new_n10910, new_n11122);
not_8  g08774(new_n11122, new_n11123);
nand_5 g08775(new_n11123, new_n11121_1, new_n11124);
xnor_4 g08776(new_n11122, new_n11121_1, new_n11125);
xnor_4 g08777(new_n11072, new_n11051, new_n11126);
xnor_4 g08778(new_n10928, new_n10913, new_n11127_1);
not_8  g08779(new_n11127_1, new_n11128);
nor_5  g08780(new_n11128, new_n11126, new_n11129);
xnor_4 g08781(new_n11128, new_n11126, new_n11130);
xnor_4 g08782(new_n11070, new_n11059, new_n11131);
xnor_4 g08783(new_n10926, new_n10916, new_n11132_1);
nor_5  g08784(new_n11132_1, new_n11131, new_n11133);
not_8  g08785(new_n11133, new_n11134_1);
not_8  g08786(new_n11132_1, new_n11135);
xnor_4 g08787(new_n11135, new_n11131, new_n11136);
xnor_4 g08788(new_n11067, new_n11064, new_n11137);
not_8  g08789(new_n11137, new_n11138_1);
not_8  g08790(new_n10924_1, new_n11139);
xnor_4 g08791(new_n5949, n13044, new_n11140);
xnor_4 g08792(new_n11140, new_n11139, new_n11141);
not_8  g08793(new_n11141, new_n11142);
nor_5  g08794(new_n11142, new_n11138_1, new_n11143);
not_8  g08795(new_n11143, new_n11144);
not_8  g08796(new_n6124, new_n11145);
nor_5  g08797(new_n6140, new_n11145, new_n11146);
nor_5  g08798(new_n6142, new_n6119, new_n11147);
nor_5  g08799(new_n11147, new_n11146, new_n11148);
not_8  g08800(new_n11148, new_n11149);
xnor_4 g08801(new_n11142, new_n11137, new_n11150);
nand_5 g08802(new_n11150, new_n11149, new_n11151);
nand_5 g08803(new_n11151, new_n11144, new_n11152);
nand_5 g08804(new_n11152, new_n11136, new_n11153);
nand_5 g08805(new_n11153, new_n11134_1, new_n11154);
nor_5  g08806(new_n11154, new_n11130, new_n11155);
nor_5  g08807(new_n11155, new_n11129, new_n11156);
nand_5 g08808(new_n11156, new_n11125, new_n11157);
nand_5 g08809(new_n11157, new_n11124, new_n11158);
not_8  g08810(new_n11158, new_n11159);
xnor_4 g08811(new_n11116, new_n11115, new_n11160);
nand_5 g08812(new_n11160, new_n11159, new_n11161);
nand_5 g08813(new_n11161, new_n11119, new_n11162);
nor_5  g08814(new_n11162, new_n11113, new_n11163);
nor_5  g08815(new_n11163, new_n11110, new_n11164);
xnor_4 g08816(new_n11104, new_n11103_1, new_n11165);
nand_5 g08817(new_n11165, new_n11164, new_n11166);
nand_5 g08818(new_n11166, new_n11107, new_n11167);
nand_5 g08819(new_n11167, new_n11101_1, new_n11168);
nand_5 g08820(new_n11168, new_n11100, new_n11169);
nor_5  g08821(new_n11169, new_n11095, new_n11170);
nor_5  g08822(new_n11170, new_n11092, new_n11171);
xnor_4 g08823(new_n11171, new_n11088, n1357);
xnor_4 g08824(new_n8471, n25240, new_n11173);
nand_5 g08825(new_n8476, new_n7647_1, new_n11174);
xnor_4 g08826(new_n8476, n10125, new_n11175);
nand_5 g08827(new_n8481, new_n7650, new_n11176);
xnor_4 g08828(new_n8481, n8067, new_n11177);
not_8  g08829(n20923, new_n11178);
nand_5 g08830(new_n8485, new_n11178, new_n11179);
xnor_4 g08831(new_n8485, n20923, new_n11180);
not_8  g08832(new_n8490, new_n11181);
nor_5  g08833(new_n11181, n18157, new_n11182_1);
not_8  g08834(new_n8958, new_n11183);
nor_5  g08835(new_n8969, new_n11183, new_n11184_1);
nor_5  g08836(new_n11184_1, new_n11182_1, new_n11185);
not_8  g08837(new_n11185, new_n11186);
nand_5 g08838(new_n11186, new_n11180, new_n11187);
nand_5 g08839(new_n11187, new_n11179, new_n11188);
nand_5 g08840(new_n11188, new_n11177, new_n11189);
nand_5 g08841(new_n11189, new_n11176, new_n11190);
nand_5 g08842(new_n11190, new_n11175, new_n11191);
nand_5 g08843(new_n11191, new_n11174, new_n11192_1);
xnor_4 g08844(new_n11192_1, new_n11173, new_n11193);
not_8  g08845(n5077, new_n11194);
not_8  g08846(n1099, new_n11195);
xnor_4 g08847(n6381, new_n11195, new_n11196);
nor_5  g08848(n14345, n2113, new_n11197);
not_8  g08849(new_n11197, new_n11198);
not_8  g08850(n2113, new_n11199);
xnor_4 g08851(n14345, new_n11199, new_n11200);
nor_5  g08852(n21134, n11356, new_n11201_1);
not_8  g08853(new_n11201_1, new_n11202);
not_8  g08854(n11356, new_n11203);
xnor_4 g08855(n21134, new_n11203, new_n11204);
nand_5 g08856(n6369, n3164, new_n11205);
not_8  g08857(new_n11205, new_n11206);
nor_5  g08858(n6369, n3164, new_n11207);
nor_5  g08859(n25797, n10611, new_n11208);
not_8  g08860(new_n11208, new_n11209);
not_8  g08861(new_n6945, new_n11210);
nor_5  g08862(new_n6957, new_n11210, new_n11211);
not_8  g08863(new_n11211, new_n11212);
nand_5 g08864(new_n11212, new_n11209, new_n11213);
nor_5  g08865(new_n11213, new_n11207, new_n11214);
nor_5  g08866(new_n11214, new_n11206, new_n11215);
nand_5 g08867(new_n11215, new_n11204, new_n11216);
nand_5 g08868(new_n11216, new_n11202, new_n11217);
nand_5 g08869(new_n11217, new_n11200, new_n11218);
nand_5 g08870(new_n11218, new_n11198, new_n11219);
xnor_4 g08871(new_n11219, new_n11196, new_n11220_1);
xnor_4 g08872(new_n11220_1, new_n11194, new_n11221);
not_8  g08873(n15546, new_n11222);
xnor_4 g08874(new_n11217, new_n11200, new_n11223_1);
not_8  g08875(new_n11223_1, new_n11224);
nor_5  g08876(new_n11224, new_n11222, new_n11225);
xnor_4 g08877(new_n11223_1, new_n11222, new_n11226);
not_8  g08878(new_n11226, new_n11227);
xnor_4 g08879(new_n11215, new_n11204, new_n11228);
nor_5  g08880(new_n11228, n26452, new_n11229);
not_8  g08881(new_n11229, new_n11230);
not_8  g08882(n19905, new_n11231);
xnor_4 g08883(n6369, new_n9683, new_n11232);
xnor_4 g08884(new_n11232, new_n11213, new_n11233);
not_8  g08885(new_n11233, new_n11234_1);
nor_5  g08886(new_n11234_1, new_n11231, new_n11235);
xnor_4 g08887(new_n11233, new_n11231, new_n11236);
not_8  g08888(new_n11236, new_n11237);
nor_5  g08889(new_n6958, new_n4359, new_n11238);
nand_5 g08890(new_n9003_1, new_n8998, new_n11239);
not_8  g08891(new_n11239, new_n11240);
nor_5  g08892(new_n11240, new_n11238, new_n11241);
nor_5  g08893(new_n11241, new_n11237, new_n11242);
nor_5  g08894(new_n11242, new_n11235, new_n11243);
not_8  g08895(n26452, new_n11244);
xnor_4 g08896(new_n11228, new_n11244, new_n11245_1);
nand_5 g08897(new_n11245_1, new_n11243, new_n11246);
nand_5 g08898(new_n11246, new_n11230, new_n11247);
nor_5  g08899(new_n11247, new_n11227, new_n11248);
nor_5  g08900(new_n11248, new_n11225, new_n11249);
xnor_4 g08901(new_n11249, new_n11221, new_n11250);
xnor_4 g08902(new_n11250, new_n11193, new_n11251);
not_8  g08903(new_n11175, new_n11252);
xnor_4 g08904(new_n11190, new_n11252, new_n11253);
xnor_4 g08905(new_n11247, new_n11226, new_n11254);
nand_5 g08906(new_n11254, new_n11253, new_n11255);
not_8  g08907(new_n11254, new_n11256);
xnor_4 g08908(new_n11256, new_n11253, new_n11257);
xnor_4 g08909(new_n11188, new_n11177, new_n11258);
not_8  g08910(new_n11258, new_n11259);
xnor_4 g08911(new_n11245_1, new_n11243, new_n11260);
nand_5 g08912(new_n11260, new_n11259, new_n11261_1);
xnor_4 g08913(new_n11260, new_n11258, new_n11262);
xnor_4 g08914(new_n11185, new_n11180, new_n11263);
not_8  g08915(new_n11263, new_n11264);
xnor_4 g08916(new_n11241, new_n11236, new_n11265);
not_8  g08917(new_n11265, new_n11266_1);
nor_5  g08918(new_n11266_1, new_n11264, new_n11267);
not_8  g08919(new_n11267, new_n11268);
xnor_4 g08920(new_n11265, new_n11264, new_n11269);
nor_5  g08921(new_n8996, new_n8970, new_n11270);
not_8  g08922(new_n9004, new_n11271);
nor_5  g08923(new_n11271, new_n8997, new_n11272);
nor_5  g08924(new_n11272, new_n11270, new_n11273_1);
nand_5 g08925(new_n11273_1, new_n11269, new_n11274);
nand_5 g08926(new_n11274, new_n11268, new_n11275_1);
nand_5 g08927(new_n11275_1, new_n11262, new_n11276);
nand_5 g08928(new_n11276, new_n11261_1, new_n11277);
nand_5 g08929(new_n11277, new_n11257, new_n11278);
nand_5 g08930(new_n11278, new_n11255, new_n11279);
xnor_4 g08931(new_n11279, new_n11251, n1371);
xnor_4 g08932(n17250, n15241, new_n11281);
not_8  g08933(new_n11281, new_n11282);
not_8  g08934(n23160, new_n11283);
nor_5  g08935(new_n11283, n7678, new_n11284);
not_8  g08936(n16524, new_n11285);
nor_5  g08937(new_n11285, n3785, new_n11286);
xnor_4 g08938(n16524, n3785, new_n11287);
not_8  g08939(new_n11287, new_n11288);
nand_5 g08940(n20250, new_n6979, new_n11289);
nand_5 g08941(new_n8159_1, n5822, new_n11290_1);
xnor_4 g08942(n15271, n5822, new_n11291);
nand_5 g08943(n26443, new_n8163, new_n11292);
nand_5 g08944(new_n6091, new_n6090, new_n11293);
nand_5 g08945(new_n11293, new_n11292, new_n11294);
nand_5 g08946(new_n11294, new_n11291, new_n11295);
nand_5 g08947(new_n11295, new_n11290_1, new_n11296);
xnor_4 g08948(n20250, n11056, new_n11297);
nand_5 g08949(new_n11297, new_n11296, new_n11298);
nand_5 g08950(new_n11298, new_n11289, new_n11299);
nor_5  g08951(new_n11299, new_n11288, new_n11300);
nor_5  g08952(new_n11300, new_n11286, new_n11301);
xnor_4 g08953(n23160, n7678, new_n11302_1);
not_8  g08954(new_n11302_1, new_n11303);
nor_5  g08955(new_n11303, new_n11301, new_n11304);
nor_5  g08956(new_n11304, new_n11284, new_n11305);
xnor_4 g08957(new_n11305, new_n11282, new_n11306);
xnor_4 g08958(new_n10270, new_n2422, new_n11307);
nor_5  g08959(new_n10275_1, n26660, new_n11308);
xnor_4 g08960(new_n10275_1, new_n8101, new_n11309);
not_8  g08961(new_n11309, new_n11310);
not_8  g08962(n3018, new_n11311);
nor_5  g08963(new_n10299, new_n11311, new_n11312);
not_8  g08964(new_n11312, new_n11313_1);
nor_5  g08965(new_n10280, n3018, new_n11314);
not_8  g08966(new_n11314, new_n11315);
nor_5  g08967(new_n10283, new_n2398, new_n11316);
not_8  g08968(new_n11316, new_n11317);
not_8  g08969(new_n10049, new_n11318);
not_8  g08970(new_n10055_1, new_n11319);
nand_5 g08971(new_n11319, new_n10050, new_n11320);
nand_5 g08972(new_n11320, new_n11318, new_n11321);
nand_5 g08973(new_n11321, new_n10046, new_n11322);
nand_5 g08974(new_n11322, new_n11317, new_n11323);
nand_5 g08975(new_n11323, new_n11315, new_n11324);
nand_5 g08976(new_n11324, new_n11313_1, new_n11325_1);
nor_5  g08977(new_n11325_1, new_n11310, new_n11326_1);
nor_5  g08978(new_n11326_1, new_n11308, new_n11327);
xnor_4 g08979(new_n11327, new_n11307, new_n11328);
xnor_4 g08980(new_n11328, new_n11306, new_n11329);
xnor_4 g08981(new_n11325_1, new_n11309, new_n11330_1);
xnor_4 g08982(new_n11303, new_n11301, new_n11331);
nor_5  g08983(new_n11331, new_n11330_1, new_n11332);
xnor_4 g08984(new_n11331, new_n11330_1, new_n11333);
xnor_4 g08985(new_n11299, new_n11287, new_n11334);
not_8  g08986(new_n11334, new_n11335);
xnor_4 g08987(new_n10280, new_n11311, new_n11336);
xnor_4 g08988(new_n11336, new_n11323, new_n11337);
nand_5 g08989(new_n11337, new_n11335, new_n11338);
xnor_4 g08990(new_n11337, new_n11334, new_n11339);
xnor_4 g08991(new_n11297, new_n11296, new_n11340);
nor_5  g08992(new_n11340, new_n10058, new_n11341);
not_8  g08993(new_n11341, new_n11342);
not_8  g08994(new_n11340, new_n11343);
xnor_4 g08995(new_n11343, new_n10058, new_n11344);
not_8  g08996(new_n11291, new_n11345);
xnor_4 g08997(new_n11294, new_n11345, new_n11346);
nor_5  g08998(new_n11346, new_n10060, new_n11347_1);
xnor_4 g08999(new_n11346, new_n10060, new_n11348_1);
nand_5 g09000(new_n6092, new_n6089, new_n11349);
not_8  g09001(new_n11349, new_n11350);
not_8  g09002(new_n6094, new_n11351);
nor_5  g09003(new_n6104_1, new_n11351, new_n11352_1);
nor_5  g09004(new_n11352_1, new_n11350, new_n11353);
nor_5  g09005(new_n11353, new_n11348_1, new_n11354);
nor_5  g09006(new_n11354, new_n11347_1, new_n11355);
nand_5 g09007(new_n11355, new_n11344, new_n11356_1);
nand_5 g09008(new_n11356_1, new_n11342, new_n11357);
nand_5 g09009(new_n11357, new_n11339, new_n11358);
nand_5 g09010(new_n11358, new_n11338, new_n11359);
nor_5  g09011(new_n11359, new_n11333, new_n11360);
nor_5  g09012(new_n11360, new_n11332, new_n11361);
xnor_4 g09013(new_n11361, new_n11329, new_n11362);
xnor_4 g09014(new_n11362, new_n5924, new_n11363);
not_8  g09015(new_n11333, new_n11364);
xnor_4 g09016(new_n11359, new_n11364, new_n11365);
nor_5  g09017(new_n11365, new_n5929, new_n11366);
not_8  g09018(new_n11366, new_n11367);
xnor_4 g09019(new_n11365, new_n5930, new_n11368);
not_8  g09020(new_n11357, new_n11369);
xnor_4 g09021(new_n11369, new_n11339, new_n11370);
nor_5  g09022(new_n11370, new_n5935, new_n11371);
xnor_4 g09023(new_n11355, new_n11344, new_n11372);
nor_5  g09024(new_n11372, new_n5941, new_n11373);
not_8  g09025(new_n11373, new_n11374);
xnor_4 g09026(new_n11372, new_n5945, new_n11375_1);
xnor_4 g09027(new_n11353, new_n11348_1, new_n11376);
nor_5  g09028(new_n11376, new_n5949, new_n11377);
and_5  g09029(new_n6086, new_n5957, new_n11378);
not_8  g09030(new_n6105_1, new_n11379_1);
nor_5  g09031(new_n11379_1, new_n6088, new_n11380);
nor_5  g09032(new_n11380, new_n11378, new_n11381);
xnor_4 g09033(new_n11376, new_n5949, new_n11382);
nor_5  g09034(new_n11382, new_n11381, new_n11383);
nor_5  g09035(new_n11383, new_n11377, new_n11384);
nand_5 g09036(new_n11384, new_n11375_1, new_n11385);
nand_5 g09037(new_n11385, new_n11374, new_n11386_1);
xnor_4 g09038(new_n11370, new_n5935, new_n11387);
nor_5  g09039(new_n11387, new_n11386_1, new_n11388);
nor_5  g09040(new_n11388, new_n11371, new_n11389);
nand_5 g09041(new_n11389, new_n11368, new_n11390);
nand_5 g09042(new_n11390, new_n11367, new_n11391_1);
xor_4  g09043(new_n11391_1, new_n11363, n1385);
xnor_4 g09044(n26808, new_n4488, new_n11393);
nand_5 g09045(n26808, n24732, new_n11394);
xnor_4 g09046(n7339, n6631, new_n11395);
xnor_4 g09047(new_n11395, new_n11394, new_n11396);
not_8  g09048(new_n11396, new_n11397);
nor_5  g09049(new_n11397, new_n11393, new_n11398_1);
not_8  g09050(new_n11398_1, new_n11399);
xnor_4 g09051(n14684, new_n9660, new_n11400);
nor_5  g09052(n7339, n6631, new_n11401);
not_8  g09053(new_n11394, new_n11402);
nor_5  g09054(new_n11395, new_n11402, new_n11403_1);
nor_5  g09055(new_n11403_1, new_n11401, new_n11404);
xnor_4 g09056(new_n11404, new_n11400, new_n11405);
not_8  g09057(new_n11405, new_n11406);
nor_5  g09058(new_n11406, new_n11399, new_n11407);
not_8  g09059(n2680, new_n11408);
xnor_4 g09060(n17035, new_n11408, new_n11409);
nor_5  g09061(n14684, n1667, new_n11410);
not_8  g09062(new_n11400, new_n11411);
nor_5  g09063(new_n11404, new_n11411, new_n11412);
nor_5  g09064(new_n11412, new_n11410, new_n11413);
xnor_4 g09065(new_n11413, new_n11409, new_n11414);
nand_5 g09066(new_n11414, new_n11407, new_n11415);
xnor_4 g09067(n19905, new_n9659, new_n11416);
nor_5  g09068(n17035, n2680, new_n11417);
not_8  g09069(new_n11409, new_n11418);
nor_5  g09070(new_n11413, new_n11418, new_n11419_1);
nor_5  g09071(new_n11419_1, new_n11417, new_n11420);
xnor_4 g09072(new_n11420, new_n11416, new_n11421);
not_8  g09073(new_n11421, new_n11422);
nor_5  g09074(new_n11422, new_n11415, new_n11423);
xnor_4 g09075(n26452, new_n9733, new_n11424_1);
nor_5  g09076(n19905, n2547, new_n11425);
not_8  g09077(new_n11416, new_n11426);
nor_5  g09078(new_n11420, new_n11426, new_n11427);
nor_5  g09079(new_n11427, new_n11425, new_n11428);
xnor_4 g09080(new_n11428, new_n11424_1, new_n11429);
nand_5 g09081(new_n11429, new_n11423, new_n11430);
xnor_4 g09082(n15546, new_n9658, new_n11431);
not_8  g09083(new_n11431, new_n11432);
nor_5  g09084(n26452, n2999, new_n11433);
not_8  g09085(new_n11424_1, new_n11434);
nor_5  g09086(new_n11428, new_n11434, new_n11435);
nor_5  g09087(new_n11435, new_n11433, new_n11436);
xnor_4 g09088(new_n11436, new_n11432, new_n11437);
nor_5  g09089(new_n11437, new_n11430, new_n11438);
xnor_4 g09090(n13914, new_n11194, new_n11439_1);
nor_5  g09091(n15546, n14702, new_n11440);
not_8  g09092(new_n11440, new_n11441);
not_8  g09093(new_n11436, new_n11442);
nand_5 g09094(new_n11442, new_n11431, new_n11443);
nand_5 g09095(new_n11443, new_n11441, new_n11444);
xnor_4 g09096(new_n11444, new_n11439_1, new_n11445);
not_8  g09097(new_n11445, new_n11446);
nand_5 g09098(new_n11446, new_n11438, new_n11447);
xnor_4 g09099(n18035, new_n9657, new_n11448);
or_5   g09100(n13914, n5077, new_n11449);
nand_5 g09101(new_n11444, new_n11439_1, new_n11450);
nand_5 g09102(new_n11450, new_n11449, new_n11451);
xnor_4 g09103(new_n11451, new_n11448, new_n11452);
nor_5  g09104(new_n11452, new_n11447, new_n11453);
xnor_4 g09105(n8827, new_n9656, new_n11454);
or_5   g09106(n18035, n3279, new_n11455_1);
nand_5 g09107(new_n11451, new_n11448, new_n11456);
nand_5 g09108(new_n11456, new_n11455_1, new_n11457);
xnor_4 g09109(new_n11457, new_n11454, new_n11458);
not_8  g09110(new_n11458, new_n11459);
xnor_4 g09111(new_n11459, new_n11453, new_n11460);
xnor_4 g09112(new_n11460, new_n8463, new_n11461);
not_8  g09113(new_n11461, new_n11462_1);
not_8  g09114(new_n8467, new_n11463);
xnor_4 g09115(new_n11452, new_n11447, new_n11464);
nand_5 g09116(new_n11464, new_n11463, new_n11465);
xnor_4 g09117(new_n11464, new_n8467, new_n11466);
xnor_4 g09118(new_n11446, new_n11438, new_n11467);
nand_5 g09119(new_n11467, new_n8471, new_n11468);
xnor_4 g09120(new_n11467, new_n8472, new_n11469);
xnor_4 g09121(new_n11437, new_n11430, new_n11470_1);
nand_5 g09122(new_n11470_1, new_n8476, new_n11471);
xnor_4 g09123(new_n11470_1, new_n8477, new_n11472_1);
xnor_4 g09124(new_n11429, new_n11423, new_n11473_1);
nand_5 g09125(new_n11473_1, new_n8481, new_n11474);
xnor_4 g09126(new_n11473_1, new_n8482, new_n11475);
xnor_4 g09127(new_n11421, new_n11415, new_n11476);
not_8  g09128(new_n11476, new_n11477);
nand_5 g09129(new_n11477, new_n8485, new_n11478);
xnor_4 g09130(new_n11476, new_n8485, new_n11479_1);
not_8  g09131(new_n11407, new_n11480);
xnor_4 g09132(new_n11414, new_n11480, new_n11481_1);
nor_5  g09133(new_n11481_1, new_n11181, new_n11482);
not_8  g09134(new_n11482, new_n11483);
xnor_4 g09135(new_n11481_1, new_n8490, new_n11484);
xnor_4 g09136(new_n11405, new_n11399, new_n11485);
nor_5  g09137(new_n11485, new_n8497, new_n11486_1);
not_8  g09138(new_n11486_1, new_n11487);
xnor_4 g09139(new_n11485, new_n8496, new_n11488);
not_8  g09140(new_n11393, new_n11489);
nor_5  g09141(new_n11489, new_n8502, new_n11490);
nor_5  g09142(new_n11490, new_n8506, new_n11491);
nor_5  g09143(new_n11395, new_n11489, new_n11492);
nor_5  g09144(new_n11492, new_n11398_1, new_n11493);
not_8  g09145(new_n11490, new_n11494);
nor_5  g09146(new_n11494, new_n8445, new_n11495);
nor_5  g09147(new_n11495, new_n11491, new_n11496_1);
not_8  g09148(new_n11496_1, new_n11497);
nor_5  g09149(new_n11497, new_n11493, new_n11498);
nor_5  g09150(new_n11498, new_n11491, new_n11499);
not_8  g09151(new_n11499, new_n11500);
nand_5 g09152(new_n11500, new_n11488, new_n11501);
nand_5 g09153(new_n11501, new_n11487, new_n11502);
nand_5 g09154(new_n11502, new_n11484, new_n11503_1);
nand_5 g09155(new_n11503_1, new_n11483, new_n11504);
nand_5 g09156(new_n11504, new_n11479_1, new_n11505);
nand_5 g09157(new_n11505, new_n11478, new_n11506_1);
nand_5 g09158(new_n11506_1, new_n11475, new_n11507);
nand_5 g09159(new_n11507, new_n11474, new_n11508);
nand_5 g09160(new_n11508, new_n11472_1, new_n11509);
nand_5 g09161(new_n11509, new_n11471, new_n11510);
nand_5 g09162(new_n11510, new_n11469, new_n11511);
nand_5 g09163(new_n11511, new_n11468, new_n11512);
nand_5 g09164(new_n11512, new_n11466, new_n11513);
nand_5 g09165(new_n11513, new_n11465, new_n11514);
xnor_4 g09166(new_n11514, new_n11462_1, new_n11515_1);
xnor_4 g09167(new_n11515_1, new_n9714, new_n11516);
not_8  g09168(new_n9719, new_n11517);
not_8  g09169(new_n11466, new_n11518);
xnor_4 g09170(new_n11512, new_n11518, new_n11519);
nand_5 g09171(new_n11519, new_n11517, new_n11520);
xnor_4 g09172(new_n11519, new_n9719, new_n11521);
not_8  g09173(new_n11469, new_n11522);
xnor_4 g09174(new_n11510, new_n11522, new_n11523);
nand_5 g09175(new_n11523, new_n9726_1, new_n11524);
xnor_4 g09176(new_n11523, new_n9724, new_n11525);
not_8  g09177(new_n9730, new_n11526);
not_8  g09178(new_n11472_1, new_n11527);
xnor_4 g09179(new_n11508, new_n11527, new_n11528);
nand_5 g09180(new_n11528, new_n11526, new_n11529);
xnor_4 g09181(new_n11528, new_n9730, new_n11530);
xnor_4 g09182(new_n11506_1, new_n11475, new_n11531);
not_8  g09183(new_n11531, new_n11532);
nand_5 g09184(new_n11532, new_n9735, new_n11533);
xnor_4 g09185(new_n11531, new_n9735, new_n11534);
not_8  g09186(new_n11479_1, new_n11535);
xnor_4 g09187(new_n11504, new_n11535, new_n11536);
nand_5 g09188(new_n11536, new_n9739, new_n11537);
xnor_4 g09189(new_n11536, new_n9742, new_n11538_1);
xnor_4 g09190(new_n11502, new_n11484, new_n11539);
nor_5  g09191(new_n11539, new_n9746, new_n11540);
not_8  g09192(new_n11540, new_n11541);
xnor_4 g09193(new_n11499, new_n11488, new_n11542);
not_8  g09194(new_n11542, new_n11543);
nor_5  g09195(new_n11543, new_n9752, new_n11544);
not_8  g09196(new_n11544, new_n11545);
xnor_4 g09197(new_n11542, new_n9752, new_n11546);
not_8  g09198(new_n9763_1, new_n11547);
xnor_4 g09199(new_n11393, new_n2569, new_n11548_1);
nand_5 g09200(new_n11548_1, new_n11547, new_n11549);
nor_5  g09201(new_n11549, new_n9760, new_n11550);
not_8  g09202(new_n11550, new_n11551);
xnor_4 g09203(new_n11549, new_n9759, new_n11552);
xnor_4 g09204(new_n11496_1, new_n11493, new_n11553);
nand_5 g09205(new_n11553, new_n11552, new_n11554);
nand_5 g09206(new_n11554, new_n11551, new_n11555);
nand_5 g09207(new_n11555, new_n11546, new_n11556);
nand_5 g09208(new_n11556, new_n11545, new_n11557);
xnor_4 g09209(new_n11539, new_n9745, new_n11558);
nand_5 g09210(new_n11558, new_n11557, new_n11559);
nand_5 g09211(new_n11559, new_n11541, new_n11560);
nand_5 g09212(new_n11560, new_n11538_1, new_n11561);
nand_5 g09213(new_n11561, new_n11537, new_n11562);
nand_5 g09214(new_n11562, new_n11534, new_n11563);
nand_5 g09215(new_n11563, new_n11533, new_n11564_1);
nand_5 g09216(new_n11564_1, new_n11530, new_n11565);
nand_5 g09217(new_n11565, new_n11529, new_n11566_1);
nand_5 g09218(new_n11566_1, new_n11525, new_n11567);
nand_5 g09219(new_n11567, new_n11524, new_n11568);
nand_5 g09220(new_n11568, new_n11521, new_n11569);
nand_5 g09221(new_n11569, new_n11520, new_n11570);
xnor_4 g09222(new_n11570, new_n11516, n1498);
not_8  g09223(n9090, new_n11572);
xnor_4 g09224(n20658, new_n11572, new_n11573);
xnor_4 g09225(new_n11573, new_n6283, new_n11574);
xnor_4 g09226(new_n11574, new_n5267, n1501);
not_8  g09227(n25094, new_n11576);
not_8  g09228(n5131, new_n11577);
nor_5  g09229(n15506, n11473, new_n11578);
nand_5 g09230(new_n11578, new_n11577, new_n11579_1);
nor_5  g09231(new_n11579_1, n21538, new_n11580_1);
nand_5 g09232(new_n11580_1, new_n11576, new_n11581);
nor_5  g09233(new_n11581, n1611, new_n11582);
xnor_4 g09234(new_n11582, n752, new_n11583);
not_8  g09235(new_n11583, new_n11584);
xnor_4 g09236(new_n11584, new_n10319, new_n11585);
not_8  g09237(n1611, new_n11586);
xnor_4 g09238(new_n11581, new_n11586, new_n11587);
not_8  g09239(new_n11587, new_n11588);
nand_5 g09240(new_n11588, new_n10325, new_n11589);
xnor_4 g09241(new_n11587, new_n10325, new_n11590);
xnor_4 g09242(new_n11580_1, n25094, new_n11591_1);
not_8  g09243(new_n11591_1, new_n11592);
nand_5 g09244(new_n11592, new_n10332, new_n11593);
xnor_4 g09245(new_n11592, new_n10331, new_n11594);
not_8  g09246(n21538, new_n11595);
xnor_4 g09247(new_n11579_1, new_n11595, new_n11596);
not_8  g09248(new_n11596, new_n11597);
nor_5  g09249(new_n11597, new_n10338, new_n11598);
xnor_4 g09250(new_n11578, n5131, new_n11599);
not_8  g09251(new_n11599, new_n11600);
nand_5 g09252(new_n11600, new_n10345_1, new_n11601);
xnor_4 g09253(new_n11600, new_n10344, new_n11602);
nand_5 g09254(new_n10353, n15506, new_n11603);
xnor_4 g09255(n15506, n11473, new_n11604);
nand_5 g09256(new_n11604, new_n11603, new_n11605);
not_8  g09257(new_n11605, new_n11606);
nor_5  g09258(new_n11603, n11473, new_n11607_1);
nor_5  g09259(new_n11607_1, new_n11606, new_n11608);
nand_5 g09260(new_n11608, new_n10350, new_n11609);
nand_5 g09261(new_n11609, new_n11605, new_n11610);
nand_5 g09262(new_n11610, new_n11602, new_n11611);
nand_5 g09263(new_n11611, new_n11601, new_n11612);
xnor_4 g09264(new_n11597, new_n10338, new_n11613);
nor_5  g09265(new_n11613, new_n11612, new_n11614);
nor_5  g09266(new_n11614, new_n11598, new_n11615_1);
nand_5 g09267(new_n11615_1, new_n11594, new_n11616);
nand_5 g09268(new_n11616, new_n11593, new_n11617);
nand_5 g09269(new_n11617, new_n11590, new_n11618);
nand_5 g09270(new_n11618, new_n11589, new_n11619);
xnor_4 g09271(new_n11619, new_n11585, new_n11620);
not_8  g09272(n3366, new_n11621);
xnor_4 g09273(n20470, new_n11621, new_n11622);
not_8  g09274(n21222, new_n11623);
not_8  g09275(n26565, new_n11624);
or_5   g09276(new_n11624, new_n11623, new_n11625);
nor_5  g09277(n26565, n21222, new_n11626);
not_8  g09278(new_n11626, new_n11627);
nor_5  g09279(n9832, n3959, new_n11628);
not_8  g09280(new_n10122, new_n11629);
nor_5  g09281(new_n10140, new_n11629, new_n11630_1);
nor_5  g09282(new_n11630_1, new_n11628, new_n11631);
nand_5 g09283(new_n11631, new_n11627, new_n11632);
nand_5 g09284(new_n11632, new_n11625, new_n11633);
xnor_4 g09285(new_n11633, new_n11622, new_n11634);
xnor_4 g09286(new_n11634, new_n11620, new_n11635);
xnor_4 g09287(new_n11617, new_n11590, new_n11636);
xnor_4 g09288(n26565, new_n11623, new_n11637);
xnor_4 g09289(new_n11637, new_n11631, new_n11638);
nor_5  g09290(new_n11638, new_n11636, new_n11639);
not_8  g09291(new_n11639, new_n11640);
not_8  g09292(new_n11638, new_n11641);
xnor_4 g09293(new_n11641, new_n11636, new_n11642);
xnor_4 g09294(new_n11615_1, new_n11594, new_n11643);
nor_5  g09295(new_n11643, new_n10141, new_n11644);
not_8  g09296(new_n11644, new_n11645);
not_8  g09297(new_n10141, new_n11646);
xnor_4 g09298(new_n11643, new_n11646, new_n11647_1);
xnor_4 g09299(new_n11596, new_n10338, new_n11648);
xnor_4 g09300(new_n11648, new_n11612, new_n11649);
nor_5  g09301(new_n11649, new_n10199, new_n11650);
not_8  g09302(new_n11650, new_n11651);
xnor_4 g09303(new_n11649, new_n10202, new_n11652);
xnor_4 g09304(new_n11610, new_n11602, new_n11653);
nand_5 g09305(new_n11653, new_n10206, new_n11654);
xnor_4 g09306(new_n11608, new_n10350, new_n11655);
nor_5  g09307(new_n11655, new_n10212, new_n11656);
not_8  g09308(n15506, new_n11657);
xnor_4 g09309(new_n10353, new_n11657, new_n11658);
nor_5  g09310(new_n11658, new_n7635, new_n11659);
not_8  g09311(new_n11659, new_n11660);
xnor_4 g09312(new_n11655, new_n10212, new_n11661);
nor_5  g09313(new_n11661, new_n11660, new_n11662);
nor_5  g09314(new_n11662, new_n11656, new_n11663);
xnor_4 g09315(new_n11653, new_n10207, new_n11664);
nand_5 g09316(new_n11664, new_n11663, new_n11665);
nand_5 g09317(new_n11665, new_n11654, new_n11666);
not_8  g09318(new_n11666, new_n11667_1);
nand_5 g09319(new_n11667_1, new_n11652, new_n11668);
nand_5 g09320(new_n11668, new_n11651, new_n11669);
nand_5 g09321(new_n11669, new_n11647_1, new_n11670);
nand_5 g09322(new_n11670, new_n11645, new_n11671);
nand_5 g09323(new_n11671, new_n11642, new_n11672);
nand_5 g09324(new_n11672, new_n11640, new_n11673);
xnor_4 g09325(new_n11673, new_n11635, n1518);
not_8  g09326(n17458, new_n11675);
or_5   g09327(new_n11675, n14826, new_n11676);
xnor_4 g09328(n17458, n14826, new_n11677);
not_8  g09329(n1222, new_n11678);
or_5   g09330(n23493, new_n11678, new_n11679);
xnor_4 g09331(n23493, n1222, new_n11680);
not_8  g09332(n25240, new_n11681);
or_5   g09333(new_n11681, n10275, new_n11682_1);
xnor_4 g09334(n25240, n10275, new_n11683);
or_5   g09335(n15146, new_n7647_1, new_n11684);
xnor_4 g09336(n15146, n10125, new_n11685);
or_5   g09337(n11579, new_n7650, new_n11686);
xnor_4 g09338(n11579, n8067, new_n11687);
nor_5  g09339(new_n11178, n21, new_n11688);
xnor_4 g09340(n20923, n21, new_n11689);
not_8  g09341(new_n11689, new_n11690);
not_8  g09342(n18157, new_n11691);
nor_5  g09343(new_n11691, n1682, new_n11692);
xnor_4 g09344(n18157, n1682, new_n11693);
nor_5  g09345(n12161, new_n10522, new_n11694);
nor_5  g09346(new_n6982, n7963, new_n11695);
nor_5  g09347(new_n10524, n5026, new_n11696);
nor_5  g09348(n10017, new_n7661, new_n11697);
not_8  g09349(n3618, new_n11698);
nor_5  g09350(n8581, new_n11698, new_n11699);
not_8  g09351(new_n11699, new_n11700);
nor_5  g09352(new_n11700, new_n11697, new_n11701);
nor_5  g09353(new_n11701, new_n11696, new_n11702);
nor_5  g09354(new_n11702, new_n11695, new_n11703);
nor_5  g09355(new_n11703, new_n11694, new_n11704);
nand_5 g09356(new_n11704, new_n11693, new_n11705);
not_8  g09357(new_n11705, new_n11706);
nor_5  g09358(new_n11706, new_n11692, new_n11707);
nor_5  g09359(new_n11707, new_n11690, new_n11708);
nor_5  g09360(new_n11708, new_n11688, new_n11709);
not_8  g09361(new_n11709, new_n11710_1);
nand_5 g09362(new_n11710_1, new_n11687, new_n11711);
nand_5 g09363(new_n11711, new_n11686, new_n11712_1);
nand_5 g09364(new_n11712_1, new_n11685, new_n11713);
nand_5 g09365(new_n11713, new_n11684, new_n11714);
nand_5 g09366(new_n11714, new_n11683, new_n11715);
nand_5 g09367(new_n11715, new_n11682_1, new_n11716);
nand_5 g09368(new_n11716, new_n11680, new_n11717);
nand_5 g09369(new_n11717, new_n11679, new_n11718);
nand_5 g09370(new_n11718, new_n11677, new_n11719);
nand_5 g09371(new_n11719, new_n11676, new_n11720);
not_8  g09372(new_n11720, new_n11721);
not_8  g09373(n19282, new_n11722);
nand_5 g09374(new_n4386, new_n2734, new_n11723);
nor_5  g09375(new_n11723, n12821, new_n11724_1);
nand_5 g09376(new_n11724_1, new_n2726, new_n11725);
nor_5  g09377(new_n11725, n7330, new_n11726);
nand_5 g09378(new_n11726, new_n2720, new_n11727);
xnor_4 g09379(new_n11727, new_n2717, new_n11728);
not_8  g09380(new_n11728, new_n11729);
nor_5  g09381(new_n11729, new_n11722, new_n11730);
nor_5  g09382(new_n11727, n2944, new_n11731);
not_8  g09383(new_n11731, new_n11732);
xnor_4 g09384(new_n11726, n767, new_n11733);
nor_5  g09385(new_n11733, n12657, new_n11734);
xnor_4 g09386(new_n11733, new_n2986, new_n11735);
not_8  g09387(new_n11735, new_n11736_1);
xnor_4 g09388(new_n11725, new_n2723, new_n11737);
nand_5 g09389(new_n11737, n17077, new_n11738);
not_8  g09390(n17077, new_n11739);
xnor_4 g09391(new_n11737, new_n11739, new_n11740);
xnor_4 g09392(new_n11724_1, n22492, new_n11741_1);
nand_5 g09393(new_n11741_1, n26510, new_n11742);
not_8  g09394(new_n11741_1, new_n11743);
xnor_4 g09395(new_n11743, n26510, new_n11744);
not_8  g09396(n12821, new_n11745);
xnor_4 g09397(new_n11723, new_n11745, new_n11746);
nand_5 g09398(new_n11746, n23068, new_n11747);
not_8  g09399(n23068, new_n11748);
not_8  g09400(new_n11746, new_n11749_1);
nand_5 g09401(new_n11749_1, new_n11748, new_n11750);
nand_5 g09402(new_n4387, n19514, new_n11751);
nand_5 g09403(new_n4408, new_n4389, new_n11752);
nand_5 g09404(new_n11752, new_n11751, new_n11753);
nand_5 g09405(new_n11753, new_n11750, new_n11754);
nand_5 g09406(new_n11754, new_n11747, new_n11755);
nand_5 g09407(new_n11755, new_n11744, new_n11756);
nand_5 g09408(new_n11756, new_n11742, new_n11757);
nand_5 g09409(new_n11757, new_n11740, new_n11758);
nand_5 g09410(new_n11758, new_n11738, new_n11759);
nor_5  g09411(new_n11759, new_n11736_1, new_n11760);
nor_5  g09412(new_n11760, new_n11734, new_n11761);
nand_5 g09413(new_n11729, new_n11722, new_n11762);
nand_5 g09414(new_n11762, new_n11761, new_n11763);
nand_5 g09415(new_n11763, new_n11732, new_n11764);
nor_5  g09416(new_n11764, new_n11730, new_n11765);
nor_5  g09417(new_n11765, new_n11721, new_n11766);
xnor_4 g09418(new_n11718, new_n11677, new_n11767);
xnor_4 g09419(new_n11728, new_n11722, new_n11768);
xnor_4 g09420(new_n11768, new_n11761, new_n11769);
nand_5 g09421(new_n11769, new_n11767, new_n11770_1);
not_8  g09422(new_n11769, new_n11771_1);
xnor_4 g09423(new_n11771_1, new_n11767, new_n11772);
xnor_4 g09424(new_n11716, new_n11680, new_n11773);
xnor_4 g09425(new_n11759, new_n11735, new_n11774);
nand_5 g09426(new_n11774, new_n11773, new_n11775_1);
not_8  g09427(new_n11774, new_n11776);
xnor_4 g09428(new_n11776, new_n11773, new_n11777);
not_8  g09429(new_n11683, new_n11778);
xnor_4 g09430(new_n11714, new_n11778, new_n11779);
not_8  g09431(new_n11779, new_n11780);
xnor_4 g09432(new_n11757, new_n11740, new_n11781);
nand_5 g09433(new_n11781, new_n11780, new_n11782);
xnor_4 g09434(new_n11781, new_n11779, new_n11783);
xnor_4 g09435(new_n11712_1, new_n11685, new_n11784);
xnor_4 g09436(new_n11755, new_n11744, new_n11785);
nand_5 g09437(new_n11785, new_n11784, new_n11786);
not_8  g09438(new_n11785, new_n11787);
xnor_4 g09439(new_n11787, new_n11784, new_n11788);
xnor_4 g09440(new_n11709, new_n11687, new_n11789);
not_8  g09441(new_n11789, new_n11790);
xnor_4 g09442(new_n11746, new_n11748, new_n11791);
xnor_4 g09443(new_n11791, new_n11753, new_n11792);
nand_5 g09444(new_n11792, new_n11790, new_n11793);
xnor_4 g09445(new_n11792, new_n11789, new_n11794);
xnor_4 g09446(new_n11707, new_n11689, new_n11795);
not_8  g09447(new_n11795, new_n11796);
nand_5 g09448(new_n11796, new_n4409_1, new_n11797);
xnor_4 g09449(new_n11704, new_n11693, new_n11798);
nand_5 g09450(new_n11798, new_n4440, new_n11799);
not_8  g09451(new_n11798, new_n11800);
xnor_4 g09452(new_n11800, new_n4440, new_n11801);
xnor_4 g09453(n12161, n7963, new_n11802);
xnor_4 g09454(new_n11802, new_n11702, new_n11803);
nand_5 g09455(new_n11803, new_n4462, new_n11804);
not_8  g09456(new_n11803, new_n11805);
xnor_4 g09457(new_n11805, new_n4462, new_n11806);
xnor_4 g09458(n8581, n3618, new_n11807);
nor_5  g09459(new_n11807, new_n4456, new_n11808);
xnor_4 g09460(n10017, n5026, new_n11809);
xnor_4 g09461(new_n11809, new_n11700, new_n11810);
not_8  g09462(new_n11810, new_n11811);
nor_5  g09463(new_n11811, new_n11808, new_n11812);
xnor_4 g09464(new_n11810, new_n11808, new_n11813);
not_8  g09465(new_n11813, new_n11814);
nor_5  g09466(new_n11814, new_n4448, new_n11815);
nor_5  g09467(new_n11815, new_n11812, new_n11816);
not_8  g09468(new_n11816, new_n11817);
nand_5 g09469(new_n11817, new_n11806, new_n11818_1);
nand_5 g09470(new_n11818_1, new_n11804, new_n11819);
nand_5 g09471(new_n11819, new_n11801, new_n11820);
nand_5 g09472(new_n11820, new_n11799, new_n11821);
xnor_4 g09473(new_n11795, new_n4409_1, new_n11822);
nand_5 g09474(new_n11822, new_n11821, new_n11823);
nand_5 g09475(new_n11823, new_n11797, new_n11824);
nand_5 g09476(new_n11824, new_n11794, new_n11825);
nand_5 g09477(new_n11825, new_n11793, new_n11826);
nand_5 g09478(new_n11826, new_n11788, new_n11827);
nand_5 g09479(new_n11827, new_n11786, new_n11828);
nand_5 g09480(new_n11828, new_n11783, new_n11829);
nand_5 g09481(new_n11829, new_n11782, new_n11830);
nand_5 g09482(new_n11830, new_n11777, new_n11831);
nand_5 g09483(new_n11831, new_n11775_1, new_n11832);
nand_5 g09484(new_n11832, new_n11772, new_n11833);
nand_5 g09485(new_n11833, new_n11770_1, new_n11834);
xnor_4 g09486(new_n11765, new_n11721, new_n11835);
nor_5  g09487(new_n11835, new_n11834, new_n11836);
nor_5  g09488(new_n11836, new_n11766, new_n11837_1);
or_5   g09489(n20040, new_n7886, new_n11838);
nand_5 g09490(new_n9272, new_n9235, new_n11839);
nand_5 g09491(new_n11839, new_n11838, new_n11840);
xnor_4 g09492(new_n11840, new_n11837_1, new_n11841_1);
xnor_4 g09493(new_n11835, new_n11834, new_n11842_1);
nand_5 g09494(new_n11842_1, new_n11840, new_n11843_1);
xnor_4 g09495(new_n11832, new_n11772, new_n11844);
not_8  g09496(new_n11844, new_n11845);
nand_5 g09497(new_n11845, new_n9273, new_n11846);
xnor_4 g09498(new_n11844, new_n9273, new_n11847);
xnor_4 g09499(new_n11830, new_n11777, new_n11848);
not_8  g09500(new_n11848, new_n11849);
nand_5 g09501(new_n11849, new_n9340, new_n11850);
xnor_4 g09502(new_n11848, new_n9340, new_n11851);
xnor_4 g09503(new_n11828, new_n11783, new_n11852);
not_8  g09504(new_n11852, new_n11853);
nand_5 g09505(new_n11853, new_n9348, new_n11854);
xnor_4 g09506(new_n11852, new_n9348, new_n11855);
xnor_4 g09507(new_n11826, new_n11788, new_n11856);
not_8  g09508(new_n11856, new_n11857);
nand_5 g09509(new_n11857, new_n9355, new_n11858);
xnor_4 g09510(new_n11856, new_n9355, new_n11859);
not_8  g09511(new_n11794, new_n11860);
xnor_4 g09512(new_n11824, new_n11860, new_n11861);
nand_5 g09513(new_n11861, new_n9360, new_n11862);
xnor_4 g09514(new_n11861, new_n9364_1, new_n11863);
xnor_4 g09515(new_n11822, new_n11821, new_n11864);
not_8  g09516(new_n11864, new_n11865);
nor_5  g09517(new_n11865, new_n9366, new_n11866);
xnor_4 g09518(new_n11819, new_n11801, new_n11867);
nor_5  g09519(new_n11867, new_n9372_1, new_n11868);
not_8  g09520(new_n11868, new_n11869);
xnor_4 g09521(new_n11867, new_n9371_1, new_n11870);
xnor_4 g09522(new_n11816, new_n11806, new_n11871);
not_8  g09523(new_n11871, new_n11872);
nor_5  g09524(new_n11872, new_n9380_1, new_n11873);
not_8  g09525(new_n11873, new_n11874);
xnor_4 g09526(new_n11807, new_n4455, new_n11875);
not_8  g09527(new_n11875, new_n11876);
nor_5  g09528(new_n11876, new_n9388, new_n11877);
and_5  g09529(new_n11877, new_n9386, new_n11878);
xnor_4 g09530(new_n11813, new_n4448, new_n11879);
not_8  g09531(new_n11879, new_n11880);
xnor_4 g09532(new_n11877, new_n9385, new_n11881);
and_5  g09533(new_n11881, new_n11880, new_n11882);
nor_5  g09534(new_n11882, new_n11878, new_n11883);
xnor_4 g09535(new_n11871, new_n9380_1, new_n11884);
nand_5 g09536(new_n11884, new_n11883, new_n11885);
nand_5 g09537(new_n11885, new_n11874, new_n11886);
nand_5 g09538(new_n11886, new_n11870, new_n11887);
nand_5 g09539(new_n11887, new_n11869, new_n11888);
not_8  g09540(new_n9366, new_n11889);
xnor_4 g09541(new_n11864, new_n11889, new_n11890);
nor_5  g09542(new_n11890, new_n11888, new_n11891);
nor_5  g09543(new_n11891, new_n11866, new_n11892);
nand_5 g09544(new_n11892, new_n11863, new_n11893);
nand_5 g09545(new_n11893, new_n11862, new_n11894);
nand_5 g09546(new_n11894, new_n11859, new_n11895);
nand_5 g09547(new_n11895, new_n11858, new_n11896);
nand_5 g09548(new_n11896, new_n11855, new_n11897);
nand_5 g09549(new_n11897, new_n11854, new_n11898_1);
nand_5 g09550(new_n11898_1, new_n11851, new_n11899);
nand_5 g09551(new_n11899, new_n11850, new_n11900);
nand_5 g09552(new_n11900, new_n11847, new_n11901);
nand_5 g09553(new_n11901, new_n11846, new_n11902);
not_8  g09554(new_n11840, new_n11903);
xnor_4 g09555(new_n11842_1, new_n11903, new_n11904);
nand_5 g09556(new_n11904, new_n11902, new_n11905_1);
nand_5 g09557(new_n11905_1, new_n11843_1, new_n11906);
xnor_4 g09558(new_n11906, new_n11841_1, n1527);
xnor_4 g09559(n25345, n23463, new_n11908);
or_5   g09560(new_n3171, n9655, new_n11909);
xnor_4 g09561(n13074, n9655, new_n11910);
not_8  g09562(n10739, new_n11911);
or_5   g09563(n13490, new_n11911, new_n11912);
xnor_4 g09564(n13490, n10739, new_n11913);
or_5   g09565(n22660, new_n2350, new_n11914);
xnor_4 g09566(n22660, n21753, new_n11915);
nor_5  g09567(new_n2353, n1777, new_n11916);
xnor_4 g09568(n21832, n1777, new_n11917);
nor_5  g09569(new_n2356, n8745, new_n11918);
not_8  g09570(new_n11918, new_n11919);
nor_5  g09571(n16223, new_n2445, new_n11920);
not_8  g09572(new_n10380, new_n11921);
nor_5  g09573(new_n10385_1, new_n11921, new_n11922);
nor_5  g09574(new_n11922, new_n11920, new_n11923);
xnor_4 g09575(n26913, n8745, new_n11924);
nand_5 g09576(new_n11924, new_n11923, new_n11925);
nand_5 g09577(new_n11925, new_n11919, new_n11926_1);
and_5  g09578(new_n11926_1, new_n11917, new_n11927);
nor_5  g09579(new_n11927, new_n11916, new_n11928);
not_8  g09580(new_n11928, new_n11929);
nand_5 g09581(new_n11929, new_n11915, new_n11930);
nand_5 g09582(new_n11930, new_n11914, new_n11931);
nand_5 g09583(new_n11931, new_n11913, new_n11932);
nand_5 g09584(new_n11932, new_n11912, new_n11933);
nand_5 g09585(new_n11933, new_n11910, new_n11934);
nand_5 g09586(new_n11934, new_n11909, new_n11935);
xnor_4 g09587(new_n11935, new_n11908, new_n11936);
xnor_4 g09588(new_n11936, new_n8341, new_n11937);
xnor_4 g09589(new_n11933, new_n11910, new_n11938);
nand_5 g09590(new_n11938, new_n8347, new_n11939);
xnor_4 g09591(new_n8259_1, new_n8205, new_n11940);
xnor_4 g09592(new_n11938, new_n11940, new_n11941);
xnor_4 g09593(new_n11931, new_n11913, new_n11942);
nand_5 g09594(new_n11942, new_n8353, new_n11943);
xnor_4 g09595(new_n11942, new_n8352, new_n11944);
xnor_4 g09596(new_n11928, new_n11915, new_n11945);
not_8  g09597(new_n11945, new_n11946);
nand_5 g09598(new_n11946, new_n8359, new_n11947);
xnor_4 g09599(new_n11945, new_n8359, new_n11948);
not_8  g09600(new_n11917, new_n11949);
xnor_4 g09601(new_n11926_1, new_n11949, new_n11950);
not_8  g09602(new_n11950, new_n11951);
nand_5 g09603(new_n11951, new_n8367, new_n11952);
xnor_4 g09604(new_n11950, new_n8367, new_n11953);
xnor_4 g09605(new_n11924, new_n11923, new_n11954);
nand_5 g09606(new_n11954, new_n8374, new_n11955);
nand_5 g09607(new_n10386, new_n8378, new_n11956);
nand_5 g09608(new_n10398, new_n10387_1, new_n11957);
nand_5 g09609(new_n11957, new_n11956, new_n11958);
xnor_4 g09610(new_n11954, new_n8370, new_n11959);
nand_5 g09611(new_n11959, new_n11958, new_n11960);
nand_5 g09612(new_n11960, new_n11955, new_n11961);
nand_5 g09613(new_n11961, new_n11953, new_n11962);
nand_5 g09614(new_n11962, new_n11952, new_n11963);
nand_5 g09615(new_n11963, new_n11948, new_n11964);
nand_5 g09616(new_n11964, new_n11947, new_n11965_1);
nand_5 g09617(new_n11965_1, new_n11944, new_n11966);
nand_5 g09618(new_n11966, new_n11943, new_n11967);
nand_5 g09619(new_n11967, new_n11941, new_n11968);
nand_5 g09620(new_n11968, new_n11939, new_n11969);
xnor_4 g09621(new_n11969, new_n11937, n1580);
xnor_4 g09622(n18962, n12315, new_n11971);
nor_5  g09623(new_n11971, new_n7856, new_n11972);
nor_5  g09624(new_n9149, n12315, new_n11973);
xnor_4 g09625(n10158, n3952, new_n11974);
xnor_4 g09626(new_n11974, new_n11973, new_n11975);
xnor_4 g09627(new_n11975, new_n11972, new_n11976);
xnor_4 g09628(new_n11976, new_n7862, n1586);
xnor_4 g09629(n19539, n1483, new_n11978);
not_8  g09630(n8194, new_n11979);
or_5   g09631(n24093, new_n11979, new_n11980_1);
xnor_4 g09632(n24093, n8194, new_n11981);
not_8  g09633(n23657, new_n11982);
or_5   g09634(new_n11982, n23035, new_n11983);
xnor_4 g09635(n23657, n23035, new_n11984);
not_8  g09636(n16911, new_n11985);
or_5   g09637(new_n11985, n7773, new_n11986);
nand_5 g09638(new_n6803, new_n6771, new_n11987);
nand_5 g09639(new_n11987, new_n11986, new_n11988);
nand_5 g09640(new_n11988, new_n11984, new_n11989);
nand_5 g09641(new_n11989, new_n11983, new_n11990);
nand_5 g09642(new_n11990, new_n11981, new_n11991);
nand_5 g09643(new_n11991, new_n11980_1, new_n11992);
xnor_4 g09644(new_n11992, new_n11978, new_n11993);
xnor_4 g09645(n25494, n1314, new_n11994);
or_5   g09646(n10117, new_n8786, new_n11995);
xnor_4 g09647(n10117, n3306, new_n11996);
or_5   g09648(new_n8735, n13460, new_n11997);
xnor_4 g09649(n22335, n13460, new_n11998);
or_5   g09650(new_n8740, n6104, new_n11999);
or_5   g09651(n4119, new_n8745_1, new_n12000_1);
not_8  g09652(new_n4874, new_n12001);
nand_5 g09653(new_n12001, new_n4849, new_n12002);
nand_5 g09654(new_n12002, new_n12000_1, new_n12003_1);
xnor_4 g09655(n24048, n6104, new_n12004);
nand_5 g09656(new_n12004, new_n12003_1, new_n12005);
nand_5 g09657(new_n12005, new_n11999, new_n12006);
nand_5 g09658(new_n12006, new_n11998, new_n12007);
nand_5 g09659(new_n12007, new_n11997, new_n12008);
nand_5 g09660(new_n12008, new_n11996, new_n12009);
nand_5 g09661(new_n12009, new_n11995, new_n12010);
xnor_4 g09662(new_n12010, new_n11994, new_n12011_1);
xnor_4 g09663(n25296, n23717, new_n12012);
not_8  g09664(n7788, new_n12013);
or_5   g09665(n20013, new_n12013, new_n12014);
xnor_4 g09666(n20013, n7788, new_n12015);
not_8  g09667(n5443, new_n12016);
or_5   g09668(new_n12016, n1320, new_n12017);
xnor_4 g09669(n5443, n1320, new_n12018);
not_8  g09670(n18584, new_n12019);
or_5   g09671(n19803, new_n12019, new_n12020);
nand_5 g09672(new_n6768, new_n6763, new_n12021);
nand_5 g09673(new_n12021, new_n12020, new_n12022);
nand_5 g09674(new_n12022, new_n12018, new_n12023);
nand_5 g09675(new_n12023, new_n12017, new_n12024);
nand_5 g09676(new_n12024, new_n12015, new_n12025);
nand_5 g09677(new_n12025, new_n12014, new_n12026);
xnor_4 g09678(new_n12026, new_n12012, new_n12027);
not_8  g09679(new_n12027, new_n12028);
xnor_4 g09680(new_n12028, new_n12011_1, new_n12029);
xnor_4 g09681(new_n12008, new_n11996, new_n12030);
not_8  g09682(new_n12030, new_n12031);
xnor_4 g09683(new_n12024, new_n12015, new_n12032);
not_8  g09684(new_n12032, new_n12033);
nand_5 g09685(new_n12033, new_n12031, new_n12034);
xnor_4 g09686(new_n12033, new_n12030, new_n12035);
xnor_4 g09687(new_n12006, new_n11998, new_n12036);
not_8  g09688(new_n12036, new_n12037);
xnor_4 g09689(new_n12022, new_n12018, new_n12038);
not_8  g09690(new_n12038, new_n12039);
nor_5  g09691(new_n12039, new_n12037, new_n12040);
xnor_4 g09692(new_n12038, new_n12036, new_n12041);
xnor_4 g09693(new_n12004, new_n12003_1, new_n12042);
not_8  g09694(new_n12042, new_n12043);
nand_5 g09695(new_n12043, new_n6770, new_n12044);
xnor_4 g09696(new_n12043, new_n6769, new_n12045);
nand_5 g09697(new_n4903, new_n4875, new_n12046);
nand_5 g09698(new_n4948, new_n4905, new_n12047);
nand_5 g09699(new_n12047, new_n12046, new_n12048);
nand_5 g09700(new_n12048, new_n12045, new_n12049);
nand_5 g09701(new_n12049, new_n12044, new_n12050);
nor_5  g09702(new_n12050, new_n12041, new_n12051);
nor_5  g09703(new_n12051, new_n12040, new_n12052);
nand_5 g09704(new_n12052, new_n12035, new_n12053);
nand_5 g09705(new_n12053, new_n12034, new_n12054);
xnor_4 g09706(new_n12054, new_n12029, new_n12055);
xnor_4 g09707(new_n12055, new_n11993, new_n12056);
not_8  g09708(new_n12056, new_n12057);
not_8  g09709(new_n11981, new_n12058);
xnor_4 g09710(new_n11990, new_n12058, new_n12059);
not_8  g09711(new_n12059, new_n12060);
xnor_4 g09712(new_n12052, new_n12035, new_n12061);
nand_5 g09713(new_n12061, new_n12060, new_n12062);
xnor_4 g09714(new_n12061, new_n12059, new_n12063);
xnor_4 g09715(new_n11988, new_n11984, new_n12064);
xnor_4 g09716(new_n12050, new_n12041, new_n12065);
not_8  g09717(new_n12065, new_n12066);
nand_5 g09718(new_n12066, new_n12064, new_n12067);
xnor_4 g09719(new_n12065, new_n12064, new_n12068);
xnor_4 g09720(new_n12048, new_n12045, new_n12069);
nand_5 g09721(new_n12069, new_n6804, new_n12070);
not_8  g09722(new_n12069, new_n12071);
xnor_4 g09723(new_n12071, new_n6804, new_n12072_1);
nand_5 g09724(new_n6855, new_n4949, new_n12073);
not_8  g09725(new_n6861_1, new_n12074);
nand_5 g09726(new_n12074, new_n4955, new_n12075);
xnor_4 g09727(new_n12074, new_n4952_1, new_n12076);
not_8  g09728(new_n4957_1, new_n12077);
nand_5 g09729(new_n6867_1, new_n12077, new_n12078);
nor_5  g09730(new_n6875, new_n4962, new_n12079);
xnor_4 g09731(new_n6877, new_n4962, new_n12080);
not_8  g09732(new_n12080, new_n12081);
nor_5  g09733(new_n6883, new_n4972_1, new_n12082);
nor_5  g09734(new_n12082, new_n6887, new_n12083);
xnor_4 g09735(new_n12082, new_n6886, new_n12084);
and_5  g09736(new_n12084, new_n4978, new_n12085);
nor_5  g09737(new_n12085, new_n12083, new_n12086);
nor_5  g09738(new_n12086, new_n12081, new_n12087);
nor_5  g09739(new_n12087, new_n12079, new_n12088);
not_8  g09740(new_n12088, new_n12089);
xnor_4 g09741(new_n6867_1, new_n4957_1, new_n12090);
nand_5 g09742(new_n12090, new_n12089, new_n12091);
nand_5 g09743(new_n12091, new_n12078, new_n12092);
nand_5 g09744(new_n12092, new_n12076, new_n12093);
nand_5 g09745(new_n12093, new_n12075, new_n12094);
xnor_4 g09746(new_n6854, new_n4949, new_n12095);
nand_5 g09747(new_n12095, new_n12094, new_n12096);
nand_5 g09748(new_n12096, new_n12073, new_n12097);
nand_5 g09749(new_n12097, new_n12072_1, new_n12098);
nand_5 g09750(new_n12098, new_n12070, new_n12099);
nand_5 g09751(new_n12099, new_n12068, new_n12100);
nand_5 g09752(new_n12100, new_n12067, new_n12101);
nand_5 g09753(new_n12101, new_n12063, new_n12102);
nand_5 g09754(new_n12102, new_n12062, new_n12103);
xnor_4 g09755(new_n12103, new_n12057, n1590);
xnor_4 g09756(new_n8075, new_n8057, n1602);
xnor_4 g09757(new_n2895, new_n2835, n1634);
xnor_4 g09758(new_n12101, new_n12063, n1636);
nor_5  g09759(n10514, n4514, new_n12108);
not_8  g09760(new_n12108, new_n12109);
not_8  g09761(n4514, new_n12110);
xnor_4 g09762(n10514, new_n12110, new_n12111);
nor_5  g09763(n18649, n3984, new_n12112);
not_8  g09764(new_n12112, new_n12113_1);
not_8  g09765(n3984, new_n12114);
xnor_4 g09766(n18649, new_n12114, new_n12115);
not_8  g09767(n6218, new_n12116);
not_8  g09768(n19652, new_n12117);
or_5   g09769(new_n12117, new_n12116, new_n12118);
not_8  g09770(new_n12118, new_n12119);
nor_5  g09771(n19652, n6218, new_n12120);
nor_5  g09772(n20470, n3366, new_n12121_1);
not_8  g09773(new_n11622, new_n12122);
nor_5  g09774(new_n11633, new_n12122, new_n12123);
nor_5  g09775(new_n12123, new_n12121_1, new_n12124);
not_8  g09776(new_n12124, new_n12125);
nor_5  g09777(new_n12125, new_n12120, new_n12126);
nor_5  g09778(new_n12126, new_n12119, new_n12127);
nand_5 g09779(new_n12127, new_n12115, new_n12128);
nand_5 g09780(new_n12128, new_n12113_1, new_n12129);
nand_5 g09781(new_n12129, new_n12111, new_n12130);
nand_5 g09782(new_n12130, new_n12109, new_n12131_1);
not_8  g09783(n20040, new_n12132);
xnor_4 g09784(n18880, new_n7886, new_n12133);
not_8  g09785(new_n12133, new_n12134);
or_5   g09786(n25475, n23697, new_n12135);
nand_5 g09787(new_n7156, new_n7115, new_n12136);
nand_5 g09788(new_n12136, new_n12135, new_n12137);
xnor_4 g09789(new_n12137, new_n12134, new_n12138);
nor_5  g09790(new_n12138, new_n12132, new_n12139);
not_8  g09791(new_n12139, new_n12140);
xnor_4 g09792(new_n12138, n20040, new_n12141);
not_8  g09793(n19531, new_n12142);
nor_5  g09794(new_n7157, new_n12142, new_n12143);
not_8  g09795(new_n12143, new_n12144);
xnor_4 g09796(new_n7157, n19531, new_n12145);
nor_5  g09797(new_n7160, n18345, new_n12146_1);
xnor_4 g09798(new_n7160, new_n2591, new_n12147);
not_8  g09799(new_n12147, new_n12148);
nor_5  g09800(new_n7165, n13190, new_n12149);
not_8  g09801(n13190, new_n12150);
xnor_4 g09802(new_n7164, new_n12150, new_n12151);
nor_5  g09803(new_n7169, new_n2599, new_n12152_1);
not_8  g09804(new_n12152_1, new_n12153_1);
not_8  g09805(new_n7171, new_n12154);
nor_5  g09806(new_n12154, new_n2603, new_n12155);
not_8  g09807(new_n12155, new_n12156);
nand_5 g09808(new_n10165_1, new_n10147, new_n12157_1);
nand_5 g09809(new_n12157_1, new_n12156, new_n12158_1);
xnor_4 g09810(new_n7169, n3460, new_n12159);
nand_5 g09811(new_n12159, new_n12158_1, new_n12160);
nand_5 g09812(new_n12160, new_n12153_1, new_n12161_1);
nor_5  g09813(new_n12161_1, new_n12151, new_n12162);
nor_5  g09814(new_n12162, new_n12149, new_n12163);
nor_5  g09815(new_n12163, new_n12148, new_n12164);
nor_5  g09816(new_n12164, new_n12146_1, new_n12165);
nand_5 g09817(new_n12165, new_n12145, new_n12166);
nand_5 g09818(new_n12166, new_n12144, new_n12167);
nand_5 g09819(new_n12167, new_n12141, new_n12168);
nand_5 g09820(new_n12168, new_n12140, new_n12169);
or_5   g09821(n18880, n2978, new_n12170);
nand_5 g09822(new_n12137, new_n12133, new_n12171);
nand_5 g09823(new_n12171, new_n12170, new_n12172);
xnor_4 g09824(new_n12172, new_n12169, new_n12173);
not_8  g09825(n17037, new_n12174);
not_8  g09826(n26191, new_n12175);
not_8  g09827(n19575, new_n12176);
nand_5 g09828(new_n10145, new_n12176, new_n12177);
nor_5  g09829(new_n12177, n26512, new_n12178);
nand_5 g09830(new_n12178, new_n12175, new_n12179_1);
nor_5  g09831(new_n12179_1, n5386, new_n12180);
nand_5 g09832(new_n12180, new_n12174, new_n12181);
nor_5  g09833(new_n12181, n7569, new_n12182);
xnor_4 g09834(new_n12182, new_n12173, new_n12183);
xnor_4 g09835(new_n12167, new_n12141, new_n12184);
not_8  g09836(n7569, new_n12185);
xnor_4 g09837(new_n12181, new_n12185, new_n12186);
not_8  g09838(new_n12186, new_n12187);
nand_5 g09839(new_n12187, new_n12184, new_n12188);
not_8  g09840(new_n12188, new_n12189);
xnor_4 g09841(new_n12187, new_n12184, new_n12190);
not_8  g09842(new_n12145, new_n12191);
xnor_4 g09843(new_n12165, new_n12191, new_n12192_1);
xnor_4 g09844(new_n12180, n17037, new_n12193);
nor_5  g09845(new_n12193, new_n12192_1, new_n12194);
xnor_4 g09846(new_n12193, new_n12192_1, new_n12195);
xnor_4 g09847(new_n12163, new_n12147, new_n12196);
not_8  g09848(new_n12196, new_n12197);
not_8  g09849(n5386, new_n12198);
xnor_4 g09850(new_n12179_1, new_n12198, new_n12199);
nor_5  g09851(new_n12199, new_n12197, new_n12200);
xnor_4 g09852(new_n12199, new_n12196, new_n12201);
not_8  g09853(new_n12201, new_n12202);
xnor_4 g09854(new_n12161_1, new_n12151, new_n12203);
xnor_4 g09855(new_n12178, n26191, new_n12204);
nor_5  g09856(new_n12204, new_n12203, new_n12205);
not_8  g09857(n26512, new_n12206);
xnor_4 g09858(new_n12177, new_n12206, new_n12207);
xnor_4 g09859(new_n7169, new_n2599, new_n12208);
xnor_4 g09860(new_n12208, new_n12158_1, new_n12209_1);
nand_5 g09861(new_n12209_1, new_n12207, new_n12210);
not_8  g09862(new_n12209_1, new_n12211);
xnor_4 g09863(new_n12211, new_n12207, new_n12212);
nor_5  g09864(new_n10167, new_n10146, new_n12213);
nor_5  g09865(new_n10195, new_n10168, new_n12214);
nor_5  g09866(new_n12214, new_n12213, new_n12215);
nand_5 g09867(new_n12215, new_n12212, new_n12216);
nand_5 g09868(new_n12216, new_n12210, new_n12217);
xnor_4 g09869(new_n12204, new_n12203, new_n12218);
nor_5  g09870(new_n12218, new_n12217, new_n12219);
nor_5  g09871(new_n12219, new_n12205, new_n12220);
nor_5  g09872(new_n12220, new_n12202, new_n12221);
nor_5  g09873(new_n12221, new_n12200, new_n12222);
nor_5  g09874(new_n12222, new_n12195, new_n12223_1);
nor_5  g09875(new_n12223_1, new_n12194, new_n12224);
nor_5  g09876(new_n12224, new_n12190, new_n12225_1);
nor_5  g09877(new_n12225_1, new_n12189, new_n12226);
xnor_4 g09878(new_n12226, new_n12183, new_n12227);
xnor_4 g09879(new_n12227, new_n12131_1, new_n12228_1);
not_8  g09880(new_n12190, new_n12229);
xnor_4 g09881(new_n12224, new_n12229, new_n12230);
xnor_4 g09882(new_n12129, new_n12111, new_n12231);
nand_5 g09883(new_n12231, new_n12230, new_n12232);
not_8  g09884(new_n12231, new_n12233);
xnor_4 g09885(new_n12233, new_n12230, new_n12234);
not_8  g09886(new_n12195, new_n12235_1);
xnor_4 g09887(new_n12222, new_n12235_1, new_n12236);
xnor_4 g09888(new_n12127, new_n12115, new_n12237);
nand_5 g09889(new_n12237, new_n12236, new_n12238);
xnor_4 g09890(new_n12222, new_n12195, new_n12239);
xnor_4 g09891(new_n12237, new_n12239, new_n12240);
xnor_4 g09892(new_n12220, new_n12201, new_n12241);
xnor_4 g09893(n19652, new_n12116, new_n12242);
xnor_4 g09894(new_n12242, new_n12124, new_n12243);
not_8  g09895(new_n12243, new_n12244);
nand_5 g09896(new_n12244, new_n12241, new_n12245);
xnor_4 g09897(new_n12243, new_n12241, new_n12246);
xnor_4 g09898(new_n12218, new_n12217, new_n12247);
nor_5  g09899(new_n12247, new_n11634, new_n12248);
not_8  g09900(new_n12248, new_n12249);
not_8  g09901(new_n11634, new_n12250);
xnor_4 g09902(new_n12247, new_n12250, new_n12251);
not_8  g09903(new_n12212, new_n12252);
xnor_4 g09904(new_n12215, new_n12252, new_n12253);
not_8  g09905(new_n12253, new_n12254);
nor_5  g09906(new_n12254, new_n11641, new_n12255);
nor_5  g09907(new_n12253, new_n11638, new_n12256);
nand_5 g09908(new_n10196, new_n10141, new_n12257);
not_8  g09909(new_n12257, new_n12258);
nor_5  g09910(new_n10223, new_n10197, new_n12259);
nor_5  g09911(new_n12259, new_n12258, new_n12260);
nor_5  g09912(new_n12260, new_n12256, new_n12261);
nor_5  g09913(new_n12261, new_n12255, new_n12262);
nand_5 g09914(new_n12262, new_n12251, new_n12263);
nand_5 g09915(new_n12263, new_n12249, new_n12264);
nand_5 g09916(new_n12264, new_n12246, new_n12265);
nand_5 g09917(new_n12265, new_n12245, new_n12266);
nand_5 g09918(new_n12266, new_n12240, new_n12267);
nand_5 g09919(new_n12267, new_n12238, new_n12268);
nand_5 g09920(new_n12268, new_n12234, new_n12269);
nand_5 g09921(new_n12269, new_n12232, new_n12270);
xnor_4 g09922(new_n12270, new_n12228_1, n1684);
not_8  g09923(n13026, new_n12272);
xnor_4 g09924(new_n6540, new_n12114, new_n12273);
nand_5 g09925(new_n6548, new_n12117, new_n12274);
xnor_4 g09926(new_n6546, new_n12117, new_n12275);
nand_5 g09927(new_n6553, new_n11621, new_n12276);
xnor_4 g09928(new_n6552, new_n11621, new_n12277);
nand_5 g09929(new_n4183, new_n11624, new_n12278);
xnor_4 g09930(new_n4183, n26565, new_n12279);
nand_5 g09931(new_n4187, new_n10121, new_n12280);
xnor_4 g09932(new_n4186_1, new_n10121, new_n12281);
not_8  g09933(n11566, new_n12282);
nand_5 g09934(new_n4192, new_n12282, new_n12283);
xnor_4 g09935(new_n4191, new_n12282, new_n12284);
not_8  g09936(n26744, new_n12285);
not_8  g09937(new_n4196, new_n12286);
nand_5 g09938(new_n12286, new_n12285, new_n12287);
xnor_4 g09939(new_n4196, new_n12285, new_n12288);
not_8  g09940(n26625, new_n12289);
nand_5 g09941(new_n4202, new_n12289, new_n12290);
nand_5 g09942(n19922, n14230, new_n12291);
xnor_4 g09943(new_n4202, n26625, new_n12292);
nand_5 g09944(new_n12292, new_n12291, new_n12293);
nand_5 g09945(new_n12293, new_n12290, new_n12294);
nand_5 g09946(new_n12294, new_n12288, new_n12295);
nand_5 g09947(new_n12295, new_n12287, new_n12296);
nand_5 g09948(new_n12296, new_n12284, new_n12297);
nand_5 g09949(new_n12297, new_n12283, new_n12298);
nand_5 g09950(new_n12298, new_n12281, new_n12299);
nand_5 g09951(new_n12299, new_n12280, new_n12300);
nand_5 g09952(new_n12300, new_n12279, new_n12301);
nand_5 g09953(new_n12301, new_n12278, new_n12302_1);
nand_5 g09954(new_n12302_1, new_n12277, new_n12303);
nand_5 g09955(new_n12303, new_n12276, new_n12304_1);
nand_5 g09956(new_n12304_1, new_n12275, new_n12305);
nand_5 g09957(new_n12305, new_n12274, new_n12306);
xnor_4 g09958(new_n12306, new_n12273, new_n12307);
nand_5 g09959(new_n12307, new_n12272, new_n12308);
xnor_4 g09960(new_n12307, n13026, new_n12309);
not_8  g09961(n2175, new_n12310);
xnor_4 g09962(new_n12304_1, new_n12275, new_n12311);
nand_5 g09963(new_n12311, new_n12310, new_n12312);
xnor_4 g09964(new_n12311, n2175, new_n12313);
not_8  g09965(n752, new_n12314);
xnor_4 g09966(new_n12302_1, new_n12277, new_n12315_1);
nand_5 g09967(new_n12315_1, new_n12314, new_n12316);
xnor_4 g09968(new_n12315_1, n752, new_n12317);
xnor_4 g09969(new_n12300, new_n12279, new_n12318);
nand_5 g09970(new_n12318, new_n11586, new_n12319);
xnor_4 g09971(new_n12298, new_n12281, new_n12320);
nand_5 g09972(new_n12320, new_n11576, new_n12321);
xnor_4 g09973(new_n12320, n25094, new_n12322);
xnor_4 g09974(new_n12296, new_n12284, new_n12323);
nand_5 g09975(new_n12323, new_n11595, new_n12324_1);
xnor_4 g09976(new_n12323, n21538, new_n12325_1);
xnor_4 g09977(new_n12294, new_n12288, new_n12326);
nand_5 g09978(new_n12326, new_n11577, new_n12327);
not_8  g09979(n11473, new_n12328);
xnor_4 g09980(new_n12292, new_n12291, new_n12329_1);
nand_5 g09981(new_n12329_1, new_n12328, new_n12330_1);
xnor_4 g09982(n19922, n14230, new_n12331);
nand_5 g09983(new_n12331, n15506, new_n12332);
xnor_4 g09984(new_n12329_1, n11473, new_n12333);
nand_5 g09985(new_n12333, new_n12332, new_n12334);
nand_5 g09986(new_n12334, new_n12330_1, new_n12335);
xnor_4 g09987(new_n12326, n5131, new_n12336);
nand_5 g09988(new_n12336, new_n12335, new_n12337);
nand_5 g09989(new_n12337, new_n12327, new_n12338);
nand_5 g09990(new_n12338, new_n12325_1, new_n12339);
nand_5 g09991(new_n12339, new_n12324_1, new_n12340);
nand_5 g09992(new_n12340, new_n12322, new_n12341_1);
nand_5 g09993(new_n12341_1, new_n12321, new_n12342);
xnor_4 g09994(new_n12318, n1611, new_n12343);
nand_5 g09995(new_n12343, new_n12342, new_n12344);
nand_5 g09996(new_n12344, new_n12319, new_n12345);
nand_5 g09997(new_n12345, new_n12317, new_n12346_1);
nand_5 g09998(new_n12346_1, new_n12316, new_n12347);
nand_5 g09999(new_n12347, new_n12313, new_n12348);
nand_5 g10000(new_n12348, new_n12312, new_n12349_1);
nand_5 g10001(new_n12349_1, new_n12309, new_n12350);
nand_5 g10002(new_n12350, new_n12308, new_n12351);
not_8  g10003(new_n12351, new_n12352);
nand_5 g10004(new_n12352, n23912, new_n12353);
xnor_4 g10005(new_n12351, n23912, new_n12354);
not_8  g10006(new_n6540, new_n12355);
nand_5 g10007(new_n12355, new_n12114, new_n12356);
nand_5 g10008(new_n12306, new_n12273, new_n12357);
nand_5 g10009(new_n12357, new_n12356, new_n12358);
xnor_4 g10010(new_n6533, n4514, new_n12359);
xnor_4 g10011(new_n12359, new_n12358, new_n12360);
not_8  g10012(new_n12360, new_n12361);
nand_5 g10013(new_n12361, new_n12354, new_n12362);
nand_5 g10014(new_n12362, new_n12353, new_n12363);
or_5   g10015(new_n6533, new_n12110, new_n12364_1);
nor_5  g10016(new_n6537, n4514, new_n12365);
nor_5  g10017(new_n12365, new_n12358, new_n12366);
nor_5  g10018(new_n12366, new_n6535, new_n12367);
nand_5 g10019(new_n12367, new_n12364_1, new_n12368);
not_8  g10020(new_n12368, new_n12369);
nor_5  g10021(new_n12369, new_n12363, new_n12370);
nand_5 g10022(new_n4664, new_n10962, new_n12371);
xnor_4 g10023(new_n4663, new_n10962, new_n12372);
nand_5 g10024(new_n4672, new_n10950, new_n12373);
xnor_4 g10025(new_n4671, new_n10950, new_n12374);
nand_5 g10026(new_n4677, new_n6648, new_n12375);
xnor_4 g10027(new_n4676, new_n6648, new_n12376);
nand_5 g10028(new_n4683, new_n10951, new_n12377);
xnor_4 g10029(new_n4682, new_n10951, new_n12378);
nor_5  g10030(new_n4133, n13677, new_n12379);
not_8  g10031(new_n12379, new_n12380_1);
nand_5 g10032(new_n4167, new_n4134_1, new_n12381);
nand_5 g10033(new_n12381, new_n12380_1, new_n12382);
nand_5 g10034(new_n12382, new_n12378, new_n12383_1);
nand_5 g10035(new_n12383_1, new_n12377, new_n12384_1);
nand_5 g10036(new_n12384_1, new_n12376, new_n12385);
nand_5 g10037(new_n12385, new_n12375, new_n12386);
nand_5 g10038(new_n12386, new_n12374, new_n12387);
nand_5 g10039(new_n12387, new_n12373, new_n12388);
nand_5 g10040(new_n12388, new_n12372, new_n12389);
nand_5 g10041(new_n12389, new_n12371, new_n12390);
nor_5  g10042(new_n12390, new_n4645, new_n12391);
xnor_4 g10043(new_n12390, new_n4645, new_n12392);
xnor_4 g10044(new_n12368, new_n12363, new_n12393);
not_8  g10045(new_n12393, new_n12394);
nand_5 g10046(new_n12394, new_n12392, new_n12395);
xnor_4 g10047(new_n12393, new_n12392, new_n12396);
not_8  g10048(new_n12372, new_n12397_1);
xnor_4 g10049(new_n12388, new_n12397_1, new_n12398_1);
xnor_4 g10050(new_n12360, new_n12354, new_n12399);
nand_5 g10051(new_n12399, new_n12398_1, new_n12400);
xnor_4 g10052(new_n12386, new_n12374, new_n12401);
not_8  g10053(new_n12401, new_n12402);
xnor_4 g10054(new_n12349_1, new_n12309, new_n12403);
nand_5 g10055(new_n12403, new_n12402, new_n12404);
xnor_4 g10056(new_n12403, new_n12401, new_n12405);
xnor_4 g10057(new_n12384_1, new_n12376, new_n12406);
not_8  g10058(new_n12406, new_n12407);
xnor_4 g10059(new_n12347, new_n12313, new_n12408_1);
nand_5 g10060(new_n12408_1, new_n12407, new_n12409);
xnor_4 g10061(new_n12408_1, new_n12406, new_n12410);
xnor_4 g10062(new_n12382, new_n12378, new_n12411);
not_8  g10063(new_n12411, new_n12412);
xnor_4 g10064(new_n12345, new_n12317, new_n12413);
nand_5 g10065(new_n12413, new_n12412, new_n12414);
xnor_4 g10066(new_n12413, new_n12411, new_n12415);
not_8  g10067(new_n4168, new_n12416);
xnor_4 g10068(new_n12343, new_n12342, new_n12417);
nand_5 g10069(new_n12417, new_n12416, new_n12418);
xnor_4 g10070(new_n12417, new_n4168, new_n12419);
xnor_4 g10071(new_n12340, new_n12322, new_n12420);
nand_5 g10072(new_n12420, new_n4260, new_n12421);
xnor_4 g10073(new_n12338, new_n12325_1, new_n12422);
nand_5 g10074(new_n12422, new_n4266_1, new_n12423);
xnor_4 g10075(new_n12422, new_n4265, new_n12424);
xnor_4 g10076(new_n12336, new_n12335, new_n12425);
nand_5 g10077(new_n12425, new_n4270, new_n12426);
not_8  g10078(new_n12332, new_n12427);
xnor_4 g10079(new_n12333, new_n12427, new_n12428);
nor_5  g10080(new_n12428, new_n4277, new_n12429);
not_8  g10081(new_n12429, new_n12430);
xnor_4 g10082(new_n12331, new_n11657, new_n12431);
nor_5  g10083(new_n12431, new_n4280, new_n12432);
not_8  g10084(new_n12432, new_n12433);
xnor_4 g10085(new_n12428, new_n4276, new_n12434);
nand_5 g10086(new_n12434, new_n12433, new_n12435);
nand_5 g10087(new_n12435, new_n12430, new_n12436);
xnor_4 g10088(new_n12425, new_n4269, new_n12437);
nand_5 g10089(new_n12437, new_n12436, new_n12438);
nand_5 g10090(new_n12438, new_n12426, new_n12439);
nand_5 g10091(new_n12439, new_n12424, new_n12440);
nand_5 g10092(new_n12440, new_n12423, new_n12441);
xnor_4 g10093(new_n12420, new_n4259, new_n12442);
nand_5 g10094(new_n12442, new_n12441, new_n12443);
nand_5 g10095(new_n12443, new_n12421, new_n12444);
nand_5 g10096(new_n12444, new_n12419, new_n12445);
nand_5 g10097(new_n12445, new_n12418, new_n12446_1);
nand_5 g10098(new_n12446_1, new_n12415, new_n12447);
nand_5 g10099(new_n12447, new_n12414, new_n12448);
nand_5 g10100(new_n12448, new_n12410, new_n12449_1);
nand_5 g10101(new_n12449_1, new_n12409, new_n12450);
nand_5 g10102(new_n12450, new_n12405, new_n12451);
nand_5 g10103(new_n12451, new_n12404, new_n12452);
not_8  g10104(new_n12398_1, new_n12453);
xnor_4 g10105(new_n12399, new_n12453, new_n12454);
nand_5 g10106(new_n12454, new_n12452, new_n12455);
nand_5 g10107(new_n12455, new_n12400, new_n12456);
nand_5 g10108(new_n12456, new_n12396, new_n12457);
nand_5 g10109(new_n12457, new_n12395, new_n12458);
xnor_4 g10110(new_n12458, new_n12391, new_n12459);
xnor_4 g10111(new_n12459, new_n12370, n1701);
xnor_4 g10112(new_n4091, new_n4059, n1703);
xnor_4 g10113(new_n4813, new_n4753, n1721);
nand_5 g10114(new_n8187, new_n4547, new_n12463);
not_8  g10115(new_n12463, new_n12464);
nor_5  g10116(new_n9528, new_n9527, new_n12465);
nor_5  g10117(new_n12465, new_n12464, new_n12466);
not_8  g10118(new_n12466, new_n12467_1);
nand_5 g10119(new_n12467_1, new_n9577, new_n12468);
nand_5 g10120(new_n9576, new_n9529, new_n12469_1);
nand_5 g10121(new_n9654, new_n9578, new_n12470);
nand_5 g10122(new_n12470, new_n12469_1, new_n12471);
nand_5 g10123(new_n12471, new_n12468, new_n12472);
nand_5 g10124(new_n12466, new_n9576, new_n12473);
nand_5 g10125(new_n12473, new_n12470, new_n12474);
nand_5 g10126(new_n12474, new_n12472, new_n12475);
not_8  g10127(new_n12475, n1760);
xnor_4 g10128(new_n4285, new_n4273, n1791);
xnor_4 g10129(new_n3489, new_n3488, n1808);
not_8  g10130(new_n8187, new_n12479);
nand_5 g10131(new_n12479, new_n8140, new_n12480);
nand_5 g10132(new_n8265, new_n8188, new_n12481);
nand_5 g10133(new_n12481, new_n12480, new_n12482);
or_5   g10134(n13494, new_n3164_1, new_n12483);
xnor_4 g10135(n13494, n4319, new_n12484);
not_8  g10136(n23463, new_n12485);
or_5   g10137(n25345, new_n12485, new_n12486);
nand_5 g10138(new_n11935, new_n11908, new_n12487);
nand_5 g10139(new_n12487, new_n12486, new_n12488);
nand_5 g10140(new_n12488, new_n12484, new_n12489);
nand_5 g10141(new_n12489, new_n12483, new_n12490);
nor_5  g10142(new_n12490, new_n12482, new_n12491);
nand_5 g10143(new_n12490, new_n8266, new_n12492);
not_8  g10144(new_n12492, new_n12493);
xnor_4 g10145(new_n12490, new_n8266, new_n12494);
xnor_4 g10146(new_n12488, new_n12484, new_n12495_1);
nor_5  g10147(new_n12495_1, new_n8335, new_n12496);
not_8  g10148(new_n12496, new_n12497);
xnor_4 g10149(new_n12495_1, new_n8334, new_n12498);
nor_5  g10150(new_n11936, new_n8342, new_n12499);
not_8  g10151(new_n12499, new_n12500);
not_8  g10152(new_n11969, new_n12501);
nand_5 g10153(new_n12501, new_n11937, new_n12502);
nand_5 g10154(new_n12502, new_n12500, new_n12503);
nand_5 g10155(new_n12503, new_n12498, new_n12504);
nand_5 g10156(new_n12504, new_n12497, new_n12505);
nor_5  g10157(new_n12505, new_n12494, new_n12506);
nor_5  g10158(new_n12506, new_n12493, new_n12507_1);
nor_5  g10159(new_n12507_1, new_n12491, new_n12508);
nand_5 g10160(new_n12490, new_n12482, new_n12509);
not_8  g10161(new_n12509, new_n12510);
nor_5  g10162(new_n12510, new_n12506, new_n12511);
nor_5  g10163(new_n12511, new_n12508, n1821);
xnor_4 g10164(new_n7336, new_n7335_1, n1832);
not_8  g10165(n2160, new_n12514);
xnor_4 g10166(n9934, new_n7613, new_n12515_1);
not_8  g10167(new_n12515_1, new_n12516_1);
or_5   g10168(n25331, n18496, new_n12517);
not_8  g10169(n18496, new_n12518);
xnor_4 g10170(n25331, new_n12518, new_n12519);
or_5   g10171(n26224, n18483, new_n12520);
xnor_4 g10172(n26224, new_n7362, new_n12521);
nor_5  g10173(n21934, n19327, new_n12522);
xnor_4 g10174(n21934, new_n3878, new_n12523);
not_8  g10175(new_n12523, new_n12524);
nor_5  g10176(n22597, n18901, new_n12525);
xnor_4 g10177(n22597, new_n7368, new_n12526);
not_8  g10178(new_n12526, new_n12527);
nor_5  g10179(n26107, n4376, new_n12528);
xnor_4 g10180(n26107, new_n7371, new_n12529);
not_8  g10181(new_n12529, new_n12530);
nor_5  g10182(n14570, n342, new_n12531);
xnor_4 g10183(n14570, new_n3899, new_n12532);
not_8  g10184(new_n12532, new_n12533);
nor_5  g10185(n26553, n23775, new_n12534);
xnor_4 g10186(n26553, new_n7379, new_n12535);
not_8  g10187(new_n12535, new_n12536);
nor_5  g10188(n8259, n4964, new_n12537);
nand_5 g10189(n11479, n7876, new_n12538);
not_8  g10190(new_n12538, new_n12539);
xnor_4 g10191(n8259, n4964, new_n12540_1);
nor_5  g10192(new_n12540_1, new_n12539, new_n12541);
nor_5  g10193(new_n12541, new_n12537, new_n12542);
nor_5  g10194(new_n12542, new_n12536, new_n12543);
nor_5  g10195(new_n12543, new_n12534, new_n12544);
nor_5  g10196(new_n12544, new_n12533, new_n12545_1);
nor_5  g10197(new_n12545_1, new_n12531, new_n12546_1);
nor_5  g10198(new_n12546_1, new_n12530, new_n12547);
nor_5  g10199(new_n12547, new_n12528, new_n12548);
nor_5  g10200(new_n12548, new_n12527, new_n12549);
nor_5  g10201(new_n12549, new_n12525, new_n12550);
nor_5  g10202(new_n12550, new_n12524, new_n12551);
nor_5  g10203(new_n12551, new_n12522, new_n12552_1);
not_8  g10204(new_n12552_1, new_n12553);
nand_5 g10205(new_n12553, new_n12521, new_n12554);
nand_5 g10206(new_n12554, new_n12520, new_n12555);
nand_5 g10207(new_n12555, new_n12519, new_n12556);
nand_5 g10208(new_n12556, new_n12517, new_n12557);
xnor_4 g10209(new_n12557, new_n12516_1, new_n12558);
xnor_4 g10210(new_n12558, new_n12514, new_n12559);
not_8  g10211(new_n12519, new_n12560);
xnor_4 g10212(new_n12555, new_n12560, new_n12561);
nor_5  g10213(new_n12561, n10763, new_n12562_1);
xnor_4 g10214(new_n12561, n10763, new_n12563);
xnor_4 g10215(new_n12552_1, new_n12521, new_n12564);
nand_5 g10216(new_n12564, n7437, new_n12565);
xnor_4 g10217(new_n12564, new_n2944_1, new_n12566_1);
xnor_4 g10218(new_n12550, new_n12523, new_n12567);
nand_5 g10219(new_n12567, n20700, new_n12568);
xnor_4 g10220(new_n12567, new_n2947, new_n12569_1);
xnor_4 g10221(new_n12548, new_n12526, new_n12570);
nand_5 g10222(new_n12570, n7099, new_n12571);
xnor_4 g10223(new_n12570, new_n2951, new_n12572);
xnor_4 g10224(new_n12546_1, new_n12529, new_n12573);
nand_5 g10225(new_n12573, n12811, new_n12574);
not_8  g10226(n12811, new_n12575);
xnor_4 g10227(new_n12573, new_n12575, new_n12576);
xnor_4 g10228(new_n12544, new_n12532, new_n12577);
nand_5 g10229(new_n12577, n1118, new_n12578);
not_8  g10230(new_n12578, new_n12579);
xnor_4 g10231(new_n12577, new_n2959, new_n12580);
not_8  g10232(new_n12580, new_n12581);
xnor_4 g10233(new_n12542, new_n12535, new_n12582);
nand_5 g10234(new_n12582, n25974, new_n12583);
not_8  g10235(n25974, new_n12584);
xnor_4 g10236(new_n12582, new_n12584, new_n12585);
not_8  g10237(n1630, new_n12586);
xnor_4 g10238(n11479, n7876, new_n12587_1);
nand_5 g10239(new_n12587_1, n1451, new_n12588);
nand_5 g10240(new_n12588, new_n12586, new_n12589);
not_8  g10241(new_n12589, new_n12590);
xnor_4 g10242(new_n12540_1, new_n12538, new_n12591);
xnor_4 g10243(new_n12588, n1630, new_n12592);
not_8  g10244(new_n12592, new_n12593_1);
nor_5  g10245(new_n12593_1, new_n12591, new_n12594);
nor_5  g10246(new_n12594, new_n12590, new_n12595);
nand_5 g10247(new_n12595, new_n12585, new_n12596);
nand_5 g10248(new_n12596, new_n12583, new_n12597);
not_8  g10249(new_n12597, new_n12598);
nor_5  g10250(new_n12598, new_n12581, new_n12599);
nor_5  g10251(new_n12599, new_n12579, new_n12600);
not_8  g10252(new_n12600, new_n12601);
nand_5 g10253(new_n12601, new_n12576, new_n12602);
nand_5 g10254(new_n12602, new_n12574, new_n12603);
nand_5 g10255(new_n12603, new_n12572, new_n12604);
nand_5 g10256(new_n12604, new_n12571, new_n12605);
nand_5 g10257(new_n12605, new_n12569_1, new_n12606);
nand_5 g10258(new_n12606, new_n12568, new_n12607_1);
nand_5 g10259(new_n12607_1, new_n12566_1, new_n12608);
nand_5 g10260(new_n12608, new_n12565, new_n12609);
nor_5  g10261(new_n12609, new_n12563, new_n12610);
nor_5  g10262(new_n12610, new_n12562_1, new_n12611);
xnor_4 g10263(new_n12611, new_n12559, new_n12612);
not_8  g10264(new_n12612, new_n12613);
not_8  g10265(n21784, new_n12614);
not_8  g10266(n5521, new_n12615);
nand_5 g10267(new_n3999, new_n6318, new_n12616);
nor_5  g10268(new_n12616, n11926, new_n12617);
nand_5 g10269(new_n12617, new_n12615, new_n12618);
xnor_4 g10270(new_n12618, new_n12614, new_n12619);
xnor_4 g10271(new_n12619, new_n7707, new_n12620_1);
xnor_4 g10272(new_n12617, n5521, new_n12621_1);
not_8  g10273(new_n12621_1, new_n12622);
nand_5 g10274(new_n12622, new_n7711, new_n12623);
xnor_4 g10275(new_n12621_1, new_n7711, new_n12624);
xnor_4 g10276(new_n12616, n11926, new_n12625);
nand_5 g10277(new_n12625, new_n7718, new_n12626_1);
xnor_4 g10278(new_n12625, new_n7718, new_n12627);
not_8  g10279(new_n12627, new_n12628);
not_8  g10280(new_n4000_1, new_n12629);
nand_5 g10281(new_n12629, new_n3992, new_n12630);
nand_5 g10282(new_n4052, new_n4001, new_n12631);
nand_5 g10283(new_n12631, new_n12630, new_n12632);
nand_5 g10284(new_n12632, new_n12628, new_n12633);
nand_5 g10285(new_n12633, new_n12626_1, new_n12634);
nand_5 g10286(new_n12634, new_n12624, new_n12635);
nand_5 g10287(new_n12635, new_n12623, new_n12636);
xnor_4 g10288(new_n12636, new_n12620_1, new_n12637);
xnor_4 g10289(new_n12637, new_n12613, new_n12638);
xnor_4 g10290(new_n12609, new_n12563, new_n12639);
xnor_4 g10291(new_n12634, new_n12624, new_n12640);
not_8  g10292(new_n12640, new_n12641);
nand_5 g10293(new_n12641, new_n12639, new_n12642);
xnor_4 g10294(new_n12640, new_n12639, new_n12643);
xnor_4 g10295(new_n12607_1, new_n12566_1, new_n12644);
not_8  g10296(new_n12644, new_n12645);
xnor_4 g10297(new_n12632, new_n12627, new_n12646);
nand_5 g10298(new_n12646, new_n12645, new_n12647);
xnor_4 g10299(new_n12646, new_n12644, new_n12648);
not_8  g10300(new_n4053, new_n12649);
xnor_4 g10301(new_n12605, new_n12569_1, new_n12650_1);
not_8  g10302(new_n12650_1, new_n12651);
nand_5 g10303(new_n12651, new_n12649, new_n12652);
xnor_4 g10304(new_n12651, new_n4053, new_n12653);
not_8  g10305(new_n12572, new_n12654_1);
xnor_4 g10306(new_n12603, new_n12654_1, new_n12655);
nand_5 g10307(new_n12655, new_n4056, new_n12656);
xnor_4 g10308(new_n12655, new_n4055, new_n12657_1);
xnor_4 g10309(new_n12600, new_n12576, new_n12658);
nand_5 g10310(new_n12658, new_n4061, new_n12659);
xnor_4 g10311(new_n12658, new_n4060, new_n12660);
xnor_4 g10312(new_n12598, new_n12580, new_n12661);
not_8  g10313(new_n12661, new_n12662);
nor_5  g10314(new_n12662, new_n4065, new_n12663);
not_8  g10315(new_n12663, new_n12664);
xnor_4 g10316(new_n12661, new_n4065, new_n12665_1);
xnor_4 g10317(new_n12595, new_n12585, new_n12666);
nor_5  g10318(new_n12666, new_n4070, new_n12667);
not_8  g10319(new_n12667, new_n12668);
xnor_4 g10320(new_n12666, new_n4071_1, new_n12669);
not_8  g10321(new_n4080, new_n12670_1);
not_8  g10322(n1451, new_n12671);
xnor_4 g10323(new_n12587_1, new_n12671, new_n12672);
nor_5  g10324(new_n12672, new_n12670_1, new_n12673);
xnor_4 g10325(new_n12592, new_n12591, new_n12674);
and_5  g10326(new_n12674, new_n12673, new_n12675);
xnor_4 g10327(new_n12674, new_n12673, new_n12676);
nor_5  g10328(new_n12676, new_n4076, new_n12677);
nor_5  g10329(new_n12677, new_n12675, new_n12678);
nand_5 g10330(new_n12678, new_n12669, new_n12679);
nand_5 g10331(new_n12679, new_n12668, new_n12680);
nand_5 g10332(new_n12680, new_n12665_1, new_n12681);
nand_5 g10333(new_n12681, new_n12664, new_n12682);
nand_5 g10334(new_n12682, new_n12660, new_n12683);
nand_5 g10335(new_n12683, new_n12659, new_n12684);
nand_5 g10336(new_n12684, new_n12657_1, new_n12685);
nand_5 g10337(new_n12685, new_n12656, new_n12686);
nand_5 g10338(new_n12686, new_n12653, new_n12687);
nand_5 g10339(new_n12687, new_n12652, new_n12688);
nand_5 g10340(new_n12688, new_n12648, new_n12689);
nand_5 g10341(new_n12689, new_n12647, new_n12690);
nand_5 g10342(new_n12690, new_n12643, new_n12691);
nand_5 g10343(new_n12691, new_n12642, new_n12692);
xnor_4 g10344(new_n12692, new_n12638, n1859);
xnor_4 g10345(new_n5483, new_n5456, n1860);
not_8  g10346(new_n12169, new_n12695);
nor_5  g10347(new_n12172, new_n12695, new_n12696);
nor_5  g10348(n21915, n15182, new_n12697);
not_8  g10349(new_n7217, new_n12698);
nor_5  g10350(new_n7249, new_n12698, new_n12699);
nor_5  g10351(new_n12699, new_n12697, new_n12700);
xnor_4 g10352(n25972, new_n6526, new_n12701);
xnor_4 g10353(new_n12701, new_n12700, new_n12702_1);
not_8  g10354(new_n12702_1, new_n12703);
nand_5 g10355(new_n12703, n10250, new_n12704);
xnor_4 g10356(new_n12702_1, n10250, new_n12705);
not_8  g10357(new_n7250, new_n12706);
nand_5 g10358(new_n12706, n7674, new_n12707_1);
xnor_4 g10359(new_n7250, n7674, new_n12708);
nand_5 g10360(new_n7253_1, n6397, new_n12709);
xnor_4 g10361(new_n7252, n6397, new_n12710);
nor_5  g10362(new_n7256_1, new_n6487, new_n12711);
xnor_4 g10363(new_n7256_1, n19196, new_n12712);
not_8  g10364(new_n12712, new_n12713);
not_8  g10365(n23586, new_n12714);
nor_5  g10366(new_n7260, new_n12714, new_n12715);
nor_5  g10367(new_n7265, n21226, new_n12716);
not_8  g10368(new_n12716, new_n12717);
xnor_4 g10369(new_n7264, n21226, new_n12718);
not_8  g10370(new_n7270, new_n12719);
nor_5  g10371(new_n12719, new_n6497, new_n12720);
xnor_4 g10372(new_n7270, new_n6497, new_n12721);
not_8  g10373(new_n4300, new_n12722);
nor_5  g10374(new_n12722, n20036, new_n12723);
nor_5  g10375(new_n4313, new_n4305, new_n12724);
nor_5  g10376(new_n4317, new_n4307, new_n12725_1);
xnor_4 g10377(new_n4313, n11192, new_n12726);
nand_5 g10378(new_n12726, new_n12725_1, new_n12727_1);
not_8  g10379(new_n12727_1, new_n12728);
nor_5  g10380(new_n12728, new_n12724, new_n12729);
xnor_4 g10381(new_n4300, n20036, new_n12730);
nand_5 g10382(new_n12730, new_n12729, new_n12731);
not_8  g10383(new_n12731, new_n12732);
nor_5  g10384(new_n12732, new_n12723, new_n12733);
nand_5 g10385(new_n12733, new_n12721, new_n12734);
not_8  g10386(new_n12734, new_n12735);
nor_5  g10387(new_n12735, new_n12720, new_n12736);
nand_5 g10388(new_n12736, new_n12718, new_n12737);
nand_5 g10389(new_n12737, new_n12717, new_n12738);
xnor_4 g10390(new_n7260, n23586, new_n12739);
not_8  g10391(new_n12739, new_n12740_1);
nor_5  g10392(new_n12740_1, new_n12738, new_n12741);
nor_5  g10393(new_n12741, new_n12715, new_n12742_1);
nor_5  g10394(new_n12742_1, new_n12713, new_n12743);
nor_5  g10395(new_n12743, new_n12711, new_n12744);
not_8  g10396(new_n12744, new_n12745);
nand_5 g10397(new_n12745, new_n12710, new_n12746_1);
nand_5 g10398(new_n12746_1, new_n12709, new_n12747);
nand_5 g10399(new_n12747, new_n12708, new_n12748);
nand_5 g10400(new_n12748, new_n12707_1, new_n12749);
nand_5 g10401(new_n12749, new_n12705, new_n12750);
nand_5 g10402(new_n12750, new_n12704, new_n12751);
not_8  g10403(n25972, new_n12752);
or_5   g10404(new_n12752, new_n6526, new_n12753);
not_8  g10405(new_n12753, new_n12754);
or_5   g10406(n25972, n8614, new_n12755);
and_5  g10407(new_n12755, new_n12700, new_n12756_1);
nor_5  g10408(new_n12756_1, new_n12754, new_n12757);
not_8  g10409(new_n12757, new_n12758);
nand_5 g10410(new_n12758, new_n12751, new_n12759);
nand_5 g10411(new_n12759, new_n12696, new_n12760);
not_8  g10412(new_n12696, new_n12761);
xnor_4 g10413(new_n12759, new_n12761, new_n12762);
xnor_4 g10414(new_n12757, new_n12751, new_n12763);
not_8  g10415(new_n12763, new_n12764);
nand_5 g10416(new_n12764, new_n12173, new_n12765);
xnor_4 g10417(new_n12763, new_n12173, new_n12766);
not_8  g10418(new_n12184, new_n12767);
xnor_4 g10419(new_n12749, new_n12705, new_n12768);
nand_5 g10420(new_n12768, new_n12767, new_n12769);
xnor_4 g10421(new_n12768, new_n12184, new_n12770);
xnor_4 g10422(new_n12747, new_n12708, new_n12771);
nand_5 g10423(new_n12771, new_n12192_1, new_n12772);
not_8  g10424(new_n12192_1, new_n12773);
xnor_4 g10425(new_n12771, new_n12773, new_n12774);
xnor_4 g10426(new_n12745, new_n12710, new_n12775);
nand_5 g10427(new_n12775, new_n12197, new_n12776);
xnor_4 g10428(new_n12775, new_n12196, new_n12777);
xnor_4 g10429(new_n12742_1, new_n12713, new_n12778);
nand_5 g10430(new_n12778, new_n12203, new_n12779);
not_8  g10431(new_n12203, new_n12780);
xnor_4 g10432(new_n12778, new_n12780, new_n12781);
xnor_4 g10433(new_n12740_1, new_n12738, new_n12782);
nand_5 g10434(new_n12782, new_n12209_1, new_n12783_1);
xnor_4 g10435(new_n12782, new_n12211, new_n12784);
not_8  g10436(new_n10167, new_n12785);
xnor_4 g10437(new_n12736, new_n12718, new_n12786);
nor_5  g10438(new_n12786, new_n12785, new_n12787);
not_8  g10439(new_n12787, new_n12788);
xnor_4 g10440(new_n12786, new_n10167, new_n12789);
not_8  g10441(new_n12789, new_n12790);
not_8  g10442(new_n10170, new_n12791);
xnor_4 g10443(new_n12733, new_n12721, new_n12792);
not_8  g10444(new_n12792, new_n12793);
nor_5  g10445(new_n12793, new_n12791, new_n12794);
xnor_4 g10446(new_n12792, new_n12791, new_n12795);
not_8  g10447(new_n12795, new_n12796);
not_8  g10448(new_n10176, new_n12797);
xnor_4 g10449(new_n12730, new_n12729, new_n12798);
nor_5  g10450(new_n12798, new_n12797, new_n12799);
xnor_4 g10451(new_n12798, new_n10176, new_n12800);
not_8  g10452(new_n12800, new_n12801_1);
xnor_4 g10453(new_n12726, new_n12725_1, new_n12802);
not_8  g10454(new_n12802, new_n12803);
nor_5  g10455(new_n12803, new_n10181, new_n12804);
xnor_4 g10456(new_n4317, n9380, new_n12805);
nor_5  g10457(new_n12805, new_n7637, new_n12806);
not_8  g10458(new_n12806, new_n12807);
xnor_4 g10459(new_n12802, new_n10181, new_n12808);
not_8  g10460(new_n12808, new_n12809);
nor_5  g10461(new_n12809, new_n12807, new_n12810);
nor_5  g10462(new_n12810, new_n12804, new_n12811_1);
nor_5  g10463(new_n12811_1, new_n12801_1, new_n12812_1);
nor_5  g10464(new_n12812_1, new_n12799, new_n12813);
nor_5  g10465(new_n12813, new_n12796, new_n12814);
nor_5  g10466(new_n12814, new_n12794, new_n12815);
nor_5  g10467(new_n12815, new_n12790, new_n12816_1);
not_8  g10468(new_n12816_1, new_n12817);
nand_5 g10469(new_n12817, new_n12788, new_n12818);
nand_5 g10470(new_n12818, new_n12784, new_n12819);
nand_5 g10471(new_n12819, new_n12783_1, new_n12820);
nand_5 g10472(new_n12820, new_n12781, new_n12821_1);
nand_5 g10473(new_n12821_1, new_n12779, new_n12822);
nand_5 g10474(new_n12822, new_n12777, new_n12823);
nand_5 g10475(new_n12823, new_n12776, new_n12824);
nand_5 g10476(new_n12824, new_n12774, new_n12825);
nand_5 g10477(new_n12825, new_n12772, new_n12826);
nand_5 g10478(new_n12826, new_n12770, new_n12827);
nand_5 g10479(new_n12827, new_n12769, new_n12828);
nand_5 g10480(new_n12828, new_n12766, new_n12829);
nand_5 g10481(new_n12829, new_n12765, new_n12830);
nand_5 g10482(new_n12830, new_n12762, new_n12831);
nand_5 g10483(new_n12831, new_n12760, n1861);
nor_5  g10484(n13714, n12593, new_n12833);
nand_5 g10485(new_n12833, new_n9310, new_n12834);
nor_5  g10486(new_n12834, n8309, new_n12835);
nand_5 g10487(new_n12835, new_n9301, new_n12836);
nor_5  g10488(new_n12836, n26054, new_n12837);
xnor_4 g10489(new_n12837, n26318, new_n12838);
xnor_4 g10490(new_n12838, new_n5627, new_n12839);
xnor_4 g10491(new_n12836, new_n9296, new_n12840);
not_8  g10492(new_n12840, new_n12841);
nand_5 g10493(new_n12841, new_n5633, new_n12842);
xnor_4 g10494(new_n12835, new_n9301, new_n12843_1);
nand_5 g10495(new_n12843_1, new_n5661, new_n12844);
xnor_4 g10496(new_n12843_1, new_n5661, new_n12845);
not_8  g10497(new_n12845, new_n12846);
not_8  g10498(new_n5636, new_n12847);
xnor_4 g10499(new_n12834, new_n9306, new_n12848);
nor_5  g10500(new_n12848, new_n12847, new_n12849);
not_8  g10501(new_n5640, new_n12850);
xnor_4 g10502(new_n12833, n19144, new_n12851);
nor_5  g10503(new_n12851, new_n12850, new_n12852);
xnor_4 g10504(new_n12851, new_n5640, new_n12853);
nand_5 g10505(new_n5645, n13714, new_n12854);
xnor_4 g10506(new_n12854, n12593, new_n12855);
not_8  g10507(new_n12855, new_n12856);
nor_5  g10508(new_n12856, new_n5642, new_n12857);
not_8  g10509(n13714, new_n12858);
nor_5  g10510(new_n5645, new_n12858, new_n12859);
nand_5 g10511(new_n12859, new_n9315, new_n12860);
not_8  g10512(new_n12860, new_n12861_1);
nor_5  g10513(new_n12861_1, new_n12857, new_n12862);
nand_5 g10514(new_n12862, new_n12853, new_n12863);
not_8  g10515(new_n12863, new_n12864_1);
nor_5  g10516(new_n12864_1, new_n12852, new_n12865_1);
xnor_4 g10517(new_n12848, new_n5636, new_n12866);
not_8  g10518(new_n12866, new_n12867);
nor_5  g10519(new_n12867, new_n12865_1, new_n12868);
nor_5  g10520(new_n12868, new_n12849, new_n12869);
not_8  g10521(new_n12869, new_n12870_1);
nand_5 g10522(new_n12870_1, new_n12846, new_n12871_1);
nand_5 g10523(new_n12871_1, new_n12844, new_n12872);
xnor_4 g10524(new_n12840, new_n5633, new_n12873_1);
nand_5 g10525(new_n12873_1, new_n12872, new_n12874);
nand_5 g10526(new_n12874, new_n12842, new_n12875_1);
xnor_4 g10527(new_n12875_1, new_n12839, new_n12876);
nand_5 g10528(new_n9114, new_n7898, new_n12877);
nor_5  g10529(new_n12877, n20179, new_n12878);
xnor_4 g10530(new_n12878, n1112, new_n12879);
xnor_4 g10531(new_n12879, new_n7722, new_n12880);
xnor_4 g10532(new_n12877, new_n7895, new_n12881);
not_8  g10533(new_n12881, new_n12882);
nor_5  g10534(new_n12882, new_n7726, new_n12883);
xnor_4 g10535(new_n12882, new_n7726, new_n12884);
not_8  g10536(new_n9115, new_n12885);
nand_5 g10537(new_n12885, new_n7730, new_n12886);
xnor_4 g10538(new_n9115, new_n7730, new_n12887);
not_8  g10539(new_n7733, new_n12888);
nor_5  g10540(new_n9117, new_n12888, new_n12889);
not_8  g10541(new_n12889, new_n12890);
xnor_4 g10542(new_n9117, new_n7733, new_n12891);
nor_5  g10543(new_n9122, new_n7737, new_n12892_1);
not_8  g10544(new_n7737, new_n12893);
not_8  g10545(new_n9122, new_n12894);
nor_5  g10546(new_n12894, new_n12893, new_n12895);
not_8  g10547(new_n9126, new_n12896);
nor_5  g10548(new_n12896, new_n7741, new_n12897);
not_8  g10549(new_n12897, new_n12898);
nor_5  g10550(new_n7744, new_n9149, new_n12899);
not_8  g10551(new_n12899, new_n12900_1);
xnor_4 g10552(new_n9126, new_n7741, new_n12901);
nand_5 g10553(new_n12901, new_n12900_1, new_n12902);
nand_5 g10554(new_n12902, new_n12898, new_n12903);
nor_5  g10555(new_n12903, new_n12895, new_n12904_1);
nor_5  g10556(new_n12904_1, new_n12892_1, new_n12905);
nand_5 g10557(new_n12905, new_n12891, new_n12906);
nand_5 g10558(new_n12906, new_n12890, new_n12907);
nand_5 g10559(new_n12907, new_n12887, new_n12908);
nand_5 g10560(new_n12908, new_n12886, new_n12909);
nor_5  g10561(new_n12909, new_n12884, new_n12910);
nor_5  g10562(new_n12910, new_n12883, new_n12911);
xnor_4 g10563(new_n12911, new_n12880, new_n12912);
xnor_4 g10564(new_n12912, new_n12876, new_n12913);
xnor_4 g10565(new_n12909, new_n12884, new_n12914);
xnor_4 g10566(new_n12873_1, new_n12872, new_n12915);
not_8  g10567(new_n12915, new_n12916);
nand_5 g10568(new_n12916, new_n12914, new_n12917_1);
xnor_4 g10569(new_n12915, new_n12914, new_n12918);
xnor_4 g10570(new_n12869, new_n12845, new_n12919);
not_8  g10571(new_n12919, new_n12920);
not_8  g10572(new_n12887, new_n12921);
xnor_4 g10573(new_n12907, new_n12921, new_n12922);
nand_5 g10574(new_n12922, new_n12920, new_n12923);
xnor_4 g10575(new_n12922, new_n12919, new_n12924);
xnor_4 g10576(new_n12866, new_n12865_1, new_n12925);
not_8  g10577(new_n12925, new_n12926);
xnor_4 g10578(new_n12905, new_n12891, new_n12927);
nor_5  g10579(new_n12927, new_n12926, new_n12928);
not_8  g10580(new_n12928, new_n12929);
xnor_4 g10581(new_n12927, new_n12925, new_n12930);
xnor_4 g10582(new_n12862, new_n12853, new_n12931);
xnor_4 g10583(new_n12894, new_n7737, new_n12932);
xnor_4 g10584(new_n12932, new_n12903, new_n12933);
nor_5  g10585(new_n12933, new_n12931, new_n12934);
not_8  g10586(new_n12934, new_n12935);
not_8  g10587(new_n12931, new_n12936);
xnor_4 g10588(new_n12933, new_n12936, new_n12937);
xnor_4 g10589(new_n12901, new_n12899, new_n12938);
not_8  g10590(new_n12938, new_n12939);
xnor_4 g10591(new_n12855, new_n5642, new_n12940);
nor_5  g10592(new_n12940, new_n12939, new_n12941_1);
xnor_4 g10593(new_n7744, n18962, new_n12942_1);
xnor_4 g10594(new_n5645, new_n12858, new_n12943);
not_8  g10595(new_n12943, new_n12944);
nand_5 g10596(new_n12944, new_n12942_1, new_n12945);
not_8  g10597(new_n12945, new_n12946);
xnor_4 g10598(new_n12940, new_n12938, new_n12947);
not_8  g10599(new_n12947, new_n12948);
nor_5  g10600(new_n12948, new_n12946, new_n12949);
nor_5  g10601(new_n12949, new_n12941_1, new_n12950);
not_8  g10602(new_n12950, new_n12951);
nand_5 g10603(new_n12951, new_n12937, new_n12952);
nand_5 g10604(new_n12952, new_n12935, new_n12953);
nand_5 g10605(new_n12953, new_n12930, new_n12954);
nand_5 g10606(new_n12954, new_n12929, new_n12955);
nand_5 g10607(new_n12955, new_n12924, new_n12956_1);
nand_5 g10608(new_n12956_1, new_n12923, new_n12957);
nand_5 g10609(new_n12957, new_n12918, new_n12958);
nand_5 g10610(new_n12958, new_n12917_1, new_n12959);
xnor_4 g10611(new_n12959, new_n12913, n1891);
xnor_4 g10612(n20169, n1949, new_n12961);
nor_5  g10613(new_n4178, n8285, new_n12962);
nor_5  g10614(n9323, new_n4171, new_n12963);
not_8  g10615(n10792, new_n12964);
nor_5  g10616(new_n12964, n6729, new_n12965);
nor_5  g10617(n10792, new_n4238, new_n12966);
nand_5 g10618(new_n2574, n19922, new_n12967);
nor_5  g10619(new_n12967, new_n12966, new_n12968);
nor_5  g10620(new_n12968, new_n12965, new_n12969);
nor_5  g10621(new_n12969, new_n12963, new_n12970);
nor_5  g10622(new_n12970, new_n12962, new_n12971);
xnor_4 g10623(new_n12971, new_n12961, new_n12972);
xnor_4 g10624(new_n12972, new_n6912, new_n12973);
xnor_4 g10625(n9323, n8285, new_n12974);
xnor_4 g10626(new_n12974, new_n12969, new_n12975);
not_8  g10627(new_n12975, new_n12976);
nor_5  g10628(new_n12976, new_n6917, new_n12977);
not_8  g10629(new_n12977, new_n12978_1);
xnor_4 g10630(new_n12976, new_n6916, new_n12979);
xnor_4 g10631(n21687, n19922, new_n12980_1);
nor_5  g10632(new_n12980_1, new_n6922, new_n12981);
xnor_4 g10633(n10792, n6729, new_n12982);
xnor_4 g10634(new_n12982, new_n12967, new_n12983);
not_8  g10635(new_n12983, new_n12984);
nor_5  g10636(new_n12984, new_n12981, new_n12985_1);
xnor_4 g10637(new_n12983, new_n12981, new_n12986);
not_8  g10638(new_n12986, new_n12987_1);
nor_5  g10639(new_n12987_1, new_n6925, new_n12988);
nor_5  g10640(new_n12988, new_n12985_1, new_n12989);
not_8  g10641(new_n12989, new_n12990);
nand_5 g10642(new_n12990, new_n12979, new_n12991);
nand_5 g10643(new_n12991, new_n12978_1, new_n12992_1);
xnor_4 g10644(new_n12992_1, new_n12973, n1925);
xnor_4 g10645(new_n8079, new_n8047, n1942);
xnor_4 g10646(new_n6756, new_n6693, n1972);
not_8  g10647(new_n9337, new_n12996);
nor_5  g10648(new_n12996, new_n9273, new_n12997);
nor_5  g10649(new_n9410, new_n9339, new_n12998);
nor_5  g10650(new_n12998, new_n12997, new_n12999);
or_5   g10651(new_n9282, n22764, new_n13000);
and_5  g10652(new_n9283, n12507, new_n13001);
nor_5  g10653(new_n9283, n12507, new_n13002);
nor_5  g10654(new_n9336, new_n13002, new_n13003);
nor_5  g10655(new_n13003, new_n13001, new_n13004);
nand_5 g10656(new_n13004, new_n13000, new_n13005_1);
nor_5  g10657(new_n13005_1, new_n11903, new_n13006);
nand_5 g10658(new_n13006, new_n12999, new_n13007);
nand_5 g10659(new_n13005_1, new_n11903, new_n13008);
nor_5  g10660(new_n13008, new_n12999, new_n13009);
not_8  g10661(new_n13009, new_n13010);
nand_5 g10662(new_n13010, new_n13007, new_n13011);
nor_5  g10663(new_n13011, new_n11721, new_n13012);
xnor_4 g10664(new_n13011, new_n11720, new_n13013);
not_8  g10665(new_n13013, new_n13014);
xnor_4 g10666(new_n13005_1, new_n11840, new_n13015);
xnor_4 g10667(new_n13015, new_n12999, new_n13016);
nand_5 g10668(new_n13016, new_n11720, new_n13017);
xnor_4 g10669(new_n13016, new_n11721, new_n13018);
nand_5 g10670(new_n11767, new_n9411, new_n13019);
nand_5 g10671(new_n11773, new_n9415, new_n13020);
xnor_4 g10672(new_n11773, new_n9414, new_n13021);
nand_5 g10673(new_n11780, new_n9420, new_n13022);
xnor_4 g10674(new_n11780, new_n9419_1, new_n13023);
nand_5 g10675(new_n11784, new_n9425, new_n13024);
xnor_4 g10676(new_n11784, new_n9424, new_n13025);
nand_5 g10677(new_n11790, new_n9431, new_n13026_1);
xnor_4 g10678(new_n11789, new_n9431, new_n13027);
nand_5 g10679(new_n11796, new_n9438, new_n13028);
xnor_4 g10680(new_n11795, new_n9438, new_n13029);
nand_5 g10681(new_n11798, new_n9441, new_n13030);
xnor_4 g10682(new_n11800, new_n9441, new_n13031);
nor_5  g10683(new_n11805, new_n9450, new_n13032);
xnor_4 g10684(new_n11805, new_n9446, new_n13033);
not_8  g10685(new_n13033, new_n13034);
nor_5  g10686(new_n11807, new_n9454, new_n13035);
nor_5  g10687(new_n13035, new_n11811, new_n13036);
not_8  g10688(new_n13036, new_n13037);
xnor_4 g10689(new_n13035, new_n11810, new_n13038);
nand_5 g10690(new_n13038, new_n9461, new_n13039);
nand_5 g10691(new_n13039, new_n13037, new_n13040);
not_8  g10692(new_n13040, new_n13041);
nor_5  g10693(new_n13041, new_n13034, new_n13042);
nor_5  g10694(new_n13042, new_n13032, new_n13043_1);
not_8  g10695(new_n13043_1, new_n13044_1);
nand_5 g10696(new_n13044_1, new_n13031, new_n13045);
nand_5 g10697(new_n13045, new_n13030, new_n13046);
nand_5 g10698(new_n13046, new_n13029, new_n13047);
nand_5 g10699(new_n13047, new_n13028, new_n13048_1);
nand_5 g10700(new_n13048_1, new_n13027, new_n13049);
nand_5 g10701(new_n13049, new_n13026_1, new_n13050);
nand_5 g10702(new_n13050, new_n13025, new_n13051);
nand_5 g10703(new_n13051, new_n13024, new_n13052);
nand_5 g10704(new_n13052, new_n13023, new_n13053);
nand_5 g10705(new_n13053, new_n13022, new_n13054_1);
nand_5 g10706(new_n13054_1, new_n13021, new_n13055);
nand_5 g10707(new_n13055, new_n13020, new_n13056);
not_8  g10708(new_n9411, new_n13057);
xnor_4 g10709(new_n11767, new_n13057, new_n13058);
nand_5 g10710(new_n13058, new_n13056, new_n13059);
nand_5 g10711(new_n13059, new_n13019, new_n13060);
nand_5 g10712(new_n13060, new_n13018, new_n13061);
nand_5 g10713(new_n13061, new_n13017, new_n13062);
nor_5  g10714(new_n13062, new_n13014, new_n13063);
nor_5  g10715(new_n13063, new_n13012, n1981);
xnor_4 g10716(new_n13058, new_n13056, n2004);
not_8  g10717(n5140, new_n13066);
or_5   g10718(n6105, new_n13066, new_n13067);
xnor_4 g10719(n6105, n5140, new_n13068);
not_8  g10720(n6204, new_n13069);
or_5   g10721(new_n13069, n3795, new_n13070);
xnor_4 g10722(n6204, n3795, new_n13071);
not_8  g10723(n3349, new_n13072);
or_5   g10724(n25464, new_n13072, new_n13073);
xnor_4 g10725(n25464, n3349, new_n13074_1);
or_5   g10726(n4590, new_n6805, new_n13075);
xnor_4 g10727(n4590, n1742, new_n13076);
or_5   g10728(n26752, new_n6815, new_n13077);
xnor_4 g10729(n26752, n4858, new_n13078);
nor_5  g10730(new_n6821, n6513, new_n13079);
xnor_4 g10731(n8244, n6513, new_n13080);
not_8  g10732(new_n13080, new_n13081);
nor_5  g10733(new_n6826_1, n3918, new_n13082_1);
xnor_4 g10734(n9493, n3918, new_n13083);
nor_5  g10735(n15167, new_n4327, new_n13084);
nor_5  g10736(new_n6831, n919, new_n13085);
not_8  g10737(n25316, new_n13086);
nor_5  g10738(new_n13086, n21095, new_n13087);
nor_5  g10739(n25316, new_n6836, new_n13088);
nor_5  g10740(new_n4342, n8656, new_n13089);
not_8  g10741(new_n13089, new_n13090);
nor_5  g10742(new_n13090, new_n13088, new_n13091);
nor_5  g10743(new_n13091, new_n13087, new_n13092);
nor_5  g10744(new_n13092, new_n13085, new_n13093);
nor_5  g10745(new_n13093, new_n13084, new_n13094);
nand_5 g10746(new_n13094, new_n13083, new_n13095);
not_8  g10747(new_n13095, new_n13096_1);
nor_5  g10748(new_n13096_1, new_n13082_1, new_n13097);
nor_5  g10749(new_n13097, new_n13081, new_n13098);
nor_5  g10750(new_n13098, new_n13079, new_n13099);
not_8  g10751(new_n13099, new_n13100);
nand_5 g10752(new_n13100, new_n13078, new_n13101);
nand_5 g10753(new_n13101, new_n13077, new_n13102);
nand_5 g10754(new_n13102, new_n13076, new_n13103);
nand_5 g10755(new_n13103, new_n13075, new_n13104);
nand_5 g10756(new_n13104, new_n13074_1, new_n13105);
nand_5 g10757(new_n13105, new_n13073, new_n13106);
nand_5 g10758(new_n13106, new_n13071, new_n13107);
nand_5 g10759(new_n13107, new_n13070, new_n13108);
nand_5 g10760(new_n13108, new_n13068, new_n13109);
nand_5 g10761(new_n13109, new_n13067, new_n13110_1);
not_8  g10762(new_n6525, new_n13111);
nor_5  g10763(new_n6533, n10018, new_n13112);
nand_5 g10764(new_n6533, n10018, new_n13113);
not_8  g10765(n2184, new_n13114);
nand_5 g10766(new_n6540, new_n13114, new_n13115);
xnor_4 g10767(new_n6540, n2184, new_n13116_1);
not_8  g10768(n3541, new_n13117);
nand_5 g10769(new_n6546, new_n13117, new_n13118);
xnor_4 g10770(new_n6546, n3541, new_n13119);
not_8  g10771(n16818, new_n13120);
nand_5 g10772(new_n6552, new_n13120, new_n13121);
xnor_4 g10773(new_n6552, n16818, new_n13122_1);
not_8  g10774(new_n4183, new_n13123);
nand_5 g10775(new_n13123, new_n6816, new_n13124);
xnor_4 g10776(new_n4183, new_n6816, new_n13125);
nor_5  g10777(new_n4187, n14576, new_n13126);
xnor_4 g10778(new_n4186_1, n14576, new_n13127);
not_8  g10779(new_n13127, new_n13128);
nor_5  g10780(new_n4191, new_n6827, new_n13129);
not_8  g10781(new_n13129, new_n13130);
xnor_4 g10782(new_n4191, n2985, new_n13131);
nor_5  g10783(new_n12286, n5605, new_n13132);
nand_5 g10784(new_n4202, n15652, new_n13133);
nor_5  g10785(n19922, new_n6880, new_n13134);
xnor_4 g10786(new_n4202, n15652, new_n13135);
not_8  g10787(new_n13135, new_n13136);
nand_5 g10788(new_n13136, new_n13134, new_n13137_1);
nand_5 g10789(new_n13137_1, new_n13133, new_n13138);
xnor_4 g10790(new_n4196, n5605, new_n13139);
not_8  g10791(new_n13139, new_n13140);
nor_5  g10792(new_n13140, new_n13138, new_n13141_1);
nor_5  g10793(new_n13141_1, new_n13132, new_n13142);
nand_5 g10794(new_n13142, new_n13131, new_n13143);
nand_5 g10795(new_n13143, new_n13130, new_n13144_1);
nor_5  g10796(new_n13144_1, new_n13128, new_n13145);
nor_5  g10797(new_n13145, new_n13126, new_n13146);
not_8  g10798(new_n13146, new_n13147);
nand_5 g10799(new_n13147, new_n13125, new_n13148);
nand_5 g10800(new_n13148, new_n13124, new_n13149);
nand_5 g10801(new_n13149, new_n13122_1, new_n13150);
nand_5 g10802(new_n13150, new_n13121, new_n13151);
nand_5 g10803(new_n13151, new_n13119, new_n13152);
nand_5 g10804(new_n13152, new_n13118, new_n13153);
nand_5 g10805(new_n13153, new_n13116_1, new_n13154);
nand_5 g10806(new_n13154, new_n13115, new_n13155);
nand_5 g10807(new_n13155, new_n13113, new_n13156);
xnor_4 g10808(new_n13156, new_n6535, new_n13157);
nor_5  g10809(new_n13157, new_n13112, new_n13158);
xnor_4 g10810(new_n13158, new_n13111, new_n13159);
not_8  g10811(n10018, new_n13160);
xnor_4 g10812(new_n6533, new_n13160, new_n13161);
xnor_4 g10813(new_n13161, new_n13155, new_n13162);
nand_5 g10814(new_n13162, new_n6575, new_n13163);
xnor_4 g10815(new_n13162, new_n6574, new_n13164);
xnor_4 g10816(new_n13153, new_n13116_1, new_n13165);
nand_5 g10817(new_n13165, new_n6582, new_n13166);
xnor_4 g10818(new_n13165, new_n6581, new_n13167);
xnor_4 g10819(new_n13151, new_n13119, new_n13168_1);
nand_5 g10820(new_n13168_1, new_n6587_1, new_n13169);
not_8  g10821(new_n6587_1, new_n13170);
xnor_4 g10822(new_n13168_1, new_n13170, new_n13171);
xnor_4 g10823(new_n13149, new_n13122_1, new_n13172);
nand_5 g10824(new_n13172, new_n6590_1, new_n13173);
xnor_4 g10825(new_n13147, new_n13125, new_n13174);
nand_5 g10826(new_n13174, new_n6593, new_n13175);
xnor_4 g10827(new_n13174, new_n6595, new_n13176);
xnor_4 g10828(new_n13144_1, new_n13127, new_n13177);
not_8  g10829(new_n13177, new_n13178);
nand_5 g10830(new_n13178, new_n6597, new_n13179);
xnor_4 g10831(new_n13177, new_n6597, new_n13180);
xnor_4 g10832(new_n13142, new_n13131, new_n13181);
nor_5  g10833(new_n13181, new_n6599, new_n13182);
not_8  g10834(new_n13182, new_n13183);
xnor_4 g10835(new_n13139, new_n13138, new_n13184);
not_8  g10836(new_n13184, new_n13185);
nor_5  g10837(new_n13185, new_n6601, new_n13186);
xnor_4 g10838(new_n13184, new_n6601, new_n13187);
not_8  g10839(new_n13187, new_n13188);
xnor_4 g10840(new_n13135, new_n13134, new_n13189);
nor_5  g10841(new_n13189, new_n6605, new_n13190_1);
xnor_4 g10842(n19922, n4939, new_n13191);
nor_5  g10843(new_n13191, new_n6609, new_n13192);
xnor_4 g10844(new_n13189, new_n6606, new_n13193);
nand_5 g10845(new_n13193, new_n13192, new_n13194);
not_8  g10846(new_n13194, new_n13195);
nor_5  g10847(new_n13195, new_n13190_1, new_n13196);
nor_5  g10848(new_n13196, new_n13188, new_n13197);
nor_5  g10849(new_n13197, new_n13186, new_n13198_1);
xnor_4 g10850(new_n13181, new_n6598, new_n13199_1);
nand_5 g10851(new_n13199_1, new_n13198_1, new_n13200);
nand_5 g10852(new_n13200, new_n13183, new_n13201);
nand_5 g10853(new_n13201, new_n13180, new_n13202);
nand_5 g10854(new_n13202, new_n13179, new_n13203);
nand_5 g10855(new_n13203, new_n13176, new_n13204_1);
nand_5 g10856(new_n13204_1, new_n13175, new_n13205);
not_8  g10857(new_n6590_1, new_n13206);
xnor_4 g10858(new_n13172, new_n13206, new_n13207);
nand_5 g10859(new_n13207, new_n13205, new_n13208);
nand_5 g10860(new_n13208, new_n13173, new_n13209_1);
nand_5 g10861(new_n13209_1, new_n13171, new_n13210);
nand_5 g10862(new_n13210, new_n13169, new_n13211);
nand_5 g10863(new_n13211, new_n13167, new_n13212);
nand_5 g10864(new_n13212, new_n13166, new_n13213);
nand_5 g10865(new_n13213, new_n13164, new_n13214);
nand_5 g10866(new_n13214, new_n13163, new_n13215);
xnor_4 g10867(new_n13215, new_n13159, new_n13216);
not_8  g10868(new_n13216, new_n13217);
nand_5 g10869(new_n13217, new_n13110_1, new_n13218);
xnor_4 g10870(new_n13216, new_n13110_1, new_n13219);
xnor_4 g10871(new_n13108, new_n13068, new_n13220);
xnor_4 g10872(new_n13213, new_n13164, new_n13221);
not_8  g10873(new_n13221, new_n13222);
nand_5 g10874(new_n13222, new_n13220, new_n13223);
xnor_4 g10875(new_n13221, new_n13220, new_n13224);
xnor_4 g10876(new_n13106, new_n13071, new_n13225);
xnor_4 g10877(new_n13211, new_n13167, new_n13226);
not_8  g10878(new_n13226, new_n13227);
nand_5 g10879(new_n13227, new_n13225, new_n13228);
xnor_4 g10880(new_n13226, new_n13225, new_n13229);
xnor_4 g10881(new_n13104, new_n13074_1, new_n13230);
xnor_4 g10882(new_n13209_1, new_n13171, new_n13231);
not_8  g10883(new_n13231, new_n13232);
nand_5 g10884(new_n13232, new_n13230, new_n13233);
xnor_4 g10885(new_n13231, new_n13230, new_n13234);
xnor_4 g10886(new_n13102, new_n13076, new_n13235);
not_8  g10887(new_n13207, new_n13236);
xnor_4 g10888(new_n13236, new_n13205, new_n13237);
nand_5 g10889(new_n13237, new_n13235, new_n13238);
not_8  g10890(new_n13235, new_n13239);
xnor_4 g10891(new_n13237, new_n13239, new_n13240);
xnor_4 g10892(new_n13099, new_n13078, new_n13241);
not_8  g10893(new_n13241, new_n13242);
not_8  g10894(new_n13176, new_n13243);
xnor_4 g10895(new_n13203, new_n13243, new_n13244);
nand_5 g10896(new_n13244, new_n13242, new_n13245);
xnor_4 g10897(new_n13244, new_n13241, new_n13246);
xnor_4 g10898(new_n13097, new_n13080, new_n13247);
not_8  g10899(new_n13247, new_n13248);
not_8  g10900(new_n13180, new_n13249);
xnor_4 g10901(new_n13201, new_n13249, new_n13250);
nand_5 g10902(new_n13250, new_n13248, new_n13251);
xnor_4 g10903(new_n13250, new_n13247, new_n13252);
xnor_4 g10904(new_n13094, new_n13083, new_n13253);
not_8  g10905(new_n13199_1, new_n13254);
xnor_4 g10906(new_n13254, new_n13198_1, new_n13255);
nand_5 g10907(new_n13255, new_n13253, new_n13256);
not_8  g10908(new_n13253, new_n13257);
xnor_4 g10909(new_n13255, new_n13257, new_n13258);
xnor_4 g10910(new_n13196, new_n13187, new_n13259);
xnor_4 g10911(n15167, n919, new_n13260);
xnor_4 g10912(new_n13260, new_n13092, new_n13261);
not_8  g10913(new_n13261, new_n13262);
nor_5  g10914(new_n13262, new_n13259, new_n13263_1);
not_8  g10915(new_n13263_1, new_n13264);
xnor_4 g10916(new_n13261, new_n13259, new_n13265);
xnor_4 g10917(new_n13191, new_n6608, new_n13266);
not_8  g10918(new_n13266, new_n13267);
xnor_4 g10919(n20385, n8656, new_n13268);
nor_5  g10920(new_n13268, new_n13267, new_n13269);
xnor_4 g10921(n25316, n21095, new_n13270_1);
xnor_4 g10922(new_n13270_1, new_n13090, new_n13271);
not_8  g10923(new_n13271, new_n13272);
nor_5  g10924(new_n13272, new_n13269, new_n13273_1);
not_8  g10925(new_n13273_1, new_n13274);
xnor_4 g10926(new_n13193, new_n13192, new_n13275);
xnor_4 g10927(new_n13271, new_n13269, new_n13276);
nand_5 g10928(new_n13276, new_n13275, new_n13277);
nand_5 g10929(new_n13277, new_n13274, new_n13278);
nand_5 g10930(new_n13278, new_n13265, new_n13279);
nand_5 g10931(new_n13279, new_n13264, new_n13280);
nand_5 g10932(new_n13280, new_n13258, new_n13281);
nand_5 g10933(new_n13281, new_n13256, new_n13282);
nand_5 g10934(new_n13282, new_n13252, new_n13283);
nand_5 g10935(new_n13283, new_n13251, new_n13284);
nand_5 g10936(new_n13284, new_n13246, new_n13285_1);
nand_5 g10937(new_n13285_1, new_n13245, new_n13286);
nand_5 g10938(new_n13286, new_n13240, new_n13287);
nand_5 g10939(new_n13287, new_n13238, new_n13288);
nand_5 g10940(new_n13288, new_n13234, new_n13289);
nand_5 g10941(new_n13289, new_n13233, new_n13290);
nand_5 g10942(new_n13290, new_n13229, new_n13291);
nand_5 g10943(new_n13291, new_n13228, new_n13292);
nand_5 g10944(new_n13292, new_n13224, new_n13293);
nand_5 g10945(new_n13293, new_n13223, new_n13294);
nand_5 g10946(new_n13294, new_n13219, new_n13295);
nand_5 g10947(new_n13295, new_n13218, new_n13296);
nor_5  g10948(new_n13158, new_n6525, new_n13297);
not_8  g10949(new_n13156, new_n13298);
nand_5 g10950(new_n13298, new_n6535, new_n13299);
nand_5 g10951(new_n13158, new_n6525, new_n13300);
not_8  g10952(new_n13215, new_n13301);
nand_5 g10953(new_n13301, new_n13300, new_n13302);
nand_5 g10954(new_n13302, new_n13299, new_n13303);
nor_5  g10955(new_n13303, new_n13297, new_n13304);
nand_5 g10956(new_n13304, new_n13296, new_n13305);
not_8  g10957(new_n13305, n2007);
xnor_4 g10958(new_n9464, new_n9451_1, n2061);
xnor_4 g10959(new_n12030, new_n7546, new_n13308);
nand_5 g10960(new_n12036, new_n7552, new_n13309);
xnor_4 g10961(new_n12036, new_n7551, new_n13310);
nand_5 g10962(new_n12042, new_n7557, new_n13311);
not_8  g10963(new_n4875, new_n13312);
nand_5 g10964(new_n7563, new_n13312, new_n13313);
xnor_4 g10965(new_n7563, new_n4875, new_n13314);
nand_5 g10966(new_n7568, new_n4907, new_n13315);
xnor_4 g10967(new_n7567, new_n4907, new_n13316);
nor_5  g10968(new_n7572_1, new_n4914, new_n13317);
not_8  g10969(new_n13317, new_n13318);
nor_5  g10970(new_n7578, new_n4922, new_n13319_1);
not_8  g10971(new_n13319_1, new_n13320);
xnor_4 g10972(new_n7577, new_n4922, new_n13321);
not_8  g10973(new_n4930, new_n13322);
nor_5  g10974(new_n7585_1, new_n4934, new_n13323);
and_5  g10975(new_n13323, new_n13322, new_n13324);
xnor_4 g10976(new_n13323, new_n4930, new_n13325);
and_5  g10977(new_n13325, new_n7592, new_n13326);
nor_5  g10978(new_n13326, new_n13324, new_n13327);
nand_5 g10979(new_n13327, new_n13321, new_n13328);
nand_5 g10980(new_n13328, new_n13320, new_n13329);
xnor_4 g10981(new_n7571, new_n4914, new_n13330);
nand_5 g10982(new_n13330, new_n13329, new_n13331);
nand_5 g10983(new_n13331, new_n13318, new_n13332);
nand_5 g10984(new_n13332, new_n13316, new_n13333_1);
nand_5 g10985(new_n13333_1, new_n13315, new_n13334);
nand_5 g10986(new_n13334, new_n13314, new_n13335);
nand_5 g10987(new_n13335, new_n13313, new_n13336);
xnor_4 g10988(new_n12042, new_n7556, new_n13337);
nand_5 g10989(new_n13337, new_n13336, new_n13338_1);
nand_5 g10990(new_n13338_1, new_n13311, new_n13339);
nand_5 g10991(new_n13339, new_n13310, new_n13340);
nand_5 g10992(new_n13340, new_n13309, new_n13341);
xnor_4 g10993(new_n13341, new_n13308, n2092);
not_8  g10994(n10650, new_n13343);
xnor_4 g10995(n22253, new_n13343, new_n13344);
not_8  g10996(new_n13344, new_n13345);
or_5   g10997(n12900, n1255, new_n13346);
not_8  g10998(n1255, new_n13347);
xnor_4 g10999(n12900, new_n13347, new_n13348);
or_5   g11000(n20411, n9512, new_n13349);
not_8  g11001(n9512, new_n13350);
xnor_4 g11002(n20411, new_n13350, new_n13351);
nor_5  g11003(n17069, n16608, new_n13352);
not_8  g11004(new_n13352, new_n13353);
xnor_4 g11005(n17069, new_n7412, new_n13354);
nor_5  g11006(n21735, n15918, new_n13355);
not_8  g11007(new_n13355, new_n13356);
not_8  g11008(n15918, new_n13357);
xnor_4 g11009(n21735, new_n13357, new_n13358);
nor_5  g11010(n24085, n17784, new_n13359);
not_8  g11011(new_n13359, new_n13360);
not_8  g11012(n17784, new_n13361);
xnor_4 g11013(n24085, new_n13361, new_n13362);
nor_5  g11014(n14323, n14071, new_n13363);
xnor_4 g11015(n14323, new_n4826, new_n13364);
not_8  g11016(new_n13364, new_n13365);
nor_5  g11017(n2886, n1738, new_n13366);
xnor_4 g11018(n2886, new_n4831, new_n13367_1);
not_8  g11019(new_n13367_1, new_n13368);
nor_5  g11020(n12152, n1040, new_n13369);
nand_5 g11021(n19107, n9090, new_n13370);
not_8  g11022(new_n13370, new_n13371);
not_8  g11023(n1040, new_n13372);
xnor_4 g11024(n12152, new_n13372, new_n13373);
not_8  g11025(new_n13373, new_n13374);
nor_5  g11026(new_n13374, new_n13371, new_n13375);
nor_5  g11027(new_n13375, new_n13369, new_n13376);
nor_5  g11028(new_n13376, new_n13368, new_n13377);
nor_5  g11029(new_n13377, new_n13366, new_n13378);
nor_5  g11030(new_n13378, new_n13365, new_n13379);
nor_5  g11031(new_n13379, new_n13363, new_n13380);
not_8  g11032(new_n13380, new_n13381);
nand_5 g11033(new_n13381, new_n13362, new_n13382);
nand_5 g11034(new_n13382, new_n13360, new_n13383);
nand_5 g11035(new_n13383, new_n13358, new_n13384);
nand_5 g11036(new_n13384, new_n13356, new_n13385);
nand_5 g11037(new_n13385, new_n13354, new_n13386);
nand_5 g11038(new_n13386, new_n13353, new_n13387);
nand_5 g11039(new_n13387, new_n13351, new_n13388);
nand_5 g11040(new_n13388, new_n13349, new_n13389);
nand_5 g11041(new_n13389, new_n13348, new_n13390);
nand_5 g11042(new_n13390, new_n13346, new_n13391);
xnor_4 g11043(new_n13391, new_n13345, new_n13392);
nand_5 g11044(new_n13392, n2272, new_n13393);
xnor_4 g11045(new_n13392, new_n7613, new_n13394);
not_8  g11046(new_n13348, new_n13395);
xnor_4 g11047(new_n13389, new_n13395, new_n13396);
nand_5 g11048(new_n13396, n25331, new_n13397);
xnor_4 g11049(new_n13396, new_n7359, new_n13398);
not_8  g11050(new_n13351, new_n13399);
xnor_4 g11051(new_n13387, new_n13399, new_n13400);
nand_5 g11052(new_n13400, n18483, new_n13401);
xnor_4 g11053(new_n13400, new_n7362, new_n13402);
not_8  g11054(new_n13354, new_n13403);
xnor_4 g11055(new_n13385, new_n13403, new_n13404);
nand_5 g11056(new_n13404, n21934, new_n13405);
xnor_4 g11057(new_n13404, new_n7365, new_n13406);
not_8  g11058(new_n13358, new_n13407_1);
xnor_4 g11059(new_n13383, new_n13407_1, new_n13408);
nand_5 g11060(new_n13408, n18901, new_n13409_1);
xnor_4 g11061(new_n13408, new_n7368, new_n13410);
xnor_4 g11062(new_n13380, new_n13362, new_n13411);
nand_5 g11063(new_n13411, n4376, new_n13412);
xnor_4 g11064(new_n13411, new_n7371, new_n13413);
xnor_4 g11065(new_n13378, new_n13364, new_n13414);
nand_5 g11066(new_n13414, n14570, new_n13415);
xnor_4 g11067(new_n13414, new_n7375, new_n13416);
xnor_4 g11068(new_n13376, new_n13367_1, new_n13417);
nand_5 g11069(new_n13417, n23775, new_n13418);
xnor_4 g11070(new_n13417, new_n7379, new_n13419_1);
xnor_4 g11071(n19107, n9090, new_n13420);
nand_5 g11072(new_n13420, n11479, new_n13421);
nand_5 g11073(new_n13421, new_n7382, new_n13422);
not_8  g11074(new_n13422, new_n13423);
xnor_4 g11075(new_n13373, new_n13371, new_n13424_1);
xnor_4 g11076(new_n13421, n8259, new_n13425);
not_8  g11077(new_n13425, new_n13426);
nor_5  g11078(new_n13426, new_n13424_1, new_n13427);
nor_5  g11079(new_n13427, new_n13423, new_n13428);
nand_5 g11080(new_n13428, new_n13419_1, new_n13429);
nand_5 g11081(new_n13429, new_n13418, new_n13430);
nand_5 g11082(new_n13430, new_n13416, new_n13431);
nand_5 g11083(new_n13431, new_n13415, new_n13432);
nand_5 g11084(new_n13432, new_n13413, new_n13433);
nand_5 g11085(new_n13433, new_n13412, new_n13434);
nand_5 g11086(new_n13434, new_n13410, new_n13435);
nand_5 g11087(new_n13435, new_n13409_1, new_n13436);
nand_5 g11088(new_n13436, new_n13406, new_n13437);
nand_5 g11089(new_n13437, new_n13405, new_n13438);
nand_5 g11090(new_n13438, new_n13402, new_n13439);
nand_5 g11091(new_n13439, new_n13401, new_n13440);
nand_5 g11092(new_n13440, new_n13398, new_n13441);
nand_5 g11093(new_n13441, new_n13397, new_n13442);
nand_5 g11094(new_n13442, new_n13394, new_n13443);
nand_5 g11095(new_n13443, new_n13393, new_n13444);
or_5   g11096(n22253, n10650, new_n13445);
nand_5 g11097(new_n13391, new_n13344, new_n13446);
nand_5 g11098(new_n13446, new_n13445, new_n13447);
nand_5 g11099(new_n13447, new_n13444, new_n13448);
not_8  g11100(n9934, new_n13449);
nor_5  g11101(n7876, n4964, new_n13450);
nand_5 g11102(new_n13450, new_n3904, new_n13451);
nor_5  g11103(new_n13451, n342, new_n13452);
nand_5 g11104(new_n13452, new_n3894, new_n13453_1);
nor_5  g11105(new_n13453_1, n22597, new_n13454);
nand_5 g11106(new_n13454, new_n3878, new_n13455);
nor_5  g11107(new_n13455, n26224, new_n13456_1);
and_5  g11108(new_n13456_1, new_n12518, new_n13457_1);
and_5  g11109(new_n13457_1, new_n13449, new_n13458);
xnor_4 g11110(new_n13457_1, n9934, new_n13459);
nor_5  g11111(n18409, n5704, new_n13460_1);
nand_5 g11112(new_n13460_1, new_n2390, new_n13461);
nor_5  g11113(new_n13461, n19911, new_n13462);
nand_5 g11114(new_n13462, new_n2406, new_n13463);
nor_5  g11115(new_n13463, n18907, new_n13464);
nand_5 g11116(new_n13464, new_n7695, new_n13465);
nor_5  g11117(new_n13465, n4256, new_n13466);
xnor_4 g11118(new_n13466, n21287, new_n13467);
not_8  g11119(new_n13467, new_n13468);
nand_5 g11120(new_n13468, new_n7450, new_n13469);
xnor_4 g11121(new_n13467, new_n7450, new_n13470);
xnor_4 g11122(new_n13465, new_n7692_1, new_n13471);
not_8  g11123(new_n13471, new_n13472);
nand_5 g11124(new_n13472, new_n7454, new_n13473);
xnor_4 g11125(new_n13471, new_n7454, new_n13474);
xnor_4 g11126(new_n13464, n22332, new_n13475);
not_8  g11127(new_n13475, new_n13476);
nand_5 g11128(new_n13476, new_n7457, new_n13477_1);
xnor_4 g11129(new_n13475, new_n7457, new_n13478);
xnor_4 g11130(new_n13463, new_n2415, new_n13479);
not_8  g11131(new_n13479, new_n13480);
nand_5 g11132(new_n13480, new_n5385, new_n13481);
xnor_4 g11133(new_n13479, new_n5385, new_n13482);
not_8  g11134(n16158, new_n13483);
xnor_4 g11135(new_n13462, n2731, new_n13484_1);
not_8  g11136(new_n13484_1, new_n13485);
nand_5 g11137(new_n13485, new_n13483, new_n13486_1);
xnor_4 g11138(new_n13484_1, new_n13483, new_n13487_1);
not_8  g11139(n5752, new_n13488);
xnor_4 g11140(new_n13461, new_n3969, new_n13489);
not_8  g11141(new_n13489, new_n13490_1);
nand_5 g11142(new_n13490_1, new_n13488, new_n13491);
xnor_4 g11143(new_n13460_1, n13708, new_n13492);
not_8  g11144(new_n13492, new_n13493);
nand_5 g11145(new_n13493, new_n4829, new_n13494_1);
xnor_4 g11146(new_n13492, new_n4829, new_n13495);
xnor_4 g11147(n18409, n5704, new_n13496);
nand_5 g11148(new_n13496, new_n4833, new_n13497);
nand_5 g11149(n22309, n5704, new_n13498);
xnor_4 g11150(new_n13496, n25073, new_n13499);
nand_5 g11151(new_n13499, new_n13498, new_n13500_1);
nand_5 g11152(new_n13500_1, new_n13497, new_n13501_1);
nand_5 g11153(new_n13501_1, new_n13495, new_n13502);
nand_5 g11154(new_n13502, new_n13494_1, new_n13503);
xnor_4 g11155(new_n13489, new_n13488, new_n13504);
nand_5 g11156(new_n13504, new_n13503, new_n13505);
nand_5 g11157(new_n13505, new_n13491, new_n13506_1);
nand_5 g11158(new_n13506_1, new_n13487_1, new_n13507);
nand_5 g11159(new_n13507, new_n13486_1, new_n13508);
nand_5 g11160(new_n13508, new_n13482, new_n13509);
nand_5 g11161(new_n13509, new_n13481, new_n13510);
nand_5 g11162(new_n13510, new_n13478, new_n13511);
nand_5 g11163(new_n13511, new_n13477_1, new_n13512);
nand_5 g11164(new_n13512, new_n13474, new_n13513);
nand_5 g11165(new_n13513, new_n13473, new_n13514);
nand_5 g11166(new_n13514, new_n13470, new_n13515);
nand_5 g11167(new_n13515, new_n13469, new_n13516);
nand_5 g11168(new_n13466, new_n7689, new_n13517);
xnor_4 g11169(new_n13517, new_n7686_1, new_n13518);
xnor_4 g11170(new_n13518, new_n7533, new_n13519);
xnor_4 g11171(new_n13519, new_n13516, new_n13520);
nand_5 g11172(new_n13520, new_n13459, new_n13521);
not_8  g11173(new_n13520, new_n13522);
xnor_4 g11174(new_n13522, new_n13459, new_n13523);
xnor_4 g11175(new_n13456_1, n18496, new_n13524);
xnor_4 g11176(new_n13514, new_n13470, new_n13525);
nand_5 g11177(new_n13525, new_n13524, new_n13526);
not_8  g11178(new_n13525, new_n13527);
xnor_4 g11179(new_n13527, new_n13524, new_n13528);
not_8  g11180(n26224, new_n13529);
xnor_4 g11181(new_n13455, new_n13529, new_n13530);
xnor_4 g11182(new_n13512, new_n13474, new_n13531);
nand_5 g11183(new_n13531, new_n13530, new_n13532);
not_8  g11184(new_n13531, new_n13533);
xnor_4 g11185(new_n13533, new_n13530, new_n13534);
xnor_4 g11186(new_n13454, n19327, new_n13535);
xnor_4 g11187(new_n13510, new_n13478, new_n13536);
nand_5 g11188(new_n13536, new_n13535, new_n13537);
not_8  g11189(new_n13536, new_n13538);
xnor_4 g11190(new_n13538, new_n13535, new_n13539);
xnor_4 g11191(new_n13453_1, new_n3888, new_n13540);
xnor_4 g11192(new_n13508, new_n13482, new_n13541);
nand_5 g11193(new_n13541, new_n13540, new_n13542);
not_8  g11194(new_n13541, new_n13543);
xnor_4 g11195(new_n13543, new_n13540, new_n13544);
xnor_4 g11196(new_n13452, n26107, new_n13545);
xnor_4 g11197(new_n13506_1, new_n13487_1, new_n13546);
nand_5 g11198(new_n13546, new_n13545, new_n13547);
not_8  g11199(new_n13546, new_n13548_1);
xnor_4 g11200(new_n13548_1, new_n13545, new_n13549_1);
xnor_4 g11201(new_n13451, new_n3899, new_n13550);
xnor_4 g11202(new_n13504, new_n13503, new_n13551_1);
nand_5 g11203(new_n13551_1, new_n13550, new_n13552);
not_8  g11204(new_n13551_1, new_n13553);
xnor_4 g11205(new_n13553, new_n13550, new_n13554);
xnor_4 g11206(new_n13501_1, new_n13495, new_n13555);
xnor_4 g11207(new_n13450, n26553, new_n13556);
nand_5 g11208(new_n13556, new_n13555, new_n13557);
xnor_4 g11209(new_n13556, new_n13555, new_n13558);
not_8  g11210(new_n13558, new_n13559);
xnor_4 g11211(n7876, new_n3909_1, new_n13560);
not_8  g11212(new_n13560, new_n13561);
xnor_4 g11213(new_n13499, new_n13498, new_n13562);
not_8  g11214(new_n13562, new_n13563);
nor_5  g11215(new_n13563, new_n13561, new_n13564);
not_8  g11216(new_n13564, new_n13565);
not_8  g11217(n5704, new_n13566);
xnor_4 g11218(n22309, new_n13566, new_n13567);
not_8  g11219(new_n13567, new_n13568);
nor_5  g11220(new_n13568, new_n3946, new_n13569);
xnor_4 g11221(new_n13562, new_n13561, new_n13570);
nand_5 g11222(new_n13570, new_n13569, new_n13571);
nand_5 g11223(new_n13571, new_n13565, new_n13572);
nand_5 g11224(new_n13572, new_n13559, new_n13573);
nand_5 g11225(new_n13573, new_n13557, new_n13574);
nand_5 g11226(new_n13574, new_n13554, new_n13575);
nand_5 g11227(new_n13575, new_n13552, new_n13576);
nand_5 g11228(new_n13576, new_n13549_1, new_n13577);
nand_5 g11229(new_n13577, new_n13547, new_n13578);
nand_5 g11230(new_n13578, new_n13544, new_n13579);
nand_5 g11231(new_n13579, new_n13542, new_n13580);
nand_5 g11232(new_n13580, new_n13539, new_n13581);
nand_5 g11233(new_n13581, new_n13537, new_n13582);
nand_5 g11234(new_n13582, new_n13534, new_n13583);
nand_5 g11235(new_n13583, new_n13532, new_n13584);
nand_5 g11236(new_n13584, new_n13528, new_n13585);
nand_5 g11237(new_n13585, new_n13526, new_n13586);
nand_5 g11238(new_n13586, new_n13523, new_n13587);
nand_5 g11239(new_n13587, new_n13521, new_n13588);
nor_5  g11240(new_n13588, new_n13458, new_n13589);
or_5   g11241(new_n13517, n26986, new_n13590);
or_5   g11242(new_n13518, n8305, new_n13591);
nand_5 g11243(new_n13518, n8305, new_n13592);
nand_5 g11244(new_n13592, new_n13516, new_n13593);
nand_5 g11245(new_n13593, new_n13591, new_n13594);
nand_5 g11246(new_n13594, new_n13590, new_n13595);
nand_5 g11247(new_n13595, new_n13589, new_n13596);
xnor_4 g11248(new_n13596, new_n13448, new_n13597);
xnor_4 g11249(new_n13447, new_n13444, new_n13598);
xnor_4 g11250(new_n13595, new_n13589, new_n13599);
nor_5  g11251(new_n13599, new_n13598, new_n13600);
xnor_4 g11252(new_n13599, new_n13598, new_n13601);
xnor_4 g11253(new_n13442, new_n13394, new_n13602_1);
not_8  g11254(new_n13602_1, new_n13603);
xnor_4 g11255(new_n13586, new_n13523, new_n13604);
nand_5 g11256(new_n13604, new_n13603, new_n13605);
xnor_4 g11257(new_n13604, new_n13602_1, new_n13606);
xnor_4 g11258(new_n13440, new_n13398, new_n13607);
not_8  g11259(new_n13607, new_n13608);
xnor_4 g11260(new_n13584, new_n13528, new_n13609);
nand_5 g11261(new_n13609, new_n13608, new_n13610);
xnor_4 g11262(new_n13609, new_n13607, new_n13611);
xnor_4 g11263(new_n13438, new_n13402, new_n13612);
not_8  g11264(new_n13612, new_n13613);
xnor_4 g11265(new_n13582, new_n13534, new_n13614);
nand_5 g11266(new_n13614, new_n13613, new_n13615);
xnor_4 g11267(new_n13614, new_n13612, new_n13616);
xnor_4 g11268(new_n13436, new_n13406, new_n13617);
not_8  g11269(new_n13617, new_n13618);
xnor_4 g11270(new_n13580, new_n13539, new_n13619);
nand_5 g11271(new_n13619, new_n13618, new_n13620);
xnor_4 g11272(new_n13619, new_n13617, new_n13621);
xnor_4 g11273(new_n13434, new_n13410, new_n13622);
not_8  g11274(new_n13622, new_n13623);
xnor_4 g11275(new_n13578, new_n13544, new_n13624);
nand_5 g11276(new_n13624, new_n13623, new_n13625);
xnor_4 g11277(new_n13624, new_n13622, new_n13626_1);
not_8  g11278(new_n13432, new_n13627);
xnor_4 g11279(new_n13627, new_n13413, new_n13628);
not_8  g11280(new_n13549_1, new_n13629);
xnor_4 g11281(new_n13576, new_n13629, new_n13630);
not_8  g11282(new_n13630, new_n13631);
nand_5 g11283(new_n13631, new_n13628, new_n13632);
xnor_4 g11284(new_n13630, new_n13628, new_n13633);
xnor_4 g11285(new_n13430, new_n13416, new_n13634);
not_8  g11286(new_n13634, new_n13635);
xnor_4 g11287(new_n13574, new_n13554, new_n13636);
nand_5 g11288(new_n13636, new_n13635, new_n13637);
xnor_4 g11289(new_n13636, new_n13634, new_n13638);
not_8  g11290(new_n13428, new_n13639);
xnor_4 g11291(new_n13639, new_n13419_1, new_n13640);
xnor_4 g11292(new_n13572, new_n13558, new_n13641);
not_8  g11293(new_n13641, new_n13642);
nand_5 g11294(new_n13642, new_n13640, new_n13643);
xnor_4 g11295(new_n13641, new_n13640, new_n13644);
xnor_4 g11296(new_n13570, new_n13569, new_n13645);
xnor_4 g11297(new_n13425, new_n13424_1, new_n13646);
not_8  g11298(new_n13646, new_n13647);
nor_5  g11299(new_n13647, new_n13645, new_n13648);
xnor_4 g11300(new_n13420, new_n7384, new_n13649);
xnor_4 g11301(new_n13567, new_n3946, new_n13650);
not_8  g11302(new_n13650, new_n13651);
nor_5  g11303(new_n13651, new_n13649, new_n13652);
not_8  g11304(new_n13652, new_n13653);
xnor_4 g11305(new_n13646, new_n13645, new_n13654);
not_8  g11306(new_n13654, new_n13655);
nor_5  g11307(new_n13655, new_n13653, new_n13656);
nor_5  g11308(new_n13656, new_n13648, new_n13657);
nand_5 g11309(new_n13657, new_n13644, new_n13658);
nand_5 g11310(new_n13658, new_n13643, new_n13659);
nand_5 g11311(new_n13659, new_n13638, new_n13660);
nand_5 g11312(new_n13660, new_n13637, new_n13661);
nand_5 g11313(new_n13661, new_n13633, new_n13662);
nand_5 g11314(new_n13662, new_n13632, new_n13663);
nand_5 g11315(new_n13663, new_n13626_1, new_n13664);
nand_5 g11316(new_n13664, new_n13625, new_n13665);
nand_5 g11317(new_n13665, new_n13621, new_n13666);
nand_5 g11318(new_n13666, new_n13620, new_n13667);
nand_5 g11319(new_n13667, new_n13616, new_n13668_1);
nand_5 g11320(new_n13668_1, new_n13615, new_n13669);
nand_5 g11321(new_n13669, new_n13611, new_n13670);
nand_5 g11322(new_n13670, new_n13610, new_n13671);
nand_5 g11323(new_n13671, new_n13606, new_n13672);
nand_5 g11324(new_n13672, new_n13605, new_n13673);
not_8  g11325(new_n13673, new_n13674);
nor_5  g11326(new_n13674, new_n13601, new_n13675);
nor_5  g11327(new_n13675, new_n13600, new_n13676);
xnor_4 g11328(new_n13676, new_n13597, n2095);
xnor_4 g11329(new_n12095, new_n12094, n2105);
not_8  g11330(new_n6410, new_n13679);
not_8  g11331(n8827, new_n13680);
not_8  g11332(n11898, new_n13681);
xnor_4 g11333(n23166, new_n13681, new_n13682);
not_8  g11334(n19941, new_n13683_1);
or_5   g11335(new_n13683_1, new_n9672, new_n13684);
not_8  g11336(new_n13684, new_n13685);
nor_5  g11337(n19941, n10577, new_n13686);
nor_5  g11338(n6381, n1099, new_n13687);
not_8  g11339(new_n13687, new_n13688);
nand_5 g11340(new_n11219, new_n11196, new_n13689);
nand_5 g11341(new_n13689, new_n13688, new_n13690);
nor_5  g11342(new_n13690, new_n13686, new_n13691);
nor_5  g11343(new_n13691, new_n13685, new_n13692);
xnor_4 g11344(new_n13692, new_n13682, new_n13693);
xnor_4 g11345(new_n13693, new_n13680, new_n13694);
xnor_4 g11346(n19941, new_n9672, new_n13695);
xnor_4 g11347(new_n13695, new_n13690, new_n13696);
nand_5 g11348(new_n13696, n18035, new_n13697);
not_8  g11349(new_n13697, new_n13698);
not_8  g11350(n18035, new_n13699);
xnor_4 g11351(new_n13696, new_n13699, new_n13700);
not_8  g11352(new_n13700, new_n13701);
nor_5  g11353(new_n11220_1, n5077, new_n13702);
not_8  g11354(new_n13702, new_n13703);
nand_5 g11355(new_n11249, new_n11221, new_n13704);
nand_5 g11356(new_n13704, new_n13703, new_n13705);
nor_5  g11357(new_n13705, new_n13701, new_n13706);
nor_5  g11358(new_n13706, new_n13698, new_n13707);
xnor_4 g11359(new_n13707, new_n13694, new_n13708_1);
xnor_4 g11360(new_n13708_1, new_n13679, new_n13709);
xnor_4 g11361(new_n13705, new_n13700, new_n13710_1);
nand_5 g11362(new_n13710_1, new_n6412, new_n13711);
not_8  g11363(new_n13710_1, new_n13712);
xnor_4 g11364(new_n13712, new_n6412, new_n13713);
nand_5 g11365(new_n11250, new_n6420, new_n13714_1);
not_8  g11366(new_n6420, new_n13715);
xnor_4 g11367(new_n11250, new_n13715, new_n13716);
nand_5 g11368(new_n11254, new_n6425, new_n13717);
xnor_4 g11369(new_n11256, new_n6425, new_n13718);
nand_5 g11370(new_n11260, new_n6432, new_n13719_1);
xnor_4 g11371(new_n11260, new_n6431_1, new_n13720);
nand_5 g11372(new_n11265, new_n6437_1, new_n13721);
xnor_4 g11373(new_n11266_1, new_n6437_1, new_n13722_1);
nor_5  g11374(new_n9004, new_n6441, new_n13723);
xnor_4 g11375(new_n11271, new_n6441, new_n13724);
not_8  g11376(new_n13724, new_n13725);
nor_5  g11377(new_n8979, new_n6448, new_n13726);
xnor_4 g11378(new_n8979, new_n6447, new_n13727);
not_8  g11379(new_n13727, new_n13728);
not_8  g11380(new_n6452, new_n13729);
nor_5  g11381(new_n8984, new_n13729, new_n13730);
nor_5  g11382(new_n8989, new_n6109, new_n13731);
not_8  g11383(new_n13731, new_n13732);
xnor_4 g11384(new_n8983, new_n13729, new_n13733);
not_8  g11385(new_n13733, new_n13734);
nor_5  g11386(new_n13734, new_n13732, new_n13735);
nor_5  g11387(new_n13735, new_n13730, new_n13736);
nor_5  g11388(new_n13736, new_n13728, new_n13737);
nor_5  g11389(new_n13737, new_n13726, new_n13738);
nor_5  g11390(new_n13738, new_n13725, new_n13739);
nor_5  g11391(new_n13739, new_n13723, new_n13740);
not_8  g11392(new_n13740, new_n13741);
nand_5 g11393(new_n13741, new_n13722_1, new_n13742);
nand_5 g11394(new_n13742, new_n13721, new_n13743);
nand_5 g11395(new_n13743, new_n13720, new_n13744);
nand_5 g11396(new_n13744, new_n13719_1, new_n13745);
nand_5 g11397(new_n13745, new_n13718, new_n13746);
nand_5 g11398(new_n13746, new_n13717, new_n13747);
nand_5 g11399(new_n13747, new_n13716, new_n13748);
nand_5 g11400(new_n13748, new_n13714_1, new_n13749);
nand_5 g11401(new_n13749, new_n13713, new_n13750);
nand_5 g11402(new_n13750, new_n13711, new_n13751);
xnor_4 g11403(new_n13751, new_n13709, n2122);
xnor_4 g11404(new_n2887_1, new_n2859, n2147);
xnor_4 g11405(new_n11162, new_n11113, n2209);
xor_4  g11406(new_n6085, new_n5960, n2214);
not_8  g11407(new_n4383, new_n13756);
xnor_4 g11408(new_n11864, new_n13756, new_n13757);
nor_5  g11409(new_n11867, new_n4471, new_n13758);
not_8  g11410(new_n13758, new_n13759);
xnor_4 g11411(new_n11867, new_n4472, new_n13760);
nor_5  g11412(new_n11871, new_n4478_1, new_n13761);
xnor_4 g11413(new_n11871, new_n4478_1, new_n13762);
nor_5  g11414(new_n11880, new_n4486, new_n13763);
nor_5  g11415(new_n11876, new_n4490, new_n13764_1);
xnor_4 g11416(new_n11879, new_n4486, new_n13765);
not_8  g11417(new_n13765, new_n13766);
nor_5  g11418(new_n13766, new_n13764_1, new_n13767);
nor_5  g11419(new_n13767, new_n13763, new_n13768);
not_8  g11420(new_n13768, new_n13769);
nor_5  g11421(new_n13769, new_n13762, new_n13770);
nor_5  g11422(new_n13770, new_n13761, new_n13771);
nand_5 g11423(new_n13771, new_n13760, new_n13772);
nand_5 g11424(new_n13772, new_n13759, new_n13773);
xnor_4 g11425(new_n13773, new_n13757, n2238);
xor_4  g11426(new_n11890, new_n11888, n2327);
xnor_4 g11427(new_n6068, new_n6030, n2343);
xnor_4 g11428(new_n11233, new_n8268, new_n13777);
nor_5  g11429(new_n6958, new_n8299, new_n13778);
not_8  g11430(new_n6959, new_n13779);
nor_5  g11431(new_n6977, new_n13779, new_n13780);
nor_5  g11432(new_n13780, new_n13778, new_n13781_1);
xnor_4 g11433(new_n13781_1, new_n13777, new_n13782);
xnor_4 g11434(n20923, new_n11285, new_n13783_1);
nor_5  g11435(n18157, n11056, new_n13784);
not_8  g11436(new_n6980, new_n13785);
nor_5  g11437(new_n6992, new_n13785, new_n13786);
nor_5  g11438(new_n13786, new_n13784, new_n13787);
xnor_4 g11439(new_n13787, new_n13783_1, new_n13788);
xnor_4 g11440(new_n13788, n3785, new_n13789);
nand_5 g11441(new_n6993, new_n4573, new_n13790);
not_8  g11442(new_n13790, new_n13791);
not_8  g11443(new_n6994, new_n13792);
nor_5  g11444(new_n7010, new_n13792, new_n13793);
nor_5  g11445(new_n13793, new_n13791, new_n13794);
xnor_4 g11446(new_n13794, new_n13789, new_n13795);
not_8  g11447(new_n13795, new_n13796);
xnor_4 g11448(new_n13796, new_n13782, new_n13797);
not_8  g11449(new_n6978, new_n13798_1);
nor_5  g11450(new_n7012, new_n13798_1, new_n13799);
not_8  g11451(new_n13799, new_n13800);
nand_5 g11452(new_n7034, new_n7013, new_n13801);
nand_5 g11453(new_n13801, new_n13800, new_n13802);
xnor_4 g11454(new_n13802, new_n13797, n2361);
xnor_4 g11455(new_n3855, new_n8890, n2363);
xnor_4 g11456(new_n4807, new_n4771, n2374);
not_8  g11457(new_n3931, new_n13806);
not_8  g11458(new_n5111, new_n13807);
xnor_4 g11459(n7305, new_n4015, new_n13808);
nor_5  g11460(n25872, n19618, new_n13809);
not_8  g11461(new_n6145, new_n13810);
nor_5  g11462(new_n6151, new_n13810, new_n13811);
nor_5  g11463(new_n13811, new_n13809, new_n13812);
xnor_4 g11464(new_n13812, new_n13808, new_n13813);
not_8  g11465(new_n13813, new_n13814);
nor_5  g11466(new_n13814, new_n5114, new_n13815);
not_8  g11467(new_n13815, new_n13816);
xnor_4 g11468(new_n13813, new_n5114, new_n13817);
nor_5  g11469(new_n6152, new_n6144, new_n13818);
nor_5  g11470(new_n6163, new_n6153, new_n13819);
nor_5  g11471(new_n13819, new_n13818, new_n13820);
nand_5 g11472(new_n13820, new_n13817, new_n13821);
nand_5 g11473(new_n13821, new_n13816, new_n13822);
xnor_4 g11474(n20826, new_n3993, new_n13823);
nor_5  g11475(n7305, n1204, new_n13824);
not_8  g11476(new_n13808, new_n13825);
nor_5  g11477(new_n13812, new_n13825, new_n13826);
nor_5  g11478(new_n13826, new_n13824, new_n13827);
xnor_4 g11479(new_n13827, new_n13823, new_n13828);
not_8  g11480(new_n13828, new_n13829);
xnor_4 g11481(new_n13829, new_n13822, new_n13830);
xnor_4 g11482(new_n13830, new_n13807, new_n13831);
xnor_4 g11483(new_n13831, new_n13806, new_n13832);
not_8  g11484(new_n3935, new_n13833);
xnor_4 g11485(new_n13820, new_n13817, new_n13834);
not_8  g11486(new_n13834, new_n13835_1);
nor_5  g11487(new_n13835_1, new_n13833, new_n13836);
not_8  g11488(new_n3939, new_n13837);
nor_5  g11489(new_n6164, new_n13837, new_n13838);
nand_5 g11490(new_n6174, new_n6165, new_n13839);
not_8  g11491(new_n13839, new_n13840);
nor_5  g11492(new_n13840, new_n13838, new_n13841);
xnor_4 g11493(new_n13834, new_n13833, new_n13842);
not_8  g11494(new_n13842, new_n13843);
nor_5  g11495(new_n13843, new_n13841, new_n13844);
nor_5  g11496(new_n13844, new_n13836, new_n13845);
xor_4  g11497(new_n13845, new_n13832, n2388);
xnor_4 g11498(n7335, new_n12514, new_n13847);
or_5   g11499(n10763, n5696, new_n13848);
nand_5 g11500(new_n5616, new_n5581, new_n13849);
nand_5 g11501(new_n13849, new_n13848, new_n13850_1);
xnor_4 g11502(new_n13850_1, new_n13847, new_n13851_1);
xnor_4 g11503(n11220, new_n3294, new_n13852);
or_5   g11504(n22379, n9967, new_n13853);
nand_5 g11505(new_n5579_1, new_n5543, new_n13854);
nand_5 g11506(new_n13854, new_n13853, new_n13855);
xnor_4 g11507(new_n13855, new_n13852, new_n13856);
xnor_4 g11508(new_n13856, new_n13851_1, new_n13857);
not_8  g11509(new_n5617, new_n13858);
nor_5  g11510(new_n13858, new_n5580, new_n13859);
not_8  g11511(new_n13859, new_n13860);
nand_5 g11512(new_n5672, new_n13860, new_n13861);
xnor_4 g11513(new_n13861, new_n13857, new_n13862);
not_8  g11514(new_n13862, new_n13863);
not_8  g11515(n7593, new_n13864);
nand_5 g11516(new_n5494, new_n3387, new_n13865);
xnor_4 g11517(new_n13865, new_n13864, new_n13866);
xnor_4 g11518(new_n13866, new_n3163, new_n13867);
or_5   g11519(new_n5495, n6485, new_n13868);
nand_5 g11520(new_n5541, new_n5496, new_n13869);
nand_5 g11521(new_n13869, new_n13868, new_n13870);
xnor_4 g11522(new_n13870, new_n13867, new_n13871);
xnor_4 g11523(new_n13871, new_n13863, new_n13872);
not_8  g11524(new_n5542, new_n13873);
nand_5 g11525(new_n5675, new_n13873, new_n13874);
nand_5 g11526(new_n5733, new_n13874, new_n13875);
xnor_4 g11527(new_n13875, new_n13872, n2440);
xnor_4 g11528(new_n12264, new_n12246, n2444);
xnor_4 g11529(new_n5348, new_n3351, n2513);
not_8  g11530(n14323, new_n13879);
xnor_4 g11531(new_n6268, new_n13879, new_n13880);
not_8  g11532(n2886, new_n13881);
nor_5  g11533(new_n6275, new_n13881, new_n13882);
not_8  g11534(new_n13882, new_n13883);
xnor_4 g11535(new_n6274, new_n13881, new_n13884);
nor_5  g11536(new_n6288, new_n13372, new_n13885);
not_8  g11537(new_n13885, new_n13886);
nand_5 g11538(n20658, n9090, new_n13887);
not_8  g11539(new_n13887, new_n13888);
xnor_4 g11540(new_n6288, n1040, new_n13889);
nand_5 g11541(new_n13889, new_n13888, new_n13890);
nand_5 g11542(new_n13890, new_n13886, new_n13891);
nand_5 g11543(new_n13891, new_n13884, new_n13892);
nand_5 g11544(new_n13892, new_n13883, new_n13893);
xnor_4 g11545(new_n13893, new_n13880, new_n13894);
xnor_4 g11546(new_n13894, n12562, new_n13895);
not_8  g11547(new_n13884, new_n13896);
xnor_4 g11548(new_n13891, new_n13896, new_n13897);
nor_5  g11549(new_n13897, n7949, new_n13898);
xnor_4 g11550(new_n13897, n7949, new_n13899);
not_8  g11551(new_n11573, new_n13900);
nor_5  g11552(new_n13900, new_n6281, new_n13901);
nor_5  g11553(new_n13901, n24374, new_n13902);
xnor_4 g11554(new_n13889, new_n13888, new_n13903);
not_8  g11555(new_n13903, new_n13904);
not_8  g11556(n24374, new_n13905);
xnor_4 g11557(new_n13901, new_n13905, new_n13906);
not_8  g11558(new_n13906, new_n13907);
nor_5  g11559(new_n13907, new_n13904, new_n13908);
nor_5  g11560(new_n13908, new_n13902, new_n13909);
nor_5  g11561(new_n13909, new_n13899, new_n13910);
nor_5  g11562(new_n13910, new_n13898, new_n13911);
xnor_4 g11563(new_n13911, new_n13895, new_n13912_1);
not_8  g11564(new_n13912_1, new_n13913);
xnor_4 g11565(new_n13913, new_n13636, new_n13914_1);
not_8  g11566(new_n13909, new_n13915);
xnor_4 g11567(new_n13915, new_n13899, new_n13916);
nand_5 g11568(new_n13916, new_n13642, new_n13917);
xnor_4 g11569(new_n13916, new_n13641, new_n13918);
xnor_4 g11570(new_n13906, new_n13904, new_n13919);
nand_5 g11571(new_n13919, new_n13645, new_n13920);
xnor_4 g11572(new_n11573, new_n6281, new_n13921);
and_5  g11573(new_n13921, new_n13650, new_n13922_1);
not_8  g11574(new_n13922_1, new_n13923_1);
xnor_4 g11575(new_n13919, new_n13645, new_n13924);
not_8  g11576(new_n13924, new_n13925);
nand_5 g11577(new_n13925, new_n13923_1, new_n13926);
nand_5 g11578(new_n13926, new_n13920, new_n13927);
nand_5 g11579(new_n13927, new_n13918, new_n13928);
nand_5 g11580(new_n13928, new_n13917, new_n13929);
xnor_4 g11581(new_n13929, new_n13914_1, n2515);
xnor_4 g11582(new_n11564_1, new_n11530, n2533);
or_5   g11583(n26986, new_n3294, new_n13932);
xnor_4 g11584(n26986, n3425, new_n13933);
or_5   g11585(n21287, new_n3295, new_n13934);
xnor_4 g11586(n21287, n9967, new_n13935);
or_5   g11587(new_n3317, n4256, new_n13936);
xnor_4 g11588(n20946, n4256, new_n13937);
or_5   g11589(n22332, new_n2430, new_n13938);
xnor_4 g11590(n22332, n7751, new_n13939);
or_5   g11591(new_n2434, n18907, new_n13940);
xnor_4 g11592(n26823, n18907, new_n13941);
nor_5  g11593(new_n2438, n2731, new_n13942);
not_8  g11594(new_n13942, new_n13943);
nor_5  g11595(new_n8932, new_n8919, new_n13944);
not_8  g11596(new_n13944, new_n13945);
nand_5 g11597(new_n13945, new_n13943, new_n13946);
nand_5 g11598(new_n13946, new_n13941, new_n13947);
nand_5 g11599(new_n13947, new_n13940, new_n13948);
nand_5 g11600(new_n13948, new_n13939, new_n13949);
nand_5 g11601(new_n13949, new_n13938, new_n13950);
nand_5 g11602(new_n13950, new_n13937, new_n13951_1);
nand_5 g11603(new_n13951_1, new_n13936, new_n13952);
nand_5 g11604(new_n13952, new_n13935, new_n13953);
nand_5 g11605(new_n13953, new_n13934, new_n13954);
nand_5 g11606(new_n13954, new_n13933, new_n13955);
nand_5 g11607(new_n13955, new_n13932, new_n13956);
not_8  g11608(new_n13956, new_n13957);
nand_5 g11609(new_n5390, new_n5384, new_n13958);
nor_5  g11610(new_n7480, new_n13958, new_n13959);
nand_5 g11611(new_n13959, new_n7475_1, new_n13960);
nor_5  g11612(new_n13960, new_n7470, new_n13961);
nand_5 g11613(new_n13961, new_n7539, new_n13962);
nor_5  g11614(new_n13962, new_n7622, new_n13963);
not_8  g11615(new_n13963, new_n13964);
not_8  g11616(new_n7624, new_n13965);
nand_5 g11617(new_n13962, new_n13965, new_n13966);
not_8  g11618(new_n13966, new_n13967);
nor_5  g11619(new_n13967, new_n13963, new_n13968);
not_8  g11620(new_n13968, new_n13969);
nand_5 g11621(new_n13969, new_n3290, new_n13970);
xnor_4 g11622(new_n13961, new_n7539, new_n13971);
nand_5 g11623(new_n13971, new_n3215, new_n13972);
xnor_4 g11624(new_n13971, new_n3216, new_n13973);
xnor_4 g11625(new_n13960, new_n7470, new_n13974);
nand_5 g11626(new_n13974, new_n3221, new_n13975);
xnor_4 g11627(new_n13974, new_n3222, new_n13976);
xnor_4 g11628(new_n13959, new_n7475_1, new_n13977);
nand_5 g11629(new_n13977, new_n3227, new_n13978);
xnor_4 g11630(new_n13977, new_n3228_1, new_n13979);
xnor_4 g11631(new_n7480, new_n13958, new_n13980);
nand_5 g11632(new_n13980, new_n3233, new_n13981);
xnor_4 g11633(new_n13980, new_n3234, new_n13982);
not_8  g11634(new_n3238, new_n13983);
nand_5 g11635(new_n5391, new_n13983, new_n13984);
nand_5 g11636(new_n5425, new_n5392, new_n13985);
nand_5 g11637(new_n13985, new_n13984, new_n13986);
nand_5 g11638(new_n13986, new_n13982, new_n13987);
nand_5 g11639(new_n13987, new_n13981, new_n13988);
nand_5 g11640(new_n13988, new_n13979, new_n13989);
nand_5 g11641(new_n13989, new_n13978, new_n13990);
nand_5 g11642(new_n13990, new_n13976, new_n13991);
nand_5 g11643(new_n13991, new_n13975, new_n13992);
nand_5 g11644(new_n13992, new_n13973, new_n13993);
nand_5 g11645(new_n13993, new_n13972, new_n13994);
nand_5 g11646(new_n13968, new_n3291, new_n13995);
nand_5 g11647(new_n13995, new_n13994, new_n13996);
nand_5 g11648(new_n13996, new_n13970, new_n13997);
nand_5 g11649(new_n13997, new_n13964, new_n13998);
xnor_4 g11650(new_n13998, new_n13957, new_n13999);
xnor_4 g11651(new_n13968, new_n3291, new_n14000);
xnor_4 g11652(new_n14000, new_n13994, new_n14001);
nand_5 g11653(new_n14001, new_n13956, new_n14002);
xnor_4 g11654(new_n14001, new_n13957, new_n14003);
xnor_4 g11655(new_n13954, new_n13933, new_n14004_1);
xnor_4 g11656(new_n13992, new_n13973, new_n14005);
not_8  g11657(new_n14005, new_n14006);
nand_5 g11658(new_n14006, new_n14004_1, new_n14007);
xnor_4 g11659(new_n14005, new_n14004_1, new_n14008);
xnor_4 g11660(new_n13952, new_n13935, new_n14009);
xnor_4 g11661(new_n13990, new_n13976, new_n14010);
not_8  g11662(new_n14010, new_n14011);
nand_5 g11663(new_n14011, new_n14009, new_n14012);
xnor_4 g11664(new_n14010, new_n14009, new_n14013);
xnor_4 g11665(new_n13950, new_n13937, new_n14014);
xnor_4 g11666(new_n13988, new_n13979, new_n14015);
not_8  g11667(new_n14015, new_n14016);
nand_5 g11668(new_n14016, new_n14014, new_n14017);
xnor_4 g11669(new_n14015, new_n14014, new_n14018);
xnor_4 g11670(new_n13948, new_n13939, new_n14019);
not_8  g11671(new_n14019, new_n14020);
xnor_4 g11672(new_n13986, new_n13982, new_n14021);
nor_5  g11673(new_n14021, new_n14020, new_n14022);
not_8  g11674(new_n14022, new_n14023);
xnor_4 g11675(new_n14021, new_n14019, new_n14024);
xnor_4 g11676(new_n13946, new_n13941, new_n14025);
nor_5  g11677(new_n14025, new_n5426, new_n14026);
xnor_4 g11678(new_n14025, new_n5426, new_n14027);
nor_5  g11679(new_n8933, new_n8917, new_n14028);
nor_5  g11680(new_n8956, new_n8934, new_n14029);
nor_5  g11681(new_n14029, new_n14028, new_n14030);
nor_5  g11682(new_n14030, new_n14027, new_n14031);
nor_5  g11683(new_n14031, new_n14026, new_n14032);
nand_5 g11684(new_n14032, new_n14024, new_n14033);
nand_5 g11685(new_n14033, new_n14023, new_n14034);
nand_5 g11686(new_n14034, new_n14018, new_n14035);
nand_5 g11687(new_n14035, new_n14017, new_n14036_1);
nand_5 g11688(new_n14036_1, new_n14013, new_n14037);
nand_5 g11689(new_n14037, new_n14012, new_n14038);
nand_5 g11690(new_n14038, new_n14008, new_n14039);
nand_5 g11691(new_n14039, new_n14007, new_n14040);
nand_5 g11692(new_n14040, new_n14003, new_n14041);
nand_5 g11693(new_n14041, new_n14002, new_n14042);
xnor_4 g11694(new_n14042, new_n13999, n2535);
nor_5  g11695(n20259, n3925, new_n14044);
nand_5 g11696(new_n14044, new_n5181, new_n14045);
nor_5  g11697(new_n14045, n7305, new_n14046);
nand_5 g11698(new_n14046, new_n5174, new_n14047);
xnor_4 g11699(new_n14047, new_n5170, new_n14048);
xnor_4 g11700(new_n14048, new_n5004, new_n14049);
xnor_4 g11701(new_n14046, n20826, new_n14050);
not_8  g11702(new_n14050, new_n14051);
nand_5 g11703(new_n14051, new_n5008, new_n14052);
xnor_4 g11704(new_n14050, new_n5008, new_n14053);
xnor_4 g11705(new_n14045, new_n5176, new_n14054);
not_8  g11706(new_n14054, new_n14055);
nand_5 g11707(new_n14055, new_n8754, new_n14056);
xnor_4 g11708(new_n14044, n25872, new_n14057);
not_8  g11709(new_n14057, new_n14058);
nand_5 g11710(new_n14058, new_n3694, new_n14059_1);
xnor_4 g11711(new_n14057, new_n3694, new_n14060);
xnor_4 g11712(n20259, n3925, new_n14061);
nand_5 g11713(new_n14061, new_n3698, new_n14062);
nand_5 g11714(n9246, n3925, new_n14063);
xnor_4 g11715(new_n14061, n16994, new_n14064);
nand_5 g11716(new_n14064, new_n14063, new_n14065);
nand_5 g11717(new_n14065, new_n14062, new_n14066);
nand_5 g11718(new_n14066, new_n14060, new_n14067);
nand_5 g11719(new_n14067, new_n14059_1, new_n14068);
xnor_4 g11720(new_n14054, new_n8754, new_n14069);
nand_5 g11721(new_n14069, new_n14068, new_n14070);
nand_5 g11722(new_n14070, new_n14056, new_n14071_1);
nand_5 g11723(new_n14071_1, new_n14053, new_n14072);
nand_5 g11724(new_n14072, new_n14052, new_n14073);
xnor_4 g11725(new_n14073, new_n14049, new_n14074);
xnor_4 g11726(new_n14074, new_n8213, new_n14075);
xnor_4 g11727(new_n14071_1, new_n14053, new_n14076);
nor_5  g11728(new_n14076, new_n8219, new_n14077);
not_8  g11729(new_n14077, new_n14078);
xnor_4 g11730(new_n14076, new_n8219, new_n14079);
not_8  g11731(new_n14079, new_n14080);
xnor_4 g11732(new_n14069, new_n14068, new_n14081_1);
nor_5  g11733(new_n14081_1, new_n8224, new_n14082);
not_8  g11734(new_n14082, new_n14083);
xnor_4 g11735(new_n14081_1, new_n8224, new_n14084);
not_8  g11736(new_n14084, new_n14085);
not_8  g11737(new_n8232, new_n14086);
xnor_4 g11738(new_n14066, new_n14060, new_n14087);
nand_5 g11739(new_n14087, new_n14086, new_n14088);
not_8  g11740(new_n14088, new_n14089);
xnor_4 g11741(new_n14087, new_n8232, new_n14090_1);
not_8  g11742(new_n14090_1, new_n14091);
xnor_4 g11743(new_n14064, new_n14063, new_n14092);
nand_5 g11744(new_n14092, new_n8240, new_n14093);
not_8  g11745(new_n14093, new_n14094);
not_8  g11746(new_n10376, new_n14095_1);
nor_5  g11747(new_n14095_1, new_n8243, new_n14096);
not_8  g11748(new_n14096, new_n14097);
xnor_4 g11749(new_n14092, new_n8240, new_n14098);
nor_5  g11750(new_n14098, new_n14097, new_n14099);
nor_5  g11751(new_n14099, new_n14094, new_n14100);
nor_5  g11752(new_n14100, new_n14091, new_n14101);
nor_5  g11753(new_n14101, new_n14089, new_n14102);
nand_5 g11754(new_n14102, new_n14085, new_n14103);
nand_5 g11755(new_n14103, new_n14083, new_n14104);
nand_5 g11756(new_n14104, new_n14080, new_n14105);
nand_5 g11757(new_n14105, new_n14078, new_n14106);
xnor_4 g11758(new_n14106, new_n14075, new_n14107_1);
not_8  g11759(new_n14107_1, new_n14108);
xnor_4 g11760(n1163, n329, new_n14109);
nor_5  g11761(new_n8803_1, n18537, new_n14110);
xnor_4 g11762(n24170, n18537, new_n14111);
not_8  g11763(new_n14111, new_n14112);
nor_5  g11764(n7057, new_n7422, new_n14113);
xnor_4 g11765(n7057, n2409, new_n14114);
nor_5  g11766(n8869, new_n5296, new_n14115);
nor_5  g11767(new_n8807, n8381, new_n14116);
nor_5  g11768(new_n5307, n10372, new_n14117);
nor_5  g11769(new_n9044, n7428, new_n14118);
not_8  g11770(new_n14118, new_n14119);
nor_5  g11771(n20235, new_n7431, new_n14120);
nor_5  g11772(new_n14120, new_n14119, new_n14121_1);
nor_5  g11773(new_n14121_1, new_n14117, new_n14122);
nor_5  g11774(new_n14122, new_n14116, new_n14123);
nor_5  g11775(new_n14123, new_n14115, new_n14124);
and_5  g11776(new_n14124, new_n14114, new_n14125);
nor_5  g11777(new_n14125, new_n14113, new_n14126_1);
nor_5  g11778(new_n14126_1, new_n14112, new_n14127);
nor_5  g11779(new_n14127, new_n14110, new_n14128);
xnor_4 g11780(new_n14128, new_n14109, new_n14129);
xnor_4 g11781(new_n14129, new_n14108, new_n14130_1);
xnor_4 g11782(new_n14126_1, new_n14111, new_n14131);
xnor_4 g11783(new_n14104, new_n14080, new_n14132);
nor_5  g11784(new_n14132, new_n14131, new_n14133);
xnor_4 g11785(new_n14132, new_n14131, new_n14134);
not_8  g11786(new_n14100, new_n14135);
nand_5 g11787(new_n14135, new_n14090_1, new_n14136_1);
nand_5 g11788(new_n14136_1, new_n14088, new_n14137);
xnor_4 g11789(new_n14137, new_n14084, new_n14138);
xnor_4 g11790(new_n14124, new_n14114, new_n14139);
not_8  g11791(new_n14139, new_n14140);
nor_5  g11792(new_n14140, new_n14138, new_n14141);
xnor_4 g11793(new_n14140, new_n14138, new_n14142);
xnor_4 g11794(new_n14100, new_n14090_1, new_n14143);
xnor_4 g11795(n8869, n8381, new_n14144);
xnor_4 g11796(new_n14144, new_n14122, new_n14145);
not_8  g11797(new_n14145, new_n14146);
nor_5  g11798(new_n14146, new_n14143, new_n14147_1);
xnor_4 g11799(new_n14146, new_n14143, new_n14148_1);
not_8  g11800(new_n10377, new_n14149);
nor_5  g11801(new_n10378, new_n14149, new_n14150);
xnor_4 g11802(n20235, n10372, new_n14151);
xnor_4 g11803(new_n14151, new_n14119, new_n14152);
not_8  g11804(new_n14152, new_n14153);
nor_5  g11805(new_n14153, new_n14150, new_n14154);
xnor_4 g11806(new_n14098, new_n14096, new_n14155);
not_8  g11807(new_n14155, new_n14156);
xnor_4 g11808(new_n14152, new_n14150, new_n14157);
nand_5 g11809(new_n14157, new_n14156, new_n14158);
not_8  g11810(new_n14158, new_n14159);
nor_5  g11811(new_n14159, new_n14154, new_n14160);
nor_5  g11812(new_n14160, new_n14148_1, new_n14161);
nor_5  g11813(new_n14161, new_n14147_1, new_n14162);
nor_5  g11814(new_n14162, new_n14142, new_n14163);
nor_5  g11815(new_n14163, new_n14141, new_n14164);
nor_5  g11816(new_n14164, new_n14134, new_n14165);
nor_5  g11817(new_n14165, new_n14133, new_n14166);
xnor_4 g11818(new_n14166, new_n14130_1, n2537);
xnor_4 g11819(new_n11746, new_n3049, new_n14168);
not_8  g11820(new_n14168, new_n14169);
nor_5  g11821(new_n4388, new_n3056, new_n14170);
xnor_4 g11822(new_n4387, new_n3056, new_n14171);
not_8  g11823(new_n14171, new_n14172);
nor_5  g11824(new_n4391, new_n3063, new_n14173);
not_8  g11825(new_n14173, new_n14174_1);
not_8  g11826(new_n4391, new_n14175);
xnor_4 g11827(new_n14175, new_n3063, new_n14176);
not_8  g11828(new_n4394, new_n14177);
nor_5  g11829(new_n14177, new_n3069, new_n14178);
xnor_4 g11830(new_n14177, new_n3068, new_n14179);
not_8  g11831(new_n4397, new_n14180);
nor_5  g11832(new_n14180, new_n3074, new_n14181);
nor_5  g11833(new_n3080, n1152, new_n14182);
xnor_4 g11834(new_n4397, new_n3074, new_n14183);
nand_5 g11835(new_n14183, new_n14182, new_n14184);
not_8  g11836(new_n14184, new_n14185);
nor_5  g11837(new_n14185, new_n14181, new_n14186);
nand_5 g11838(new_n14186, new_n14179, new_n14187);
not_8  g11839(new_n14187, new_n14188);
nor_5  g11840(new_n14188, new_n14178, new_n14189);
nand_5 g11841(new_n14189, new_n14176, new_n14190_1);
nand_5 g11842(new_n14190_1, new_n14174_1, new_n14191);
nor_5  g11843(new_n14191, new_n14172, new_n14192);
nor_5  g11844(new_n14192, new_n14170, new_n14193);
xnor_4 g11845(new_n14193, new_n14169, new_n14194);
xnor_4 g11846(new_n14194, new_n12209_1, new_n14195);
xnor_4 g11847(new_n14191, new_n14171, new_n14196);
nor_5  g11848(new_n14196, new_n10167, new_n14197);
xnor_4 g11849(new_n14196, new_n12785, new_n14198);
not_8  g11850(new_n14198, new_n14199);
xnor_4 g11851(new_n14189, new_n14176, new_n14200);
nor_5  g11852(new_n14200, new_n10170, new_n14201);
xnor_4 g11853(new_n14200, new_n12791, new_n14202);
not_8  g11854(new_n14202, new_n14203);
xnor_4 g11855(new_n14186, new_n14179, new_n14204);
nor_5  g11856(new_n14204, new_n12797, new_n14205);
xnor_4 g11857(new_n14204, new_n12797, new_n14206);
xnor_4 g11858(new_n14183, new_n14182, new_n14207);
nor_5  g11859(new_n14207, new_n10182, new_n14208);
xnor_4 g11860(new_n3079, n1152, new_n14209);
nor_5  g11861(new_n14209, new_n7637, new_n14210);
xnor_4 g11862(new_n14207, new_n10181, new_n14211_1);
not_8  g11863(new_n14211_1, new_n14212);
nor_5  g11864(new_n14212, new_n14210, new_n14213);
nor_5  g11865(new_n14213, new_n14208, new_n14214);
not_8  g11866(new_n14214, new_n14215);
nor_5  g11867(new_n14215, new_n14206, new_n14216);
nor_5  g11868(new_n14216, new_n14205, new_n14217);
not_8  g11869(new_n14217, new_n14218);
nor_5  g11870(new_n14218, new_n14203, new_n14219);
nor_5  g11871(new_n14219, new_n14201, new_n14220);
nor_5  g11872(new_n14220, new_n14199, new_n14221);
nor_5  g11873(new_n14221, new_n14197, new_n14222_1);
not_8  g11874(new_n14222_1, new_n14223);
xnor_4 g11875(new_n14223, new_n14195, n2553);
xnor_4 g11876(new_n12682, new_n12660, n2555);
not_8  g11877(n12892, new_n14226);
xnor_4 g11878(new_n11393, new_n14226, new_n14227);
not_8  g11879(new_n14227, new_n14228);
nor_5  g11880(new_n14228, new_n10669, new_n14229);
not_8  g11881(new_n14229, new_n14230_1);
nor_5  g11882(new_n11489, new_n14226, new_n14231);
xnor_4 g11883(new_n11396, n12209, new_n14232);
xnor_4 g11884(new_n14232, new_n14231, new_n14233);
xnor_4 g11885(new_n14233, new_n10673, new_n14234);
xnor_4 g11886(new_n14234, new_n14230_1, n2560);
or_5   g11887(n26180, n10650, new_n14236);
xnor_4 g11888(n26180, new_n13343, new_n14237);
or_5   g11889(n24004, n12900, new_n14238);
not_8  g11890(n12900, new_n14239);
xnor_4 g11891(n24004, new_n14239, new_n14240);
or_5   g11892(n20411, n12871, new_n14241);
xnor_4 g11893(n20411, new_n3614, new_n14242);
nor_5  g11894(n23304, n17069, new_n14243);
not_8  g11895(new_n14243, new_n14244);
not_8  g11896(n17069, new_n14245);
xnor_4 g11897(n23304, new_n14245, new_n14246);
nor_5  g11898(n19361, n15918, new_n14247);
xnor_4 g11899(n19361, new_n13357, new_n14248);
not_8  g11900(new_n14248, new_n14249);
nor_5  g11901(n17784, n1437, new_n14250);
xnor_4 g11902(n17784, new_n3629, new_n14251);
not_8  g11903(new_n14251, new_n14252);
nor_5  g11904(n14323, n4722, new_n14253);
xnor_4 g11905(n14323, new_n3637, new_n14254);
not_8  g11906(new_n14254, new_n14255);
nor_5  g11907(n14633, n2886, new_n14256);
xnor_4 g11908(n14633, new_n13881, new_n14257);
not_8  g11909(new_n14257, new_n14258);
nor_5  g11910(n8721, n1040, new_n14259);
nand_5 g11911(n18578, n9090, new_n14260);
not_8  g11912(new_n14260, new_n14261);
xnor_4 g11913(n8721, new_n13372, new_n14262);
not_8  g11914(new_n14262, new_n14263);
nor_5  g11915(new_n14263, new_n14261, new_n14264);
nor_5  g11916(new_n14264, new_n14259, new_n14265);
nor_5  g11917(new_n14265, new_n14258, new_n14266);
nor_5  g11918(new_n14266, new_n14256, new_n14267_1);
nor_5  g11919(new_n14267_1, new_n14255, new_n14268);
nor_5  g11920(new_n14268, new_n14253, new_n14269);
nor_5  g11921(new_n14269, new_n14252, new_n14270);
nor_5  g11922(new_n14270, new_n14250, new_n14271_1);
nor_5  g11923(new_n14271_1, new_n14249, new_n14272);
nor_5  g11924(new_n14272, new_n14247, new_n14273);
not_8  g11925(new_n14273, new_n14274);
nand_5 g11926(new_n14274, new_n14246, new_n14275_1);
nand_5 g11927(new_n14275_1, new_n14244, new_n14276);
nand_5 g11928(new_n14276, new_n14242, new_n14277_1);
nand_5 g11929(new_n14277_1, new_n14241, new_n14278);
nand_5 g11930(new_n14278, new_n14240, new_n14279);
nand_5 g11931(new_n14279, new_n14238, new_n14280);
nand_5 g11932(new_n14280, new_n14237, new_n14281);
nand_5 g11933(new_n14281, new_n14236, new_n14282);
nor_5  g11934(n9259, n6456, new_n14283);
not_8  g11935(new_n14283, new_n14284);
nand_5 g11936(new_n6235, new_n6189_1, new_n14285);
nand_5 g11937(new_n14285, new_n14284, new_n14286);
not_8  g11938(new_n14286, new_n14287);
nand_5 g11939(new_n14287, new_n14282, new_n14288);
xnor_4 g11940(new_n14286, new_n14282, new_n14289);
not_8  g11941(new_n14237, new_n14290);
xnor_4 g11942(new_n14280, new_n14290, new_n14291);
nand_5 g11943(new_n14291, new_n6236, new_n14292);
xnor_4 g11944(new_n14280, new_n14237, new_n14293);
xnor_4 g11945(new_n14293, new_n6236, new_n14294_1);
not_8  g11946(new_n14240, new_n14295);
xnor_4 g11947(new_n14278, new_n14295, new_n14296);
nand_5 g11948(new_n14296, new_n6240, new_n14297);
xnor_4 g11949(new_n14278, new_n14240, new_n14298);
xnor_4 g11950(new_n14298, new_n6240, new_n14299);
not_8  g11951(new_n14242, new_n14300);
xnor_4 g11952(new_n14276, new_n14300, new_n14301);
nand_5 g11953(new_n14301, new_n6247, new_n14302);
xnor_4 g11954(new_n14301, new_n6246, new_n14303);
xnor_4 g11955(new_n14273, new_n14246, new_n14304);
nand_5 g11956(new_n14304, new_n6253, new_n14305);
xnor_4 g11957(new_n14304, new_n6252, new_n14306);
xnor_4 g11958(new_n14271_1, new_n14248, new_n14307);
nand_5 g11959(new_n14307, new_n6259, new_n14308);
xnor_4 g11960(new_n14307, new_n6258, new_n14309);
not_8  g11961(new_n6263, new_n14310_1);
xnor_4 g11962(new_n14269, new_n14251, new_n14311);
nor_5  g11963(new_n14311, new_n14310_1, new_n14312);
xnor_4 g11964(new_n14311, new_n6263, new_n14313);
not_8  g11965(new_n14313, new_n14314);
not_8  g11966(new_n6269, new_n14315);
xnor_4 g11967(new_n14267_1, new_n14254, new_n14316);
nor_5  g11968(new_n14316, new_n14315, new_n14317);
xnor_4 g11969(new_n14316, new_n6269, new_n14318);
not_8  g11970(new_n14318, new_n14319);
xnor_4 g11971(new_n14265, new_n14257, new_n14320);
nor_5  g11972(new_n14320, new_n6277, new_n14321);
xnor_4 g11973(new_n14320, new_n6276_1, new_n14322);
not_8  g11974(new_n14322, new_n14323_1);
xnor_4 g11975(n18578, new_n11572, new_n14324);
nor_5  g11976(new_n14324, new_n6283, new_n14325);
nor_5  g11977(new_n14325, new_n6286, new_n14326_1);
xnor_4 g11978(new_n14262, new_n14261, new_n14327);
not_8  g11979(new_n14326_1, new_n14328);
not_8  g11980(new_n6218_1, new_n14329);
nand_5 g11981(new_n14325, new_n14329, new_n14330);
nand_5 g11982(new_n14330, new_n14328, new_n14331);
nor_5  g11983(new_n14331, new_n14327, new_n14332);
nor_5  g11984(new_n14332, new_n14326_1, new_n14333);
nor_5  g11985(new_n14333, new_n14323_1, new_n14334);
nor_5  g11986(new_n14334, new_n14321, new_n14335);
nor_5  g11987(new_n14335, new_n14319, new_n14336);
nor_5  g11988(new_n14336, new_n14317, new_n14337);
nor_5  g11989(new_n14337, new_n14314, new_n14338);
nor_5  g11990(new_n14338, new_n14312, new_n14339);
nand_5 g11991(new_n14339, new_n14309, new_n14340);
nand_5 g11992(new_n14340, new_n14308, new_n14341);
nand_5 g11993(new_n14341, new_n14306, new_n14342_1);
nand_5 g11994(new_n14342_1, new_n14305, new_n14343);
nand_5 g11995(new_n14343, new_n14303, new_n14344);
nand_5 g11996(new_n14344, new_n14302, new_n14345_1);
nand_5 g11997(new_n14345_1, new_n14299, new_n14346);
nand_5 g11998(new_n14346, new_n14297, new_n14347);
nand_5 g11999(new_n14347, new_n14294_1, new_n14348);
nand_5 g12000(new_n14348, new_n14292, new_n14349);
nand_5 g12001(new_n14349, new_n14289, new_n14350);
nand_5 g12002(new_n14350, new_n14288, new_n14351);
not_8  g12003(new_n14351, new_n14352);
xnor_4 g12004(new_n14349, new_n14289, new_n14353_1);
not_8  g12005(new_n14353_1, new_n14354);
not_8  g12006(n2743, new_n14355);
or_5   g12007(n3506, new_n14355, new_n14356);
nand_5 g12008(new_n3721, new_n3674, new_n14357);
nand_5 g12009(new_n14357, new_n14356, new_n14358);
not_8  g12010(new_n14358, new_n14359);
nand_5 g12011(new_n14359, new_n14354, new_n14360);
xnor_4 g12012(new_n14359, new_n14353_1, new_n14361);
not_8  g12013(new_n3722, new_n14362);
xnor_4 g12014(new_n14347, new_n14294_1, new_n14363);
not_8  g12015(new_n14363, new_n14364_1);
nand_5 g12016(new_n14364_1, new_n14362, new_n14365);
xnor_4 g12017(new_n14363, new_n14362, new_n14366);
xnor_4 g12018(new_n14345_1, new_n14299, new_n14367);
not_8  g12019(new_n14367, new_n14368);
nand_5 g12020(new_n14368, new_n3739, new_n14369);
xnor_4 g12021(new_n14367, new_n3739, new_n14370);
not_8  g12022(new_n3745, new_n14371);
xnor_4 g12023(new_n14343, new_n14303, new_n14372);
not_8  g12024(new_n14372, new_n14373);
nand_5 g12025(new_n14373, new_n14371, new_n14374);
xnor_4 g12026(new_n14372, new_n14371, new_n14375_1);
not_8  g12027(new_n3751, new_n14376);
not_8  g12028(new_n14306, new_n14377);
xnor_4 g12029(new_n14341, new_n14377, new_n14378);
nand_5 g12030(new_n14378, new_n14376, new_n14379);
xnor_4 g12031(new_n14378, new_n3751, new_n14380);
not_8  g12032(new_n3756, new_n14381);
not_8  g12033(new_n14309, new_n14382);
xnor_4 g12034(new_n14339, new_n14382, new_n14383);
nand_5 g12035(new_n14383, new_n14381, new_n14384);
xnor_4 g12036(new_n14383, new_n3756, new_n14385);
xnor_4 g12037(new_n14337, new_n14314, new_n14386);
nand_5 g12038(new_n14386, new_n3764, new_n14387);
xnor_4 g12039(new_n14386, new_n3765, new_n14388);
xnor_4 g12040(new_n14335, new_n14318, new_n14389);
nor_5  g12041(new_n14389, new_n3771, new_n14390);
xnor_4 g12042(new_n14389, new_n3771, new_n14391);
xnor_4 g12043(new_n14333, new_n14322, new_n14392);
nor_5  g12044(new_n14392, new_n3776, new_n14393);
xnor_4 g12045(new_n14392, new_n3776, new_n14394);
xnor_4 g12046(new_n14331, new_n14327, new_n14395);
not_8  g12047(new_n14395, new_n14396);
nor_5  g12048(new_n14396, new_n3783, new_n14397);
xnor_4 g12049(new_n14324, new_n6282, new_n14398);
not_8  g12050(new_n14398, new_n14399);
nor_5  g12051(new_n14399, new_n3785_1, new_n14400);
not_8  g12052(new_n14400, new_n14401);
xnor_4 g12053(new_n14395, new_n3783, new_n14402);
not_8  g12054(new_n14402, new_n14403);
nor_5  g12055(new_n14403, new_n14401, new_n14404);
nor_5  g12056(new_n14404, new_n14397, new_n14405);
nor_5  g12057(new_n14405, new_n14394, new_n14406);
nor_5  g12058(new_n14406, new_n14393, new_n14407);
nor_5  g12059(new_n14407, new_n14391, new_n14408);
nor_5  g12060(new_n14408, new_n14390, new_n14409);
not_8  g12061(new_n14409, new_n14410);
nand_5 g12062(new_n14410, new_n14388, new_n14411);
nand_5 g12063(new_n14411, new_n14387, new_n14412_1);
nand_5 g12064(new_n14412_1, new_n14385, new_n14413);
nand_5 g12065(new_n14413, new_n14384, new_n14414_1);
nand_5 g12066(new_n14414_1, new_n14380, new_n14415);
nand_5 g12067(new_n14415, new_n14379, new_n14416);
nand_5 g12068(new_n14416, new_n14375_1, new_n14417);
nand_5 g12069(new_n14417, new_n14374, new_n14418);
nand_5 g12070(new_n14418, new_n14370, new_n14419);
nand_5 g12071(new_n14419, new_n14369, new_n14420);
nand_5 g12072(new_n14420, new_n14366, new_n14421);
nand_5 g12073(new_n14421, new_n14365, new_n14422);
nand_5 g12074(new_n14422, new_n14361, new_n14423);
nand_5 g12075(new_n14423, new_n14360, new_n14424);
xnor_4 g12076(new_n14424, new_n14352, n2561);
xor_4  g12077(new_n8949, new_n8947, n2573);
xnor_4 g12078(n18558, n10411, new_n14427);
nor_5  g12079(new_n2705, n7149, new_n14428);
nor_5  g12080(n16971, new_n2742, new_n14429);
nor_5  g12081(n14148, new_n2801, new_n14430);
nor_5  g12082(new_n2919, n11503, new_n14431);
nor_5  g12083(new_n10717, n1152, new_n14432);
not_8  g12084(new_n14432, new_n14433);
nor_5  g12085(new_n14433, new_n14431, new_n14434);
nor_5  g12086(new_n14434, new_n14430, new_n14435);
nor_5  g12087(new_n14435, new_n14429, new_n14436);
nor_5  g12088(new_n14436, new_n14428, new_n14437);
xnor_4 g12089(new_n14437, new_n14427, new_n14438);
nor_5  g12090(n7963, new_n10521, new_n14439);
nor_5  g12091(new_n10522, n6590, new_n14440_1);
nor_5  g12092(new_n10525_1, n10017, new_n14441);
nor_5  g12093(n20349, new_n10524, new_n14442);
nand_5 g12094(n15936, new_n11698, new_n14443);
nor_5  g12095(new_n14443, new_n14442, new_n14444);
nor_5  g12096(new_n14444, new_n14441, new_n14445);
nor_5  g12097(new_n14445, new_n14440_1, new_n14446);
nor_5  g12098(new_n14446, new_n14439, new_n14447);
xnor_4 g12099(new_n14447, new_n10574, new_n14448);
xnor_4 g12100(new_n14448, new_n14438, new_n14449);
xnor_4 g12101(n16971, n7149, new_n14450);
xnor_4 g12102(new_n14450, new_n14435, new_n14451);
xnor_4 g12103(new_n14445, new_n10579, new_n14452);
nor_5  g12104(new_n14452, new_n14451, new_n14453);
not_8  g12105(new_n14452, new_n14454);
xnor_4 g12106(new_n14454, new_n14451, new_n14455);
xnor_4 g12107(n18151, n1152, new_n14456);
nor_5  g12108(new_n14456, new_n10587, new_n14457_1);
xnor_4 g12109(n14148, n11503, new_n14458);
xnor_4 g12110(new_n14458, new_n14433, new_n14459);
not_8  g12111(new_n14459, new_n14460);
nor_5  g12112(new_n14460, new_n14457_1, new_n14461);
xnor_4 g12113(new_n14459, new_n14457_1, new_n14462);
not_8  g12114(new_n14462, new_n14463);
xnor_4 g12115(new_n14443, new_n10583, new_n14464_1);
nor_5  g12116(new_n14464_1, new_n14463, new_n14465);
nor_5  g12117(new_n14465, new_n14461, new_n14466);
nand_5 g12118(new_n14466, new_n14455, new_n14467);
not_8  g12119(new_n14467, new_n14468);
nor_5  g12120(new_n14468, new_n14453, new_n14469);
xnor_4 g12121(new_n14469, new_n14449, new_n14470);
xnor_4 g12122(n19515, n17035, new_n14471_1);
not_8  g12123(n22588, new_n14472);
nor_5  g12124(new_n14472, n14684, new_n14473);
nor_5  g12125(n22588, new_n4353, new_n14474);
not_8  g12126(n12209, new_n14475_1);
nor_5  g12127(new_n14475_1, n6631, new_n14476);
nor_5  g12128(n12209, new_n8975, new_n14477);
nand_5 g12129(new_n4488, n12892, new_n14478);
nor_5  g12130(new_n14478, new_n14477, new_n14479);
nor_5  g12131(new_n14479, new_n14476, new_n14480);
nor_5  g12132(new_n14480, new_n14474, new_n14481);
nor_5  g12133(new_n14481, new_n14473, new_n14482);
xnor_4 g12134(new_n14482, new_n14471_1, new_n14483);
xnor_4 g12135(new_n14483, new_n14470, new_n14484);
xnor_4 g12136(new_n14466, new_n14455, new_n14485);
not_8  g12137(new_n14485, new_n14486);
xnor_4 g12138(n22588, n14684, new_n14487);
xnor_4 g12139(new_n14487, new_n14480, new_n14488);
not_8  g12140(new_n14488, new_n14489);
nor_5  g12141(new_n14489, new_n14486, new_n14490);
xnor_4 g12142(n24732, n12892, new_n14491);
not_8  g12143(new_n10587, new_n14492);
xnor_4 g12144(new_n14456, new_n14492, new_n14493);
not_8  g12145(new_n14493, new_n14494);
nor_5  g12146(new_n14494, new_n14491, new_n14495);
xnor_4 g12147(n12209, n6631, new_n14496);
xnor_4 g12148(new_n14496, new_n14478, new_n14497);
not_8  g12149(new_n14497, new_n14498);
nor_5  g12150(new_n14498, new_n14495, new_n14499);
xnor_4 g12151(new_n14497, new_n14495, new_n14500);
not_8  g12152(new_n14500, new_n14501);
xnor_4 g12153(new_n14464_1, new_n14462, new_n14502);
not_8  g12154(new_n14502, new_n14503);
nor_5  g12155(new_n14503, new_n14501, new_n14504);
nor_5  g12156(new_n14504, new_n14499, new_n14505);
xnor_4 g12157(new_n14489, new_n14485, new_n14506);
not_8  g12158(new_n14506, new_n14507);
nor_5  g12159(new_n14507, new_n14505, new_n14508);
nor_5  g12160(new_n14508, new_n14490, new_n14509);
not_8  g12161(new_n14509, new_n14510_1);
xnor_4 g12162(new_n14510_1, new_n14484, n2578);
not_8  g12163(new_n8331, new_n14512);
nor_5  g12164(new_n12482, new_n14512, new_n14513);
xnor_4 g12165(new_n12482, new_n8331, new_n14514);
not_8  g12166(new_n14514, new_n14515);
nor_5  g12167(new_n8331, new_n8266, new_n14516);
nor_5  g12168(new_n8414, new_n8332, new_n14517);
nor_5  g12169(new_n14517, new_n14516, new_n14518);
nor_5  g12170(new_n14518, new_n14515, new_n14519);
nor_5  g12171(new_n14519, new_n14513, n2582);
xor_4  g12172(new_n4495, new_n4480, n2602);
nor_5  g12173(n22201, n2420, new_n14522);
nand_5 g12174(new_n14522, new_n8601, new_n14523);
nor_5  g12175(new_n14523, n21078, new_n14524);
nand_5 g12176(new_n14524, new_n8593, new_n14525);
xnor_4 g12177(new_n14525, new_n8589, new_n14526);
not_8  g12178(new_n14526, new_n14527);
xnor_4 g12179(new_n14527, new_n4133, new_n14528);
xnor_4 g12180(new_n14524, n12546, new_n14529);
not_8  g12181(new_n14529, new_n14530);
nand_5 g12182(new_n14530, new_n4692, new_n14531);
xnor_4 g12183(new_n14523, new_n8597, new_n14532);
not_8  g12184(new_n14532, new_n14533);
nand_5 g12185(new_n14533, new_n4140, new_n14534);
xnor_4 g12186(new_n14533, new_n4139, new_n14535);
xnor_4 g12187(new_n14522, new_n8601, new_n14536);
nor_5  g12188(new_n14536, new_n4146_1, new_n14537);
xnor_4 g12189(new_n14536, new_n4146_1, new_n14538);
xnor_4 g12190(new_n8612, n2420, new_n14539);
nor_5  g12191(new_n14539, new_n4151_1, new_n14540);
not_8  g12192(new_n14540, new_n14541_1);
nor_5  g12193(new_n4154, new_n8612, new_n14542);
not_8  g12194(new_n14542, new_n14543);
xnor_4 g12195(new_n14539, new_n4152_1, new_n14544);
nand_5 g12196(new_n14544, new_n14543, new_n14545);
nand_5 g12197(new_n14545, new_n14541_1, new_n14546_1);
nor_5  g12198(new_n14546_1, new_n14538, new_n14547_1);
nor_5  g12199(new_n14547_1, new_n14537, new_n14548);
nand_5 g12200(new_n14548, new_n14535, new_n14549);
nand_5 g12201(new_n14549, new_n14534, new_n14550);
xnor_4 g12202(new_n14530, new_n4135, new_n14551);
nand_5 g12203(new_n14551, new_n14550, new_n14552);
nand_5 g12204(new_n14552, new_n14531, new_n14553);
xnor_4 g12205(new_n14553, new_n14528, new_n14554);
xnor_4 g12206(new_n8590, new_n4564, new_n14555);
nand_5 g12207(new_n8594_1, new_n4568, new_n14556);
xnor_4 g12208(new_n8594_1, n3785, new_n14557);
nand_5 g12209(new_n8598, new_n4573, new_n14558);
xnor_4 g12210(new_n8598, n20250, new_n14559);
nor_5  g12211(new_n8603, new_n4577, new_n14560);
nor_5  g12212(new_n8605, n5822, new_n14561);
nor_5  g12213(new_n8609, n26443, new_n14562);
nor_5  g12214(new_n2571, new_n2568, new_n14563);
xnor_4 g12215(new_n8608_1, n26443, new_n14564);
not_8  g12216(new_n14564, new_n14565);
nor_5  g12217(new_n14565, new_n14563, new_n14566);
nor_5  g12218(new_n14566, new_n14562, new_n14567);
not_8  g12219(new_n14567, new_n14568);
nor_5  g12220(new_n14568, new_n14561, new_n14569);
nor_5  g12221(new_n14569, new_n14560, new_n14570_1);
nand_5 g12222(new_n14570_1, new_n14559, new_n14571);
nand_5 g12223(new_n14571, new_n14558, new_n14572);
nand_5 g12224(new_n14572, new_n14557, new_n14573);
nand_5 g12225(new_n14573, new_n14556, new_n14574);
xnor_4 g12226(new_n14574, new_n14555, new_n14575_1);
xnor_4 g12227(new_n14575_1, new_n14554, new_n14576_1);
xnor_4 g12228(new_n14572, new_n14557, new_n14577);
not_8  g12229(new_n14577, new_n14578);
not_8  g12230(new_n14551, new_n14579);
xnor_4 g12231(new_n14579, new_n14550, new_n14580);
nand_5 g12232(new_n14580, new_n14578, new_n14581);
xnor_4 g12233(new_n14580, new_n14577, new_n14582);
xnor_4 g12234(new_n14548, new_n14535, new_n14583);
not_8  g12235(new_n14583, new_n14584);
not_8  g12236(new_n14559, new_n14585);
xnor_4 g12237(new_n14570_1, new_n14585, new_n14586);
nand_5 g12238(new_n14586, new_n14584, new_n14587);
xnor_4 g12239(new_n14586, new_n14583, new_n14588);
xnor_4 g12240(new_n14546_1, new_n14538, new_n14589);
xnor_4 g12241(new_n8603, n5822, new_n14590);
xnor_4 g12242(new_n14590, new_n14568, new_n14591);
not_8  g12243(new_n14591, new_n14592);
nor_5  g12244(new_n14592, new_n14589, new_n14593_1);
xnor_4 g12245(new_n14544, new_n14543, new_n14594);
xnor_4 g12246(new_n14564, new_n14563, new_n14595);
not_8  g12247(new_n14595, new_n14596);
nor_5  g12248(new_n14596, new_n14594, new_n14597);
not_8  g12249(new_n14597, new_n14598);
xnor_4 g12250(new_n2571, n1681, new_n14599);
not_8  g12251(new_n14599, new_n14600);
xnor_4 g12252(new_n2581, new_n8612, new_n14601);
not_8  g12253(new_n14601, new_n14602);
nor_5  g12254(new_n14602, new_n14600, new_n14603_1);
not_8  g12255(new_n14603_1, new_n14604);
xnor_4 g12256(new_n14595, new_n14594, new_n14605);
nand_5 g12257(new_n14605, new_n14604, new_n14606);
nand_5 g12258(new_n14606, new_n14598, new_n14607);
xnor_4 g12259(new_n14592, new_n14589, new_n14608);
nor_5  g12260(new_n14608, new_n14607, new_n14609);
nor_5  g12261(new_n14609, new_n14593_1, new_n14610);
nand_5 g12262(new_n14610, new_n14588, new_n14611);
nand_5 g12263(new_n14611, new_n14587, new_n14612);
nand_5 g12264(new_n14612, new_n14582, new_n14613);
nand_5 g12265(new_n14613, new_n14581, new_n14614);
xnor_4 g12266(new_n14614, new_n14576_1, n2619);
nor_5  g12267(new_n6238, n12900, new_n14616);
xnor_4 g12268(new_n6238, new_n14239, new_n14617);
not_8  g12269(new_n14617, new_n14618);
nor_5  g12270(new_n6244, n20411, new_n14619);
xnor_4 g12271(new_n6245_1, n20411, new_n14620);
not_8  g12272(new_n14620, new_n14621);
nor_5  g12273(new_n6250, n17069, new_n14622);
xnor_4 g12274(new_n6250, new_n14245, new_n14623);
not_8  g12275(new_n14623, new_n14624);
nor_5  g12276(new_n6256_1, n15918, new_n14625);
nor_5  g12277(new_n6262, n17784, new_n14626);
xnor_4 g12278(new_n6262, new_n13361, new_n14627);
not_8  g12279(new_n14627, new_n14628);
nor_5  g12280(new_n6272, new_n13879, new_n14629);
not_8  g12281(new_n14629, new_n14630);
nand_5 g12282(new_n13893, new_n13880, new_n14631);
nand_5 g12283(new_n14631, new_n14630, new_n14632);
nor_5  g12284(new_n14632, new_n14628, new_n14633_1);
nor_5  g12285(new_n14633_1, new_n14626, new_n14634);
xnor_4 g12286(new_n6256_1, new_n13357, new_n14635);
not_8  g12287(new_n14635, new_n14636_1);
nor_5  g12288(new_n14636_1, new_n14634, new_n14637);
nor_5  g12289(new_n14637, new_n14625, new_n14638);
nor_5  g12290(new_n14638, new_n14624, new_n14639);
nor_5  g12291(new_n14639, new_n14622, new_n14640);
nor_5  g12292(new_n14640, new_n14621, new_n14641);
nor_5  g12293(new_n14641, new_n14619, new_n14642);
nor_5  g12294(new_n14642, new_n14618, new_n14643);
nor_5  g12295(new_n14643, new_n14616, new_n14644);
xnor_4 g12296(new_n6186, n10650, new_n14645);
xnor_4 g12297(new_n14645, new_n14644, new_n14646);
not_8  g12298(new_n14646, new_n14647);
nor_5  g12299(new_n14647, n6456, new_n14648);
not_8  g12300(new_n14648, new_n14649);
xnor_4 g12301(new_n14646, n6456, new_n14650);
xnor_4 g12302(new_n14642, new_n14618, new_n14651);
nor_5  g12303(new_n14651, n4085, new_n14652);
not_8  g12304(new_n14652, new_n14653);
xnor_4 g12305(new_n14651, new_n6191, new_n14654);
xnor_4 g12306(new_n14640, new_n14621, new_n14655);
nor_5  g12307(new_n14655, n26725, new_n14656);
not_8  g12308(new_n14656, new_n14657);
xnor_4 g12309(new_n14655, n26725, new_n14658);
xnor_4 g12310(new_n14638, new_n14623, new_n14659);
not_8  g12311(new_n14659, new_n14660);
nor_5  g12312(new_n14660, n11980, new_n14661);
xnor_4 g12313(new_n14659, new_n6196, new_n14662);
xnor_4 g12314(new_n14635, new_n14634, new_n14663);
not_8  g12315(new_n14663, new_n14664);
nor_5  g12316(new_n14664, n3253, new_n14665);
xnor_4 g12317(new_n14663, new_n6200, new_n14666);
xnor_4 g12318(new_n14632, new_n14627, new_n14667);
nor_5  g12319(new_n14667, new_n6204_1, new_n14668);
not_8  g12320(new_n14668, new_n14669);
xnor_4 g12321(new_n14667, n7759, new_n14670);
nor_5  g12322(new_n13894, new_n6208, new_n14671);
not_8  g12323(new_n14671, new_n14672);
nand_5 g12324(new_n13911, new_n13895, new_n14673);
nand_5 g12325(new_n14673, new_n14672, new_n14674);
nand_5 g12326(new_n14674, new_n14670, new_n14675);
nand_5 g12327(new_n14675, new_n14669, new_n14676);
nor_5  g12328(new_n14676, new_n14666, new_n14677);
nor_5  g12329(new_n14677, new_n14665, new_n14678);
nor_5  g12330(new_n14678, new_n14662, new_n14679);
nor_5  g12331(new_n14679, new_n14661, new_n14680_1);
nor_5  g12332(new_n14680_1, new_n14658, new_n14681);
not_8  g12333(new_n14681, new_n14682);
nand_5 g12334(new_n14682, new_n14657, new_n14683);
nand_5 g12335(new_n14683, new_n14654, new_n14684_1);
nand_5 g12336(new_n14684_1, new_n14653, new_n14685);
nand_5 g12337(new_n14685, new_n14650, new_n14686);
nand_5 g12338(new_n14686, new_n14649, new_n14687);
not_8  g12339(new_n14644, new_n14688);
nor_5  g12340(new_n6187, n10650, new_n14689);
nor_5  g12341(new_n14689, new_n14688, new_n14690);
nor_5  g12342(new_n6185, n2979, new_n14691);
nor_5  g12343(new_n6186, new_n13343, new_n14692_1);
nor_5  g12344(new_n14692_1, new_n14691, new_n14693);
not_8  g12345(new_n14693, new_n14694);
nor_5  g12346(new_n14694, new_n14690, new_n14695);
not_8  g12347(new_n14695, new_n14696);
nor_5  g12348(new_n14696, new_n14687, new_n14697);
not_8  g12349(new_n14697, new_n14698);
nand_5 g12350(new_n14698, new_n13596, new_n14699);
xnor_4 g12351(new_n14697, new_n13596, new_n14700);
not_8  g12352(new_n13599, new_n14701_1);
xnor_4 g12353(new_n14695, new_n14687, new_n14702_1);
not_8  g12354(new_n14702_1, new_n14703);
nand_5 g12355(new_n14703, new_n14701_1, new_n14704_1);
xnor_4 g12356(new_n14703, new_n13599, new_n14705);
xnor_4 g12357(new_n14685, new_n14650, new_n14706);
not_8  g12358(new_n14706, new_n14707);
nand_5 g12359(new_n14707, new_n13604, new_n14708);
xnor_4 g12360(new_n14706, new_n13604, new_n14709);
xnor_4 g12361(new_n14683, new_n14654, new_n14710);
not_8  g12362(new_n14710, new_n14711);
nand_5 g12363(new_n14711, new_n13609, new_n14712);
xnor_4 g12364(new_n14710, new_n13609, new_n14713);
xnor_4 g12365(new_n14680_1, new_n14658, new_n14714);
not_8  g12366(new_n14714, new_n14715);
nand_5 g12367(new_n14715, new_n13614, new_n14716);
xnor_4 g12368(new_n14714, new_n13614, new_n14717);
xnor_4 g12369(new_n14678, new_n14662, new_n14718);
not_8  g12370(new_n14718, new_n14719);
nand_5 g12371(new_n14719, new_n13619, new_n14720);
xnor_4 g12372(new_n14718, new_n13619, new_n14721);
xnor_4 g12373(new_n14676, new_n14666, new_n14722);
not_8  g12374(new_n14722, new_n14723);
nand_5 g12375(new_n14723, new_n13624, new_n14724);
xnor_4 g12376(new_n14722, new_n13624, new_n14725);
xnor_4 g12377(new_n14674, new_n14670, new_n14726);
nand_5 g12378(new_n14726, new_n13631, new_n14727);
xnor_4 g12379(new_n14726, new_n13630, new_n14728);
nand_5 g12380(new_n13912_1, new_n13636, new_n14729);
nand_5 g12381(new_n13929, new_n13914_1, new_n14730);
nand_5 g12382(new_n14730, new_n14729, new_n14731);
nand_5 g12383(new_n14731, new_n14728, new_n14732);
nand_5 g12384(new_n14732, new_n14727, new_n14733);
nand_5 g12385(new_n14733, new_n14725, new_n14734_1);
nand_5 g12386(new_n14734_1, new_n14724, new_n14735);
nand_5 g12387(new_n14735, new_n14721, new_n14736);
nand_5 g12388(new_n14736, new_n14720, new_n14737);
nand_5 g12389(new_n14737, new_n14717, new_n14738);
nand_5 g12390(new_n14738, new_n14716, new_n14739);
nand_5 g12391(new_n14739, new_n14713, new_n14740);
nand_5 g12392(new_n14740, new_n14712, new_n14741);
nand_5 g12393(new_n14741, new_n14709, new_n14742);
nand_5 g12394(new_n14742, new_n14708, new_n14743);
nand_5 g12395(new_n14743, new_n14705, new_n14744);
nand_5 g12396(new_n14744, new_n14704_1, new_n14745);
nand_5 g12397(new_n14745, new_n14700, new_n14746_1);
nand_5 g12398(new_n14746_1, new_n14699, new_n14747);
not_8  g12399(new_n14747, n2661);
xnor_4 g12400(new_n11884, new_n11883, n2693);
xnor_4 g12401(new_n14438, new_n12888, new_n14750);
not_8  g12402(new_n14451, new_n14751);
nand_5 g12403(new_n14751, new_n12893, new_n14752);
xnor_4 g12404(new_n14451, new_n12893, new_n14753);
nand_5 g12405(new_n14460, new_n7741, new_n14754);
nor_5  g12406(new_n14456, new_n7744, new_n14755);
xnor_4 g12407(new_n14459, new_n7741, new_n14756);
nand_5 g12408(new_n14756, new_n14755, new_n14757);
nand_5 g12409(new_n14757, new_n14754, new_n14758);
nand_5 g12410(new_n14758, new_n14753, new_n14759);
nand_5 g12411(new_n14759, new_n14752, new_n14760);
xnor_4 g12412(new_n14760, new_n14750, new_n14761);
xnor_4 g12413(n8309, n4665, new_n14762);
nor_5  g12414(new_n9310, n19005, new_n14763_1);
nor_5  g12415(n19144, new_n2917, new_n14764);
nor_5  g12416(new_n9315, n4326, new_n14765);
not_8  g12417(new_n14765, new_n14766);
nor_5  g12418(n12593, new_n2921, new_n14767);
not_8  g12419(new_n14767, new_n14768);
nor_5  g12420(new_n12858, n5438, new_n14769);
nand_5 g12421(new_n14769, new_n14768, new_n14770);
nand_5 g12422(new_n14770, new_n14766, new_n14771);
not_8  g12423(new_n14771, new_n14772_1);
nor_5  g12424(new_n14772_1, new_n14764, new_n14773);
nor_5  g12425(new_n14773, new_n14763_1, new_n14774);
xnor_4 g12426(new_n14774, new_n14762, new_n14775);
not_8  g12427(new_n14775, new_n14776);
xnor_4 g12428(new_n14776, new_n14761, new_n14777);
xnor_4 g12429(new_n14758, new_n14753, new_n14778);
xnor_4 g12430(n19144, n19005, new_n14779);
xnor_4 g12431(new_n14779, new_n14772_1, new_n14780);
nand_5 g12432(new_n14780, new_n14778, new_n14781);
xnor_4 g12433(new_n14780, new_n14778, new_n14782);
not_8  g12434(new_n14782, new_n14783);
xnor_4 g12435(n13714, n5438, new_n14784);
xnor_4 g12436(new_n14456, new_n7854, new_n14785);
not_8  g12437(new_n14785, new_n14786);
nor_5  g12438(new_n14786, new_n14784, new_n14787);
xnor_4 g12439(n12593, n4326, new_n14788);
xnor_4 g12440(new_n14788, new_n14769, new_n14789);
nor_5  g12441(new_n14789, new_n14787, new_n14790_1);
xnor_4 g12442(new_n14756, new_n14755, new_n14791);
not_8  g12443(new_n14791, new_n14792);
xnor_4 g12444(new_n14789, new_n14787, new_n14793);
nor_5  g12445(new_n14793, new_n14792, new_n14794);
nor_5  g12446(new_n14794, new_n14790_1, new_n14795);
not_8  g12447(new_n14795, new_n14796);
nand_5 g12448(new_n14796, new_n14783, new_n14797);
nand_5 g12449(new_n14797, new_n14781, new_n14798);
xnor_4 g12450(new_n14798, new_n14777, n2703);
xnor_4 g12451(new_n13738, new_n13725, n2706);
nor_5  g12452(n3320, new_n6478, new_n14801_1);
xnor_4 g12453(n3320, n1831, new_n14802);
not_8  g12454(new_n14802, new_n14803);
not_8  g12455(n13137, new_n14804);
nor_5  g12456(new_n14804, n1288, new_n14805);
xnor_4 g12457(n13137, n1288, new_n14806);
not_8  g12458(new_n14806, new_n14807);
not_8  g12459(n18452, new_n14808);
nor_5  g12460(new_n14808, n1752, new_n14809);
xnor_4 g12461(n18452, n1752, new_n14810);
not_8  g12462(new_n14810, new_n14811);
not_8  g12463(n21317, new_n14812);
nor_5  g12464(new_n14812, n13110, new_n14813);
xnor_4 g12465(n21317, n13110, new_n14814);
not_8  g12466(new_n14814, new_n14815);
nor_5  g12467(n25694, new_n4169, new_n14816);
xnor_4 g12468(n25694, n12398, new_n14817);
not_8  g12469(new_n14817, new_n14818);
nor_5  g12470(new_n4170, n15424, new_n14819_1);
xnor_4 g12471(n19789, n15424, new_n14820);
nor_5  g12472(n20169, new_n4190, new_n14821);
not_8  g12473(new_n12961, new_n14822);
nor_5  g12474(new_n12971, new_n14822, new_n14823);
nor_5  g12475(new_n14823, new_n14821, new_n14824);
and_5  g12476(new_n14824, new_n14820, new_n14825);
nor_5  g12477(new_n14825, new_n14819_1, new_n14826_1);
nor_5  g12478(new_n14826_1, new_n14818, new_n14827_1);
nor_5  g12479(new_n14827_1, new_n14816, new_n14828);
nor_5  g12480(new_n14828, new_n14815, new_n14829);
nor_5  g12481(new_n14829, new_n14813, new_n14830);
nor_5  g12482(new_n14830, new_n14811, new_n14831);
nor_5  g12483(new_n14831, new_n14809, new_n14832);
nor_5  g12484(new_n14832, new_n14807, new_n14833);
nor_5  g12485(new_n14833, new_n14805, new_n14834);
nor_5  g12486(new_n14834, new_n14803, new_n14835);
nor_5  g12487(new_n14835, new_n14801_1, new_n14836);
not_8  g12488(new_n14836, new_n14837);
not_8  g12489(n1483, new_n14838);
or_5   g12490(n19539, new_n14838, new_n14839_1);
nand_5 g12491(new_n11992, new_n11978, new_n14840);
nand_5 g12492(new_n14840, new_n14839_1, new_n14841);
not_8  g12493(new_n14841, new_n14842);
not_8  g12494(new_n11993, new_n14843);
nand_5 g12495(new_n6812, new_n13120, new_n14844);
nor_5  g12496(new_n14844, n3541, new_n14845);
xnor_4 g12497(new_n14845, n2184, new_n14846);
not_8  g12498(new_n14846, new_n14847);
nand_5 g12499(new_n14847, new_n13069, new_n14848);
xnor_4 g12500(new_n14846, new_n13069, new_n14849_1);
xnor_4 g12501(new_n14844, new_n13117, new_n14850);
not_8  g12502(new_n14850, new_n14851);
nor_5  g12503(new_n14851, new_n13072, new_n14852);
nor_5  g12504(new_n14850, n3349, new_n14853);
not_8  g12505(new_n6813, new_n14854);
nor_5  g12506(new_n14854, new_n6805, new_n14855);
nor_5  g12507(new_n6813, n1742, new_n14856);
nor_5  g12508(new_n6851, new_n14856, new_n14857);
nor_5  g12509(new_n14857, new_n14855, new_n14858);
nor_5  g12510(new_n14858, new_n14853, new_n14859);
nor_5  g12511(new_n14859, new_n14852, new_n14860);
nand_5 g12512(new_n14860, new_n14849_1, new_n14861);
nand_5 g12513(new_n14861, new_n14848, new_n14862);
nand_5 g12514(new_n14845, new_n13114, new_n14863);
xnor_4 g12515(new_n14863, new_n13160, new_n14864);
xnor_4 g12516(new_n14864, new_n13066, new_n14865);
xnor_4 g12517(new_n14865, new_n14862, new_n14866);
nor_5  g12518(new_n14866, new_n14843, new_n14867);
xnor_4 g12519(new_n14866, new_n14843, new_n14868);
xnor_4 g12520(new_n14860, new_n14849_1, new_n14869);
nor_5  g12521(new_n14869, new_n12059, new_n14870);
xnor_4 g12522(new_n14869, new_n12059, new_n14871);
not_8  g12523(new_n12064, new_n14872);
xnor_4 g12524(new_n14850, new_n13072, new_n14873);
xnor_4 g12525(new_n14873, new_n14858, new_n14874);
nand_5 g12526(new_n14874, new_n14872, new_n14875);
xnor_4 g12527(new_n14874, new_n12064, new_n14876);
not_8  g12528(new_n6852, new_n14877);
nor_5  g12529(new_n14877, new_n6804, new_n14878);
not_8  g12530(new_n14878, new_n14879);
nand_5 g12531(new_n6901, new_n6853_1, new_n14880);
nand_5 g12532(new_n14880, new_n14879, new_n14881);
nand_5 g12533(new_n14881, new_n14876, new_n14882);
nand_5 g12534(new_n14882, new_n14875, new_n14883);
nor_5  g12535(new_n14883, new_n14871, new_n14884);
nor_5  g12536(new_n14884, new_n14870, new_n14885);
nor_5  g12537(new_n14885, new_n14868, new_n14886);
nor_5  g12538(new_n14886, new_n14867, new_n14887);
not_8  g12539(new_n14887, new_n14888);
or_5   g12540(new_n14863, n10018, new_n14889);
or_5   g12541(new_n14864, n5140, new_n14890);
nand_5 g12542(new_n14864, n5140, new_n14891_1);
nand_5 g12543(new_n14891_1, new_n14862, new_n14892);
nand_5 g12544(new_n14892, new_n14890, new_n14893);
nand_5 g12545(new_n14893, new_n14889, new_n14894);
not_8  g12546(new_n14894, new_n14895);
nor_5  g12547(new_n14895, new_n14888, new_n14896);
nand_5 g12548(new_n14896, new_n14842, new_n14897);
nor_5  g12549(new_n14894, new_n14887, new_n14898);
nand_5 g12550(new_n14898, new_n14841, new_n14899_1);
nand_5 g12551(new_n14899_1, new_n14897, new_n14900);
xnor_4 g12552(new_n14900, new_n14837, new_n14901);
xnor_4 g12553(new_n14895, new_n14887, new_n14902);
xnor_4 g12554(new_n14902, new_n14841, new_n14903);
nor_5  g12555(new_n14903, new_n14837, new_n14904);
not_8  g12556(new_n14903, new_n14905);
nor_5  g12557(new_n14905, new_n14836, new_n14906);
xnor_4 g12558(new_n14834, new_n14802, new_n14907);
xnor_4 g12559(new_n14885, new_n14868, new_n14908);
nor_5  g12560(new_n14908, new_n14907, new_n14909);
not_8  g12561(new_n14909, new_n14910);
not_8  g12562(new_n14908, new_n14911);
xnor_4 g12563(new_n14911, new_n14907, new_n14912);
xnor_4 g12564(new_n14832, new_n14807, new_n14913);
xnor_4 g12565(new_n14883, new_n14871, new_n14914);
not_8  g12566(new_n14914, new_n14915);
nand_5 g12567(new_n14915, new_n14913, new_n14916);
xnor_4 g12568(new_n14914, new_n14913, new_n14917);
xnor_4 g12569(new_n14830, new_n14810, new_n14918);
not_8  g12570(new_n14918, new_n14919);
xnor_4 g12571(new_n14881, new_n14876, new_n14920);
nand_5 g12572(new_n14920, new_n14919, new_n14921);
xnor_4 g12573(new_n14920, new_n14918, new_n14922);
xnor_4 g12574(new_n14828, new_n14814, new_n14923);
not_8  g12575(new_n14923, new_n14924);
nand_5 g12576(new_n14924, new_n6902, new_n14925);
xnor_4 g12577(new_n14826_1, new_n14817, new_n14926);
not_8  g12578(new_n14926, new_n14927);
nand_5 g12579(new_n14927, new_n6904, new_n14928);
xnor_4 g12580(new_n14926, new_n6904, new_n14929);
xnor_4 g12581(new_n14824, new_n14820, new_n14930);
nand_5 g12582(new_n14930, new_n6908, new_n14931_1);
xnor_4 g12583(new_n14930, new_n6907, new_n14932);
nand_5 g12584(new_n12972, new_n6913, new_n14933);
nand_5 g12585(new_n12992_1, new_n12973, new_n14934);
nand_5 g12586(new_n14934, new_n14933, new_n14935);
nand_5 g12587(new_n14935, new_n14932, new_n14936);
nand_5 g12588(new_n14936, new_n14931_1, new_n14937);
nand_5 g12589(new_n14937, new_n14929, new_n14938);
nand_5 g12590(new_n14938, new_n14928, new_n14939);
xnor_4 g12591(new_n14923, new_n6902, new_n14940);
nand_5 g12592(new_n14940, new_n14939, new_n14941);
nand_5 g12593(new_n14941, new_n14925, new_n14942);
nand_5 g12594(new_n14942, new_n14922, new_n14943);
nand_5 g12595(new_n14943, new_n14921, new_n14944_1);
nand_5 g12596(new_n14944_1, new_n14917, new_n14945);
nand_5 g12597(new_n14945, new_n14916, new_n14946);
nand_5 g12598(new_n14946, new_n14912, new_n14947);
nand_5 g12599(new_n14947, new_n14910, new_n14948);
nor_5  g12600(new_n14948, new_n14906, new_n14949);
nor_5  g12601(new_n14949, new_n14904, new_n14950);
xnor_4 g12602(new_n14950, new_n14901, n2711);
xnor_4 g12603(n10611, n2680, new_n14952);
nor_5  g12604(n2783, new_n9660, new_n14953);
nor_5  g12605(new_n6947, n1667, new_n14954_1);
nor_5  g12606(n15490, new_n9755, new_n14955);
nor_5  g12607(new_n9693, n7339, new_n14956);
nand_5 g12608(n26808, new_n6967_1, new_n14957);
nor_5  g12609(new_n14957, new_n14956, new_n14958);
nor_5  g12610(new_n14958, new_n14955, new_n14959);
nor_5  g12611(new_n14959, new_n14954_1, new_n14960);
nor_5  g12612(new_n14960, new_n14953, new_n14961);
xnor_4 g12613(new_n14961, new_n14952, new_n14962);
xnor_4 g12614(new_n14962, new_n9613, new_n14963);
xnor_4 g12615(n2783, n1667, new_n14964);
xnor_4 g12616(new_n14964, new_n14959, new_n14965);
not_8  g12617(new_n14965, new_n14966);
nor_5  g12618(new_n14966, new_n9617, new_n14967);
not_8  g12619(new_n14967, new_n14968);
xnor_4 g12620(new_n14965, new_n9617, new_n14969);
not_8  g12621(new_n14969, new_n14970);
xnor_4 g12622(n26808, n18, new_n14971);
nor_5  g12623(new_n14971, new_n9626_1, new_n14972);
xnor_4 g12624(n15490, n7339, new_n14973);
xnor_4 g12625(new_n14973, new_n14957, new_n14974);
not_8  g12626(new_n14974, new_n14975);
nor_5  g12627(new_n14975, new_n14972, new_n14976);
xnor_4 g12628(new_n14974, new_n14972, new_n14977_1);
not_8  g12629(new_n14977_1, new_n14978);
nor_5  g12630(new_n14978, new_n9632, new_n14979);
nor_5  g12631(new_n14979, new_n14976, new_n14980);
nor_5  g12632(new_n14980, new_n14970, new_n14981);
not_8  g12633(new_n14981, new_n14982);
nand_5 g12634(new_n14982, new_n14968, new_n14983);
xnor_4 g12635(new_n14983, new_n14963, n2761);
xnor_4 g12636(n25120, new_n6308_1, new_n14985);
or_5   g12637(n8363, n2816, new_n14986);
xnor_4 g12638(n8363, new_n6359, new_n14987);
or_5   g12639(n20359, n14680, new_n14988);
not_8  g12640(n14680, new_n14989_1);
xnor_4 g12641(n20359, new_n14989_1, new_n14990);
nor_5  g12642(n17250, n4409, new_n14991);
not_8  g12643(new_n14991, new_n14992);
not_8  g12644(new_n9937, new_n14993);
nand_5 g12645(new_n14993, new_n9910, new_n14994);
nand_5 g12646(new_n14994, new_n14992, new_n14995);
nand_5 g12647(new_n14995, new_n14990, new_n14996);
nand_5 g12648(new_n14996, new_n14988, new_n14997);
nand_5 g12649(new_n14997, new_n14987, new_n14998);
nand_5 g12650(new_n14998, new_n14986, new_n14999);
xnor_4 g12651(new_n14999, new_n14985, new_n15000);
nor_5  g12652(new_n15000, n17458, new_n15001);
xnor_4 g12653(new_n15000, new_n11675, new_n15002_1);
not_8  g12654(new_n15002_1, new_n15003);
not_8  g12655(new_n14987, new_n15004_1);
xnor_4 g12656(new_n14997, new_n15004_1, new_n15005);
nor_5  g12657(new_n15005, new_n11678, new_n15006);
not_8  g12658(new_n15006, new_n15007);
xnor_4 g12659(new_n14995, new_n14990, new_n15008);
nor_5  g12660(new_n15008, n25240, new_n15009);
not_8  g12661(new_n15009, new_n15010);
xnor_4 g12662(new_n15008, new_n11681, new_n15011_1);
nor_5  g12663(new_n9938_1, new_n7647_1, new_n15012);
xnor_4 g12664(new_n9938_1, new_n7647_1, new_n15013);
nor_5  g12665(new_n9941, new_n7650, new_n15014);
xnor_4 g12666(new_n9941, new_n7650, new_n15015);
nor_5  g12667(new_n9946_1, new_n11178, new_n15016);
xnor_4 g12668(new_n9945, n20923, new_n15017);
nor_5  g12669(new_n9950, new_n11691, new_n15018);
xnor_4 g12670(new_n9950, new_n11691, new_n15019_1);
nor_5  g12671(new_n9954, new_n6982, new_n15020);
nor_5  g12672(new_n9957, n5026, new_n15021);
not_8  g12673(new_n15021, new_n15022);
nor_5  g12674(new_n9961, new_n7664, new_n15023);
not_8  g12675(new_n15023, new_n15024);
xnor_4 g12676(new_n9956, n5026, new_n15025);
nand_5 g12677(new_n15025, new_n15024, new_n15026);
nand_5 g12678(new_n15026, new_n15022, new_n15027);
xnor_4 g12679(new_n9954, new_n6982, new_n15028);
nor_5  g12680(new_n15028, new_n15027, new_n15029);
nor_5  g12681(new_n15029, new_n15020, new_n15030);
nor_5  g12682(new_n15030, new_n15019_1, new_n15031_1);
nor_5  g12683(new_n15031_1, new_n15018, new_n15032);
nor_5  g12684(new_n15032, new_n15017, new_n15033_1);
nor_5  g12685(new_n15033_1, new_n15016, new_n15034);
nor_5  g12686(new_n15034, new_n15015, new_n15035);
nor_5  g12687(new_n15035, new_n15014, new_n15036);
nor_5  g12688(new_n15036, new_n15013, new_n15037);
nor_5  g12689(new_n15037, new_n15012, new_n15038);
nand_5 g12690(new_n15038, new_n15011_1, new_n15039);
nand_5 g12691(new_n15039, new_n15010, new_n15040);
not_8  g12692(new_n15040, new_n15041);
xnor_4 g12693(new_n15005, n1222, new_n15042);
nand_5 g12694(new_n15042, new_n15041, new_n15043);
nand_5 g12695(new_n15043, new_n15007, new_n15044);
nor_5  g12696(new_n15044, new_n15003, new_n15045);
nor_5  g12697(new_n15045, new_n15001, new_n15046);
nor_5  g12698(n25120, n8526, new_n15047);
not_8  g12699(new_n15047, new_n15048);
nand_5 g12700(new_n14999, new_n14985, new_n15049);
nand_5 g12701(new_n15049, new_n15048, new_n15050);
not_8  g12702(new_n15050, new_n15051);
nand_5 g12703(new_n15051, new_n15046, new_n15052_1);
nand_5 g12704(new_n3885, new_n11199, new_n15053_1);
nor_5  g12705(new_n15053_1, n1099, new_n15054);
nand_5 g12706(new_n15054, new_n13683_1, new_n15055);
xnor_4 g12707(new_n15055, new_n13681, new_n15056);
not_8  g12708(new_n15056, new_n15057);
nand_5 g12709(new_n15057, new_n5089, new_n15058);
xnor_4 g12710(new_n15057, new_n5088, new_n15059);
xnor_4 g12711(new_n15054, n19941, new_n15060);
not_8  g12712(new_n15060, new_n15061);
nand_5 g12713(new_n15061, new_n5094, new_n15062);
xnor_4 g12714(new_n15061, new_n5093, new_n15063);
xnor_4 g12715(new_n15053_1, new_n11195, new_n15064);
not_8  g12716(new_n15064, new_n15065);
nand_5 g12717(new_n15065, new_n5097, new_n15066);
xnor_4 g12718(new_n15064, new_n5097, new_n15067);
not_8  g12719(new_n3886, new_n15068);
nand_5 g12720(new_n5102, new_n15068, new_n15069);
xnor_4 g12721(new_n5101_1, new_n15068, new_n15070);
nand_5 g12722(new_n5107, new_n3891_1, new_n15071);
xnor_4 g12723(new_n5106, new_n3891_1, new_n15072);
nor_5  g12724(new_n13807, new_n3895, new_n15073);
not_8  g12725(new_n15073, new_n15074);
xnor_4 g12726(new_n5111, new_n3895, new_n15075);
nor_5  g12727(new_n5114, new_n3901, new_n15076);
not_8  g12728(new_n15076, new_n15077_1);
xnor_4 g12729(new_n5114, new_n3902, new_n15078);
nor_5  g12730(new_n5118, new_n3905, new_n15079);
not_8  g12731(new_n15079, new_n15080);
xnor_4 g12732(new_n5118, new_n3906, new_n15081);
nor_5  g12733(new_n6157, n25435, new_n15082_1);
nand_5 g12734(new_n15082_1, new_n4368, new_n15083);
not_8  g12735(new_n15083, new_n15084);
not_8  g12736(new_n3910, new_n15085);
not_8  g12737(new_n15082_1, new_n15086);
nand_5 g12738(new_n15086, new_n15085, new_n15087);
nand_5 g12739(new_n15087, new_n15083, new_n15088);
nor_5  g12740(new_n15088, new_n5122, new_n15089);
nor_5  g12741(new_n15089, new_n15084, new_n15090);
not_8  g12742(new_n15090, new_n15091);
nand_5 g12743(new_n15091, new_n15081, new_n15092);
nand_5 g12744(new_n15092, new_n15080, new_n15093);
nand_5 g12745(new_n15093, new_n15078, new_n15094_1);
nand_5 g12746(new_n15094_1, new_n15077_1, new_n15095);
nand_5 g12747(new_n15095, new_n15075, new_n15096);
nand_5 g12748(new_n15096, new_n15074, new_n15097);
nand_5 g12749(new_n15097, new_n15072, new_n15098);
nand_5 g12750(new_n15098, new_n15071, new_n15099);
nand_5 g12751(new_n15099, new_n15070, new_n15100);
nand_5 g12752(new_n15100, new_n15069, new_n15101);
nand_5 g12753(new_n15101, new_n15067, new_n15102);
nand_5 g12754(new_n15102, new_n15066, new_n15103);
nand_5 g12755(new_n15103, new_n15063, new_n15104);
nand_5 g12756(new_n15104, new_n15062, new_n15105);
nand_5 g12757(new_n15105, new_n15059, new_n15106);
nand_5 g12758(new_n15106, new_n15058, new_n15107);
not_8  g12759(new_n15107, new_n15108);
nor_5  g12760(new_n15055, n11898, new_n15109);
nand_5 g12761(new_n15109, new_n5151, new_n15110);
not_8  g12762(new_n15110, new_n15111);
nand_5 g12763(new_n15111, new_n15108, new_n15112);
nor_5  g12764(new_n15109, new_n5151, new_n15113);
nand_5 g12765(new_n15113, new_n15107, new_n15114);
nand_5 g12766(new_n15114, new_n15112, new_n15115);
nor_5  g12767(new_n15115, new_n15052_1, new_n15116);
nand_5 g12768(new_n15115, new_n15052_1, new_n15117);
xnor_4 g12769(new_n15050, new_n15046, new_n15118_1);
not_8  g12770(new_n5151, new_n15119);
xnor_4 g12771(new_n15109, new_n15119, new_n15120);
xnor_4 g12772(new_n15120, new_n15108, new_n15121);
nor_5  g12773(new_n15121, new_n15118_1, new_n15122);
xnor_4 g12774(new_n15121, new_n15118_1, new_n15123);
xnor_4 g12775(new_n15044, new_n15002_1, new_n15124);
xnor_4 g12776(new_n15105, new_n15059, new_n15125);
not_8  g12777(new_n15125, new_n15126);
nand_5 g12778(new_n15126, new_n15124, new_n15127);
xnor_4 g12779(new_n15125, new_n15124, new_n15128_1);
xnor_4 g12780(new_n15103, new_n15063, new_n15129);
not_8  g12781(new_n15129, new_n15130);
xnor_4 g12782(new_n15042, new_n15041, new_n15131);
nand_5 g12783(new_n15131, new_n15130, new_n15132);
xnor_4 g12784(new_n15131, new_n15129, new_n15133);
not_8  g12785(new_n15011_1, new_n15134);
xnor_4 g12786(new_n15038, new_n15134, new_n15135);
xnor_4 g12787(new_n15101, new_n15067, new_n15136);
not_8  g12788(new_n15136, new_n15137);
nand_5 g12789(new_n15137, new_n15135, new_n15138);
xnor_4 g12790(new_n15136, new_n15135, new_n15139_1);
xnor_4 g12791(new_n15099, new_n15070, new_n15140);
not_8  g12792(new_n15140, new_n15141);
xnor_4 g12793(new_n15036, new_n15013, new_n15142);
nand_5 g12794(new_n15142, new_n15141, new_n15143);
xnor_4 g12795(new_n15142, new_n15140, new_n15144);
not_8  g12796(new_n15072, new_n15145_1);
xnor_4 g12797(new_n15097, new_n15145_1, new_n15146_1);
xnor_4 g12798(new_n15034, new_n15015, new_n15147);
nand_5 g12799(new_n15147, new_n15146_1, new_n15148);
not_8  g12800(new_n15147, new_n15149);
xnor_4 g12801(new_n15149, new_n15146_1, new_n15150);
xnor_4 g12802(new_n15095, new_n15075, new_n15151);
not_8  g12803(new_n15151, new_n15152);
xnor_4 g12804(new_n15032, new_n15017, new_n15153);
nand_5 g12805(new_n15153, new_n15152, new_n15154);
xnor_4 g12806(new_n15153, new_n15151, new_n15155);
xnor_4 g12807(new_n15093, new_n15078, new_n15156);
xnor_4 g12808(new_n15030, new_n15019_1, new_n15157);
not_8  g12809(new_n15157, new_n15158);
nor_5  g12810(new_n15158, new_n15156, new_n15159);
not_8  g12811(new_n15159, new_n15160);
xnor_4 g12812(new_n15157, new_n15156, new_n15161);
xnor_4 g12813(new_n15091, new_n15081, new_n15162);
not_8  g12814(new_n15162, new_n15163);
xnor_4 g12815(new_n15028, new_n15027, new_n15164);
nor_5  g12816(new_n15164, new_n15163, new_n15165_1);
xnor_4 g12817(new_n15164, new_n15163, new_n15166);
xnor_4 g12818(new_n15025, new_n15023, new_n15167_1);
not_8  g12819(new_n15167_1, new_n15168);
xnor_4 g12820(new_n15088, new_n6154, new_n15169);
not_8  g12821(new_n15169, new_n15170);
nor_5  g12822(new_n15170, new_n15168, new_n15171);
not_8  g12823(new_n15171, new_n15172);
xnor_4 g12824(new_n9960, new_n7664, new_n15173);
xnor_4 g12825(new_n5126, n25435, new_n15174);
not_8  g12826(new_n15174, new_n15175);
nand_5 g12827(new_n15175, new_n15173, new_n15176_1);
xnor_4 g12828(new_n15169, new_n15168, new_n15177);
nand_5 g12829(new_n15177, new_n15176_1, new_n15178);
nand_5 g12830(new_n15178, new_n15172, new_n15179);
nor_5  g12831(new_n15179, new_n15166, new_n15180_1);
nor_5  g12832(new_n15180_1, new_n15165_1, new_n15181);
nand_5 g12833(new_n15181, new_n15161, new_n15182_1);
nand_5 g12834(new_n15182_1, new_n15160, new_n15183);
nand_5 g12835(new_n15183, new_n15155, new_n15184);
nand_5 g12836(new_n15184, new_n15154, new_n15185);
nand_5 g12837(new_n15185, new_n15150, new_n15186);
nand_5 g12838(new_n15186, new_n15148, new_n15187);
nand_5 g12839(new_n15187, new_n15144, new_n15188);
nand_5 g12840(new_n15188, new_n15143, new_n15189);
nand_5 g12841(new_n15189, new_n15139_1, new_n15190);
nand_5 g12842(new_n15190, new_n15138, new_n15191);
nand_5 g12843(new_n15191, new_n15133, new_n15192);
nand_5 g12844(new_n15192, new_n15132, new_n15193);
nand_5 g12845(new_n15193, new_n15128_1, new_n15194);
nand_5 g12846(new_n15194, new_n15127, new_n15195);
not_8  g12847(new_n15195, new_n15196);
nor_5  g12848(new_n15196, new_n15123, new_n15197);
nor_5  g12849(new_n15197, new_n15122, new_n15198);
nand_5 g12850(new_n15198, new_n15117, new_n15199);
nand_5 g12851(new_n15199, new_n15112, new_n15200);
nor_5  g12852(new_n15200, new_n15116, n2774);
nor_5  g12853(new_n10026, n20478, new_n15202);
nand_5 g12854(new_n15202, new_n8152, new_n15203);
nor_5  g12855(new_n15203, n2421, new_n15204);
nand_5 g12856(new_n15204, new_n8147, new_n15205_1);
nor_5  g12857(new_n15205_1, n5031, new_n15206);
xnor_4 g12858(new_n15206, n2145, new_n15207);
xnor_4 g12859(new_n15207, new_n5158_1, new_n15208);
xnor_4 g12860(new_n15205_1, new_n6315, new_n15209);
nor_5  g12861(new_n15209, n2659, new_n15210);
not_8  g12862(new_n15210, new_n15211);
xnor_4 g12863(new_n15209, new_n5162, new_n15212);
xnor_4 g12864(new_n15204, n11044, new_n15213);
nor_5  g12865(new_n15213, n24327, new_n15214);
xnor_4 g12866(new_n15213, new_n5166, new_n15215);
not_8  g12867(new_n15215, new_n15216);
xnor_4 g12868(new_n15203, new_n6322, new_n15217);
nor_5  g12869(new_n15217, n22198, new_n15218);
xnor_4 g12870(new_n15202, n987, new_n15219);
nand_5 g12871(new_n15219, n20826, new_n15220);
xnor_4 g12872(new_n15219, new_n5174, new_n15221);
nand_5 g12873(new_n10027, n7305, new_n15222);
nand_5 g12874(new_n10041, new_n10028, new_n15223);
nand_5 g12875(new_n15223, new_n15222, new_n15224);
nand_5 g12876(new_n15224, new_n15221, new_n15225);
nand_5 g12877(new_n15225, new_n15220, new_n15226);
xnor_4 g12878(new_n15217, new_n5170, new_n15227);
not_8  g12879(new_n15227, new_n15228);
nor_5  g12880(new_n15228, new_n15226, new_n15229);
nor_5  g12881(new_n15229, new_n15218, new_n15230_1);
nor_5  g12882(new_n15230_1, new_n15216, new_n15231);
nor_5  g12883(new_n15231, new_n15214, new_n15232);
not_8  g12884(new_n15232, new_n15233);
nand_5 g12885(new_n15233, new_n15212, new_n15234);
nand_5 g12886(new_n15234, new_n15211, new_n15235);
xnor_4 g12887(new_n15235, new_n15208, new_n15236);
xnor_4 g12888(new_n15236, new_n3610, new_n15237);
xnor_4 g12889(new_n15232, new_n15212, new_n15238);
nor_5  g12890(new_n15238, new_n3616, new_n15239);
not_8  g12891(new_n15239, new_n15240);
xnor_4 g12892(new_n15230_1, new_n15216, new_n15241_1);
nor_5  g12893(new_n15241_1, new_n3620, new_n15242);
xnor_4 g12894(new_n15241_1, new_n3620, new_n15243);
xnor_4 g12895(new_n15227, new_n15226, new_n15244);
not_8  g12896(new_n15244, new_n15245);
nor_5  g12897(new_n15245, new_n3625, new_n15246);
xnor_4 g12898(new_n15244, new_n3625, new_n15247);
not_8  g12899(new_n15247, new_n15248);
xnor_4 g12900(new_n15224, new_n15221, new_n15249);
not_8  g12901(new_n15249, new_n15250);
nor_5  g12902(new_n15250, new_n3630, new_n15251);
xnor_4 g12903(new_n15250, new_n3630, new_n15252);
not_8  g12904(new_n10042, new_n15253);
nand_5 g12905(new_n15253, new_n3634, new_n15254);
xnor_4 g12906(new_n10042, new_n3634, new_n15255_1);
nor_5  g12907(new_n10062, new_n3641, new_n15256);
not_8  g12908(new_n15256, new_n15257);
xnor_4 g12909(new_n10062, new_n3640, new_n15258_1);
nor_5  g12910(new_n10067, new_n3647, new_n15259);
not_8  g12911(new_n15259, new_n15260);
nor_5  g12912(new_n10071, new_n3652, new_n15261);
xnor_4 g12913(new_n10067, new_n3646, new_n15262);
nand_5 g12914(new_n15262, new_n15261, new_n15263);
nand_5 g12915(new_n15263, new_n15260, new_n15264);
nand_5 g12916(new_n15264, new_n15258_1, new_n15265);
nand_5 g12917(new_n15265, new_n15257, new_n15266);
nand_5 g12918(new_n15266, new_n15255_1, new_n15267);
nand_5 g12919(new_n15267, new_n15254, new_n15268);
nor_5  g12920(new_n15268, new_n15252, new_n15269);
nor_5  g12921(new_n15269, new_n15251, new_n15270);
nor_5  g12922(new_n15270, new_n15248, new_n15271_1);
nor_5  g12923(new_n15271_1, new_n15246, new_n15272);
nor_5  g12924(new_n15272, new_n15243, new_n15273);
nor_5  g12925(new_n15273, new_n15242, new_n15274);
xnor_4 g12926(new_n15238, new_n3615, new_n15275_1);
nand_5 g12927(new_n15275_1, new_n15274, new_n15276);
nand_5 g12928(new_n15276, new_n15240, new_n15277);
xnor_4 g12929(new_n15277, new_n15237, new_n15278);
xnor_4 g12930(new_n3741, new_n3675, new_n15279);
nor_5  g12931(new_n3748, new_n3678, new_n15280);
nor_5  g12932(new_n3747, n13719, new_n15281);
or_5   g12933(new_n3752, n442, new_n15282);
xnor_4 g12934(new_n3752, new_n3681, new_n15283);
nand_5 g12935(new_n3759, new_n3684, new_n15284);
xnor_4 g12936(new_n3758_1, new_n3684, new_n15285);
nand_5 g12937(new_n3763, new_n3687, new_n15286);
xnor_4 g12938(new_n3762, new_n3687, new_n15287);
nand_5 g12939(new_n3770, new_n3691, new_n15288);
nand_5 g12940(new_n3774, new_n3696, new_n15289_1);
xnor_4 g12941(new_n3773, new_n3696, new_n15290);
nand_5 g12942(new_n3781_1, new_n3700, new_n15291);
not_8  g12943(new_n15291, new_n15292);
nand_5 g12944(n21993, n7139, new_n15293);
not_8  g12945(new_n15293, new_n15294);
xnor_4 g12946(new_n3780, new_n3700, new_n15295);
not_8  g12947(new_n15295, new_n15296);
nor_5  g12948(new_n15296, new_n15294, new_n15297);
nor_5  g12949(new_n15297, new_n15292, new_n15298);
not_8  g12950(new_n15298, new_n15299);
nand_5 g12951(new_n15299, new_n15290, new_n15300_1);
nand_5 g12952(new_n15300_1, new_n15289_1, new_n15301);
xnor_4 g12953(new_n3769, new_n3691, new_n15302);
nand_5 g12954(new_n15302, new_n15301, new_n15303);
nand_5 g12955(new_n15303, new_n15288, new_n15304);
nand_5 g12956(new_n15304, new_n15287, new_n15305);
nand_5 g12957(new_n15305, new_n15286, new_n15306);
nand_5 g12958(new_n15306, new_n15285, new_n15307_1);
nand_5 g12959(new_n15307_1, new_n15284, new_n15308);
nand_5 g12960(new_n15308, new_n15283, new_n15309);
nand_5 g12961(new_n15309, new_n15282, new_n15310);
nor_5  g12962(new_n15310, new_n15281, new_n15311);
nor_5  g12963(new_n15311, new_n15280, new_n15312);
xnor_4 g12964(new_n15312, new_n15279, new_n15313);
xnor_4 g12965(new_n15313, new_n15278, new_n15314);
xnor_4 g12966(new_n15275_1, new_n15274, new_n15315);
not_8  g12967(new_n15315, new_n15316);
xnor_4 g12968(new_n3747, new_n3678, new_n15317);
xnor_4 g12969(new_n15317, new_n15310, new_n15318);
nand_5 g12970(new_n15318, new_n15316, new_n15319);
xnor_4 g12971(new_n15318, new_n15315, new_n15320);
xnor_4 g12972(new_n15308, new_n15283, new_n15321);
xnor_4 g12973(new_n15272, new_n15243, new_n15322);
nor_5  g12974(new_n15322, new_n15321, new_n15323);
xnor_4 g12975(new_n15322, new_n15321, new_n15324);
xnor_4 g12976(new_n15306, new_n15285, new_n15325);
xnor_4 g12977(new_n15270, new_n15247, new_n15326);
not_8  g12978(new_n15326, new_n15327_1);
nor_5  g12979(new_n15327_1, new_n15325, new_n15328);
xnor_4 g12980(new_n15327_1, new_n15325, new_n15329);
xnor_4 g12981(new_n15304, new_n15287, new_n15330);
not_8  g12982(new_n15330, new_n15331);
xnor_4 g12983(new_n15268, new_n15252, new_n15332_1);
not_8  g12984(new_n15332_1, new_n15333);
nor_5  g12985(new_n15333, new_n15331, new_n15334);
not_8  g12986(new_n15334, new_n15335);
xnor_4 g12987(new_n15302, new_n15301, new_n15336);
not_8  g12988(new_n15336, new_n15337);
xnor_4 g12989(new_n15266, new_n15255_1, new_n15338);
nor_5  g12990(new_n15338, new_n15337, new_n15339);
not_8  g12991(new_n15339, new_n15340);
xnor_4 g12992(new_n15338, new_n15336, new_n15341);
xnor_4 g12993(new_n15298, new_n15290, new_n15342);
xnor_4 g12994(new_n15264, new_n15258_1, new_n15343);
nor_5  g12995(new_n15343, new_n15342, new_n15344);
not_8  g12996(new_n15344, new_n15345_1);
xnor_4 g12997(new_n15343, new_n15342, new_n15346);
not_8  g12998(new_n15346, new_n15347);
xnor_4 g12999(new_n15262, new_n15261, new_n15348);
not_8  g13000(new_n15348, new_n15349);
nor_5  g13001(new_n15349, new_n15295, new_n15350);
xnor_4 g13002(new_n15295, new_n15294, new_n15351);
nor_5  g13003(new_n15351, new_n15348, new_n15352);
xnor_4 g13004(n21993, new_n3702, new_n15353_1);
xnor_4 g13005(new_n10070, new_n3652, new_n15354);
nand_5 g13006(new_n15354, new_n15353_1, new_n15355);
not_8  g13007(new_n15355, new_n15356);
nor_5  g13008(new_n15356, new_n15352, new_n15357);
nor_5  g13009(new_n15357, new_n15350, new_n15358);
nand_5 g13010(new_n15358, new_n15347, new_n15359);
nand_5 g13011(new_n15359, new_n15345_1, new_n15360);
nand_5 g13012(new_n15360, new_n15341, new_n15361);
nand_5 g13013(new_n15361, new_n15340, new_n15362);
xnor_4 g13014(new_n15332_1, new_n15331, new_n15363);
nand_5 g13015(new_n15363, new_n15362, new_n15364);
nand_5 g13016(new_n15364, new_n15335, new_n15365);
nor_5  g13017(new_n15365, new_n15329, new_n15366_1);
nor_5  g13018(new_n15366_1, new_n15328, new_n15367);
nor_5  g13019(new_n15367, new_n15324, new_n15368);
nor_5  g13020(new_n15368, new_n15323, new_n15369);
nand_5 g13021(new_n15369, new_n15320, new_n15370);
nand_5 g13022(new_n15370, new_n15319, new_n15371);
xnor_4 g13023(new_n15371, new_n15314, n2779);
not_8  g13024(n25751, new_n15373);
nand_5 g13025(new_n10966, new_n15373, new_n15374);
xnor_4 g13026(new_n10965, new_n15373, new_n15375);
not_8  g13027(n26053, new_n15376);
nand_5 g13028(new_n10970, new_n15376, new_n15377);
xnor_4 g13029(new_n10969, new_n15376, new_n15378_1);
not_8  g13030(n7917, new_n15379);
not_8  g13031(new_n10973, new_n15380);
nand_5 g13032(new_n15380, new_n15379, new_n15381);
xnor_4 g13033(new_n10973, new_n15379, new_n15382_1);
not_8  g13034(n17302, new_n15383);
not_8  g13035(new_n10977, new_n15384);
nand_5 g13036(new_n15384, new_n15383, new_n15385);
xnor_4 g13037(new_n10977, new_n15383, new_n15386);
not_8  g13038(n2013, new_n15387);
not_8  g13039(new_n10980, new_n15388);
nand_5 g13040(new_n15388, new_n15387, new_n15389);
xnor_4 g13041(new_n10980, new_n15387, new_n15390);
not_8  g13042(n23755, new_n15391);
nand_5 g13043(new_n10985, new_n15391, new_n15392);
not_8  g13044(n19163, new_n15393);
nand_5 g13045(new_n10989, new_n15393, new_n15394);
xnor_4 g13046(new_n10988, new_n15393, new_n15395);
not_8  g13047(n22358, new_n15396);
nand_5 g13048(new_n6126, new_n15396, new_n15397);
nand_5 g13049(n25926, n9646, new_n15398);
xnor_4 g13050(new_n6126, n22358, new_n15399);
nand_5 g13051(new_n15399, new_n15398, new_n15400);
nand_5 g13052(new_n15400, new_n15397, new_n15401);
nand_5 g13053(new_n15401, new_n15395, new_n15402);
nand_5 g13054(new_n15402, new_n15394, new_n15403);
xnor_4 g13055(new_n10984, new_n15391, new_n15404);
nand_5 g13056(new_n15404, new_n15403, new_n15405);
nand_5 g13057(new_n15405, new_n15392, new_n15406);
nand_5 g13058(new_n15406, new_n15390, new_n15407_1);
nand_5 g13059(new_n15407_1, new_n15389, new_n15408);
nand_5 g13060(new_n15408, new_n15386, new_n15409);
nand_5 g13061(new_n15409, new_n15385, new_n15410);
nand_5 g13062(new_n15410, new_n15382_1, new_n15411);
nand_5 g13063(new_n15411, new_n15381, new_n15412);
nand_5 g13064(new_n15412, new_n15378_1, new_n15413);
nand_5 g13065(new_n15413, new_n15377, new_n15414);
nand_5 g13066(new_n15414, new_n15375, new_n15415);
nand_5 g13067(new_n15415, new_n15374, new_n15416);
not_8  g13068(n25586, new_n15417);
xnor_4 g13069(new_n10963, new_n15417, new_n15418);
xnor_4 g13070(new_n15418, new_n15416, new_n15419);
xnor_4 g13071(new_n15419, n4514, new_n15420);
xnor_4 g13072(new_n15414, new_n15375, new_n15421);
nand_5 g13073(new_n15421, new_n12114, new_n15422);
xnor_4 g13074(new_n15421, n3984, new_n15423);
xnor_4 g13075(new_n15412, new_n15378_1, new_n15424_1);
nand_5 g13076(new_n15424_1, new_n12117, new_n15425);
xnor_4 g13077(new_n15424_1, n19652, new_n15426);
xnor_4 g13078(new_n15410, new_n15382_1, new_n15427);
nand_5 g13079(new_n15427, new_n11621, new_n15428_1);
xnor_4 g13080(new_n15408, new_n15386, new_n15429);
nand_5 g13081(new_n15429, new_n11624, new_n15430);
xnor_4 g13082(new_n15429, n26565, new_n15431);
xnor_4 g13083(new_n15406, new_n15390, new_n15432);
nand_5 g13084(new_n15432, new_n10121, new_n15433);
xnor_4 g13085(new_n15432, n3959, new_n15434);
xnor_4 g13086(new_n15404, new_n15403, new_n15435_1);
nand_5 g13087(new_n15435_1, new_n12282, new_n15436);
xnor_4 g13088(new_n15435_1, n11566, new_n15437);
xnor_4 g13089(new_n15401, new_n15395, new_n15438_1);
nand_5 g13090(new_n15438_1, new_n12285, new_n15439);
xnor_4 g13091(new_n15399, new_n15398, new_n15440);
nand_5 g13092(new_n15440, new_n12289, new_n15441);
nand_5 g13093(new_n6941, n14230, new_n15442);
xnor_4 g13094(new_n15440, n26625, new_n15443);
nand_5 g13095(new_n15443, new_n15442, new_n15444);
nand_5 g13096(new_n15444, new_n15441, new_n15445);
xnor_4 g13097(new_n15438_1, n26744, new_n15446);
nand_5 g13098(new_n15446, new_n15445, new_n15447);
nand_5 g13099(new_n15447, new_n15439, new_n15448);
nand_5 g13100(new_n15448, new_n15437, new_n15449);
nand_5 g13101(new_n15449, new_n15436, new_n15450);
nand_5 g13102(new_n15450, new_n15434, new_n15451);
nand_5 g13103(new_n15451, new_n15433, new_n15452);
nand_5 g13104(new_n15452, new_n15431, new_n15453);
nand_5 g13105(new_n15453, new_n15430, new_n15454);
xnor_4 g13106(new_n15427, n3366, new_n15455);
nand_5 g13107(new_n15455, new_n15454, new_n15456);
nand_5 g13108(new_n15456, new_n15428_1, new_n15457);
nand_5 g13109(new_n15457, new_n15426, new_n15458);
nand_5 g13110(new_n15458, new_n15425, new_n15459);
nand_5 g13111(new_n15459, new_n15423, new_n15460);
nand_5 g13112(new_n15460, new_n15422, new_n15461);
xnor_4 g13113(new_n15461, new_n15420, new_n15462);
nand_5 g13114(new_n15462, new_n11097, new_n15463);
xnor_4 g13115(new_n15462, new_n11096, new_n15464);
xnor_4 g13116(new_n15459, new_n15423, new_n15465_1);
nand_5 g13117(new_n15465_1, new_n11105, new_n15466);
xnor_4 g13118(new_n15465_1, new_n11104, new_n15467_1);
xnor_4 g13119(new_n15457, new_n15426, new_n15468);
nand_5 g13120(new_n15468, new_n11111, new_n15469);
xnor_4 g13121(new_n15468, new_n11109, new_n15470_1);
xnor_4 g13122(new_n15455, new_n15454, new_n15471);
nand_5 g13123(new_n15471, new_n11117, new_n15472);
xnor_4 g13124(new_n15471, new_n11116, new_n15473);
xnor_4 g13125(new_n15452, new_n15431, new_n15474);
nand_5 g13126(new_n15474, new_n11123, new_n15475);
xnor_4 g13127(new_n15474, new_n11122, new_n15476);
xnor_4 g13128(new_n15450, new_n15434, new_n15477_1);
nand_5 g13129(new_n15477_1, new_n11128, new_n15478);
xnor_4 g13130(new_n15477_1, new_n11127_1, new_n15479);
xnor_4 g13131(new_n15448, new_n15437, new_n15480);
nand_5 g13132(new_n15480, new_n11135, new_n15481_1);
xnor_4 g13133(new_n15480, new_n11132_1, new_n15482);
not_8  g13134(new_n15446, new_n15483);
xnor_4 g13135(new_n15483, new_n15445, new_n15484);
not_8  g13136(new_n15484, new_n15485);
nand_5 g13137(new_n15485, new_n11141, new_n15486);
xnor_4 g13138(new_n15484, new_n11141, new_n15487);
not_8  g13139(new_n15442, new_n15488);
xnor_4 g13140(new_n15443, new_n15488, new_n15489);
nor_5  g13141(new_n15489, new_n6123, new_n15490_1);
not_8  g13142(new_n15490_1, new_n15491);
nor_5  g13143(new_n6942, new_n6118, new_n15492);
not_8  g13144(new_n15492, new_n15493);
nand_5 g13145(new_n15489, new_n11145, new_n15494);
nand_5 g13146(new_n15494, new_n15493, new_n15495);
nand_5 g13147(new_n15495, new_n15491, new_n15496_1);
nand_5 g13148(new_n15496_1, new_n15487, new_n15497);
nand_5 g13149(new_n15497, new_n15486, new_n15498);
nand_5 g13150(new_n15498, new_n15482, new_n15499);
nand_5 g13151(new_n15499, new_n15481_1, new_n15500);
nand_5 g13152(new_n15500, new_n15479, new_n15501_1);
nand_5 g13153(new_n15501_1, new_n15478, new_n15502);
nand_5 g13154(new_n15502, new_n15476, new_n15503);
nand_5 g13155(new_n15503, new_n15475, new_n15504);
nand_5 g13156(new_n15504, new_n15473, new_n15505);
nand_5 g13157(new_n15505, new_n15472, new_n15506_1);
nand_5 g13158(new_n15506_1, new_n15470_1, new_n15507);
nand_5 g13159(new_n15507, new_n15469, new_n15508_1);
nand_5 g13160(new_n15508_1, new_n15467_1, new_n15509);
nand_5 g13161(new_n15509, new_n15466, new_n15510);
nand_5 g13162(new_n15510, new_n15464, new_n15511);
nand_5 g13163(new_n15511, new_n15463, new_n15512);
xnor_4 g13164(new_n15512, new_n11093, new_n15513);
nor_5  g13165(new_n15419, new_n12110, new_n15514);
not_8  g13166(new_n15420, new_n15515);
nor_5  g13167(new_n15461, new_n15515, new_n15516);
nor_5  g13168(new_n15516, new_n15514, new_n15517);
nor_5  g13169(new_n10963, n25586, new_n15518);
nor_5  g13170(new_n15518, new_n15416, new_n15519);
not_8  g13171(new_n10963, new_n15520);
nor_5  g13172(new_n15520, new_n15417, new_n15521);
or_5   g13173(new_n15521, new_n10960, new_n15522);
nor_5  g13174(new_n15522, new_n15519, new_n15523);
xnor_4 g13175(new_n15523, new_n15517, new_n15524);
xnor_4 g13176(new_n15524, new_n15513, n2826);
nand_5 g13177(new_n6574, n5140, new_n15526);
xnor_4 g13178(new_n6574, new_n13066, new_n15527);
nand_5 g13179(new_n6581, n6204, new_n15528);
xnor_4 g13180(new_n6581, new_n13069, new_n15529);
nand_5 g13181(new_n13170, n3349, new_n15530);
xnor_4 g13182(new_n6587_1, n3349, new_n15531);
nand_5 g13183(new_n13206, n1742, new_n15532);
xnor_4 g13184(new_n6590_1, n1742, new_n15533);
nor_5  g13185(new_n6593, new_n6815, new_n15534);
not_8  g13186(new_n15534, new_n15535);
and_5  g13187(new_n6597, new_n6821, new_n15536);
xnor_4 g13188(new_n6597, n8244, new_n15537);
nor_5  g13189(new_n6598, new_n6826_1, new_n15538);
xnor_4 g13190(new_n6598, n9493, new_n15539_1);
not_8  g13191(new_n6601, new_n15540);
nor_5  g13192(new_n15540, n15167, new_n15541);
nor_5  g13193(new_n6605, new_n6836, new_n15542);
not_8  g13194(new_n15542, new_n15543);
not_8  g13195(n8656, new_n15544);
nor_5  g13196(new_n6609, new_n15544, new_n15545);
xnor_4 g13197(new_n6605, n21095, new_n15546_1);
nand_5 g13198(new_n15546_1, new_n15545, new_n15547);
nand_5 g13199(new_n15547, new_n15543, new_n15548);
xnor_4 g13200(new_n6601, n15167, new_n15549);
not_8  g13201(new_n15549, new_n15550);
nor_5  g13202(new_n15550, new_n15548, new_n15551);
nor_5  g13203(new_n15551, new_n15541, new_n15552);
nand_5 g13204(new_n15552, new_n15539_1, new_n15553);
not_8  g13205(new_n15553, new_n15554);
nor_5  g13206(new_n15554, new_n15538, new_n15555_1);
nand_5 g13207(new_n15555_1, new_n15537, new_n15556);
not_8  g13208(new_n15556, new_n15557);
nor_5  g13209(new_n15557, new_n15536, new_n15558_1);
xnor_4 g13210(new_n6593, n4858, new_n15559_1);
nand_5 g13211(new_n15559_1, new_n15558_1, new_n15560);
nand_5 g13212(new_n15560, new_n15535, new_n15561);
nand_5 g13213(new_n15561, new_n15533, new_n15562);
nand_5 g13214(new_n15562, new_n15532, new_n15563);
nand_5 g13215(new_n15563, new_n15531, new_n15564);
nand_5 g13216(new_n15564, new_n15530, new_n15565);
nand_5 g13217(new_n15565, new_n15529, new_n15566);
nand_5 g13218(new_n15566, new_n15528, new_n15567);
nand_5 g13219(new_n15567, new_n15527, new_n15568);
nand_5 g13220(new_n15568, new_n15526, new_n15569);
nand_5 g13221(new_n15569, new_n13111, new_n15570_1);
not_8  g13222(n25365, new_n15571);
nor_5  g13223(new_n2634, new_n15571, new_n15572);
not_8  g13224(new_n2635, new_n15573_1);
nor_5  g13225(new_n2700, new_n15573_1, new_n15574);
nor_5  g13226(new_n15574, new_n15572, new_n15575);
or_5   g13227(n20040, n9396, new_n15576);
nand_5 g13228(new_n2633, new_n2585, new_n15577);
nand_5 g13229(new_n15577, new_n15576, new_n15578);
nor_5  g13230(new_n15578, new_n15575, new_n15579);
not_8  g13231(new_n15579, new_n15580);
xnor_4 g13232(new_n15580, new_n15570_1, new_n15581);
xnor_4 g13233(new_n15569, new_n13111, new_n15582);
xnor_4 g13234(new_n15578, new_n15575, new_n15583);
not_8  g13235(new_n15583, new_n15584);
nand_5 g13236(new_n15584, new_n15582, new_n15585);
xnor_4 g13237(new_n15583, new_n15582, new_n15586);
xnor_4 g13238(new_n15567, new_n15527, new_n15587);
nand_5 g13239(new_n15587, new_n2701, new_n15588_1);
xnor_4 g13240(new_n15587, new_n2702, new_n15589);
xnor_4 g13241(new_n15565, new_n15529, new_n15590_1);
nand_5 g13242(new_n15590_1, new_n2831, new_n15591);
xnor_4 g13243(new_n15590_1, new_n2832, new_n15592);
xnor_4 g13244(new_n15563, new_n15531, new_n15593);
nand_5 g13245(new_n15593, new_n2838, new_n15594);
xnor_4 g13246(new_n15593, new_n2837, new_n15595);
xnor_4 g13247(new_n15561, new_n15533, new_n15596);
nand_5 g13248(new_n15596, new_n2843, new_n15597);
xnor_4 g13249(new_n15596, new_n2847, new_n15598_1);
not_8  g13250(new_n2850, new_n15599);
xnor_4 g13251(new_n15559_1, new_n15558_1, new_n15600);
nand_5 g13252(new_n15600, new_n15599, new_n15601);
xnor_4 g13253(new_n15600, new_n2850, new_n15602_1);
xnor_4 g13254(new_n15555_1, new_n15537, new_n15603);
not_8  g13255(new_n15603, new_n15604);
nand_5 g13256(new_n15604, new_n2854, new_n15605);
xnor_4 g13257(new_n15603, new_n2854, new_n15606);
xnor_4 g13258(new_n15552, new_n15539_1, new_n15607);
not_8  g13259(new_n15607, new_n15608);
nor_5  g13260(new_n15608, new_n2864, new_n15609);
xnor_4 g13261(new_n15608, new_n2861, new_n15610);
not_8  g13262(new_n15610, new_n15611);
xnor_4 g13263(new_n15549, new_n15548, new_n15612);
and_5  g13264(new_n15612, new_n2867, new_n15613);
xnor_4 g13265(new_n15612, new_n2869, new_n15614_1);
not_8  g13266(new_n15614_1, new_n15615);
xnor_4 g13267(new_n15546_1, new_n15545, new_n15616);
and_5  g13268(new_n15616, new_n2880, new_n15617);
xnor_4 g13269(new_n6608, new_n15544, new_n15618);
nor_5  g13270(new_n15618, new_n2876, new_n15619);
not_8  g13271(new_n15619, new_n15620);
xnor_4 g13272(new_n15616, new_n2873, new_n15621);
not_8  g13273(new_n15621, new_n15622);
nor_5  g13274(new_n15622, new_n15620, new_n15623);
nor_5  g13275(new_n15623, new_n15617, new_n15624);
nor_5  g13276(new_n15624, new_n15615, new_n15625);
nor_5  g13277(new_n15625, new_n15613, new_n15626);
nor_5  g13278(new_n15626, new_n15611, new_n15627);
nor_5  g13279(new_n15627, new_n15609, new_n15628);
not_8  g13280(new_n15628, new_n15629);
nand_5 g13281(new_n15629, new_n15606, new_n15630);
nand_5 g13282(new_n15630, new_n15605, new_n15631);
nand_5 g13283(new_n15631, new_n15602_1, new_n15632);
nand_5 g13284(new_n15632, new_n15601, new_n15633);
nand_5 g13285(new_n15633, new_n15598_1, new_n15634);
nand_5 g13286(new_n15634, new_n15597, new_n15635);
nand_5 g13287(new_n15635, new_n15595, new_n15636_1);
nand_5 g13288(new_n15636_1, new_n15594, new_n15637);
nand_5 g13289(new_n15637, new_n15592, new_n15638);
nand_5 g13290(new_n15638, new_n15591, new_n15639);
nand_5 g13291(new_n15639, new_n15589, new_n15640);
nand_5 g13292(new_n15640, new_n15588_1, new_n15641);
nand_5 g13293(new_n15641, new_n15586, new_n15642);
nand_5 g13294(new_n15642, new_n15585, new_n15643);
xnor_4 g13295(new_n15643, new_n15581, n2853);
xnor_4 g13296(n7099, n2035, new_n15645);
nor_5  g13297(new_n12575, n5213, new_n15646);
not_8  g13298(new_n15646, new_n15647);
xnor_4 g13299(n12811, n5213, new_n15648);
nor_5  g13300(n4665, new_n2959, new_n15649);
xnor_4 g13301(n4665, n1118, new_n15650);
nor_5  g13302(n25974, new_n2917, new_n15651);
nor_5  g13303(new_n12584, n19005, new_n15652_1);
nor_5  g13304(new_n2921, n1630, new_n15653);
nor_5  g13305(n4326, new_n12586, new_n15654);
nand_5 g13306(n5438, new_n12671, new_n15655);
nor_5  g13307(new_n15655, new_n15654, new_n15656);
nor_5  g13308(new_n15656, new_n15653, new_n15657);
nor_5  g13309(new_n15657, new_n15652_1, new_n15658);
nor_5  g13310(new_n15658, new_n15651, new_n15659);
and_5  g13311(new_n15659, new_n15650, new_n15660);
nor_5  g13312(new_n15660, new_n15649, new_n15661);
not_8  g13313(new_n15661, new_n15662_1);
nand_5 g13314(new_n15662_1, new_n15648, new_n15663);
nand_5 g13315(new_n15663, new_n15647, new_n15664);
xnor_4 g13316(new_n15664, new_n15645, new_n15665);
not_8  g13317(new_n11792, new_n15666);
nand_5 g13318(new_n4414, new_n6373, new_n15667);
xnor_4 g13319(new_n15667, new_n9912, new_n15668);
xnor_4 g13320(new_n15668, new_n4003, new_n15669);
nand_5 g13321(new_n4415, n626, new_n15670);
nand_5 g13322(new_n4437, new_n4416, new_n15671);
nand_5 g13323(new_n15671, new_n15670, new_n15672);
xnor_4 g13324(new_n15672, new_n15669, new_n15673);
xnor_4 g13325(new_n15673, new_n15666, new_n15674);
not_8  g13326(new_n4438, new_n15675);
nand_5 g13327(new_n15675, new_n4410, new_n15676);
nand_5 g13328(new_n4468, new_n4439, new_n15677);
nand_5 g13329(new_n15677, new_n15676, new_n15678);
xnor_4 g13330(new_n15678, new_n15674, new_n15679);
xnor_4 g13331(new_n15679, new_n15665, new_n15680);
xnor_4 g13332(new_n15661, new_n15648, new_n15681);
not_8  g13333(new_n15681, new_n15682);
nand_5 g13334(new_n15682, new_n4469, new_n15683);
xnor_4 g13335(new_n15659, new_n15650, new_n15684);
nand_5 g13336(new_n15684, new_n4473, new_n15685);
not_8  g13337(new_n15684, new_n15686);
xnor_4 g13338(new_n15686, new_n4473, new_n15687);
xnor_4 g13339(n25974, n19005, new_n15688);
xnor_4 g13340(new_n15688, new_n15657, new_n15689);
nand_5 g13341(new_n15689, new_n4477, new_n15690);
xnor_4 g13342(new_n15689, new_n4476_1, new_n15691);
xnor_4 g13343(n5438, n1451, new_n15692);
nor_5  g13344(new_n15692, new_n4491, new_n15693);
xnor_4 g13345(n4326, n1630, new_n15694);
xnor_4 g13346(new_n15694, new_n15655, new_n15695);
not_8  g13347(new_n15695, new_n15696);
and_5  g13348(new_n15696, new_n15693, new_n15697);
xnor_4 g13349(new_n15695, new_n15693, new_n15698);
not_8  g13350(new_n15698, new_n15699);
nor_5  g13351(new_n15699, new_n4481, new_n15700);
nor_5  g13352(new_n15700, new_n15697, new_n15701);
nand_5 g13353(new_n15701, new_n15691, new_n15702);
nand_5 g13354(new_n15702, new_n15690, new_n15703);
nand_5 g13355(new_n15703, new_n15687, new_n15704);
nand_5 g13356(new_n15704, new_n15685, new_n15705);
xnor_4 g13357(new_n15681, new_n4469, new_n15706);
nand_5 g13358(new_n15706, new_n15705, new_n15707);
nand_5 g13359(new_n15707, new_n15683, new_n15708);
xor_4  g13360(new_n15708, new_n15680, n2860);
xnor_4 g13361(new_n14737, new_n14717, n2887);
nor_5  g13362(new_n15667, n3570, new_n15711);
nand_5 g13363(new_n15711, new_n9909, new_n15712);
nor_5  g13364(new_n15712, n20359, new_n15713);
nand_5 g13365(new_n15713, new_n6359, new_n15714);
xnor_4 g13366(new_n15714, new_n6308_1, new_n15715);
not_8  g13367(new_n15715, new_n15716_1);
nand_5 g13368(new_n15716_1, new_n12614, new_n15717);
xnor_4 g13369(new_n15713, n2816, new_n15718);
nand_5 g13370(new_n15718, n5521, new_n15719);
not_8  g13371(new_n15718, new_n15720);
nand_5 g13372(new_n15720, new_n12615, new_n15721);
xnor_4 g13373(new_n15712, new_n7644, new_n15722);
nor_5  g13374(new_n15722, n11926, new_n15723);
xnor_4 g13375(new_n15722, n11926, new_n15724);
xnor_4 g13376(new_n15711, n4409, new_n15725);
nand_5 g13377(new_n15725, n4325, new_n15726);
not_8  g13378(new_n15725, new_n15727);
nand_5 g13379(new_n15727, new_n6318, new_n15728);
nand_5 g13380(new_n15668, n5337, new_n15729);
not_8  g13381(new_n15668, new_n15730);
nand_5 g13382(new_n15730, new_n4003, new_n15731);
nand_5 g13383(new_n15672, new_n15731, new_n15732);
nand_5 g13384(new_n15732, new_n15729, new_n15733);
nand_5 g13385(new_n15733, new_n15728, new_n15734);
nand_5 g13386(new_n15734, new_n15726, new_n15735);
nor_5  g13387(new_n15735, new_n15724, new_n15736);
nor_5  g13388(new_n15736, new_n15723, new_n15737);
nand_5 g13389(new_n15737, new_n15721, new_n15738);
nand_5 g13390(new_n15738, new_n15719, new_n15739);
nand_5 g13391(new_n15739, new_n15717, new_n15740);
nor_5  g13392(new_n15714, n8526, new_n15741);
nor_5  g13393(new_n15716_1, new_n12614, new_n15742);
nor_5  g13394(new_n15742, new_n15741, new_n15743_1);
nand_5 g13395(new_n15743_1, new_n15740, new_n15744);
xnor_4 g13396(new_n15744, new_n11765, new_n15745);
xnor_4 g13397(new_n15715, new_n12614, new_n15746);
xnor_4 g13398(new_n15746, new_n15739, new_n15747);
nor_5  g13399(new_n15747, new_n11769, new_n15748);
not_8  g13400(new_n15748, new_n15749_1);
xnor_4 g13401(new_n15747, new_n11771_1, new_n15750);
xnor_4 g13402(new_n15718, new_n12615, new_n15751);
xnor_4 g13403(new_n15751, new_n15737, new_n15752);
not_8  g13404(new_n15752, new_n15753);
nor_5  g13405(new_n15753, new_n11776, new_n15754);
xnor_4 g13406(new_n15752, new_n11774, new_n15755);
not_8  g13407(new_n11781, new_n15756);
xnor_4 g13408(new_n15735, new_n15724, new_n15757);
nor_5  g13409(new_n15757, new_n15756, new_n15758);
xnor_4 g13410(new_n15725, new_n6318, new_n15759);
xnor_4 g13411(new_n15759, new_n15733, new_n15760);
not_8  g13412(new_n15760, new_n15761_1);
nand_5 g13413(new_n15761_1, new_n11787, new_n15762_1);
xnor_4 g13414(new_n15760, new_n11787, new_n15763);
not_8  g13415(new_n15673, new_n15764);
nand_5 g13416(new_n15764, new_n15666, new_n15765);
nand_5 g13417(new_n15678, new_n15674, new_n15766_1);
nand_5 g13418(new_n15766_1, new_n15765, new_n15767);
nand_5 g13419(new_n15767, new_n15763, new_n15768);
nand_5 g13420(new_n15768, new_n15762_1, new_n15769);
xnor_4 g13421(new_n15757, new_n11781, new_n15770);
not_8  g13422(new_n15770, new_n15771);
nor_5  g13423(new_n15771, new_n15769, new_n15772);
nor_5  g13424(new_n15772, new_n15758, new_n15773);
nor_5  g13425(new_n15773, new_n15755, new_n15774);
nor_5  g13426(new_n15774, new_n15754, new_n15775);
nand_5 g13427(new_n15775, new_n15750, new_n15776);
nand_5 g13428(new_n15776, new_n15749_1, new_n15777);
xnor_4 g13429(new_n15777, new_n15745, new_n15778);
nand_5 g13430(new_n4356, new_n11231, new_n15779);
nor_5  g13431(new_n15779, n26452, new_n15780_1);
nand_5 g13432(new_n15780_1, new_n11222, new_n15781);
nor_5  g13433(new_n15781, n5077, new_n15782);
nand_5 g13434(new_n15782, new_n13699, new_n15783);
or_5   g13435(new_n15783, n8827, new_n15784);
xnor_4 g13436(new_n15783, new_n13680, new_n15785);
or_5   g13437(new_n15785, n11898, new_n15786);
xnor_4 g13438(new_n15782, n18035, new_n15787);
or_5   g13439(new_n15787, n19941, new_n15788);
xnor_4 g13440(new_n15787, new_n13683_1, new_n15789);
xnor_4 g13441(new_n15781, new_n11194, new_n15790);
or_5   g13442(new_n15790, n1099, new_n15791);
xnor_4 g13443(new_n15790, new_n11195, new_n15792);
xnor_4 g13444(new_n15780_1, n15546, new_n15793_1);
or_5   g13445(new_n15793_1, n2113, new_n15794);
xnor_4 g13446(new_n15779, new_n11244, new_n15795);
not_8  g13447(new_n15795, new_n15796);
nand_5 g13448(new_n15796, new_n3889, new_n15797);
xnor_4 g13449(new_n15795, new_n3889, new_n15798);
not_8  g13450(new_n4357, new_n15799);
nand_5 g13451(new_n15799, new_n3879, new_n15800);
nand_5 g13452(new_n4382, new_n4358, new_n15801);
nand_5 g13453(new_n15801, new_n15800, new_n15802);
nand_5 g13454(new_n15802, new_n15798, new_n15803);
nand_5 g13455(new_n15803, new_n15797, new_n15804);
xnor_4 g13456(new_n15793_1, new_n11199, new_n15805);
nand_5 g13457(new_n15805, new_n15804, new_n15806);
nand_5 g13458(new_n15806, new_n15794, new_n15807);
nand_5 g13459(new_n15807, new_n15792, new_n15808);
nand_5 g13460(new_n15808, new_n15791, new_n15809);
nand_5 g13461(new_n15809, new_n15789, new_n15810);
nand_5 g13462(new_n15810, new_n15788, new_n15811);
nand_5 g13463(new_n15785, n11898, new_n15812_1);
nand_5 g13464(new_n15812_1, new_n15811, new_n15813);
nand_5 g13465(new_n15813, new_n15786, new_n15814);
nand_5 g13466(new_n15814, new_n15784, new_n15815_1);
xnor_4 g13467(new_n15815_1, new_n15778, new_n15816_1);
not_8  g13468(new_n15816_1, new_n15817);
xnor_4 g13469(new_n15775, new_n15750, new_n15818);
xnor_4 g13470(new_n15785, new_n13681, new_n15819);
xnor_4 g13471(new_n15819, new_n15811, new_n15820);
not_8  g13472(new_n15820, new_n15821);
nand_5 g13473(new_n15821, new_n15818, new_n15822);
xnor_4 g13474(new_n15820, new_n15818, new_n15823);
xnor_4 g13475(new_n15809, new_n15789, new_n15824);
not_8  g13476(new_n15824, new_n15825);
xnor_4 g13477(new_n15773, new_n15755, new_n15826);
not_8  g13478(new_n15826, new_n15827);
nand_5 g13479(new_n15827, new_n15825, new_n15828);
xnor_4 g13480(new_n15827, new_n15824, new_n15829);
xnor_4 g13481(new_n15807, new_n15792, new_n15830);
not_8  g13482(new_n15830, new_n15831_1);
xnor_4 g13483(new_n15770, new_n15769, new_n15832);
nand_5 g13484(new_n15832, new_n15831_1, new_n15833);
xnor_4 g13485(new_n15832, new_n15830, new_n15834);
xnor_4 g13486(new_n15767, new_n15763, new_n15835);
xnor_4 g13487(new_n15805, new_n15804, new_n15836);
not_8  g13488(new_n15836, new_n15837);
nand_5 g13489(new_n15837, new_n15835, new_n15838);
xnor_4 g13490(new_n15836, new_n15835, new_n15839);
xnor_4 g13491(new_n15802, new_n15798, new_n15840);
not_8  g13492(new_n15840, new_n15841);
nand_5 g13493(new_n15841, new_n15679, new_n15842);
xnor_4 g13494(new_n15840, new_n15679, new_n15843);
nand_5 g13495(new_n4469, new_n13756, new_n15844);
nand_5 g13496(new_n4499, new_n4470, new_n15845);
nand_5 g13497(new_n15845, new_n15844, new_n15846_1);
nand_5 g13498(new_n15846_1, new_n15843, new_n15847);
nand_5 g13499(new_n15847, new_n15842, new_n15848);
nand_5 g13500(new_n15848, new_n15839, new_n15849);
nand_5 g13501(new_n15849, new_n15838, new_n15850);
nand_5 g13502(new_n15850, new_n15834, new_n15851);
nand_5 g13503(new_n15851, new_n15833, new_n15852);
nand_5 g13504(new_n15852, new_n15829, new_n15853);
nand_5 g13505(new_n15853, new_n15828, new_n15854);
nand_5 g13506(new_n15854, new_n15823, new_n15855);
nand_5 g13507(new_n15855, new_n15822, new_n15856);
xnor_4 g13508(new_n15856, new_n15817, n2929);
xnor_4 g13509(n22793, n767, new_n15858);
not_8  g13510(new_n15858, new_n15859_1);
nor_5  g13511(n8439, new_n2723, new_n15860);
xnor_4 g13512(n8439, n7330, new_n15861);
not_8  g13513(new_n15861, new_n15862);
nor_5  g13514(n25523, new_n2726, new_n15863);
xnor_4 g13515(n25523, n22492, new_n15864);
not_8  g13516(new_n15864, new_n15865);
nor_5  g13517(new_n11745, n5579, new_n15866);
xnor_4 g13518(n12821, n5579, new_n15867);
not_8  g13519(new_n15867, new_n15868);
nor_5  g13520(n23430, new_n2734, new_n15869_1);
xnor_4 g13521(n23430, n3468, new_n15870);
nor_5  g13522(n18558, new_n2792, new_n15871);
not_8  g13523(new_n14427, new_n15872);
nor_5  g13524(new_n14437, new_n15872, new_n15873);
nor_5  g13525(new_n15873, new_n15871, new_n15874);
nand_5 g13526(new_n15874, new_n15870, new_n15875);
not_8  g13527(new_n15875, new_n15876);
nor_5  g13528(new_n15876, new_n15869_1, new_n15877);
nor_5  g13529(new_n15877, new_n15868, new_n15878);
nor_5  g13530(new_n15878, new_n15866, new_n15879);
nor_5  g13531(new_n15879, new_n15865, new_n15880);
nor_5  g13532(new_n15880, new_n15863, new_n15881);
nor_5  g13533(new_n15881, new_n15862, new_n15882);
nor_5  g13534(new_n15882, new_n15860, new_n15883);
xnor_4 g13535(new_n15883, new_n15859_1, new_n15884_1);
xnor_4 g13536(new_n15884_1, new_n7713, new_n15885_1);
xnor_4 g13537(new_n15881, new_n15861, new_n15886);
nand_5 g13538(new_n15886, new_n7716, new_n15887);
xnor_4 g13539(new_n15886, new_n7717, new_n15888);
xnor_4 g13540(new_n15879, new_n15864, new_n15889_1);
nor_5  g13541(new_n15889_1, new_n7722, new_n15890);
xnor_4 g13542(new_n15889_1, new_n7723, new_n15891);
not_8  g13543(new_n15891, new_n15892);
xnor_4 g13544(new_n15877, new_n15867, new_n15893);
nor_5  g13545(new_n15893, new_n7728, new_n15894);
xnor_4 g13546(new_n15893, new_n7726, new_n15895);
not_8  g13547(new_n15895, new_n15896);
not_8  g13548(new_n7730, new_n15897);
xnor_4 g13549(new_n15874, new_n15870, new_n15898);
not_8  g13550(new_n15898, new_n15899);
nand_5 g13551(new_n15899, new_n15897, new_n15900);
xnor_4 g13552(new_n15898, new_n15897, new_n15901);
not_8  g13553(new_n14438, new_n15902);
nand_5 g13554(new_n15902, new_n12888, new_n15903);
nand_5 g13555(new_n14760, new_n14750, new_n15904);
nand_5 g13556(new_n15904, new_n15903, new_n15905);
nand_5 g13557(new_n15905, new_n15901, new_n15906);
nand_5 g13558(new_n15906, new_n15900, new_n15907);
nor_5  g13559(new_n15907, new_n15896, new_n15908);
nor_5  g13560(new_n15908, new_n15894, new_n15909);
nor_5  g13561(new_n15909, new_n15892, new_n15910);
nor_5  g13562(new_n15910, new_n15890, new_n15911);
nand_5 g13563(new_n15911, new_n15888, new_n15912);
nand_5 g13564(new_n15912, new_n15887, new_n15913);
xnor_4 g13565(new_n15913, new_n15885_1, new_n15914);
xnor_4 g13566(n22379, n15077, new_n15915);
nor_5  g13567(n3710, new_n2900, new_n15916);
xnor_4 g13568(n3710, n1662, new_n15917_1);
not_8  g13569(new_n15917_1, new_n15918_1);
nor_5  g13570(n26318, new_n2903, new_n15919);
xnor_4 g13571(n26318, n12875, new_n15920);
not_8  g13572(new_n15920, new_n15921);
nor_5  g13573(n26054, new_n2906, new_n15922_1);
xnor_4 g13574(n26054, n2035, new_n15923);
not_8  g13575(new_n15923, new_n15924);
nor_5  g13576(n19081, new_n2909, new_n15925);
nor_5  g13577(new_n9301, n5213, new_n15926);
nor_5  g13578(new_n9306, n4665, new_n15927);
not_8  g13579(new_n14762, new_n15928);
nor_5  g13580(new_n14774, new_n15928, new_n15929);
nor_5  g13581(new_n15929, new_n15927, new_n15930);
not_8  g13582(new_n15930, new_n15931);
nor_5  g13583(new_n15931, new_n15926, new_n15932);
nor_5  g13584(new_n15932, new_n15925, new_n15933);
nor_5  g13585(new_n15933, new_n15924, new_n15934);
nor_5  g13586(new_n15934, new_n15922_1, new_n15935);
nor_5  g13587(new_n15935, new_n15921, new_n15936_1);
nor_5  g13588(new_n15936_1, new_n15919, new_n15937);
nor_5  g13589(new_n15937, new_n15918_1, new_n15938);
nor_5  g13590(new_n15938, new_n15916, new_n15939);
xnor_4 g13591(new_n15939, new_n15915, new_n15940);
xnor_4 g13592(new_n15940, new_n15914, new_n15941);
xnor_4 g13593(new_n15937, new_n15917_1, new_n15942);
not_8  g13594(new_n15942, new_n15943);
xnor_4 g13595(new_n15911, new_n15888, new_n15944);
nand_5 g13596(new_n15944, new_n15943, new_n15945);
xnor_4 g13597(new_n15944, new_n15942, new_n15946);
xnor_4 g13598(new_n15935, new_n15920, new_n15947_1);
not_8  g13599(new_n15947_1, new_n15948);
xnor_4 g13600(new_n15909, new_n15891, new_n15949);
nand_5 g13601(new_n15949, new_n15948, new_n15950);
xnor_4 g13602(new_n15949, new_n15947_1, new_n15951);
xnor_4 g13603(new_n15933, new_n15923, new_n15952);
not_8  g13604(new_n15952, new_n15953);
xnor_4 g13605(new_n15907, new_n15895, new_n15954);
nand_5 g13606(new_n15954, new_n15953, new_n15955);
xnor_4 g13607(new_n15905, new_n15901, new_n15956_1);
xnor_4 g13608(n19081, n5213, new_n15957);
xnor_4 g13609(new_n15957, new_n15930, new_n15958_1);
nand_5 g13610(new_n15958_1, new_n15956_1, new_n15959);
not_8  g13611(new_n15956_1, new_n15960);
xnor_4 g13612(new_n15958_1, new_n15960, new_n15961);
nand_5 g13613(new_n14775, new_n14761, new_n15962);
nand_5 g13614(new_n14798, new_n14777, new_n15963);
nand_5 g13615(new_n15963, new_n15962, new_n15964);
nand_5 g13616(new_n15964, new_n15961, new_n15965);
nand_5 g13617(new_n15965, new_n15959, new_n15966);
xnor_4 g13618(new_n15954, new_n15952, new_n15967_1);
nand_5 g13619(new_n15967_1, new_n15966, new_n15968);
nand_5 g13620(new_n15968, new_n15955, new_n15969);
nand_5 g13621(new_n15969, new_n15951, new_n15970);
nand_5 g13622(new_n15970, new_n15950, new_n15971);
nand_5 g13623(new_n15971, new_n15946, new_n15972);
nand_5 g13624(new_n15972, new_n15945, new_n15973);
xnor_4 g13625(new_n15973, new_n15941, n2948);
xor_4  g13626(new_n15360, new_n15341, n2961);
xnor_4 g13627(new_n12097, new_n12072_1, n2971);
xnor_4 g13628(new_n2560_1, new_n2537_1, n3010);
xnor_4 g13629(new_n7106, new_n7094, n3017);
xnor_4 g13630(new_n12466, new_n9576, new_n15979_1);
xnor_4 g13631(new_n15979_1, new_n12471, n3020);
xnor_4 g13632(new_n6465_1, new_n6439, n3067);
xnor_4 g13633(n23541, new_n7636, new_n15982);
xnor_4 g13634(n27134, n4588, new_n15983);
xnor_4 g13635(new_n15983, new_n15982, new_n15984);
xnor_4 g13636(new_n15984, new_n10587, n3076);
nor_5  g13637(n15490, n18, new_n15986_1);
nand_5 g13638(new_n15986_1, new_n6947, new_n15987);
xnor_4 g13639(new_n15987, new_n6944, new_n15988);
xnor_4 g13640(new_n15988, new_n8299, new_n15989);
xnor_4 g13641(new_n15986_1, n2783, new_n15990);
not_8  g13642(new_n15990, new_n15991);
nor_5  g13643(new_n15991, new_n6960, new_n15992);
xnor_4 g13644(new_n15990, n19680, new_n15993);
not_8  g13645(n2809, new_n15994);
xnor_4 g13646(n15490, n18, new_n15995);
nand_5 g13647(new_n15995, new_n15994, new_n15996);
nand_5 g13648(n15508, n18, new_n15997);
xnor_4 g13649(new_n15995, n2809, new_n15998);
nand_5 g13650(new_n15998, new_n15997, new_n15999);
nand_5 g13651(new_n15999, new_n15996, new_n16000);
nor_5  g13652(new_n16000, new_n15993, new_n16001);
nor_5  g13653(new_n16001, new_n15992, new_n16002);
xnor_4 g13654(new_n16002, new_n15989, new_n16003);
xnor_4 g13655(new_n16003, new_n11372, new_n16004);
xnor_4 g13656(new_n16000, new_n15993, new_n16005);
nor_5  g13657(new_n16005, new_n11376, new_n16006);
xnor_4 g13658(new_n16005, new_n11376, new_n16007);
nor_5  g13659(new_n15998, new_n6105_1, new_n16008);
not_8  g13660(new_n16008, new_n16009);
xnor_4 g13661(new_n15998, new_n15997, new_n16010);
nand_5 g13662(new_n16010, new_n6105_1, new_n16011);
xnor_4 g13663(n15508, new_n6967_1, new_n16012);
not_8  g13664(new_n16012, new_n16013_1);
nor_5  g13665(new_n16013_1, new_n6085, new_n16014);
not_8  g13666(new_n16014, new_n16015);
nand_5 g13667(new_n16015, new_n16011, new_n16016);
nand_5 g13668(new_n16016, new_n16009, new_n16017);
nor_5  g13669(new_n16017, new_n16007, new_n16018);
nor_5  g13670(new_n16018, new_n16006, new_n16019);
xor_4  g13671(new_n16019, new_n16004, n3089);
xor_4  g13672(new_n5469, new_n5468, n3125);
xnor_4 g13673(n21839, new_n11722, new_n16022);
or_5   g13674(n27089, n12657, new_n16023);
nand_5 g13675(new_n3030_1, new_n2987, new_n16024);
nand_5 g13676(new_n16024, new_n16023, new_n16025);
xnor_4 g13677(new_n16025, new_n16022, new_n16026);
and_5  g13678(new_n16026, new_n11729, new_n16027);
xnor_4 g13679(new_n16026, new_n11728, new_n16028);
not_8  g13680(new_n16028, new_n16029_1);
nor_5  g13681(new_n11733, new_n3031, new_n16030);
nor_5  g13682(new_n11737, new_n3037, new_n16031);
xnor_4 g13683(new_n11737, new_n3035, new_n16032);
not_8  g13684(new_n16032, new_n16033);
nor_5  g13685(new_n11743, new_n3042, new_n16034);
not_8  g13686(new_n16034, new_n16035);
xnor_4 g13687(new_n11741_1, new_n3042, new_n16036);
nor_5  g13688(new_n11749_1, new_n3049, new_n16037);
nor_5  g13689(new_n14193, new_n14169, new_n16038);
nor_5  g13690(new_n16038, new_n16037, new_n16039);
not_8  g13691(new_n16039, new_n16040);
nand_5 g13692(new_n16040, new_n16036, new_n16041);
nand_5 g13693(new_n16041, new_n16035, new_n16042);
nor_5  g13694(new_n16042, new_n16033, new_n16043);
nor_5  g13695(new_n16043, new_n16031, new_n16044);
xnor_4 g13696(new_n11733, new_n3032, new_n16045);
not_8  g13697(new_n16045, new_n16046);
nor_5  g13698(new_n16046, new_n16044, new_n16047);
nor_5  g13699(new_n16047, new_n16030, new_n16048);
nor_5  g13700(new_n16048, new_n16029_1, new_n16049);
nor_5  g13701(new_n16049, new_n16027, new_n16050);
not_8  g13702(new_n16050, new_n16051);
or_5   g13703(n21839, n19282, new_n16052);
nand_5 g13704(new_n16025, new_n16022, new_n16053);
nand_5 g13705(new_n16053, new_n16052, new_n16054);
nand_5 g13706(new_n16054, new_n11731, new_n16055);
nor_5  g13707(new_n16055, new_n16051, new_n16056);
not_8  g13708(new_n16054, new_n16057);
nand_5 g13709(new_n16057, new_n11732, new_n16058);
nor_5  g13710(new_n16058, new_n16050, new_n16059);
nor_5  g13711(new_n16059, new_n16056, new_n16060_1);
xnor_4 g13712(new_n16060_1, new_n12761, new_n16061);
not_8  g13713(new_n12173, new_n16062_1);
xnor_4 g13714(new_n16054, new_n11732, new_n16063);
xnor_4 g13715(new_n16063, new_n16050, new_n16064);
not_8  g13716(new_n16064, new_n16065);
nand_5 g13717(new_n16065, new_n16062_1, new_n16066);
xnor_4 g13718(new_n16064, new_n16062_1, new_n16067);
xnor_4 g13719(new_n16048, new_n16028, new_n16068_1);
nand_5 g13720(new_n16068_1, new_n12184, new_n16069);
xnor_4 g13721(new_n16068_1, new_n12767, new_n16070);
xnor_4 g13722(new_n16045, new_n16044, new_n16071);
nand_5 g13723(new_n16071, new_n12773, new_n16072);
xnor_4 g13724(new_n16071, new_n12192_1, new_n16073);
xnor_4 g13725(new_n16042, new_n16032, new_n16074);
nand_5 g13726(new_n16074, new_n12196, new_n16075);
xnor_4 g13727(new_n16074, new_n12197, new_n16076);
xnor_4 g13728(new_n16040, new_n16036, new_n16077);
nand_5 g13729(new_n16077, new_n12780, new_n16078);
xnor_4 g13730(new_n16077, new_n12203, new_n16079);
nand_5 g13731(new_n14194, new_n12211, new_n16080_1);
nand_5 g13732(new_n14223, new_n14195, new_n16081);
nand_5 g13733(new_n16081, new_n16080_1, new_n16082);
nand_5 g13734(new_n16082, new_n16079, new_n16083);
nand_5 g13735(new_n16083, new_n16078, new_n16084);
nand_5 g13736(new_n16084, new_n16076, new_n16085);
nand_5 g13737(new_n16085, new_n16075, new_n16086);
nand_5 g13738(new_n16086, new_n16073, new_n16087);
nand_5 g13739(new_n16087, new_n16072, new_n16088);
nand_5 g13740(new_n16088, new_n16070, new_n16089);
nand_5 g13741(new_n16089, new_n16069, new_n16090);
nand_5 g13742(new_n16090, new_n16067, new_n16091);
nand_5 g13743(new_n16091, new_n16066, new_n16092);
xnor_4 g13744(new_n16092, new_n16061, n3126);
xnor_4 g13745(new_n12822, new_n12777, n3208);
xnor_4 g13746(new_n15177, new_n15176_1, n3219);
xnor_4 g13747(new_n15624, new_n15615, n3235);
xnor_4 g13748(new_n11963, new_n11948, n3244);
or_5   g13749(new_n8425, n5532, new_n16098_1);
not_8  g13750(n11579, new_n16099);
nor_5  g13751(new_n16099, n3962, new_n16100);
nor_5  g13752(n23513, new_n8432_1, new_n16101);
nand_5 g13753(new_n14447, new_n10575, new_n16102);
not_8  g13754(new_n16102, new_n16103);
nor_5  g13755(n6427, new_n8436, new_n16104);
nor_5  g13756(new_n16104, new_n16103, new_n16105);
nor_5  g13757(new_n16105, new_n10517, new_n16106);
nor_5  g13758(new_n16106, new_n16101, new_n16107);
nor_5  g13759(new_n16107, new_n10539, new_n16108);
nor_5  g13760(new_n16108, new_n16100, new_n16109);
not_8  g13761(new_n16109, new_n16110_1);
nand_5 g13762(new_n16110_1, new_n10542, new_n16111);
nand_5 g13763(new_n16111, new_n16098_1, new_n16112);
xnor_4 g13764(new_n16112, new_n10547, new_n16113);
xnor_4 g13765(new_n16113, new_n15886, new_n16114);
not_8  g13766(new_n15889_1, new_n16115);
xnor_4 g13767(new_n16109, new_n10542, new_n16116);
not_8  g13768(new_n16116, new_n16117);
nand_5 g13769(new_n16117, new_n16115, new_n16118);
xnor_4 g13770(new_n16117, new_n15889_1, new_n16119);
xnor_4 g13771(new_n16107, new_n10538, new_n16120);
nor_5  g13772(new_n16120, new_n15893, new_n16121);
not_8  g13773(new_n16121, new_n16122);
not_8  g13774(new_n16120, new_n16123);
xnor_4 g13775(new_n16123, new_n15893, new_n16124);
xnor_4 g13776(new_n16105, new_n10516, new_n16125);
nor_5  g13777(new_n16125, new_n15899, new_n16126);
not_8  g13778(new_n16126, new_n16127);
xnor_4 g13779(new_n16125, new_n15898, new_n16128);
not_8  g13780(new_n14448, new_n16129);
nor_5  g13781(new_n16129, new_n14438, new_n16130);
not_8  g13782(new_n14449, new_n16131);
nor_5  g13783(new_n14469, new_n16131, new_n16132);
nor_5  g13784(new_n16132, new_n16130, new_n16133);
nand_5 g13785(new_n16133, new_n16128, new_n16134);
nand_5 g13786(new_n16134, new_n16127, new_n16135);
nand_5 g13787(new_n16135, new_n16124, new_n16136);
nand_5 g13788(new_n16136, new_n16122, new_n16137);
nand_5 g13789(new_n16137, new_n16119, new_n16138);
nand_5 g13790(new_n16138, new_n16118, new_n16139);
xnor_4 g13791(new_n16139, new_n16114, new_n16140);
not_8  g13792(n26483, new_n16141);
nor_5  g13793(n23541, n16247, new_n16142_1);
nand_5 g13794(new_n16142_1, new_n2669, new_n16143);
nor_5  g13795(new_n16143, n15979, new_n16144);
nand_5 g13796(new_n16144, new_n16141, new_n16145);
nor_5  g13797(new_n16145, n24768, new_n16146);
nand_5 g13798(new_n16146, new_n2647, new_n16147);
xnor_4 g13799(new_n16147, new_n2642, new_n16148);
xnor_4 g13800(new_n16148, new_n2591, new_n16149);
xnor_4 g13801(new_n16146, n8687, new_n16150);
not_8  g13802(new_n16150, new_n16151);
nand_5 g13803(new_n16151, new_n12150, new_n16152);
xnor_4 g13804(new_n16150, new_n12150, new_n16153);
xnor_4 g13805(new_n16145, n24768, new_n16154);
nand_5 g13806(new_n16154, new_n2599, new_n16155);
xnor_4 g13807(new_n16154, n3460, new_n16156);
xnor_4 g13808(new_n16144, n26483, new_n16157);
not_8  g13809(new_n16157, new_n16158_1);
nand_5 g13810(new_n16158_1, new_n2603, new_n16159);
xnor_4 g13811(new_n16157, new_n2603, new_n16160);
xnor_4 g13812(new_n16143, new_n2664, new_n16161);
not_8  g13813(new_n16161, new_n16162);
nand_5 g13814(new_n16162, new_n10148, new_n16163);
xnor_4 g13815(new_n16142_1, n8638, new_n16164);
not_8  g13816(new_n16164, new_n16165);
nand_5 g13817(new_n16165, new_n2610, new_n16166);
xnor_4 g13818(new_n16164, new_n2610, new_n16167_1);
xnor_4 g13819(n23541, n16247, new_n16168);
nand_5 g13820(new_n16168, new_n9252, new_n16169);
nand_5 g13821(n23541, n19234, new_n16170);
xnor_4 g13822(new_n16168, n1136, new_n16171);
nand_5 g13823(new_n16171, new_n16170, new_n16172);
nand_5 g13824(new_n16172, new_n16169, new_n16173);
nand_5 g13825(new_n16173, new_n16167_1, new_n16174);
nand_5 g13826(new_n16174, new_n16166, new_n16175);
xnor_4 g13827(new_n16161, new_n10148, new_n16176);
nand_5 g13828(new_n16176, new_n16175, new_n16177);
nand_5 g13829(new_n16177, new_n16163, new_n16178);
nand_5 g13830(new_n16178, new_n16160, new_n16179);
nand_5 g13831(new_n16179, new_n16159, new_n16180);
nand_5 g13832(new_n16180, new_n16156, new_n16181);
nand_5 g13833(new_n16181, new_n16155, new_n16182);
nand_5 g13834(new_n16182, new_n16153, new_n16183);
nand_5 g13835(new_n16183, new_n16152, new_n16184);
xnor_4 g13836(new_n16184, new_n16149, new_n16185_1);
xnor_4 g13837(new_n16185_1, new_n16140, new_n16186);
xnor_4 g13838(new_n16182, new_n16153, new_n16187);
not_8  g13839(new_n16187, new_n16188);
xnor_4 g13840(new_n16137, new_n16119, new_n16189);
not_8  g13841(new_n16189, new_n16190);
nand_5 g13842(new_n16190, new_n16188, new_n16191);
not_8  g13843(new_n16156, new_n16192);
xnor_4 g13844(new_n16180, new_n16192, new_n16193);
not_8  g13845(new_n16124, new_n16194);
xnor_4 g13846(new_n16135, new_n16194, new_n16195);
nand_5 g13847(new_n16195, new_n16193, new_n16196_1);
not_8  g13848(new_n16193, new_n16197);
xnor_4 g13849(new_n16195, new_n16197, new_n16198);
xnor_4 g13850(new_n16178, new_n16160, new_n16199);
not_8  g13851(new_n16199, new_n16200);
not_8  g13852(new_n16128, new_n16201);
xnor_4 g13853(new_n16133, new_n16201, new_n16202);
nand_5 g13854(new_n16202, new_n16200, new_n16203);
not_8  g13855(new_n14470, new_n16204);
xnor_4 g13856(new_n16176, new_n16175, new_n16205);
not_8  g13857(new_n16205, new_n16206_1);
nand_5 g13858(new_n16206_1, new_n16204, new_n16207);
xnor_4 g13859(new_n16206_1, new_n14470, new_n16208);
not_8  g13860(new_n16167_1, new_n16209);
xnor_4 g13861(new_n16173, new_n16209, new_n16210);
nor_5  g13862(new_n16210, new_n14485, new_n16211);
xnor_4 g13863(new_n16210, new_n14486, new_n16212);
not_8  g13864(new_n16212, new_n16213);
xnor_4 g13865(new_n16171, new_n16170, new_n16214);
nor_5  g13866(new_n16214, new_n14503, new_n16215_1);
not_8  g13867(new_n15982, new_n16216);
nor_5  g13868(new_n16216, new_n14494, new_n16217_1);
xnor_4 g13869(new_n16214, new_n14502, new_n16218_1);
not_8  g13870(new_n16218_1, new_n16219_1);
nor_5  g13871(new_n16219_1, new_n16217_1, new_n16220);
nor_5  g13872(new_n16220, new_n16215_1, new_n16221);
not_8  g13873(new_n16221, new_n16222);
nor_5  g13874(new_n16222, new_n16213, new_n16223_1);
nor_5  g13875(new_n16223_1, new_n16211, new_n16224);
nand_5 g13876(new_n16224, new_n16208, new_n16225);
nand_5 g13877(new_n16225, new_n16207, new_n16226);
xnor_4 g13878(new_n16202, new_n16199, new_n16227);
nand_5 g13879(new_n16227, new_n16226, new_n16228);
nand_5 g13880(new_n16228, new_n16203, new_n16229);
nand_5 g13881(new_n16229, new_n16198, new_n16230_1);
nand_5 g13882(new_n16230_1, new_n16196_1, new_n16231);
xnor_4 g13883(new_n16189, new_n16188, new_n16232);
nand_5 g13884(new_n16232, new_n16231, new_n16233);
nand_5 g13885(new_n16233, new_n16191, new_n16234);
xnor_4 g13886(new_n16234, new_n16186, n3263);
xnor_4 g13887(new_n13046, new_n13029, n3289);
not_8  g13888(n18537, new_n16237);
xnor_4 g13889(n21832, new_n2955, new_n16238);
nand_5 g13890(n26913, n12956, new_n16239);
nor_5  g13891(n26913, n12956, new_n16240);
not_8  g13892(new_n16240, new_n16241);
nor_5  g13893(n18295, n16223, new_n16242);
nor_5  g13894(new_n5304, new_n5297, new_n16243_1);
nor_5  g13895(new_n16243_1, new_n16242, new_n16244);
nand_5 g13896(new_n16244, new_n16241, new_n16245);
nand_5 g13897(new_n16245, new_n16239, new_n16246);
xnor_4 g13898(new_n16246, new_n16238, new_n16247_1);
xnor_4 g13899(new_n16247_1, new_n16237, new_n16248);
not_8  g13900(new_n16248, new_n16249);
xnor_4 g13901(n26913, new_n9546, new_n16250);
not_8  g13902(new_n16250, new_n16251);
xnor_4 g13903(new_n16251, new_n16244, new_n16252);
not_8  g13904(new_n16252, new_n16253);
nor_5  g13905(new_n16253, n7057, new_n16254);
xnor_4 g13906(new_n16252, n7057, new_n16255);
not_8  g13907(new_n16255, new_n16256);
nor_5  g13908(new_n5305, n8381, new_n16257);
not_8  g13909(new_n5306, new_n16258);
nor_5  g13910(new_n5316, new_n16258, new_n16259);
nor_5  g13911(new_n16259, new_n16257, new_n16260);
nor_5  g13912(new_n16260, new_n16256, new_n16261);
nor_5  g13913(new_n16261, new_n16254, new_n16262);
xnor_4 g13914(new_n16262, new_n16249, new_n16263);
not_8  g13915(new_n16263, new_n16264);
xnor_4 g13916(new_n15249, n21649, new_n16265);
nand_5 g13917(new_n10042, new_n5432, new_n16266);
xnor_4 g13918(new_n10042, n18274, new_n16267);
nand_5 g13919(new_n10062, new_n5436, new_n16268);
nor_5  g13920(new_n10068, n23842, new_n16269);
not_8  g13921(new_n16269, new_n16270);
not_8  g13922(n21654, new_n16271);
nor_5  g13923(new_n10071, new_n16271, new_n16272);
not_8  g13924(new_n16272, new_n16273);
xnor_4 g13925(new_n10067, n23842, new_n16274);
nand_5 g13926(new_n16274, new_n16273, new_n16275_1);
nand_5 g13927(new_n16275_1, new_n16270, new_n16276);
xnor_4 g13928(new_n10062, n3828, new_n16277);
nand_5 g13929(new_n16277, new_n16276, new_n16278);
nand_5 g13930(new_n16278, new_n16268, new_n16279_1);
nand_5 g13931(new_n16279_1, new_n16267, new_n16280);
nand_5 g13932(new_n16280, new_n16266, new_n16281);
xnor_4 g13933(new_n16281, new_n16265, new_n16282);
xnor_4 g13934(new_n16282, new_n16264, new_n16283);
xnor_4 g13935(new_n16260, new_n16255, new_n16284);
xnor_4 g13936(new_n16279_1, new_n16267, new_n16285);
not_8  g13937(new_n16285, new_n16286);
nand_5 g13938(new_n16286, new_n16284, new_n16287);
xnor_4 g13939(new_n16285, new_n16284, new_n16288);
not_8  g13940(new_n16277, new_n16289);
xnor_4 g13941(new_n16289, new_n16276, new_n16290);
nand_5 g13942(new_n16290, new_n5317, new_n16291);
xnor_4 g13943(new_n16274, new_n16273, new_n16292);
not_8  g13944(new_n16292, new_n16293);
nand_5 g13945(new_n16293, new_n5343, new_n16294);
not_8  g13946(new_n5347, new_n16295);
xnor_4 g13947(new_n10070, new_n16271, new_n16296);
nand_5 g13948(new_n16296, new_n16295, new_n16297);
xnor_4 g13949(new_n16292, new_n5343, new_n16298);
nand_5 g13950(new_n16298, new_n16297, new_n16299);
nand_5 g13951(new_n16299, new_n16294, new_n16300);
not_8  g13952(new_n5317, new_n16301);
xnor_4 g13953(new_n16290, new_n16301, new_n16302);
nand_5 g13954(new_n16302, new_n16300, new_n16303);
nand_5 g13955(new_n16303, new_n16291, new_n16304);
nand_5 g13956(new_n16304, new_n16288, new_n16305);
nand_5 g13957(new_n16305, new_n16287, new_n16306);
xnor_4 g13958(new_n16306, new_n16283, n3301);
xnor_4 g13959(new_n11421, n3030, new_n16308);
not_8  g13960(n19515, new_n16309);
nor_5  g13961(new_n11414, new_n16309, new_n16310);
xnor_4 g13962(new_n11414, n19515, new_n16311);
not_8  g13963(new_n16311, new_n16312);
nor_5  g13964(new_n11405, new_n14472, new_n16313);
xnor_4 g13965(new_n11405, n22588, new_n16314);
nor_5  g13966(new_n11397, n12209, new_n16315);
not_8  g13967(new_n14232, new_n16316);
nor_5  g13968(new_n16316, new_n14231, new_n16317);
nor_5  g13969(new_n16317, new_n16315, new_n16318);
nand_5 g13970(new_n16318, new_n16314, new_n16319);
not_8  g13971(new_n16319, new_n16320);
nor_5  g13972(new_n16320, new_n16313, new_n16321);
nor_5  g13973(new_n16321, new_n16312, new_n16322_1);
nor_5  g13974(new_n16322_1, new_n16310, new_n16323);
xnor_4 g13975(new_n16323, new_n16308, new_n16324);
xnor_4 g13976(new_n16324, new_n10648, new_n16325);
xnor_4 g13977(new_n16321, new_n16311, new_n16326);
not_8  g13978(new_n16326, new_n16327_1);
nor_5  g13979(new_n16327_1, new_n10654, new_n16328);
xnor_4 g13980(new_n16326, new_n10655, new_n16329);
xnor_4 g13981(new_n16318, new_n16314, new_n16330);
nor_5  g13982(new_n16330, new_n10660, new_n16331);
xnor_4 g13983(new_n16330, new_n10660, new_n16332);
nor_5  g13984(new_n14233, new_n10673, new_n16333);
nor_5  g13985(new_n14234, new_n14230_1, new_n16334);
nor_5  g13986(new_n16334, new_n16333, new_n16335);
nor_5  g13987(new_n16335, new_n16332, new_n16336);
nor_5  g13988(new_n16336, new_n16331, new_n16337);
nor_5  g13989(new_n16337, new_n16329, new_n16338);
nor_5  g13990(new_n16338, new_n16328, new_n16339);
xor_4  g13991(new_n16339, new_n16325, n3316);
xnor_4 g13992(new_n14217, new_n14202, n3332);
not_8  g13993(new_n8463, new_n16342);
nand_5 g13994(new_n16342, new_n11675, new_n16343);
xnor_4 g13995(new_n8463, new_n11675, new_n16344);
nand_5 g13996(new_n11463, new_n11678, new_n16345);
xnor_4 g13997(new_n8467, new_n11678, new_n16346);
nand_5 g13998(new_n8471, new_n11681, new_n16347);
nand_5 g13999(new_n11192_1, new_n11173, new_n16348);
nand_5 g14000(new_n16348, new_n16347, new_n16349);
nand_5 g14001(new_n16349, new_n16346, new_n16350_1);
nand_5 g14002(new_n16350_1, new_n16345, new_n16351);
nand_5 g14003(new_n16351, new_n16344, new_n16352);
nand_5 g14004(new_n16352, new_n16343, new_n16353);
nor_5  g14005(new_n16353, new_n8528, new_n16354);
and_5  g14006(new_n13693, n8827, new_n16355);
not_8  g14007(new_n13694, new_n16356);
nor_5  g14008(new_n13707, new_n16356, new_n16357);
nor_5  g14009(new_n16357, new_n16355, new_n16358);
nor_5  g14010(n23166, n11898, new_n16359);
and_5  g14011(new_n13692, new_n13682, new_n16360);
nor_5  g14012(new_n16360, new_n16359, new_n16361);
not_8  g14013(new_n16361, new_n16362);
nor_5  g14014(new_n16362, new_n16358, new_n16363);
xnor_4 g14015(new_n16363, new_n16354, new_n16364);
xnor_4 g14016(new_n16353, new_n8529, new_n16365);
not_8  g14017(new_n16365, new_n16366);
xnor_4 g14018(new_n16361, new_n16358, new_n16367_1);
nand_5 g14019(new_n16367_1, new_n16366, new_n16368);
xnor_4 g14020(new_n16367_1, new_n16365, new_n16369);
not_8  g14021(new_n16344, new_n16370);
xnor_4 g14022(new_n16351, new_n16370, new_n16371);
nor_5  g14023(new_n16371, new_n13708_1, new_n16372);
xnor_4 g14024(new_n16371, new_n13708_1, new_n16373);
not_8  g14025(new_n16346, new_n16374);
xnor_4 g14026(new_n16349, new_n16374, new_n16375);
nand_5 g14027(new_n16375, new_n13710_1, new_n16376_1);
not_8  g14028(new_n11193, new_n16377);
nand_5 g14029(new_n11250, new_n16377, new_n16378);
nand_5 g14030(new_n11279, new_n11251, new_n16379_1);
nand_5 g14031(new_n16379_1, new_n16378, new_n16380);
xnor_4 g14032(new_n16375, new_n13712, new_n16381);
nand_5 g14033(new_n16381, new_n16380, new_n16382);
nand_5 g14034(new_n16382, new_n16376_1, new_n16383);
nor_5  g14035(new_n16383, new_n16373, new_n16384);
nor_5  g14036(new_n16384, new_n16372, new_n16385);
nand_5 g14037(new_n16385, new_n16369, new_n16386);
nand_5 g14038(new_n16386, new_n16368, new_n16387);
xnor_4 g14039(new_n16387, new_n16364, n3340);
xnor_4 g14040(n13851, n5077, new_n16389);
not_8  g14041(new_n16389, new_n16390);
nor_5  g14042(n24937, new_n11222, new_n16391);
xnor_4 g14043(n24937, n15546, new_n16392);
not_8  g14044(new_n16392, new_n16393);
nor_5  g14045(new_n11244, n5098, new_n16394);
xnor_4 g14046(n26452, n5098, new_n16395);
not_8  g14047(new_n16395, new_n16396_1);
nor_5  g14048(new_n11231, n3030, new_n16397);
xnor_4 g14049(n19905, n3030, new_n16398_1);
nor_5  g14050(new_n16309, n17035, new_n16399);
not_8  g14051(new_n14471_1, new_n16400);
nor_5  g14052(new_n14482, new_n16400, new_n16401);
nor_5  g14053(new_n16401, new_n16399, new_n16402);
and_5  g14054(new_n16402, new_n16398_1, new_n16403);
nor_5  g14055(new_n16403, new_n16397, new_n16404);
nor_5  g14056(new_n16404, new_n16396_1, new_n16405);
nor_5  g14057(new_n16405, new_n16394, new_n16406_1);
nor_5  g14058(new_n16406_1, new_n16393, new_n16407_1);
nor_5  g14059(new_n16407_1, new_n16391, new_n16408);
xnor_4 g14060(new_n16408, new_n16390, new_n16409);
xnor_4 g14061(new_n16409, new_n16140, new_n16410);
xnor_4 g14062(new_n16406_1, new_n16392, new_n16411);
not_8  g14063(new_n16411, new_n16412);
nand_5 g14064(new_n16412, new_n16190, new_n16413);
xnor_4 g14065(new_n16411, new_n16190, new_n16414);
xnor_4 g14066(new_n16404, new_n16395, new_n16415);
not_8  g14067(new_n16415, new_n16416);
nand_5 g14068(new_n16416, new_n16195, new_n16417);
xnor_4 g14069(new_n16415, new_n16195, new_n16418);
xnor_4 g14070(new_n16402, new_n16398_1, new_n16419_1);
nor_5  g14071(new_n16419_1, new_n16202, new_n16420);
xnor_4 g14072(new_n16419_1, new_n16202, new_n16421);
not_8  g14073(new_n14483, new_n16422);
nor_5  g14074(new_n16422, new_n14470, new_n16423);
not_8  g14075(new_n16423, new_n16424_1);
nand_5 g14076(new_n14510_1, new_n14484, new_n16425);
nand_5 g14077(new_n16425, new_n16424_1, new_n16426);
nor_5  g14078(new_n16426, new_n16421, new_n16427);
nor_5  g14079(new_n16427, new_n16420, new_n16428_1);
nand_5 g14080(new_n16428_1, new_n16418, new_n16429);
nand_5 g14081(new_n16429, new_n16417, new_n16430);
nand_5 g14082(new_n16430, new_n16414, new_n16431);
nand_5 g14083(new_n16431, new_n16413, new_n16432);
xor_4  g14084(new_n16432, new_n16410, n3343);
nor_5  g14085(new_n16147, n19270, new_n16434);
nand_5 g14086(new_n16434, new_n2636, new_n16435);
or_5   g14087(new_n16435, n25365, new_n16436);
xnor_4 g14088(new_n16435, new_n15571, new_n16437);
or_5   g14089(new_n16437, n20040, new_n16438);
xnor_4 g14090(new_n16434, n14704, new_n16439_1);
not_8  g14091(new_n16439_1, new_n16440_1);
nand_5 g14092(new_n16440_1, new_n12142, new_n16441);
xnor_4 g14093(new_n16439_1, new_n12142, new_n16442);
not_8  g14094(new_n16148, new_n16443);
nand_5 g14095(new_n16443, new_n2591, new_n16444);
nand_5 g14096(new_n16184, new_n16149, new_n16445_1);
nand_5 g14097(new_n16445_1, new_n16444, new_n16446);
nand_5 g14098(new_n16446, new_n16442, new_n16447);
nand_5 g14099(new_n16447, new_n16441, new_n16448);
nand_5 g14100(new_n16437, n20040, new_n16449);
nand_5 g14101(new_n16449, new_n16448, new_n16450);
nand_5 g14102(new_n16450, new_n16438, new_n16451);
nand_5 g14103(new_n16451, new_n16436, new_n16452);
not_8  g14104(new_n16452, new_n16453);
not_8  g14105(new_n14864, new_n16454);
xnor_4 g14106(new_n16437, new_n12132, new_n16455);
xnor_4 g14107(new_n16455, new_n16448, new_n16456);
not_8  g14108(new_n16456, new_n16457);
nor_5  g14109(new_n16457, new_n16454, new_n16458);
nand_5 g14110(new_n16457, new_n16454, new_n16459);
xnor_4 g14111(new_n16446, new_n16442, new_n16460_1);
nand_5 g14112(new_n16460_1, new_n14846, new_n16461);
xnor_4 g14113(new_n16460_1, new_n14847, new_n16462);
nand_5 g14114(new_n16185_1, new_n14850, new_n16463);
xnor_4 g14115(new_n16185_1, new_n14851, new_n16464);
nand_5 g14116(new_n16187, new_n6813, new_n16465);
xnor_4 g14117(new_n16187, new_n14854, new_n16466);
nand_5 g14118(new_n16197, new_n6817, new_n16467);
nor_5  g14119(new_n16200, new_n6823, new_n16468);
not_8  g14120(new_n16468, new_n16469);
xnor_4 g14121(new_n16199, new_n6823, new_n16470);
nor_5  g14122(new_n16205, new_n6828, new_n16471);
xnor_4 g14123(new_n16205, new_n6829, new_n16472);
not_8  g14124(new_n16472, new_n16473);
nor_5  g14125(new_n16210, new_n6833, new_n16474);
not_8  g14126(new_n16474, new_n16475);
xnor_4 g14127(new_n16210, new_n6832, new_n16476_1);
not_8  g14128(new_n6837, new_n16477);
nor_5  g14129(new_n16214, new_n16477, new_n16478);
nor_5  g14130(new_n16216, new_n6880, new_n16479);
xnor_4 g14131(new_n16214, new_n16477, new_n16480);
nor_5  g14132(new_n16480, new_n16479, new_n16481_1);
nor_5  g14133(new_n16481_1, new_n16478, new_n16482_1);
nand_5 g14134(new_n16482_1, new_n16476_1, new_n16483);
nand_5 g14135(new_n16483, new_n16475, new_n16484);
nor_5  g14136(new_n16484, new_n16473, new_n16485);
nor_5  g14137(new_n16485, new_n16471, new_n16486);
nand_5 g14138(new_n16486, new_n16470, new_n16487);
nand_5 g14139(new_n16487, new_n16469, new_n16488);
xnor_4 g14140(new_n16193, new_n6817, new_n16489);
nand_5 g14141(new_n16489, new_n16488, new_n16490);
nand_5 g14142(new_n16490, new_n16467, new_n16491);
nand_5 g14143(new_n16491, new_n16466, new_n16492);
nand_5 g14144(new_n16492, new_n16465, new_n16493_1);
nand_5 g14145(new_n16493_1, new_n16464, new_n16494);
nand_5 g14146(new_n16494, new_n16463, new_n16495);
nand_5 g14147(new_n16495, new_n16462, new_n16496);
nand_5 g14148(new_n16496, new_n16461, new_n16497);
nand_5 g14149(new_n16497, new_n16459, new_n16498);
nand_5 g14150(new_n16498, new_n14889, new_n16499);
nor_5  g14151(new_n16499, new_n16458, new_n16500);
xnor_4 g14152(new_n16500, new_n16453, new_n16501);
not_8  g14153(new_n16501, new_n16502_1);
not_8  g14154(n10250, new_n16503);
not_8  g14155(new_n13220, new_n16504);
nand_5 g14156(new_n16504, new_n16503, new_n16505);
xnor_4 g14157(new_n13220, new_n16503, new_n16506_1);
not_8  g14158(new_n13225, new_n16507_1);
nand_5 g14159(new_n16507_1, new_n6481, new_n16508);
xnor_4 g14160(new_n13225, new_n6481, new_n16509);
not_8  g14161(new_n13230, new_n16510);
nand_5 g14162(new_n16510, new_n6484, new_n16511);
xnor_4 g14163(new_n13230, new_n6484, new_n16512);
nand_5 g14164(new_n13239, new_n6487, new_n16513);
xnor_4 g14165(new_n13235, new_n6487, new_n16514);
nand_5 g14166(new_n13241, new_n12714, new_n16515);
xnor_4 g14167(new_n13241, n23586, new_n16516_1);
not_8  g14168(n21226, new_n16517_1);
nand_5 g14169(new_n13247, new_n16517_1, new_n16518);
xnor_4 g14170(new_n13247, n21226, new_n16519);
nand_5 g14171(new_n13257, new_n6497, new_n16520);
xnor_4 g14172(new_n13253, new_n6497, new_n16521_1);
nand_5 g14173(new_n13262, new_n9210, new_n16522);
xnor_4 g14174(new_n13261, new_n9210, new_n16523);
nor_5  g14175(new_n13272, new_n4305, new_n16524_1);
nor_5  g14176(new_n13268, n9380, new_n16525);
xnor_4 g14177(new_n13271, new_n4305, new_n16526);
not_8  g14178(new_n16526, new_n16527_1);
nor_5  g14179(new_n16527_1, new_n16525, new_n16528);
nor_5  g14180(new_n16528, new_n16524_1, new_n16529);
nand_5 g14181(new_n16529, new_n16523, new_n16530);
nand_5 g14182(new_n16530, new_n16522, new_n16531);
nand_5 g14183(new_n16531, new_n16521_1, new_n16532);
nand_5 g14184(new_n16532, new_n16520, new_n16533);
nand_5 g14185(new_n16533, new_n16519, new_n16534);
nand_5 g14186(new_n16534, new_n16518, new_n16535);
nand_5 g14187(new_n16535, new_n16516_1, new_n16536);
nand_5 g14188(new_n16536, new_n16515, new_n16537);
nand_5 g14189(new_n16537, new_n16514, new_n16538);
nand_5 g14190(new_n16538, new_n16513, new_n16539);
nand_5 g14191(new_n16539, new_n16512, new_n16540);
nand_5 g14192(new_n16540, new_n16511, new_n16541);
nand_5 g14193(new_n16541, new_n16509, new_n16542);
nand_5 g14194(new_n16542, new_n16508, new_n16543);
nand_5 g14195(new_n16543, new_n16506_1, new_n16544_1);
nand_5 g14196(new_n16544_1, new_n16505, new_n16545);
xnor_4 g14197(new_n16545, new_n13110_1, new_n16546);
nor_5  g14198(new_n16546, new_n16502_1, new_n16547);
xnor_4 g14199(new_n16543, new_n16506_1, new_n16548);
not_8  g14200(new_n16548, new_n16549);
xnor_4 g14201(new_n16456, new_n16454, new_n16550);
xnor_4 g14202(new_n16550, new_n16497, new_n16551);
nand_5 g14203(new_n16551, new_n16549, new_n16552);
xnor_4 g14204(new_n16551, new_n16548, new_n16553);
xnor_4 g14205(new_n16541, new_n16509, new_n16554_1);
not_8  g14206(new_n16554_1, new_n16555);
xnor_4 g14207(new_n16495, new_n16462, new_n16556);
nand_5 g14208(new_n16556, new_n16555, new_n16557);
xnor_4 g14209(new_n16556, new_n16554_1, new_n16558);
xnor_4 g14210(new_n16539, new_n16512, new_n16559);
not_8  g14211(new_n16559, new_n16560);
xnor_4 g14212(new_n16493_1, new_n16464, new_n16561);
nand_5 g14213(new_n16561, new_n16560, new_n16562);
xnor_4 g14214(new_n16561, new_n16559, new_n16563);
xnor_4 g14215(new_n16537, new_n16514, new_n16564);
not_8  g14216(new_n16564, new_n16565);
xnor_4 g14217(new_n16491, new_n16466, new_n16566);
nand_5 g14218(new_n16566, new_n16565, new_n16567);
xnor_4 g14219(new_n16566, new_n16564, new_n16568);
xnor_4 g14220(new_n16535, new_n16516_1, new_n16569);
not_8  g14221(new_n16569, new_n16570);
xnor_4 g14222(new_n16489, new_n16488, new_n16571);
nand_5 g14223(new_n16571, new_n16570, new_n16572);
xnor_4 g14224(new_n16571, new_n16569, new_n16573);
xnor_4 g14225(new_n16533, new_n16519, new_n16574);
not_8  g14226(new_n16574, new_n16575);
xnor_4 g14227(new_n16486, new_n16470, new_n16576);
nand_5 g14228(new_n16576, new_n16575, new_n16577);
xnor_4 g14229(new_n16576, new_n16574, new_n16578);
not_8  g14230(new_n16521_1, new_n16579);
xnor_4 g14231(new_n16531, new_n16579, new_n16580);
xnor_4 g14232(new_n16484, new_n16472, new_n16581);
nand_5 g14233(new_n16581, new_n16580, new_n16582);
not_8  g14234(new_n16581, new_n16583_1);
xnor_4 g14235(new_n16583_1, new_n16580, new_n16584_1);
xnor_4 g14236(new_n16529, new_n16523, new_n16585);
not_8  g14237(new_n16585, new_n16586);
xnor_4 g14238(new_n16482_1, new_n16476_1, new_n16587);
nand_5 g14239(new_n16587, new_n16586, new_n16588);
xnor_4 g14240(new_n16480, new_n16479, new_n16589_1);
not_8  g14241(new_n16589_1, new_n16590);
xnor_4 g14242(new_n16526, new_n16525, new_n16591);
not_8  g14243(new_n16591, new_n16592);
nor_5  g14244(new_n16592, new_n16590, new_n16593);
xnor_4 g14245(new_n15982, new_n6880, new_n16594);
not_8  g14246(new_n16594, new_n16595);
xnor_4 g14247(new_n13268, new_n4307, new_n16596_1);
nor_5  g14248(new_n16596_1, new_n16595, new_n16597);
not_8  g14249(new_n16597, new_n16598);
xnor_4 g14250(new_n16591, new_n16589_1, new_n16599);
nor_5  g14251(new_n16599, new_n16598, new_n16600);
nor_5  g14252(new_n16600, new_n16593, new_n16601);
xnor_4 g14253(new_n16587, new_n16585, new_n16602);
nand_5 g14254(new_n16602, new_n16601, new_n16603);
nand_5 g14255(new_n16603, new_n16588, new_n16604);
nand_5 g14256(new_n16604, new_n16584_1, new_n16605);
nand_5 g14257(new_n16605, new_n16582, new_n16606);
nand_5 g14258(new_n16606, new_n16578, new_n16607);
nand_5 g14259(new_n16607, new_n16577, new_n16608_1);
nand_5 g14260(new_n16608_1, new_n16573, new_n16609);
nand_5 g14261(new_n16609, new_n16572, new_n16610);
nand_5 g14262(new_n16610, new_n16568, new_n16611);
nand_5 g14263(new_n16611, new_n16567, new_n16612);
nand_5 g14264(new_n16612, new_n16563, new_n16613);
nand_5 g14265(new_n16613, new_n16562, new_n16614);
nand_5 g14266(new_n16614, new_n16558, new_n16615);
nand_5 g14267(new_n16615, new_n16557, new_n16616);
nand_5 g14268(new_n16616, new_n16553, new_n16617_1);
nand_5 g14269(new_n16617_1, new_n16552, new_n16618);
xnor_4 g14270(new_n16546, new_n16501, new_n16619);
nand_5 g14271(new_n16619, new_n16618, new_n16620);
not_8  g14272(new_n16620, new_n16621);
nor_5  g14273(new_n16621, new_n16547, new_n16622);
not_8  g14274(new_n16622, new_n16623);
nand_5 g14275(new_n16500, new_n16452, new_n16624);
not_8  g14276(new_n16545, new_n16625);
nand_5 g14277(new_n16625, new_n13110_1, new_n16626);
xnor_4 g14278(new_n16626, new_n16624, new_n16627);
xnor_4 g14279(new_n16627, new_n16623, n3390);
xnor_4 g14280(new_n6927, new_n6925, n3426);
xnor_4 g14281(new_n4971, new_n4969, n3451);
xnor_4 g14282(new_n12953, new_n12930, n3459);
xnor_4 g14283(n6773, n583, new_n16632);
xnor_4 g14284(new_n16632, new_n2574, new_n16633);
nor_5  g14285(new_n16633, new_n14602, new_n16634);
not_8  g14286(new_n16634, new_n16635);
nand_5 g14287(new_n16632, n21687, new_n16636);
nand_5 g14288(new_n16636, new_n4238, new_n16637);
nand_5 g14289(n21687, n6729, new_n16638);
not_8  g14290(new_n16638, new_n16639);
nand_5 g14291(new_n16632, new_n16639, new_n16640_1);
nand_5 g14292(new_n16640_1, new_n16637, new_n16641);
nand_5 g14293(n6773, n583, new_n16642);
not_8  g14294(new_n16642, new_n16643);
xnor_4 g14295(n22173, new_n4201, new_n16644);
xnor_4 g14296(new_n16644, new_n16643, new_n16645);
xnor_4 g14297(new_n16645, new_n16641, new_n16646);
xnor_4 g14298(new_n16646, new_n14594, new_n16647);
xnor_4 g14299(new_n16647, new_n16635, n3502);
xnor_4 g14300(new_n11566_1, new_n11525, n3516);
not_8  g14301(n25126, new_n16650);
nor_5  g14302(n24129, n22274, new_n16651);
nand_5 g14303(new_n16651, new_n4301, new_n16652);
nor_5  g14304(new_n16652, n19608, new_n16653);
nand_5 g14305(new_n16653, new_n16650, new_n16654);
nor_5  g14306(new_n16654, n10712, new_n16655);
xnor_4 g14307(new_n16655, n18145, new_n16656_1);
xnor_4 g14308(new_n16656_1, n15761, new_n16657);
not_8  g14309(n10712, new_n16658);
xnor_4 g14310(new_n16654, new_n16658, new_n16659);
not_8  g14311(new_n16659, new_n16660);
nand_5 g14312(new_n16660, n11201, new_n16661);
xnor_4 g14313(new_n16659, n11201, new_n16662);
xnor_4 g14314(new_n16653, n25126, new_n16663);
not_8  g14315(new_n16663, new_n16664);
nand_5 g14316(new_n16664, n18690, new_n16665);
xnor_4 g14317(new_n16663, n18690, new_n16666);
not_8  g14318(n19608, new_n16667);
xnor_4 g14319(new_n16652, new_n16667, new_n16668);
not_8  g14320(new_n16668, new_n16669);
nand_5 g14321(new_n16669, n12153, new_n16670);
xnor_4 g14322(new_n16668, n12153, new_n16671);
xnor_4 g14323(new_n16651, n1689, new_n16672);
not_8  g14324(new_n16672, new_n16673);
nand_5 g14325(new_n16673, n13044, new_n16674_1);
xnor_4 g14326(new_n16672, n13044, new_n16675);
xnor_4 g14327(n24129, n22274, new_n16676);
nand_5 g14328(new_n16676, n18745, new_n16677);
nor_5  g14329(n24129, new_n6120, new_n16678);
xnor_4 g14330(new_n16676, new_n6122, new_n16679);
nand_5 g14331(new_n16679, new_n16678, new_n16680);
nand_5 g14332(new_n16680, new_n16677, new_n16681);
nand_5 g14333(new_n16681, new_n16675, new_n16682_1);
nand_5 g14334(new_n16682_1, new_n16674_1, new_n16683);
nand_5 g14335(new_n16683, new_n16671, new_n16684_1);
nand_5 g14336(new_n16684_1, new_n16670, new_n16685);
nand_5 g14337(new_n16685, new_n16666, new_n16686);
nand_5 g14338(new_n16686, new_n16665, new_n16687);
nand_5 g14339(new_n16687, new_n16662, new_n16688_1);
nand_5 g14340(new_n16688_1, new_n16661, new_n16689);
xnor_4 g14341(new_n16689, new_n16657, new_n16690);
xnor_4 g14342(new_n16690, new_n7256_1, new_n16691);
xnor_4 g14343(new_n16687, new_n16662, new_n16692);
not_8  g14344(new_n16692, new_n16693);
nand_5 g14345(new_n16693, new_n7260, new_n16694);
xnor_4 g14346(new_n16692, new_n7260, new_n16695);
xnor_4 g14347(new_n16685, new_n16666, new_n16696);
not_8  g14348(new_n16696, new_n16697);
nand_5 g14349(new_n16697, new_n7264, new_n16698);
xnor_4 g14350(new_n16696, new_n7264, new_n16699);
xnor_4 g14351(new_n16683, new_n16671, new_n16700);
nor_5  g14352(new_n16700, new_n7270, new_n16701);
not_8  g14353(new_n16701, new_n16702);
xnor_4 g14354(new_n16700, new_n12719, new_n16703);
xnor_4 g14355(new_n16681, new_n16675, new_n16704);
not_8  g14356(new_n16704, new_n16705);
nor_5  g14357(new_n16705, new_n4300, new_n16706);
xnor_4 g14358(new_n16704, new_n4300, new_n16707);
not_8  g14359(new_n16707, new_n16708);
xnor_4 g14360(new_n16679, new_n16678, new_n16709);
nand_5 g14361(new_n16709, new_n7275, new_n16710);
xnor_4 g14362(n24129, n16167, new_n16711);
nor_5  g14363(new_n16711, new_n4317, new_n16712);
xnor_4 g14364(new_n16709, new_n4313, new_n16713);
nand_5 g14365(new_n16713, new_n16712, new_n16714);
nand_5 g14366(new_n16714, new_n16710, new_n16715);
not_8  g14367(new_n16715, new_n16716);
nor_5  g14368(new_n16716, new_n16708, new_n16717);
nor_5  g14369(new_n16717, new_n16706, new_n16718);
nand_5 g14370(new_n16718, new_n16703, new_n16719);
nand_5 g14371(new_n16719, new_n16702, new_n16720);
nand_5 g14372(new_n16720, new_n16699, new_n16721);
nand_5 g14373(new_n16721, new_n16698, new_n16722_1);
nand_5 g14374(new_n16722_1, new_n16695, new_n16723);
nand_5 g14375(new_n16723, new_n16694, new_n16724);
xnor_4 g14376(new_n16724, new_n16691, new_n16725);
xnor_4 g14377(new_n16725, new_n11038, new_n16726);
xnor_4 g14378(new_n16722_1, new_n16695, new_n16727);
not_8  g14379(new_n16727, new_n16728);
nand_5 g14380(new_n16728, new_n11043, new_n16729);
xnor_4 g14381(new_n16727, new_n11043, new_n16730);
not_8  g14382(new_n16699, new_n16731);
xnor_4 g14383(new_n16720, new_n16731, new_n16732);
nand_5 g14384(new_n16732, new_n11049, new_n16733_1);
xnor_4 g14385(new_n16732, new_n11048, new_n16734);
not_8  g14386(new_n16703, new_n16735);
xnor_4 g14387(new_n16718, new_n16735, new_n16736);
nand_5 g14388(new_n16736, new_n11057, new_n16737);
xnor_4 g14389(new_n16716, new_n16707, new_n16738);
not_8  g14390(new_n16738, new_n16739);
nand_5 g14391(new_n16739, new_n11060, new_n16740);
xnor_4 g14392(new_n16738, new_n11060, new_n16741);
xnor_4 g14393(new_n16713, new_n16712, new_n16742);
nand_5 g14394(new_n16742, new_n6128, new_n16743_1);
xnor_4 g14395(new_n16711, new_n4318, new_n16744);
not_8  g14396(new_n16744, new_n16745);
nor_5  g14397(new_n16745, new_n6114, new_n16746);
not_8  g14398(new_n16746, new_n16747);
xnor_4 g14399(new_n16742, new_n11065, new_n16748);
nand_5 g14400(new_n16748, new_n16747, new_n16749);
nand_5 g14401(new_n16749, new_n16743_1, new_n16750);
nand_5 g14402(new_n16750, new_n16741, new_n16751);
nand_5 g14403(new_n16751, new_n16740, new_n16752);
xnor_4 g14404(new_n16736, new_n11056_1, new_n16753);
nand_5 g14405(new_n16753, new_n16752, new_n16754);
nand_5 g14406(new_n16754, new_n16737, new_n16755);
nand_5 g14407(new_n16755, new_n16734, new_n16756);
nand_5 g14408(new_n16756, new_n16733_1, new_n16757);
nand_5 g14409(new_n16757, new_n16730, new_n16758);
nand_5 g14410(new_n16758, new_n16729, new_n16759);
xnor_4 g14411(new_n16759, new_n16726, n3528);
xnor_4 g14412(new_n9652, new_n9584, n3555);
nor_5  g14413(new_n2766, new_n2716, new_n16762);
nor_5  g14414(new_n2828, new_n2767, new_n16763);
nor_5  g14415(new_n16763, new_n16762, new_n16764);
not_8  g14416(new_n16764, new_n16765);
not_8  g14417(new_n2714, new_n16766);
nor_5  g14418(new_n16766, n13951, new_n16767);
nand_5 g14419(new_n10760, new_n16767, new_n16768);
not_8  g14420(new_n16768, new_n16769);
nand_5 g14421(new_n16769, new_n16765, new_n16770);
nor_5  g14422(new_n10760, new_n16767, new_n16771);
nand_5 g14423(new_n16771, new_n16764, new_n16772);
nand_5 g14424(new_n16772, new_n16770, new_n16773);
nand_5 g14425(new_n16773, new_n15580, new_n16774);
xnor_4 g14426(new_n16773, new_n15579, new_n16775);
not_8  g14427(new_n10760, new_n16776);
xnor_4 g14428(new_n16776, new_n16767, new_n16777);
xnor_4 g14429(new_n16777, new_n16765, new_n16778);
not_8  g14430(new_n16778, new_n16779);
nand_5 g14431(new_n16779, new_n15583, new_n16780);
xnor_4 g14432(new_n16778, new_n15583, new_n16781);
not_8  g14433(new_n2829, new_n16782);
nand_5 g14434(new_n16782, new_n2702, new_n16783);
nand_5 g14435(new_n2897, new_n2830, new_n16784);
nand_5 g14436(new_n16784, new_n16783, new_n16785);
nand_5 g14437(new_n16785, new_n16781, new_n16786);
nand_5 g14438(new_n16786, new_n16780, new_n16787);
nand_5 g14439(new_n16787, new_n16775, new_n16788);
nand_5 g14440(new_n16788, new_n16774, new_n16789);
nand_5 g14441(new_n16789, new_n16770, new_n16790);
not_8  g14442(new_n16790, n3561);
xnor_4 g14443(n16439, n14680, new_n16792);
not_8  g14444(new_n16792, new_n16793);
and_5  g14445(n17250, new_n4560, new_n16794);
nor_5  g14446(new_n11305, new_n11282, new_n16795);
nor_5  g14447(new_n16795, new_n16794, new_n16796);
xnor_4 g14448(new_n16796, new_n16793, new_n16797);
xnor_4 g14449(new_n10266, new_n7935, new_n16798_1);
nor_5  g14450(new_n10270, n13783, new_n16799);
not_8  g14451(new_n11307, new_n16800);
nor_5  g14452(new_n11327, new_n16800, new_n16801);
nor_5  g14453(new_n16801, new_n16799, new_n16802);
xnor_4 g14454(new_n16802, new_n16798_1, new_n16803);
xnor_4 g14455(new_n16803, new_n16797, new_n16804);
nor_5  g14456(new_n11328, new_n11306, new_n16805);
nor_5  g14457(new_n11361, new_n11329, new_n16806);
nor_5  g14458(new_n16806, new_n16805, new_n16807);
xnor_4 g14459(new_n16807, new_n16804, new_n16808);
xnor_4 g14460(new_n16808, new_n5919, new_n16809);
nor_5  g14461(new_n11362, new_n5924, new_n16810);
nor_5  g14462(new_n11391_1, new_n11363, new_n16811);
nor_5  g14463(new_n16811, new_n16810, new_n16812_1);
xor_4  g14464(new_n16812_1, new_n16809, n3563);
xnor_4 g14465(new_n6459, new_n6457_1, n3617);
xnor_4 g14466(n22253, n8305, new_n16815);
or_5   g14467(n12861, new_n13347, new_n16816);
xnor_4 g14468(n12861, n1255, new_n16817);
or_5   g14469(n13333, new_n13350, new_n16818_1);
xnor_4 g14470(n13333, n9512, new_n16819);
or_5   g14471(new_n7412, n2210, new_n16820);
nand_5 g14472(n21735, new_n5385, new_n16821);
nand_5 g14473(new_n4847, new_n4821, new_n16822);
nand_5 g14474(new_n16822, new_n16821, new_n16823);
xnor_4 g14475(n16608, n2210, new_n16824_1);
nand_5 g14476(new_n16824_1, new_n16823, new_n16825);
nand_5 g14477(new_n16825, new_n16820, new_n16826);
nand_5 g14478(new_n16826, new_n16819, new_n16827);
nand_5 g14479(new_n16827, new_n16818_1, new_n16828);
nand_5 g14480(new_n16828, new_n16817, new_n16829);
nand_5 g14481(new_n16829, new_n16816, new_n16830);
xnor_4 g14482(new_n16830, new_n16815, new_n16831);
xnor_4 g14483(new_n16831, new_n12055, new_n16832);
not_8  g14484(new_n16832, new_n16833);
xnor_4 g14485(new_n16828, new_n16817, new_n16834_1);
nand_5 g14486(new_n16834_1, new_n12061, new_n16835);
xnor_4 g14487(new_n16834_1, new_n12061, new_n16836);
not_8  g14488(new_n16836, new_n16837_1);
not_8  g14489(new_n16819, new_n16838);
xnor_4 g14490(new_n16826, new_n16838, new_n16839);
nor_5  g14491(new_n16839, new_n12065, new_n16840);
not_8  g14492(new_n16840, new_n16841_1);
xnor_4 g14493(new_n16824_1, new_n16823, new_n16842);
nor_5  g14494(new_n16842, new_n12069, new_n16843);
xnor_4 g14495(new_n16842, new_n12069, new_n16844);
nor_5  g14496(new_n4949, new_n4848, new_n16845);
nor_5  g14497(new_n4989, new_n4950, new_n16846);
nor_5  g14498(new_n16846, new_n16845, new_n16847);
nor_5  g14499(new_n16847, new_n16844, new_n16848);
nor_5  g14500(new_n16848, new_n16843, new_n16849);
xnor_4 g14501(new_n16839, new_n12066, new_n16850);
nand_5 g14502(new_n16850, new_n16849, new_n16851);
nand_5 g14503(new_n16851, new_n16841_1, new_n16852);
nand_5 g14504(new_n16852, new_n16837_1, new_n16853);
nand_5 g14505(new_n16853, new_n16835, new_n16854);
xnor_4 g14506(new_n16854, new_n16833, n3642);
not_8  g14507(n3324, new_n16856);
xnor_4 g14508(n16544, new_n3164_1, new_n16857);
nor_5  g14509(n23463, n6814, new_n16858);
xnor_4 g14510(n23463, new_n2941, new_n16859);
not_8  g14511(new_n16859, new_n16860);
nor_5  g14512(n19701, n13074, new_n16861);
xnor_4 g14513(n19701, new_n3171, new_n16862);
not_8  g14514(new_n16862, new_n16863);
nor_5  g14515(n23529, n10739, new_n16864);
xnor_4 g14516(n23529, new_n11911, new_n16865);
not_8  g14517(new_n16865, new_n16866);
nor_5  g14518(n24620, n21753, new_n16867);
xnor_4 g14519(n24620, new_n2350, new_n16868);
not_8  g14520(new_n16868, new_n16869);
nor_5  g14521(n21832, n5211, new_n16870);
not_8  g14522(new_n16238, new_n16871);
nor_5  g14523(new_n16246, new_n16871, new_n16872);
nor_5  g14524(new_n16872, new_n16870, new_n16873);
nor_5  g14525(new_n16873, new_n16869, new_n16874);
nor_5  g14526(new_n16874, new_n16867, new_n16875);
nor_5  g14527(new_n16875, new_n16866, new_n16876);
nor_5  g14528(new_n16876, new_n16864, new_n16877);
nor_5  g14529(new_n16877, new_n16863, new_n16878);
nor_5  g14530(new_n16878, new_n16861, new_n16879);
nor_5  g14531(new_n16879, new_n16860, new_n16880);
nor_5  g14532(new_n16880, new_n16858, new_n16881);
xnor_4 g14533(new_n16881, new_n16857, new_n16882);
xnor_4 g14534(new_n16882, new_n16856, new_n16883);
not_8  g14535(n17911, new_n16884);
xnor_4 g14536(new_n16879, new_n16859, new_n16885_1);
not_8  g14537(new_n16885_1, new_n16886);
nand_5 g14538(new_n16886, new_n16884, new_n16887);
xnor_4 g14539(new_n16885_1, new_n16884, new_n16888);
not_8  g14540(n21997, new_n16889);
xnor_4 g14541(new_n16877, new_n16862, new_n16890);
not_8  g14542(new_n16890, new_n16891);
nand_5 g14543(new_n16891, new_n16889, new_n16892);
xnor_4 g14544(new_n16890, new_n16889, new_n16893);
not_8  g14545(n25119, new_n16894);
xnor_4 g14546(new_n16875, new_n16865, new_n16895);
not_8  g14547(new_n16895, new_n16896);
nand_5 g14548(new_n16896, new_n16894, new_n16897);
xnor_4 g14549(new_n16895, new_n16894, new_n16898);
xnor_4 g14550(new_n16873, new_n16868, new_n16899);
not_8  g14551(new_n16899, new_n16900);
nor_5  g14552(new_n16900, new_n9035, new_n16901);
nor_5  g14553(new_n16247_1, n18537, new_n16902);
not_8  g14554(new_n16902, new_n16903);
not_8  g14555(new_n16262, new_n16904);
nand_5 g14556(new_n16904, new_n16248, new_n16905_1);
nand_5 g14557(new_n16905_1, new_n16903, new_n16906);
xnor_4 g14558(new_n16899, new_n9035, new_n16907);
not_8  g14559(new_n16907, new_n16908);
nor_5  g14560(new_n16908, new_n16906, new_n16909);
nor_5  g14561(new_n16909, new_n16901, new_n16910);
nand_5 g14562(new_n16910, new_n16898, new_n16911_1);
nand_5 g14563(new_n16911_1, new_n16897, new_n16912);
nand_5 g14564(new_n16912, new_n16893, new_n16913);
nand_5 g14565(new_n16913, new_n16892, new_n16914);
nand_5 g14566(new_n16914, new_n16888, new_n16915);
nand_5 g14567(new_n16915, new_n16887, new_n16916);
xnor_4 g14568(new_n16916, new_n16883, new_n16917);
not_8  g14569(new_n16917, new_n16918);
xnor_4 g14570(n23250, n16507, new_n16919);
not_8  g14571(n11455, new_n16920);
or_5   g14572(n22470, new_n16920, new_n16921);
xnor_4 g14573(n22470, n11455, new_n16922);
not_8  g14574(n3945, new_n16923);
or_5   g14575(n19116, new_n16923, new_n16924);
xnor_4 g14576(n19116, n3945, new_n16925);
not_8  g14577(n5255, new_n16926);
nor_5  g14578(n6861, new_n16926, new_n16927);
not_8  g14579(new_n16927, new_n16928);
xnor_4 g14580(n6861, n5255, new_n16929);
nor_5  g14581(new_n5428, n19357, new_n16930);
xnor_4 g14582(n21649, n19357, new_n16931);
not_8  g14583(new_n16931, new_n16932);
nor_5  g14584(new_n5432, n2328, new_n16933);
nand_5 g14585(n15053, new_n5436, new_n16934);
nand_5 g14586(new_n5335, new_n5331, new_n16935);
nand_5 g14587(new_n16935, new_n16934, new_n16936);
xnor_4 g14588(n18274, n2328, new_n16937);
not_8  g14589(new_n16937, new_n16938);
nor_5  g14590(new_n16938, new_n16936, new_n16939);
nor_5  g14591(new_n16939, new_n16933, new_n16940);
nor_5  g14592(new_n16940, new_n16932, new_n16941);
nor_5  g14593(new_n16941, new_n16930, new_n16942);
not_8  g14594(new_n16942, new_n16943);
nand_5 g14595(new_n16943, new_n16929, new_n16944);
nand_5 g14596(new_n16944, new_n16928, new_n16945);
nand_5 g14597(new_n16945, new_n16925, new_n16946);
nand_5 g14598(new_n16946, new_n16924, new_n16947);
nand_5 g14599(new_n16947, new_n16922, new_n16948);
nand_5 g14600(new_n16948, new_n16921, new_n16949);
xnor_4 g14601(new_n16949, new_n16919, new_n16950);
not_8  g14602(new_n16950, new_n16951_1);
nor_5  g14603(new_n16951_1, n4967, new_n16952);
not_8  g14604(n4967, new_n16953);
xnor_4 g14605(new_n16950, new_n16953, new_n16954_1);
xnor_4 g14606(new_n16947, new_n16922, new_n16955);
not_8  g14607(new_n16955, new_n16956);
nor_5  g14608(new_n16956, n15602, new_n16957);
xnor_4 g14609(new_n16945, new_n16925, new_n16958);
not_8  g14610(new_n16958, new_n16959);
nand_5 g14611(new_n16959, n8694, new_n16960);
xnor_4 g14612(new_n16942, new_n16929, new_n16961);
nor_5  g14613(new_n16961, n12380, new_n16962);
not_8  g14614(n12380, new_n16963);
xnor_4 g14615(new_n16961, new_n16963, new_n16964);
not_8  g14616(new_n16964, new_n16965);
xnor_4 g14617(new_n16940, new_n16931, new_n16966);
nor_5  g14618(new_n16966, n8943, new_n16967);
not_8  g14619(n8943, new_n16968_1);
xnor_4 g14620(new_n16966, new_n16968_1, new_n16969);
not_8  g14621(new_n16969, new_n16970);
not_8  g14622(n8255, new_n16971_1);
xnor_4 g14623(new_n16937, new_n16936, new_n16972);
not_8  g14624(new_n16972, new_n16973);
nor_5  g14625(new_n16973, new_n16971_1, new_n16974);
not_8  g14626(new_n16974, new_n16975);
not_8  g14627(n11184, new_n16976);
not_8  g14628(new_n5336, new_n16977);
nor_5  g14629(new_n16977, new_n16976, new_n16978);
not_8  g14630(new_n16978, new_n16979);
not_8  g14631(new_n5337_1, new_n16980);
nand_5 g14632(new_n16980, new_n5330_1, new_n16981);
nand_5 g14633(new_n16981, new_n16979, new_n16982);
xnor_4 g14634(new_n16972, n8255, new_n16983);
not_8  g14635(new_n16983, new_n16984);
nand_5 g14636(new_n16984, new_n16982, new_n16985);
nand_5 g14637(new_n16985, new_n16975, new_n16986);
nor_5  g14638(new_n16986, new_n16970, new_n16987);
nor_5  g14639(new_n16987, new_n16967, new_n16988_1);
nor_5  g14640(new_n16988_1, new_n16965, new_n16989_1);
nor_5  g14641(new_n16989_1, new_n16962, new_n16990);
xnor_4 g14642(new_n16958, n8694, new_n16991);
nand_5 g14643(new_n16991, new_n16990, new_n16992);
nand_5 g14644(new_n16992, new_n16960, new_n16993);
not_8  g14645(n15602, new_n16994_1);
xnor_4 g14646(new_n16955, new_n16994_1, new_n16995);
nor_5  g14647(new_n16995, new_n16993, new_n16996);
nor_5  g14648(new_n16996, new_n16957, new_n16997);
nor_5  g14649(new_n16997, new_n16954_1, new_n16998);
nor_5  g14650(new_n16998, new_n16952, new_n16999);
not_8  g14651(n13419, new_n17000);
xnor_4 g14652(n6659, n5101, new_n17001);
not_8  g14653(n23250, new_n17002);
or_5   g14654(new_n17002, n16507, new_n17003);
nand_5 g14655(new_n16949, new_n16919, new_n17004);
nand_5 g14656(new_n17004, new_n17003, new_n17005);
xnor_4 g14657(new_n17005, new_n17001, new_n17006_1);
xnor_4 g14658(new_n17006_1, new_n17000, new_n17007);
not_8  g14659(new_n17007, new_n17008);
xnor_4 g14660(new_n17008, new_n16999, new_n17009);
xnor_4 g14661(new_n17009, new_n16918, new_n17010);
xnor_4 g14662(new_n16914, new_n16888, new_n17011);
not_8  g14663(new_n17011, new_n17012);
not_8  g14664(new_n16954_1, new_n17013);
xnor_4 g14665(new_n16997, new_n17013, new_n17014);
nand_5 g14666(new_n17014, new_n17012, new_n17015);
xnor_4 g14667(new_n17014, new_n17011, new_n17016);
not_8  g14668(new_n16893, new_n17017);
xnor_4 g14669(new_n16912, new_n17017, new_n17018);
xnor_4 g14670(new_n16995, new_n16993, new_n17019);
not_8  g14671(new_n17019, new_n17020);
nand_5 g14672(new_n17020, new_n17018, new_n17021);
xnor_4 g14673(new_n17019, new_n17018, new_n17022);
xnor_4 g14674(new_n16910, new_n16898, new_n17023);
not_8  g14675(new_n17023, new_n17024);
xnor_4 g14676(new_n16991, new_n16990, new_n17025);
nand_5 g14677(new_n17025, new_n17024, new_n17026);
xnor_4 g14678(new_n17025, new_n17023, new_n17027);
xnor_4 g14679(new_n16988_1, new_n16964, new_n17028);
xnor_4 g14680(new_n16907, new_n16906, new_n17029);
not_8  g14681(new_n17029, new_n17030);
nand_5 g14682(new_n17030, new_n17028, new_n17031);
xnor_4 g14683(new_n17029, new_n17028, new_n17032);
xnor_4 g14684(new_n16986, new_n16969, new_n17033);
nand_5 g14685(new_n17033, new_n16264, new_n17034);
xnor_4 g14686(new_n17033, new_n16263, new_n17035_1);
not_8  g14687(new_n16284, new_n17036);
xnor_4 g14688(new_n16983, new_n16982, new_n17037_1);
nor_5  g14689(new_n17037_1, new_n17036, new_n17038);
not_8  g14690(new_n17038, new_n17039);
xnor_4 g14691(new_n17037_1, new_n16284, new_n17040);
nor_5  g14692(new_n5338, new_n16301, new_n17041);
not_8  g14693(new_n17041, new_n17042);
nand_5 g14694(new_n5354, new_n5339, new_n17043);
nand_5 g14695(new_n17043, new_n17042, new_n17044);
nand_5 g14696(new_n17044, new_n17040, new_n17045);
nand_5 g14697(new_n17045, new_n17039, new_n17046);
nand_5 g14698(new_n17046, new_n17035_1, new_n17047);
nand_5 g14699(new_n17047, new_n17034, new_n17048);
nand_5 g14700(new_n17048, new_n17032, new_n17049);
nand_5 g14701(new_n17049, new_n17031, new_n17050);
nand_5 g14702(new_n17050, new_n17027, new_n17051);
nand_5 g14703(new_n17051, new_n17026, new_n17052);
nand_5 g14704(new_n17052, new_n17022, new_n17053);
nand_5 g14705(new_n17053, new_n17021, new_n17054);
nand_5 g14706(new_n17054, new_n17016, new_n17055);
nand_5 g14707(new_n17055, new_n17015, new_n17056);
not_8  g14708(new_n17056, new_n17057);
xnor_4 g14709(new_n17057, new_n17010, n3649);
nor_5  g14710(n26625, n14230, new_n17059);
nand_5 g14711(new_n17059, new_n12285, new_n17060);
nor_5  g14712(new_n17060, n11566, new_n17061);
nand_5 g14713(new_n17061, new_n10121, new_n17062);
nor_5  g14714(new_n17062, n26565, new_n17063);
xnor_4 g14715(new_n17063, n3366, new_n17064);
xnor_4 g14716(new_n17064, n26191, new_n17065);
xnor_4 g14717(new_n17062, new_n11624, new_n17066);
nand_5 g14718(new_n17066, new_n12206, new_n17067);
xnor_4 g14719(new_n17066, n26512, new_n17068_1);
xnor_4 g14720(new_n17061, n3959, new_n17069_1);
nand_5 g14721(new_n17069_1, new_n12176, new_n17070_1);
xnor_4 g14722(new_n17069_1, n19575, new_n17071);
xnor_4 g14723(new_n17060, new_n12282, new_n17072);
nand_5 g14724(new_n17072, new_n10171, new_n17073);
xnor_4 g14725(new_n17072, n15378, new_n17074);
xnor_4 g14726(new_n17059, n26744, new_n17075_1);
nand_5 g14727(new_n17075_1, new_n10142, new_n17076);
not_8  g14728(new_n17076, new_n17077_1);
xnor_4 g14729(n26625, n14230, new_n17078);
nand_5 g14730(new_n17078, n22591, new_n17079);
nor_5  g14731(new_n10184, n14230, new_n17080);
xnor_4 g14732(new_n17078, new_n10183, new_n17081);
nand_5 g14733(new_n17081, new_n17080, new_n17082);
nand_5 g14734(new_n17082, new_n17079, new_n17083);
xnor_4 g14735(new_n17075_1, n17095, new_n17084_1);
not_8  g14736(new_n17084_1, new_n17085);
nor_5  g14737(new_n17085, new_n17083, new_n17086);
nor_5  g14738(new_n17086, new_n17077_1, new_n17087);
not_8  g14739(new_n17087, new_n17088);
nand_5 g14740(new_n17088, new_n17074, new_n17089);
nand_5 g14741(new_n17089, new_n17073, new_n17090_1);
nand_5 g14742(new_n17090_1, new_n17071, new_n17091);
nand_5 g14743(new_n17091, new_n17070_1, new_n17092);
nand_5 g14744(new_n17092, new_n17068_1, new_n17093);
nand_5 g14745(new_n17093, new_n17067, new_n17094);
xnor_4 g14746(new_n17094, new_n17065, new_n17095_1);
xnor_4 g14747(new_n17095_1, n7917, new_n17096);
not_8  g14748(new_n17096, new_n17097);
xnor_4 g14749(new_n17092, new_n17068_1, new_n17098);
nor_5  g14750(new_n17098, n17302, new_n17099);
xnor_4 g14751(new_n17098, n17302, new_n17100);
xnor_4 g14752(new_n17090_1, new_n17071, new_n17101);
nand_5 g14753(new_n17101, n2013, new_n17102);
xnor_4 g14754(new_n17101, new_n15387, new_n17103);
xnor_4 g14755(new_n17087, new_n17074, new_n17104_1);
nor_5  g14756(new_n17104_1, new_n15391, new_n17105);
not_8  g14757(new_n17105, new_n17106_1);
xnor_4 g14758(new_n17104_1, n23755, new_n17107);
xnor_4 g14759(new_n17084_1, new_n17083, new_n17108);
nor_5  g14760(new_n17108, new_n15393, new_n17109);
not_8  g14761(new_n17109, new_n17110);
xnor_4 g14762(new_n17108, n19163, new_n17111);
xnor_4 g14763(new_n17081, new_n17080, new_n17112);
nor_5  g14764(new_n17112, new_n15396, new_n17113);
nand_5 g14765(new_n17112, new_n15396, new_n17114);
xnor_4 g14766(n26167, n14230, new_n17115);
nand_5 g14767(new_n17115, n9646, new_n17116);
not_8  g14768(new_n17116, new_n17117);
nand_5 g14769(new_n17117, new_n17114, new_n17118);
not_8  g14770(new_n17118, new_n17119_1);
nor_5  g14771(new_n17119_1, new_n17113, new_n17120);
not_8  g14772(new_n17120, new_n17121);
nand_5 g14773(new_n17121, new_n17111, new_n17122);
nand_5 g14774(new_n17122, new_n17110, new_n17123);
nand_5 g14775(new_n17123, new_n17107, new_n17124);
nand_5 g14776(new_n17124, new_n17106_1, new_n17125);
nand_5 g14777(new_n17125, new_n17103, new_n17126);
nand_5 g14778(new_n17126, new_n17102, new_n17127);
nor_5  g14779(new_n17127, new_n17100, new_n17128);
nor_5  g14780(new_n17128, new_n17099, new_n17129);
xnor_4 g14781(new_n17129, new_n17097, new_n17130_1);
xnor_4 g14782(new_n17130_1, new_n7305_1, new_n17131);
xnor_4 g14783(new_n17127, new_n17100, new_n17132);
nand_5 g14784(new_n17132, new_n7310, new_n17133);
xnor_4 g14785(new_n17132, new_n7308_1, new_n17134);
not_8  g14786(new_n17125, new_n17135);
xnor_4 g14787(new_n17135, new_n17103, new_n17136);
nand_5 g14788(new_n17136, new_n7313_1, new_n17137);
xnor_4 g14789(new_n17136, new_n7312, new_n17138_1);
xnor_4 g14790(new_n17123, new_n17107, new_n17139);
not_8  g14791(new_n17139, new_n17140);
nand_5 g14792(new_n17140, new_n7319, new_n17141);
xnor_4 g14793(new_n17139, new_n7319, new_n17142);
xnor_4 g14794(new_n17120, new_n17111, new_n17143);
not_8  g14795(new_n17143, new_n17144);
nor_5  g14796(new_n17144, new_n7327, new_n17145);
not_8  g14797(new_n17145, new_n17146);
xnor_4 g14798(new_n17143, new_n7327, new_n17147);
xnor_4 g14799(new_n17112, n22358, new_n17148);
xnor_4 g14800(new_n17148, new_n17116, new_n17149);
nor_5  g14801(new_n17149, new_n7332, new_n17150);
xnor_4 g14802(new_n17115, n9646, new_n17151);
not_8  g14803(new_n17151, new_n17152);
nor_5  g14804(new_n17152, new_n7335_1, new_n17153);
not_8  g14805(new_n17153, new_n17154);
xnor_4 g14806(new_n17149, new_n7339_1, new_n17155);
not_8  g14807(new_n17155, new_n17156);
nor_5  g14808(new_n17156, new_n17154, new_n17157);
nor_5  g14809(new_n17157, new_n17150, new_n17158);
nand_5 g14810(new_n17158, new_n17147, new_n17159);
nand_5 g14811(new_n17159, new_n17146, new_n17160);
nand_5 g14812(new_n17160, new_n17142, new_n17161);
nand_5 g14813(new_n17161, new_n17141, new_n17162);
nand_5 g14814(new_n17162, new_n17138_1, new_n17163_1);
nand_5 g14815(new_n17163_1, new_n17137, new_n17164);
nand_5 g14816(new_n17164, new_n17134, new_n17165);
nand_5 g14817(new_n17165, new_n17133, new_n17166);
xnor_4 g14818(new_n17166, new_n17131, n3665);
xnor_4 g14819(new_n6117, new_n6116, n3679);
nor_5  g14820(n16521, n7139, new_n17169);
nand_5 g14821(new_n17169, new_n3696, new_n17170);
nor_5  g14822(new_n17170, n604, new_n17171);
nand_5 g14823(new_n17171, new_n3687, new_n17172);
nor_5  g14824(new_n17172, n9172, new_n17173);
nand_5 g14825(new_n17173, new_n3681, new_n17174);
nor_5  g14826(new_n17174, n13719, new_n17175);
xnor_4 g14827(new_n17175, n7026, new_n17176);
xnor_4 g14828(new_n17176, new_n6240, new_n17177);
xnor_4 g14829(new_n17174, new_n3678, new_n17178);
not_8  g14830(new_n17178, new_n17179);
nor_5  g14831(new_n17179, new_n6247, new_n17180);
xnor_4 g14832(new_n17178, new_n6246, new_n17181);
xnor_4 g14833(new_n17173, n442, new_n17182);
nor_5  g14834(new_n17182, new_n6252, new_n17183);
not_8  g14835(new_n17183, new_n17184);
xnor_4 g14836(new_n17182, new_n6253, new_n17185);
xnor_4 g14837(new_n17172, new_n3684, new_n17186);
nor_5  g14838(new_n17186, new_n6258, new_n17187);
not_8  g14839(new_n17187, new_n17188);
xnor_4 g14840(new_n17186, new_n6258, new_n17189);
not_8  g14841(new_n17189, new_n17190);
xnor_4 g14842(new_n17171, n4913, new_n17191);
nor_5  g14843(new_n17191, new_n6263, new_n17192);
not_8  g14844(new_n17192, new_n17193);
xnor_4 g14845(new_n17191, new_n6263, new_n17194);
not_8  g14846(new_n17194, new_n17195);
xnor_4 g14847(new_n17170, new_n3691, new_n17196);
nor_5  g14848(new_n17196, new_n6269, new_n17197);
xnor_4 g14849(new_n17196, new_n6269, new_n17198);
xnor_4 g14850(new_n17169, n16824, new_n17199);
nor_5  g14851(new_n17199, new_n6276_1, new_n17200);
xnor_4 g14852(new_n17199, new_n6276_1, new_n17201);
nand_5 g14853(new_n17169, new_n6282, new_n17202_1);
not_8  g14854(new_n17202_1, new_n17203);
nand_5 g14855(new_n6283, new_n3702, new_n17204);
xnor_4 g14856(new_n17204, new_n3700, new_n17205);
nor_5  g14857(new_n17205, new_n6453, new_n17206);
nor_5  g14858(new_n17206, new_n17203, new_n17207);
nor_5  g14859(new_n17207, new_n17201, new_n17208);
nor_5  g14860(new_n17208, new_n17200, new_n17209);
nor_5  g14861(new_n17209, new_n17198, new_n17210);
nor_5  g14862(new_n17210, new_n17197, new_n17211);
not_8  g14863(new_n17211, new_n17212);
nand_5 g14864(new_n17212, new_n17195, new_n17213);
nand_5 g14865(new_n17213, new_n17193, new_n17214);
nand_5 g14866(new_n17214, new_n17190, new_n17215);
nand_5 g14867(new_n17215, new_n17188, new_n17216);
nand_5 g14868(new_n17216, new_n17185, new_n17217);
nand_5 g14869(new_n17217, new_n17184, new_n17218);
nor_5  g14870(new_n17218, new_n17181, new_n17219_1);
nor_5  g14871(new_n17219_1, new_n17180, new_n17220);
xnor_4 g14872(new_n17220, new_n17177, new_n17221);
xnor_4 g14873(new_n6357, n2858, new_n17222);
nand_5 g14874(new_n6362, n2659, new_n17223);
xnor_4 g14875(new_n6361, n2659, new_n17224);
nand_5 g14876(new_n6366, n24327, new_n17225);
nand_5 g14877(new_n9031, new_n9006, new_n17226);
nand_5 g14878(new_n17226, new_n17225, new_n17227);
nand_5 g14879(new_n17227, new_n17224, new_n17228);
nand_5 g14880(new_n17228, new_n17223, new_n17229);
xnor_4 g14881(new_n17229, new_n17222, new_n17230);
not_8  g14882(new_n17230, new_n17231);
xnor_4 g14883(new_n17231, new_n17221, new_n17232_1);
xnor_4 g14884(new_n17227, new_n17224, new_n17233);
xnor_4 g14885(new_n17218, new_n17181, new_n17234);
nand_5 g14886(new_n17234, new_n17233, new_n17235);
not_8  g14887(new_n17233, new_n17236_1);
xnor_4 g14888(new_n17234, new_n17236_1, new_n17237);
xnor_4 g14889(new_n17216, new_n17185, new_n17238);
not_8  g14890(new_n17238, new_n17239);
nand_5 g14891(new_n17239, new_n9032_1, new_n17240);
xnor_4 g14892(new_n17238, new_n9032_1, new_n17241);
xnor_4 g14893(new_n17214, new_n17189, new_n17242);
nand_5 g14894(new_n17242, new_n9064, new_n17243_1);
xnor_4 g14895(new_n17242, new_n9065, new_n17244);
xnor_4 g14896(new_n17211, new_n17195, new_n17245);
nand_5 g14897(new_n17245, new_n9071, new_n17246);
not_8  g14898(new_n9071, new_n17247);
xnor_4 g14899(new_n17245, new_n17247, new_n17248);
not_8  g14900(new_n17198, new_n17249);
xnor_4 g14901(new_n17209, new_n17249, new_n17250_1);
not_8  g14902(new_n17250_1, new_n17251_1);
nor_5  g14903(new_n17251_1, new_n9078, new_n17252);
not_8  g14904(new_n17252, new_n17253);
xnor_4 g14905(new_n17250_1, new_n9078, new_n17254);
xnor_4 g14906(new_n17207, new_n17201, new_n17255);
not_8  g14907(new_n17255, new_n17256);
nor_5  g14908(new_n17256, new_n9082, new_n17257);
xnor_4 g14909(new_n17256, new_n9082, new_n17258);
xnor_4 g14910(new_n17205, new_n6286, new_n17259);
not_8  g14911(new_n17259, new_n17260);
nor_5  g14912(new_n17260, new_n9088, new_n17261);
not_8  g14913(new_n17261, new_n17262);
xnor_4 g14914(new_n6282, new_n3702, new_n17263_1);
nand_5 g14915(new_n17263_1, new_n9091, new_n17264);
xnor_4 g14916(new_n17259, new_n9088, new_n17265);
nand_5 g14917(new_n17265, new_n17264, new_n17266);
nand_5 g14918(new_n17266, new_n17262, new_n17267);
nor_5  g14919(new_n17267, new_n17258, new_n17268);
nor_5  g14920(new_n17268, new_n17257, new_n17269);
nand_5 g14921(new_n17269, new_n17254, new_n17270);
nand_5 g14922(new_n17270, new_n17253, new_n17271);
nand_5 g14923(new_n17271, new_n17248, new_n17272);
nand_5 g14924(new_n17272, new_n17246, new_n17273);
nand_5 g14925(new_n17273, new_n17244, new_n17274);
nand_5 g14926(new_n17274, new_n17243_1, new_n17275);
nand_5 g14927(new_n17275, new_n17241, new_n17276);
nand_5 g14928(new_n17276, new_n17240, new_n17277);
nand_5 g14929(new_n17277, new_n17237, new_n17278);
nand_5 g14930(new_n17278, new_n17235, new_n17279);
xnor_4 g14931(new_n17279, new_n17232_1, n3725);
not_8  g14932(new_n15744, new_n17281);
or_5   g14933(n11220, n3425, new_n17282);
nand_5 g14934(new_n13855, new_n13852, new_n17283);
nand_5 g14935(new_n17283, new_n17282, new_n17284);
or_5   g14936(n7335, n2160, new_n17285_1);
nand_5 g14937(new_n13850_1, new_n13847, new_n17286);
nand_5 g14938(new_n17286, new_n17285_1, new_n17287);
xnor_4 g14939(new_n17287, new_n17284, new_n17288);
not_8  g14940(new_n13851_1, new_n17289);
nor_5  g14941(new_n13856, new_n17289, new_n17290);
not_8  g14942(new_n17290, new_n17291);
nand_5 g14943(new_n13861, new_n13857, new_n17292);
nand_5 g14944(new_n17292, new_n17291, new_n17293);
xnor_4 g14945(new_n17293, new_n17288, new_n17294);
xnor_4 g14946(new_n17294, new_n17281, new_n17295);
nand_5 g14947(new_n15747, new_n13862, new_n17296);
xnor_4 g14948(new_n15747, new_n13863, new_n17297);
not_8  g14949(new_n5675, new_n17298);
nor_5  g14950(new_n15752, new_n17298, new_n17299);
xnor_4 g14951(new_n15753, new_n5675, new_n17300);
not_8  g14952(new_n15757, new_n17301);
nor_5  g14953(new_n17301, new_n5678, new_n17302_1);
nor_5  g14954(new_n15761_1, new_n5683, new_n17303);
not_8  g14955(new_n17303, new_n17304);
xnor_4 g14956(new_n15760, new_n5683, new_n17305);
nor_5  g14957(new_n15764, new_n5687_1, new_n17306);
not_8  g14958(new_n17306, new_n17307);
xnor_4 g14959(new_n15673, new_n5687_1, new_n17308);
nor_5  g14960(new_n5693, new_n15675, new_n17309);
not_8  g14961(new_n17309, new_n17310);
nor_5  g14962(new_n5697, new_n4442, new_n17311);
xnor_4 g14963(new_n5697, new_n4442, new_n17312);
nor_5  g14964(new_n5706, new_n4446, new_n17313);
xnor_4 g14965(new_n5706, new_n4446, new_n17314);
nor_5  g14966(new_n5712, new_n4449, new_n17315);
nor_5  g14967(new_n5710, new_n4430, new_n17316);
nor_5  g14968(new_n5717, new_n4454, new_n17317);
not_8  g14969(new_n17317, new_n17318);
nor_5  g14970(new_n17318, new_n17316, new_n17319);
nor_5  g14971(new_n17319, new_n17315, new_n17320_1);
nor_5  g14972(new_n17320_1, new_n17314, new_n17321);
nor_5  g14973(new_n17321, new_n17313, new_n17322);
nor_5  g14974(new_n17322, new_n17312, new_n17323);
nor_5  g14975(new_n17323, new_n17311, new_n17324);
xnor_4 g14976(new_n5692, new_n15675, new_n17325);
nand_5 g14977(new_n17325, new_n17324, new_n17326);
nand_5 g14978(new_n17326, new_n17310, new_n17327);
nand_5 g14979(new_n17327, new_n17308, new_n17328);
nand_5 g14980(new_n17328, new_n17307, new_n17329);
nand_5 g14981(new_n17329, new_n17305, new_n17330);
nand_5 g14982(new_n17330, new_n17304, new_n17331);
xnor_4 g14983(new_n17301, new_n5678, new_n17332);
nor_5  g14984(new_n17332, new_n17331, new_n17333);
nor_5  g14985(new_n17333, new_n17302_1, new_n17334);
nor_5  g14986(new_n17334, new_n17300, new_n17335);
nor_5  g14987(new_n17335, new_n17299, new_n17336);
nand_5 g14988(new_n17336, new_n17297, new_n17337_1);
nand_5 g14989(new_n17337_1, new_n17296, new_n17338);
xnor_4 g14990(new_n17338, new_n17295, n3733);
not_8  g14991(new_n11437, new_n17340);
xnor_4 g14992(new_n17340, n24937, new_n17341);
not_8  g14993(new_n17341, new_n17342);
not_8  g14994(new_n11429, new_n17343);
nand_5 g14995(new_n17343, n5098, new_n17344_1);
xnor_4 g14996(new_n11429, n5098, new_n17345);
not_8  g14997(n3030, new_n17346);
nor_5  g14998(new_n11421, new_n17346, new_n17347);
not_8  g14999(new_n16308, new_n17348);
nor_5  g15000(new_n16323, new_n17348, new_n17349);
nor_5  g15001(new_n17349, new_n17347, new_n17350);
not_8  g15002(new_n17350, new_n17351_1);
nand_5 g15003(new_n17351_1, new_n17345, new_n17352);
nand_5 g15004(new_n17352, new_n17344_1, new_n17353);
xnor_4 g15005(new_n17353, new_n17342, new_n17354);
xnor_4 g15006(new_n17354, new_n10638, new_n17355);
xnor_4 g15007(new_n17350, new_n17345, new_n17356);
not_8  g15008(new_n17356, new_n17357);
nand_5 g15009(new_n17357, new_n10643, new_n17358);
xnor_4 g15010(new_n17356, new_n10643, new_n17359_1);
not_8  g15011(new_n16324, new_n17360);
nand_5 g15012(new_n17360, new_n10648, new_n17361);
nand_5 g15013(new_n16339, new_n16325, new_n17362);
nand_5 g15014(new_n17362, new_n17361, new_n17363);
nand_5 g15015(new_n17363, new_n17359_1, new_n17364);
nand_5 g15016(new_n17364, new_n17358, new_n17365);
xor_4  g15017(new_n17365, new_n17355, n3755);
xnor_4 g15018(new_n9644, new_n9605, n3758);
not_8  g15019(n2570, new_n17368);
not_8  g15020(n19033, new_n17369);
not_8  g15021(n18145, new_n17370);
nand_5 g15022(new_n16655, new_n17370, new_n17371);
nor_5  g15023(new_n17371, n655, new_n17372);
nand_5 g15024(new_n17372, new_n17369, new_n17373);
xnor_4 g15025(new_n17373, new_n17368, new_n17374);
xnor_4 g15026(new_n17374, n14692, new_n17375);
xnor_4 g15027(new_n17372, n19033, new_n17376);
not_8  g15028(new_n17376, new_n17377);
nand_5 g15029(new_n17377, n4100, new_n17378);
xnor_4 g15030(new_n17376, n4100, new_n17379);
not_8  g15031(n655, new_n17380);
xnor_4 g15032(new_n17371, new_n17380, new_n17381);
not_8  g15033(new_n17381, new_n17382);
nand_5 g15034(new_n17382, n21957, new_n17383);
xnor_4 g15035(new_n17381, n21957, new_n17384);
not_8  g15036(new_n16656_1, new_n17385);
nand_5 g15037(new_n17385, n15761, new_n17386);
nand_5 g15038(new_n16689, new_n16657, new_n17387_1);
nand_5 g15039(new_n17387_1, new_n17386, new_n17388);
nand_5 g15040(new_n17388, new_n17384, new_n17389);
nand_5 g15041(new_n17389, new_n17383, new_n17390);
nand_5 g15042(new_n17390, new_n17379, new_n17391_1);
nand_5 g15043(new_n17391_1, new_n17378, new_n17392_1);
xnor_4 g15044(new_n17392_1, new_n17375, new_n17393);
not_8  g15045(new_n17393, new_n17394);
nand_5 g15046(new_n17394, new_n12702_1, new_n17395);
xnor_4 g15047(new_n17393, new_n12702_1, new_n17396);
xnor_4 g15048(new_n17390, new_n17379, new_n17397);
not_8  g15049(new_n17397, new_n17398);
nand_5 g15050(new_n17398, new_n7250, new_n17399);
xnor_4 g15051(new_n17397, new_n7250, new_n17400);
xnor_4 g15052(new_n17388, new_n17384, new_n17401);
not_8  g15053(new_n17401, new_n17402);
nand_5 g15054(new_n17402, new_n7252, new_n17403);
xnor_4 g15055(new_n17401, new_n7252, new_n17404);
not_8  g15056(new_n16690, new_n17405);
nand_5 g15057(new_n17405, new_n7256_1, new_n17406);
nand_5 g15058(new_n16724, new_n16691, new_n17407);
nand_5 g15059(new_n17407, new_n17406, new_n17408);
nand_5 g15060(new_n17408, new_n17404, new_n17409);
nand_5 g15061(new_n17409, new_n17403, new_n17410);
nand_5 g15062(new_n17410, new_n17400, new_n17411);
nand_5 g15063(new_n17411, new_n17399, new_n17412);
nand_5 g15064(new_n17412, new_n17396, new_n17413);
nand_5 g15065(new_n17413, new_n17395, new_n17414);
nor_5  g15066(new_n17373, n2570, new_n17415);
or_5   g15067(new_n17374, new_n10896, new_n17416);
nand_5 g15068(new_n17392_1, new_n17375, new_n17417);
nand_5 g15069(new_n17417, new_n17416, new_n17418);
xnor_4 g15070(new_n17418, new_n17415, new_n17419);
xnor_4 g15071(new_n17419, new_n12757, new_n17420);
xnor_4 g15072(new_n17420, new_n17414, new_n17421_1);
not_8  g15073(new_n17421_1, new_n17422);
nand_5 g15074(new_n17422, new_n11016, new_n17423);
xnor_4 g15075(new_n17421_1, new_n11016, new_n17424);
xnor_4 g15076(new_n17412, new_n17396, new_n17425);
not_8  g15077(new_n17425, new_n17426);
nand_5 g15078(new_n17426, new_n11022, new_n17427);
xnor_4 g15079(new_n17425, new_n11022, new_n17428);
xnor_4 g15080(new_n17410, new_n17400, new_n17429);
not_8  g15081(new_n17429, new_n17430);
nand_5 g15082(new_n17430, new_n11027, new_n17431);
xnor_4 g15083(new_n17429, new_n11027, new_n17432_1);
xnor_4 g15084(new_n17408, new_n17404, new_n17433);
not_8  g15085(new_n17433, new_n17434);
nand_5 g15086(new_n17434, new_n11032, new_n17435);
xnor_4 g15087(new_n17433, new_n11032, new_n17436_1);
not_8  g15088(new_n16725, new_n17437);
nor_5  g15089(new_n17437, new_n11038, new_n17438);
not_8  g15090(new_n16726, new_n17439);
nor_5  g15091(new_n16759, new_n17439, new_n17440_1);
nor_5  g15092(new_n17440_1, new_n17438, new_n17441);
nand_5 g15093(new_n17441, new_n17436_1, new_n17442);
nand_5 g15094(new_n17442, new_n17435, new_n17443);
nand_5 g15095(new_n17443, new_n17432_1, new_n17444);
nand_5 g15096(new_n17444, new_n17431, new_n17445);
nand_5 g15097(new_n17445, new_n17428, new_n17446);
nand_5 g15098(new_n17446, new_n17427, new_n17447);
nand_5 g15099(new_n17447, new_n17424, new_n17448);
nand_5 g15100(new_n17448, new_n17423, new_n17449);
not_8  g15101(new_n17419, new_n17450_1);
nor_5  g15102(new_n17450_1, new_n12757, new_n17451);
not_8  g15103(new_n17418, new_n17452);
nand_5 g15104(new_n17452, new_n17415, new_n17453);
not_8  g15105(new_n17414, new_n17454);
nand_5 g15106(new_n17450_1, new_n12757, new_n17455);
nand_5 g15107(new_n17455, new_n17454, new_n17456);
nand_5 g15108(new_n17456, new_n17453, new_n17457);
nor_5  g15109(new_n17457, new_n17451, new_n17458_1);
xnor_4 g15110(new_n17458_1, new_n17449, n3760);
xnor_4 g15111(new_n4089_1, new_n4064, n3781);
xnor_4 g15112(new_n14412_1, new_n14385, n3794);
not_8  g15113(new_n11574, new_n17462);
nor_5  g15114(new_n17462, new_n5267, new_n17463);
nor_5  g15115(new_n17463, new_n5273_1, new_n17464);
nand_5 g15116(new_n17463, new_n5020_1, new_n17465);
not_8  g15117(new_n17465, new_n17466_1);
nor_5  g15118(new_n17466_1, new_n17464, new_n17467);
nor_5  g15119(new_n13900, new_n6283, new_n17468);
not_8  g15120(new_n17468, new_n17469);
nor_5  g15121(new_n6283, new_n6218_1, new_n17470);
nor_5  g15122(new_n6286, new_n6282, new_n17471);
nor_5  g15123(new_n17471, new_n17470, new_n17472);
xnor_4 g15124(new_n17472, new_n13903, new_n17473);
xnor_4 g15125(new_n17473, new_n17469, new_n17474);
xor_4  g15126(new_n17474, new_n17467, n3842);
xnor_4 g15127(new_n13038, new_n9461, n3850);
xnor_4 g15128(new_n15698, new_n4481, n3869);
not_8  g15129(n19584, new_n17478);
xnor_4 g15130(n21749, new_n4327, new_n17479);
nor_5  g15131(n25316, n7769, new_n17480);
nand_5 g15132(n21138, n20385, new_n17481);
xnor_4 g15133(n25316, new_n10133, new_n17482);
nand_5 g15134(new_n17482, new_n17481, new_n17483);
not_8  g15135(new_n17483, new_n17484);
nor_5  g15136(new_n17484, new_n17480, new_n17485);
xnor_4 g15137(new_n17485, new_n17479, new_n17486);
xnor_4 g15138(new_n17486, new_n17478, new_n17487);
not_8  g15139(n5060, new_n17488);
xnor_4 g15140(n21138, n20385, new_n17489);
nand_5 g15141(new_n17489, n15332, new_n17490);
nand_5 g15142(new_n17490, new_n17488, new_n17491);
not_8  g15143(new_n17491, new_n17492);
not_8  g15144(new_n17481, new_n17493_1);
xnor_4 g15145(new_n17482, new_n17493_1, new_n17494);
xnor_4 g15146(new_n17490, new_n17488, new_n17495);
nor_5  g15147(new_n17495, new_n17494, new_n17496);
nor_5  g15148(new_n17496, new_n17492, new_n17497);
xnor_4 g15149(new_n17497, new_n17487, new_n17498);
xnor_4 g15150(new_n17498, new_n16587, new_n17499);
xnor_4 g15151(new_n17495, new_n17494, new_n17500_1);
nand_5 g15152(new_n17500_1, new_n16590, new_n17501);
not_8  g15153(n15332, new_n17502);
xnor_4 g15154(new_n17489, new_n17502, new_n17503);
nor_5  g15155(new_n17503, new_n16595, new_n17504);
not_8  g15156(new_n17504, new_n17505);
xnor_4 g15157(new_n17500_1, new_n16589_1, new_n17506);
nand_5 g15158(new_n17506, new_n17505, new_n17507);
nand_5 g15159(new_n17507, new_n17501, new_n17508);
xnor_4 g15160(new_n17508, new_n17499, n3871);
xor_4  g15161(new_n17267, new_n17258, n3891);
xnor_4 g15162(n10250, n2570, new_n17511);
or_5   g15163(n19033, new_n6481, new_n17512);
xnor_4 g15164(n19033, n7674, new_n17513);
or_5   g15165(new_n6484, n655, new_n17514);
xnor_4 g15166(n6397, n655, new_n17515);
or_5   g15167(new_n6487, n18145, new_n17516);
xnor_4 g15168(n19196, n18145, new_n17517);
or_5   g15169(new_n12714, n10712, new_n17518);
xnor_4 g15170(n23586, n10712, new_n17519);
nor_5  g15171(n25126, new_n16517_1, new_n17520);
xnor_4 g15172(n25126, n21226, new_n17521);
not_8  g15173(new_n17521, new_n17522);
nor_5  g15174(n19608, new_n6497, new_n17523);
nor_5  g15175(n20036, new_n4301, new_n17524_1);
nor_5  g15176(new_n4310, new_n4302, new_n17525);
nor_5  g15177(new_n17525, new_n17524_1, new_n17526);
xnor_4 g15178(n19608, n4426, new_n17527);
nand_5 g15179(new_n17527, new_n17526, new_n17528);
not_8  g15180(new_n17528, new_n17529_1);
nor_5  g15181(new_n17529_1, new_n17523, new_n17530);
nor_5  g15182(new_n17530, new_n17522, new_n17531);
nor_5  g15183(new_n17531, new_n17520, new_n17532);
not_8  g15184(new_n17532, new_n17533);
nand_5 g15185(new_n17533, new_n17519, new_n17534);
nand_5 g15186(new_n17534, new_n17518, new_n17535);
nand_5 g15187(new_n17535, new_n17517, new_n17536);
nand_5 g15188(new_n17536, new_n17516, new_n17537);
nand_5 g15189(new_n17537, new_n17515, new_n17538);
nand_5 g15190(new_n17538, new_n17514, new_n17539);
nand_5 g15191(new_n17539, new_n17513, new_n17540);
nand_5 g15192(new_n17540, new_n17512, new_n17541);
xnor_4 g15193(new_n17541, new_n17511, new_n17542);
xnor_4 g15194(new_n17542, new_n12703, new_n17543);
xnor_4 g15195(new_n17539, new_n17513, new_n17544);
nand_5 g15196(new_n17544, new_n7250, new_n17545);
xnor_4 g15197(new_n17544, new_n12706, new_n17546);
xnor_4 g15198(new_n17537, new_n17515, new_n17547);
nand_5 g15199(new_n17547, new_n7252, new_n17548);
xnor_4 g15200(new_n17547, new_n7253_1, new_n17549);
xnor_4 g15201(new_n17535, new_n17517, new_n17550);
nand_5 g15202(new_n17550, new_n7256_1, new_n17551);
xnor_4 g15203(new_n17550, new_n7256_1, new_n17552);
not_8  g15204(new_n17552, new_n17553);
xnor_4 g15205(new_n17533, new_n17519, new_n17554);
nand_5 g15206(new_n17554, new_n7260, new_n17555);
xnor_4 g15207(new_n17554, new_n7260, new_n17556);
not_8  g15208(new_n17556, new_n17557_1);
xnor_4 g15209(new_n17530, new_n17521, new_n17558);
not_8  g15210(new_n17558, new_n17559);
nand_5 g15211(new_n17559, new_n7264, new_n17560);
xnor_4 g15212(new_n17558, new_n7264, new_n17561);
xnor_4 g15213(new_n17527, new_n17526, new_n17562);
nand_5 g15214(new_n17562, new_n12719, new_n17563);
xnor_4 g15215(new_n17562, new_n7270, new_n17564);
nor_5  g15216(new_n4311, new_n12722, new_n17565);
not_8  g15217(new_n17565, new_n17566);
nand_5 g15218(new_n4324, new_n4312, new_n17567);
nand_5 g15219(new_n17567, new_n17566, new_n17568);
nand_5 g15220(new_n17568, new_n17564, new_n17569);
nand_5 g15221(new_n17569, new_n17563, new_n17570);
nand_5 g15222(new_n17570, new_n17561, new_n17571);
nand_5 g15223(new_n17571, new_n17560, new_n17572);
nand_5 g15224(new_n17572, new_n17557_1, new_n17573);
nand_5 g15225(new_n17573, new_n17555, new_n17574);
nand_5 g15226(new_n17574, new_n17553, new_n17575);
nand_5 g15227(new_n17575, new_n17551, new_n17576);
nand_5 g15228(new_n17576, new_n17549, new_n17577);
nand_5 g15229(new_n17577, new_n17548, new_n17578);
nand_5 g15230(new_n17578, new_n17546, new_n17579);
nand_5 g15231(new_n17579, new_n17545, new_n17580);
xnor_4 g15232(new_n17580, new_n17543, new_n17581);
xnor_4 g15233(new_n17581, new_n6688, new_n17582);
not_8  g15234(new_n17546, new_n17583_1);
xnor_4 g15235(new_n17578, new_n17583_1, new_n17584);
nand_5 g15236(new_n17584, new_n6697, new_n17585);
xnor_4 g15237(new_n17584, new_n6696, new_n17586);
not_8  g15238(new_n17549, new_n17587);
xnor_4 g15239(new_n17576, new_n17587, new_n17588);
nand_5 g15240(new_n17588, new_n6703, new_n17589);
xnor_4 g15241(new_n17588, new_n6702, new_n17590);
xnor_4 g15242(new_n17574, new_n17552, new_n17591);
nand_5 g15243(new_n17591, new_n6707_1, new_n17592_1);
xnor_4 g15244(new_n17591, new_n6706_1, new_n17593);
xnor_4 g15245(new_n17572, new_n17556, new_n17594);
nand_5 g15246(new_n17594, new_n6714, new_n17595);
xnor_4 g15247(new_n17594, new_n6713, new_n17596);
xnor_4 g15248(new_n17570, new_n17561, new_n17597);
not_8  g15249(new_n17597, new_n17598);
nand_5 g15250(new_n17598, new_n6719, new_n17599);
xnor_4 g15251(new_n17597, new_n6719, new_n17600);
xnor_4 g15252(new_n17568, new_n17564, new_n17601);
nor_5  g15253(new_n17601, new_n6724, new_n17602);
xnor_4 g15254(new_n17601, new_n6727, new_n17603);
not_8  g15255(new_n17603, new_n17604);
nor_5  g15256(new_n4334, new_n4325_1, new_n17605);
nor_5  g15257(new_n4351, new_n4336, new_n17606);
nor_5  g15258(new_n17606, new_n17605, new_n17607);
nor_5  g15259(new_n17607, new_n17604, new_n17608);
nor_5  g15260(new_n17608, new_n17602, new_n17609);
not_8  g15261(new_n17609, new_n17610);
nand_5 g15262(new_n17610, new_n17600, new_n17611);
nand_5 g15263(new_n17611, new_n17599, new_n17612);
nand_5 g15264(new_n17612, new_n17596, new_n17613);
nand_5 g15265(new_n17613, new_n17595, new_n17614);
nand_5 g15266(new_n17614, new_n17593, new_n17615);
nand_5 g15267(new_n17615, new_n17592_1, new_n17616);
nand_5 g15268(new_n17616, new_n17590, new_n17617);
nand_5 g15269(new_n17617, new_n17589, new_n17618);
nand_5 g15270(new_n17618, new_n17586, new_n17619);
nand_5 g15271(new_n17619, new_n17585, new_n17620);
xnor_4 g15272(new_n17620, new_n17582, n3932);
xnor_4 g15273(new_n4083, new_n4082, n3934);
xnor_4 g15274(new_n4283, new_n4282, n3971);
nor_5  g15275(n8581, n5026, new_n17624);
nand_5 g15276(new_n17624, new_n6982, new_n17625);
nor_5  g15277(new_n17625, n18157, new_n17626);
nand_5 g15278(new_n17626, new_n11178, new_n17627);
nor_5  g15279(new_n17627, n8067, new_n17628);
nand_5 g15280(new_n17628, new_n7647_1, new_n17629);
nor_5  g15281(new_n17629, n25240, new_n17630);
xnor_4 g15282(new_n17630, n1222, new_n17631);
xnor_4 g15283(new_n17631, new_n9341, new_n17632);
xnor_4 g15284(new_n17629, new_n11681, new_n17633);
not_8  g15285(new_n17633, new_n17634);
nand_5 g15286(new_n17634, new_n9349, new_n17635);
xnor_4 g15287(new_n17633, new_n9349, new_n17636);
xnor_4 g15288(new_n17628, n10125, new_n17637);
and_5  g15289(new_n17637, n26318, new_n17638_1);
nor_5  g15290(new_n17637, n26318, new_n17639);
xnor_4 g15291(new_n17627, new_n7650, new_n17640);
not_8  g15292(new_n17640, new_n17641);
nand_5 g15293(new_n17641, new_n9296, new_n17642);
xnor_4 g15294(new_n17640, new_n9296, new_n17643);
xnor_4 g15295(new_n17626, n20923, new_n17644);
not_8  g15296(new_n17644, new_n17645);
nand_5 g15297(new_n17645, new_n9301, new_n17646);
xnor_4 g15298(new_n17644, new_n9301, new_n17647);
xnor_4 g15299(new_n17625, new_n11691, new_n17648);
not_8  g15300(new_n17648, new_n17649);
nand_5 g15301(new_n17649, new_n9306, new_n17650);
xnor_4 g15302(new_n17624, n12161, new_n17651);
not_8  g15303(new_n17651, new_n17652);
nand_5 g15304(new_n17652, new_n9310, new_n17653);
xnor_4 g15305(new_n17651, new_n9310, new_n17654);
xnor_4 g15306(n8581, n5026, new_n17655);
nand_5 g15307(new_n17655, new_n9315, new_n17656);
nand_5 g15308(n13714, n8581, new_n17657);
xnor_4 g15309(new_n17655, n12593, new_n17658);
nand_5 g15310(new_n17658, new_n17657, new_n17659);
nand_5 g15311(new_n17659, new_n17656, new_n17660);
nand_5 g15312(new_n17660, new_n17654, new_n17661);
nand_5 g15313(new_n17661, new_n17653, new_n17662);
xnor_4 g15314(new_n17648, new_n9306, new_n17663);
nand_5 g15315(new_n17663, new_n17662, new_n17664_1);
nand_5 g15316(new_n17664_1, new_n17650, new_n17665);
nand_5 g15317(new_n17665, new_n17647, new_n17666);
nand_5 g15318(new_n17666, new_n17646, new_n17667);
nand_5 g15319(new_n17667, new_n17643, new_n17668);
nand_5 g15320(new_n17668, new_n17642, new_n17669);
nor_5  g15321(new_n17669, new_n17639, new_n17670);
nor_5  g15322(new_n17670, new_n17638_1, new_n17671);
nand_5 g15323(new_n17671, new_n17636, new_n17672);
nand_5 g15324(new_n17672, new_n17635, new_n17673);
xnor_4 g15325(new_n17673, new_n17632, new_n17674);
xnor_4 g15326(new_n17674, new_n5906, new_n17675);
xnor_4 g15327(new_n17671, new_n17636, new_n17676);
nand_5 g15328(new_n17676, n23913, new_n17677);
xnor_4 g15329(new_n17676, new_n5851, new_n17678);
xnor_4 g15330(new_n17637, new_n9291, new_n17679);
xnor_4 g15331(new_n17679, new_n17669, new_n17680);
nand_5 g15332(new_n17680, n22554, new_n17681);
xnor_4 g15333(new_n17680, new_n5836, new_n17682);
xnor_4 g15334(new_n17667, new_n17643, new_n17683);
nand_5 g15335(new_n17683, n20429, new_n17684);
xnor_4 g15336(new_n17683, new_n5862, new_n17685);
xnor_4 g15337(new_n17665, new_n17647, new_n17686);
nand_5 g15338(new_n17686, n3909, new_n17687_1);
xnor_4 g15339(new_n17686, new_n5837, new_n17688);
xnor_4 g15340(new_n17663, new_n17662, new_n17689);
nand_5 g15341(new_n17689, n23974, new_n17690);
xnor_4 g15342(new_n17689, new_n5873, new_n17691);
xnor_4 g15343(new_n17660, new_n17654, new_n17692);
nand_5 g15344(new_n17692, n2146, new_n17693);
xnor_4 g15345(new_n17692, new_n5838, new_n17694);
xnor_4 g15346(new_n17658, new_n17657, new_n17695);
nand_5 g15347(new_n17695, n22173, new_n17696);
xnor_4 g15348(n13714, new_n7664, new_n17697);
not_8  g15349(new_n17697, new_n17698);
nor_5  g15350(new_n17698, new_n5961, new_n17699);
xnor_4 g15351(new_n17695, new_n8553, new_n17700);
nand_5 g15352(new_n17700, new_n17699, new_n17701);
nand_5 g15353(new_n17701, new_n17696, new_n17702);
nand_5 g15354(new_n17702, new_n17694, new_n17703);
nand_5 g15355(new_n17703, new_n17693, new_n17704);
nand_5 g15356(new_n17704, new_n17691, new_n17705);
nand_5 g15357(new_n17705, new_n17690, new_n17706);
nand_5 g15358(new_n17706, new_n17688, new_n17707);
nand_5 g15359(new_n17707, new_n17687_1, new_n17708);
nand_5 g15360(new_n17708, new_n17685, new_n17709);
nand_5 g15361(new_n17709, new_n17684, new_n17710);
nand_5 g15362(new_n17710, new_n17682, new_n17711);
nand_5 g15363(new_n17711, new_n17681, new_n17712);
nand_5 g15364(new_n17712, new_n17678, new_n17713);
nand_5 g15365(new_n17713, new_n17677, new_n17714);
xnor_4 g15366(new_n17714, new_n17675, new_n17715);
xnor_4 g15367(new_n17715, new_n8647, new_n17716);
not_8  g15368(new_n17678, new_n17717);
xnor_4 g15369(new_n17712, new_n17717, new_n17718);
not_8  g15370(new_n17718, new_n17719);
nand_5 g15371(new_n17719, new_n8654, new_n17720);
xnor_4 g15372(new_n17718, new_n8654, new_n17721_1);
xnor_4 g15373(new_n17710, new_n17682, new_n17722);
nand_5 g15374(new_n17722, new_n8660, new_n17723);
xnor_4 g15375(new_n17722, new_n8659, new_n17724);
xnor_4 g15376(new_n17708, new_n17685, new_n17725);
nand_5 g15377(new_n17725, new_n8666, new_n17726);
xnor_4 g15378(new_n17725, new_n8665, new_n17727);
not_8  g15379(new_n17688, new_n17728);
xnor_4 g15380(new_n17706, new_n17728, new_n17729);
not_8  g15381(new_n17729, new_n17730);
nand_5 g15382(new_n17730, new_n8672, new_n17731);
xnor_4 g15383(new_n17729, new_n8672, new_n17732);
xnor_4 g15384(new_n17704, new_n17691, new_n17733);
nand_5 g15385(new_n17733, new_n8681, new_n17734);
xnor_4 g15386(new_n17733, new_n8677, new_n17735_1);
not_8  g15387(new_n17694, new_n17736);
xnor_4 g15388(new_n17702, new_n17736, new_n17737);
not_8  g15389(new_n17737, new_n17738_1);
nand_5 g15390(new_n17738_1, new_n8688, new_n17739);
xnor_4 g15391(new_n17700, new_n17699, new_n17740);
nand_5 g15392(new_n17740, new_n8691, new_n17741);
xnor_4 g15393(new_n17697, new_n5961, new_n17742);
nand_5 g15394(new_n17742, new_n8693, new_n17743);
not_8  g15395(new_n8691, new_n17744);
xnor_4 g15396(new_n17740, new_n17744, new_n17745);
nand_5 g15397(new_n17745, new_n17743, new_n17746_1);
nand_5 g15398(new_n17746_1, new_n17741, new_n17747);
xnor_4 g15399(new_n17737, new_n8688, new_n17748);
nand_5 g15400(new_n17748, new_n17747, new_n17749_1);
nand_5 g15401(new_n17749_1, new_n17739, new_n17750);
nand_5 g15402(new_n17750, new_n17735_1, new_n17751);
nand_5 g15403(new_n17751, new_n17734, new_n17752);
nand_5 g15404(new_n17752, new_n17732, new_n17753);
nand_5 g15405(new_n17753, new_n17731, new_n17754);
nand_5 g15406(new_n17754, new_n17727, new_n17755);
nand_5 g15407(new_n17755, new_n17726, new_n17756);
nand_5 g15408(new_n17756, new_n17724, new_n17757);
nand_5 g15409(new_n17757, new_n17723, new_n17758);
nand_5 g15410(new_n17758, new_n17721_1, new_n17759);
nand_5 g15411(new_n17759, new_n17720, new_n17760);
xnor_4 g15412(new_n17760, new_n17716, n3983);
not_8  g15413(new_n7024, new_n17762);
xnor_4 g15414(n13714, n583, new_n17763);
xnor_4 g15415(new_n17763, n6611, new_n17764);
nor_5  g15416(new_n17764, new_n17762, new_n17765);
nor_5  g15417(new_n17763, new_n9555, new_n17766);
nand_5 g15418(n13714, n583, new_n17767);
xnor_4 g15419(n22173, n12593, new_n17768);
xnor_4 g15420(new_n17768, new_n17767, new_n17769);
xnor_4 g15421(new_n17769, new_n5882_1, new_n17770);
not_8  g15422(new_n17770, new_n17771);
xnor_4 g15423(new_n17771, new_n17766, new_n17772);
xnor_4 g15424(new_n17772, new_n17765, new_n17773);
xor_4  g15425(new_n17773, new_n7021, n4000);
xnor_4 g15426(n26823, n20179, new_n17775);
nor_5  g15427(n19228, new_n2438, new_n17776);
xnor_4 g15428(n19228, n4812, new_n17777);
not_8  g15429(new_n17777, new_n17778);
nor_5  g15430(new_n2442, n15539, new_n17779);
xnor_4 g15431(n24278, n15539, new_n17780);
not_8  g15432(new_n17780, new_n17781);
nor_5  g15433(new_n2446, n8052, new_n17782);
nor_5  g15434(n24618, new_n7136, new_n17783);
nand_5 g15435(n10158, new_n3348, new_n17784_1);
nand_5 g15436(new_n11974, new_n11973, new_n17785);
nand_5 g15437(new_n17785, new_n17784_1, new_n17786);
nor_5  g15438(new_n17786, new_n17783, new_n17787);
nor_5  g15439(new_n17787, new_n17782, new_n17788);
nor_5  g15440(new_n17788, new_n17781, new_n17789);
nor_5  g15441(new_n17789, new_n17779, new_n17790);
nor_5  g15442(new_n17790, new_n17778, new_n17791);
nor_5  g15443(new_n17791, new_n17776, new_n17792);
xnor_4 g15444(new_n17792, new_n17775, new_n17793);
xnor_4 g15445(new_n17793, new_n7833, new_n17794);
xnor_4 g15446(new_n17790, new_n17777, new_n17795);
not_8  g15447(new_n17795, new_n17796);
nand_5 g15448(new_n17796, new_n7839, new_n17797);
xnor_4 g15449(new_n17795, new_n7839, new_n17798);
xnor_4 g15450(new_n17788, new_n17780, new_n17799);
not_8  g15451(new_n17799, new_n17800);
nand_5 g15452(new_n17800, new_n7843, new_n17801);
xnor_4 g15453(n24618, n8052, new_n17802);
xnor_4 g15454(new_n17802, new_n17786, new_n17803);
nor_5  g15455(new_n17803, new_n7846, new_n17804);
not_8  g15456(new_n17804, new_n17805);
xnor_4 g15457(new_n17803, new_n7846, new_n17806);
not_8  g15458(new_n17806, new_n17807);
and_5  g15459(new_n11975, new_n11972, new_n17808);
not_8  g15460(new_n7862, new_n17809);
nor_5  g15461(new_n11976, new_n17809, new_n17810);
nor_5  g15462(new_n17810, new_n17808, new_n17811);
nand_5 g15463(new_n17811, new_n17807, new_n17812);
nand_5 g15464(new_n17812, new_n17805, new_n17813);
xnor_4 g15465(new_n17800, new_n7842, new_n17814);
nand_5 g15466(new_n17814, new_n17813, new_n17815);
nand_5 g15467(new_n17815, new_n17801, new_n17816);
nand_5 g15468(new_n17816, new_n17798, new_n17817);
nand_5 g15469(new_n17817, new_n17797, new_n17818);
xnor_4 g15470(new_n17818, new_n17794, n4010);
xnor_4 g15471(n11220, n2160, new_n17820_1);
not_8  g15472(n10763, new_n17821);
or_5   g15473(n22379, new_n17821, new_n17822);
xnor_4 g15474(n22379, n10763, new_n17823);
or_5   g15475(new_n2944_1, n1662, new_n17824);
xnor_4 g15476(n7437, n1662, new_n17825);
or_5   g15477(new_n2947, n12875, new_n17826);
or_5   g15478(new_n2951, n2035, new_n17827);
nand_5 g15479(new_n15664, new_n15645, new_n17828);
nand_5 g15480(new_n17828, new_n17827, new_n17829);
xnor_4 g15481(n20700, n12875, new_n17830);
nand_5 g15482(new_n17830, new_n17829, new_n17831);
nand_5 g15483(new_n17831, new_n17826, new_n17832);
nand_5 g15484(new_n17832, new_n17825, new_n17833);
nand_5 g15485(new_n17833, new_n17824, new_n17834);
nand_5 g15486(new_n17834, new_n17823, new_n17835);
nand_5 g15487(new_n17835, new_n17822, new_n17836);
xnor_4 g15488(new_n17836, new_n17820_1, new_n17837);
xnor_4 g15489(new_n17837, new_n15818, new_n17838);
not_8  g15490(new_n17838, new_n17839);
xnor_4 g15491(new_n17834, new_n17823, new_n17840);
nand_5 g15492(new_n17840, new_n15827, new_n17841);
xnor_4 g15493(new_n17840, new_n15826, new_n17842);
xnor_4 g15494(new_n17832, new_n17825, new_n17843);
nand_5 g15495(new_n17843, new_n15832, new_n17844);
xnor_4 g15496(new_n17830, new_n17829, new_n17845);
nor_5  g15497(new_n17845, new_n15835, new_n17846);
xnor_4 g15498(new_n17845, new_n15835, new_n17847);
nor_5  g15499(new_n15679, new_n15665, new_n17848);
nor_5  g15500(new_n15708, new_n15680, new_n17849);
nor_5  g15501(new_n17849, new_n17848, new_n17850);
nor_5  g15502(new_n17850, new_n17847, new_n17851);
nor_5  g15503(new_n17851, new_n17846, new_n17852);
not_8  g15504(new_n15832, new_n17853);
xnor_4 g15505(new_n17843, new_n17853, new_n17854);
nand_5 g15506(new_n17854, new_n17852, new_n17855_1);
nand_5 g15507(new_n17855_1, new_n17844, new_n17856);
nand_5 g15508(new_n17856, new_n17842, new_n17857);
nand_5 g15509(new_n17857, new_n17841, new_n17858);
xnor_4 g15510(new_n17858, new_n17839, n4014);
xnor_4 g15511(new_n15060, new_n12518, new_n17860);
nand_5 g15512(new_n15065, new_n13529, new_n17861);
xnor_4 g15513(new_n15064, new_n13529, new_n17862);
nand_5 g15514(new_n15068, new_n3878, new_n17863);
nand_5 g15515(new_n3924, new_n3887, new_n17864);
nand_5 g15516(new_n17864, new_n17863, new_n17865);
nand_5 g15517(new_n17865, new_n17862, new_n17866);
nand_5 g15518(new_n17866, new_n17861, new_n17867);
xnor_4 g15519(new_n17867, new_n17860, new_n17868);
xnor_4 g15520(new_n17868, new_n5046_1, new_n17869);
xnor_4 g15521(new_n17865, new_n17862, new_n17870);
nand_5 g15522(new_n17870, n20409, new_n17871);
xnor_4 g15523(new_n17870, new_n6243, new_n17872);
nand_5 g15524(new_n3925_1, n25749, new_n17873);
nand_5 g15525(new_n3961, new_n3926, new_n17874);
nand_5 g15526(new_n17874, new_n17873, new_n17875);
nand_5 g15527(new_n17875, new_n17872, new_n17876);
nand_5 g15528(new_n17876, new_n17871, new_n17877_1);
xnor_4 g15529(new_n17877_1, new_n17869, new_n17878);
xnor_4 g15530(new_n17878, new_n12640, new_n17879);
xnor_4 g15531(new_n17875, new_n17872, new_n17880);
nand_5 g15532(new_n17880, new_n12646, new_n17881);
not_8  g15533(new_n12646, new_n17882);
xnor_4 g15534(new_n17880, new_n17882, new_n17883);
nand_5 g15535(new_n12649, new_n3962_1, new_n17884);
nand_5 g15536(new_n4093, new_n4054, new_n17885);
nand_5 g15537(new_n17885, new_n17884, new_n17886);
nand_5 g15538(new_n17886, new_n17883, new_n17887);
nand_5 g15539(new_n17887, new_n17881, new_n17888);
xnor_4 g15540(new_n17888, new_n17879, n4071);
xnor_4 g15541(new_n13736, new_n13728, n4088);
or_5   g15542(new_n13865, n7593, new_n17891);
or_5   g15543(new_n13866, n5025, new_n17892);
nand_5 g15544(new_n13866, n5025, new_n17893);
nand_5 g15545(new_n13870, new_n17893, new_n17894);
nand_5 g15546(new_n17894, new_n17892, new_n17895);
nand_5 g15547(new_n17895, new_n17891, new_n17896);
not_8  g15548(new_n17284, new_n17897);
and_5  g15549(new_n17287, new_n17897, new_n17898);
nor_5  g15550(new_n17287, new_n17897, new_n17899);
nor_5  g15551(new_n17293, new_n17899, new_n17900);
nor_5  g15552(new_n17900, new_n17898, new_n17901);
not_8  g15553(new_n17901, new_n17902);
nor_5  g15554(new_n17902, new_n17896, new_n17903);
not_8  g15555(new_n17294, new_n17904);
not_8  g15556(new_n17896, new_n17905);
nor_5  g15557(new_n17905, new_n17904, new_n17906);
nor_5  g15558(new_n17896, new_n17294, new_n17907);
nand_5 g15559(new_n13871, new_n13863, new_n17908);
xnor_4 g15560(new_n13871, new_n13862, new_n17909);
nand_5 g15561(new_n13875, new_n17909, new_n17910);
nand_5 g15562(new_n17910, new_n17908, new_n17911_1);
nor_5  g15563(new_n17911_1, new_n17907, new_n17912_1);
nor_5  g15564(new_n17912_1, new_n17906, new_n17913);
nor_5  g15565(new_n17913, new_n17903, new_n17914);
nor_5  g15566(new_n17901, new_n17905, new_n17915);
nor_5  g15567(new_n17915, new_n17912_1, new_n17916);
nor_5  g15568(new_n17916, new_n17914, n4089);
nand_5 g15569(new_n12878, new_n7122, new_n17918);
xnor_4 g15570(new_n17918, new_n7118, new_n17919);
xnor_4 g15571(new_n17919, new_n3390_1, new_n17920);
nor_5  g15572(new_n12879, n5302, new_n17921);
not_8  g15573(new_n17921, new_n17922);
xnor_4 g15574(new_n12879, new_n3393, new_n17923);
nor_5  g15575(new_n12882, new_n5504, new_n17924);
nor_5  g15576(new_n12881, n25738, new_n17925);
nor_5  g15577(new_n9115, n21471, new_n17926);
not_8  g15578(new_n17926, new_n17927_1);
nand_5 g15579(new_n9135, new_n9116, new_n17928);
nand_5 g15580(new_n17928, new_n17927_1, new_n17929);
nor_5  g15581(new_n17929, new_n17925, new_n17930);
nor_5  g15582(new_n17930, new_n17924, new_n17931_1);
nand_5 g15583(new_n17931_1, new_n17923, new_n17932);
nand_5 g15584(new_n17932, new_n17922, new_n17933);
xnor_4 g15585(new_n17933, new_n17920, new_n17934);
xnor_4 g15586(new_n17934, new_n7219, new_n17935);
xnor_4 g15587(new_n17931_1, new_n17923, new_n17936);
nor_5  g15588(new_n17936, n1293, new_n17937);
not_8  g15589(new_n17937, new_n17938);
xnor_4 g15590(new_n17936, new_n7223, new_n17939);
xnor_4 g15591(new_n12881, new_n5504, new_n17940);
xnor_4 g15592(new_n17940, new_n17929, new_n17941);
nand_5 g15593(new_n17941, n19042, new_n17942);
not_8  g15594(new_n17942, new_n17943);
not_8  g15595(new_n9136, new_n17944);
nor_5  g15596(new_n17944, new_n9111, new_n17945);
nor_5  g15597(new_n9168, new_n9138, new_n17946);
nor_5  g15598(new_n17946, new_n17945, new_n17947);
xnor_4 g15599(new_n17941, new_n7227, new_n17948_1);
not_8  g15600(new_n17948_1, new_n17949);
nor_5  g15601(new_n17949, new_n17947, new_n17950);
nor_5  g15602(new_n17950, new_n17943, new_n17951);
nand_5 g15603(new_n17951, new_n17939, new_n17952);
nand_5 g15604(new_n17952, new_n17938, new_n17953);
xnor_4 g15605(new_n17953, new_n17935, new_n17954_1);
xnor_4 g15606(new_n8004, n11736, new_n17955);
nand_5 g15607(new_n2464, n23200, new_n17956_1);
xnor_4 g15608(new_n2464, n23200, new_n17957);
not_8  g15609(new_n17957, new_n17958);
nand_5 g15610(new_n2470, n17959, new_n17959_1);
xnor_4 g15611(new_n2470, new_n5749, new_n17960);
nand_5 g15612(new_n2476, n7566, new_n17961);
nand_5 g15613(new_n7054, new_n7040, new_n17962);
nand_5 g15614(new_n17962, new_n17961, new_n17963_1);
nand_5 g15615(new_n17963_1, new_n17960, new_n17964);
nand_5 g15616(new_n17964, new_n17959_1, new_n17965);
nand_5 g15617(new_n17965, new_n17958, new_n17966);
nand_5 g15618(new_n17966, new_n17956_1, new_n17967);
xnor_4 g15619(new_n17967, new_n17955, new_n17968_1);
xnor_4 g15620(new_n17968_1, new_n17954_1, new_n17969);
not_8  g15621(new_n17939, new_n17970);
not_8  g15622(new_n17945, new_n17971);
not_8  g15623(new_n9168, new_n17972);
nand_5 g15624(new_n17972, new_n9137, new_n17973);
nand_5 g15625(new_n17973, new_n17971, new_n17974);
nand_5 g15626(new_n17948_1, new_n17974, new_n17975);
nand_5 g15627(new_n17975, new_n17942, new_n17976_1);
xnor_4 g15628(new_n17976_1, new_n17970, new_n17977);
not_8  g15629(new_n17977, new_n17978);
xnor_4 g15630(new_n17965, new_n17957, new_n17979);
not_8  g15631(new_n17979, new_n17980);
nand_5 g15632(new_n17980, new_n17978, new_n17981);
xnor_4 g15633(new_n17980, new_n17977, new_n17982);
xnor_4 g15634(new_n17963_1, new_n17960, new_n17983);
xnor_4 g15635(new_n17948_1, new_n17947, new_n17984);
not_8  g15636(new_n17984, new_n17985);
nand_5 g15637(new_n17985, new_n17983, new_n17986);
nand_5 g15638(new_n9169, new_n7055, new_n17987);
nand_5 g15639(new_n9193, new_n9170, new_n17988);
nand_5 g15640(new_n17988, new_n17987, new_n17989);
xnor_4 g15641(new_n17984, new_n17983, new_n17990);
nand_5 g15642(new_n17990, new_n17989, new_n17991);
nand_5 g15643(new_n17991, new_n17986, new_n17992);
nand_5 g15644(new_n17992, new_n17982, new_n17993);
nand_5 g15645(new_n17993, new_n17981, new_n17994);
xnor_4 g15646(new_n17994, new_n17969, n4103);
nand_5 g15647(new_n15744, new_n13595, new_n17996);
not_8  g15648(new_n17996, new_n17997);
xnor_4 g15649(new_n15744, new_n13595, new_n17998_1);
nand_5 g15650(new_n15747, new_n13522, new_n17999);
nand_5 g15651(new_n15752, new_n13527, new_n18000);
xnor_4 g15652(new_n15752, new_n13525, new_n18001);
nand_5 g15653(new_n17301, new_n13533, new_n18002);
xnor_4 g15654(new_n15757, new_n13533, new_n18003);
nand_5 g15655(new_n15760, new_n13538, new_n18004);
xnor_4 g15656(new_n15760, new_n13536, new_n18005);
nand_5 g15657(new_n15673, new_n13543, new_n18006);
nand_5 g15658(new_n13548_1, new_n4438, new_n18007);
xnor_4 g15659(new_n13546, new_n4438, new_n18008);
nor_5  g15660(new_n13553, new_n4442, new_n18009);
xnor_4 g15661(new_n13553, new_n4442, new_n18010);
nor_5  g15662(new_n13555, new_n4447, new_n18011);
not_8  g15663(new_n18011, new_n18012);
xnor_4 g15664(new_n13555, new_n4446, new_n18013);
nor_5  g15665(new_n13562, new_n4450, new_n18014);
not_8  g15666(new_n18014, new_n18015);
nor_5  g15667(new_n13568, new_n4454, new_n18016);
not_8  g15668(new_n18016, new_n18017);
xnor_4 g15669(new_n13562, new_n4449, new_n18018);
nand_5 g15670(new_n18018, new_n18017, new_n18019);
nand_5 g15671(new_n18019, new_n18015, new_n18020);
nand_5 g15672(new_n18020, new_n18013, new_n18021);
nand_5 g15673(new_n18021, new_n18012, new_n18022);
nor_5  g15674(new_n18022, new_n18010, new_n18023);
nor_5  g15675(new_n18023, new_n18009, new_n18024);
nand_5 g15676(new_n18024, new_n18008, new_n18025_1);
nand_5 g15677(new_n18025_1, new_n18007, new_n18026);
xnor_4 g15678(new_n15673, new_n13541, new_n18027);
nand_5 g15679(new_n18027, new_n18026, new_n18028);
nand_5 g15680(new_n18028, new_n18006, new_n18029);
nand_5 g15681(new_n18029, new_n18005, new_n18030);
nand_5 g15682(new_n18030, new_n18004, new_n18031);
nand_5 g15683(new_n18031, new_n18003, new_n18032);
nand_5 g15684(new_n18032, new_n18002, new_n18033);
nand_5 g15685(new_n18033, new_n18001, new_n18034);
nand_5 g15686(new_n18034, new_n18000, new_n18035_1);
xnor_4 g15687(new_n15747, new_n13520, new_n18036);
nand_5 g15688(new_n18036, new_n18035_1, new_n18037);
nand_5 g15689(new_n18037, new_n17999, new_n18038);
nor_5  g15690(new_n18038, new_n17998_1, new_n18039);
nor_5  g15691(new_n18039, new_n17997, new_n18040);
not_8  g15692(new_n18040, new_n18041);
nor_5  g15693(new_n6186, new_n6188, new_n18042);
not_8  g15694(new_n18042, new_n18043_1);
nor_5  g15695(new_n6187, n6456, new_n18044);
or_5   g15696(new_n6238, n4085, new_n18045_1);
xnor_4 g15697(new_n6238, new_n6191, new_n18046);
or_5   g15698(new_n6244, n26725, new_n18047);
xnor_4 g15699(new_n6245_1, n26725, new_n18048);
or_5   g15700(new_n6250, n11980, new_n18049);
xnor_4 g15701(new_n6250, new_n6196, new_n18050);
or_5   g15702(new_n6256_1, n3253, new_n18051);
xnor_4 g15703(new_n6256_1, new_n6200, new_n18052);
nand_5 g15704(new_n6266, new_n6204_1, new_n18053);
xnor_4 g15705(new_n6262, new_n6204_1, new_n18054);
nand_5 g15706(new_n6272, new_n6208, new_n18055);
nand_5 g15707(new_n6275, new_n6212, new_n18056);
xnor_4 g15708(new_n6274, new_n6212, new_n18057);
nand_5 g15709(new_n6288, new_n13905, new_n18058);
not_8  g15710(new_n18058, new_n18059_1);
nand_5 g15711(n20658, n14575, new_n18060);
not_8  g15712(new_n18060, new_n18061_1);
xnor_4 g15713(new_n6288, n24374, new_n18062);
not_8  g15714(new_n18062, new_n18063);
nor_5  g15715(new_n18063, new_n18061_1, new_n18064);
nor_5  g15716(new_n18064, new_n18059_1, new_n18065);
not_8  g15717(new_n18065, new_n18066);
nand_5 g15718(new_n18066, new_n18057, new_n18067);
nand_5 g15719(new_n18067, new_n18056, new_n18068);
xnor_4 g15720(new_n6268, new_n6208, new_n18069);
nand_5 g15721(new_n18069, new_n18068, new_n18070);
nand_5 g15722(new_n18070, new_n18055, new_n18071_1);
nand_5 g15723(new_n18071_1, new_n18054, new_n18072);
nand_5 g15724(new_n18072, new_n18053, new_n18073);
nand_5 g15725(new_n18073, new_n18052, new_n18074);
nand_5 g15726(new_n18074, new_n18051, new_n18075);
nand_5 g15727(new_n18075, new_n18050, new_n18076);
nand_5 g15728(new_n18076, new_n18049, new_n18077);
nand_5 g15729(new_n18077, new_n18048, new_n18078);
nand_5 g15730(new_n18078, new_n18047, new_n18079);
nand_5 g15731(new_n18079, new_n18046, new_n18080);
nand_5 g15732(new_n18080, new_n18045_1, new_n18081);
nor_5  g15733(new_n18081, new_n18044, new_n18082);
nor_5  g15734(new_n18082, new_n14691, new_n18083);
nand_5 g15735(new_n18083, new_n18043_1, new_n18084);
not_8  g15736(new_n18084, new_n18085);
nand_5 g15737(new_n18085, new_n18041, new_n18086);
xnor_4 g15738(new_n18038, new_n17998_1, new_n18087);
nand_5 g15739(new_n18087, new_n18084, new_n18088);
xnor_4 g15740(new_n18087, new_n18085, new_n18089);
not_8  g15741(new_n18036, new_n18090);
xnor_4 g15742(new_n18090, new_n18035_1, new_n18091);
xnor_4 g15743(new_n6186, n6456, new_n18092);
xnor_4 g15744(new_n18092, new_n18081, new_n18093);
not_8  g15745(new_n18093, new_n18094);
nand_5 g15746(new_n18094, new_n18091, new_n18095);
xnor_4 g15747(new_n18093, new_n18091, new_n18096);
xnor_4 g15748(new_n18079, new_n18046, new_n18097);
not_8  g15749(new_n18097, new_n18098);
not_8  g15750(new_n18001, new_n18099);
xnor_4 g15751(new_n18033, new_n18099, new_n18100);
nand_5 g15752(new_n18100, new_n18098, new_n18101);
xnor_4 g15753(new_n18100, new_n18097, new_n18102);
xnor_4 g15754(new_n18077, new_n18048, new_n18103);
not_8  g15755(new_n18103, new_n18104);
not_8  g15756(new_n18003, new_n18105_1);
xnor_4 g15757(new_n18031, new_n18105_1, new_n18106);
nand_5 g15758(new_n18106, new_n18104, new_n18107);
xnor_4 g15759(new_n18106, new_n18103, new_n18108);
xnor_4 g15760(new_n18075, new_n18050, new_n18109);
not_8  g15761(new_n18109, new_n18110);
not_8  g15762(new_n18005, new_n18111);
xnor_4 g15763(new_n18029, new_n18111, new_n18112);
nand_5 g15764(new_n18112, new_n18110, new_n18113);
xnor_4 g15765(new_n18112, new_n18109, new_n18114);
xnor_4 g15766(new_n18073, new_n18052, new_n18115);
not_8  g15767(new_n18115, new_n18116);
not_8  g15768(new_n18027, new_n18117);
xnor_4 g15769(new_n18117, new_n18026, new_n18118);
nand_5 g15770(new_n18118, new_n18116, new_n18119);
xnor_4 g15771(new_n18118, new_n18115, new_n18120);
not_8  g15772(new_n18054, new_n18121);
xnor_4 g15773(new_n18071_1, new_n18121, new_n18122);
xnor_4 g15774(new_n18024, new_n18008, new_n18123);
not_8  g15775(new_n18123, new_n18124);
nand_5 g15776(new_n18124, new_n18122, new_n18125);
xnor_4 g15777(new_n18123, new_n18122, new_n18126);
xnor_4 g15778(new_n18022, new_n18010, new_n18127);
not_8  g15779(new_n18127, new_n18128);
xnor_4 g15780(new_n18069, new_n18068, new_n18129);
nor_5  g15781(new_n18129, new_n18128, new_n18130);
not_8  g15782(new_n18130, new_n18131);
xnor_4 g15783(new_n18129, new_n18127, new_n18132);
xnor_4 g15784(new_n18065, new_n18057, new_n18133);
not_8  g15785(new_n18020, new_n18134);
xnor_4 g15786(new_n18134, new_n18013, new_n18135);
nor_5  g15787(new_n18135, new_n18133, new_n18136);
xnor_4 g15788(new_n18135, new_n18133, new_n18137);
xnor_4 g15789(new_n18018, new_n18016, new_n18138);
not_8  g15790(new_n18138, new_n18139);
nor_5  g15791(new_n18139, new_n18062, new_n18140);
not_8  g15792(new_n18140, new_n18141);
xnor_4 g15793(new_n18062, new_n18061_1, new_n18142);
nor_5  g15794(new_n18142, new_n18138, new_n18143_1);
not_8  g15795(new_n18143_1, new_n18144);
xnor_4 g15796(n20658, new_n6281, new_n18145_1);
xnor_4 g15797(new_n13567, new_n4454, new_n18146);
and_5  g15798(new_n18146, new_n18145_1, new_n18147);
not_8  g15799(new_n18147, new_n18148);
nand_5 g15800(new_n18148, new_n18144, new_n18149);
nand_5 g15801(new_n18149, new_n18141, new_n18150);
nor_5  g15802(new_n18150, new_n18137, new_n18151_1);
nor_5  g15803(new_n18151_1, new_n18136, new_n18152_1);
nand_5 g15804(new_n18152_1, new_n18132, new_n18153);
nand_5 g15805(new_n18153, new_n18131, new_n18154);
nand_5 g15806(new_n18154, new_n18126, new_n18155);
nand_5 g15807(new_n18155, new_n18125, new_n18156);
nand_5 g15808(new_n18156, new_n18120, new_n18157_1);
nand_5 g15809(new_n18157_1, new_n18119, new_n18158);
nand_5 g15810(new_n18158, new_n18114, new_n18159);
nand_5 g15811(new_n18159, new_n18113, new_n18160);
nand_5 g15812(new_n18160, new_n18108, new_n18161);
nand_5 g15813(new_n18161, new_n18107, new_n18162);
nand_5 g15814(new_n18162, new_n18102, new_n18163);
nand_5 g15815(new_n18163, new_n18101, new_n18164);
nand_5 g15816(new_n18164, new_n18096, new_n18165);
nand_5 g15817(new_n18165, new_n18095, new_n18166);
nand_5 g15818(new_n18166, new_n18089, new_n18167);
nand_5 g15819(new_n18167, new_n18088, new_n18168);
nand_5 g15820(new_n18168, new_n18086, new_n18169);
nand_5 g15821(new_n18084, new_n18040, new_n18170);
nand_5 g15822(new_n18170, new_n18167, new_n18171_1);
nand_5 g15823(new_n18171_1, new_n18169, new_n18172);
not_8  g15824(new_n18172, n4123);
xnor_4 g15825(new_n14132, new_n8365, new_n18174);
not_8  g15826(new_n14138, new_n18175);
nand_5 g15827(new_n18175, new_n8375, new_n18176);
xnor_4 g15828(new_n14138, new_n8375, new_n18177);
not_8  g15829(new_n14143, new_n18178);
nand_5 g15830(new_n18178, new_n8396, new_n18179);
xnor_4 g15831(new_n14143, new_n8396, new_n18180);
not_8  g15832(new_n8381_1, new_n18181);
nor_5  g15833(new_n14156, new_n18181, new_n18182);
nor_5  g15834(new_n14149, new_n8384, new_n18183);
not_8  g15835(new_n18183, new_n18184);
xnor_4 g15836(new_n14155, new_n8381_1, new_n18185);
nor_5  g15837(new_n18185, new_n18184, new_n18186);
nor_5  g15838(new_n18186, new_n18182, new_n18187);
nand_5 g15839(new_n18187, new_n18180, new_n18188);
nand_5 g15840(new_n18188, new_n18179, new_n18189);
nand_5 g15841(new_n18189, new_n18177, new_n18190);
nand_5 g15842(new_n18190, new_n18176, new_n18191);
xnor_4 g15843(new_n18191, new_n18174, n4134);
xnor_4 g15844(new_n9650, new_n9589, n4146);
xnor_4 g15845(new_n16326, new_n15158, new_n18194);
not_8  g15846(new_n16330, new_n18195);
nor_5  g15847(new_n18195, new_n15164, new_n18196);
xnor_4 g15848(new_n18195, new_n15164, new_n18197);
nor_5  g15849(new_n15168, new_n14233, new_n18198);
nor_5  g15850(new_n15173, new_n14228, new_n18199);
not_8  g15851(new_n18199, new_n18200);
xnor_4 g15852(new_n15167_1, new_n14233, new_n18201);
not_8  g15853(new_n18201, new_n18202);
nor_5  g15854(new_n18202, new_n18200, new_n18203);
nor_5  g15855(new_n18203, new_n18198, new_n18204);
not_8  g15856(new_n18204, new_n18205);
nor_5  g15857(new_n18205, new_n18197, new_n18206);
nor_5  g15858(new_n18206, new_n18196, new_n18207);
xnor_4 g15859(new_n18207, new_n18194, n4150);
xnor_4 g15860(new_n13330, new_n13329, n4151);
xnor_4 g15861(new_n13671, new_n13606, n4152);
xnor_4 g15862(new_n6469, new_n6427_1, n4153);
or_5   g15863(new_n12752, n10250, new_n18212);
nand_5 g15864(new_n9233, new_n9195, new_n18213);
nand_5 g15865(new_n18213, new_n18212, new_n18214);
xnor_4 g15866(new_n18214, new_n13011, new_n18215);
nor_5  g15867(new_n18214, new_n13016, new_n18216);
not_8  g15868(new_n13016, new_n18217);
not_8  g15869(new_n18214, new_n18218);
nor_5  g15870(new_n18218, new_n18217, new_n18219);
nor_5  g15871(new_n9411, new_n9234, new_n18220);
nor_5  g15872(new_n9478, new_n9412, new_n18221);
nor_5  g15873(new_n18221, new_n18220, new_n18222);
nor_5  g15874(new_n18222, new_n18219, new_n18223);
nor_5  g15875(new_n18223, new_n18216, new_n18224);
xnor_4 g15876(new_n18224, new_n18215, n4165);
xnor_4 g15877(new_n12268, new_n12234, n4172);
xnor_4 g15878(new_n12084, new_n4978, n4173);
xnor_4 g15879(new_n6934, new_n6910, n4176);
xnor_4 g15880(new_n9634, new_n9632, n4186);
xnor_4 g15881(new_n17754, new_n17727, n4204);
not_8  g15882(new_n12172, new_n18231);
not_8  g15883(new_n12138, new_n18232_1);
nand_5 g15884(new_n18232_1, n13494, new_n18233);
xnor_4 g15885(new_n12138, n13494, new_n18234);
not_8  g15886(new_n7157, new_n18235);
nand_5 g15887(new_n18235, n25345, new_n18236);
nand_5 g15888(new_n7214, new_n7158, new_n18237);
nand_5 g15889(new_n18237, new_n18236, new_n18238_1);
nand_5 g15890(new_n18238_1, new_n18234, new_n18239);
nand_5 g15891(new_n18239, new_n18233, new_n18240);
nand_5 g15892(new_n18240, new_n18231, new_n18241_1);
not_8  g15893(new_n18241_1, new_n18242);
nand_5 g15894(new_n17063, new_n11621, new_n18243);
nor_5  g15895(new_n18243, n19652, new_n18244);
xnor_4 g15896(new_n18244, n3984, new_n18245);
nand_5 g15897(new_n18245, new_n12174, new_n18246);
xnor_4 g15898(new_n18245, n17037, new_n18247);
xnor_4 g15899(new_n18243, new_n12117, new_n18248);
nor_5  g15900(new_n18248, new_n12198, new_n18249);
nand_5 g15901(new_n17064, new_n12175, new_n18250);
nand_5 g15902(new_n17094, new_n17065, new_n18251);
nand_5 g15903(new_n18251, new_n18250, new_n18252);
xnor_4 g15904(new_n18248, new_n12198, new_n18253);
nor_5  g15905(new_n18253, new_n18252, new_n18254_1);
nor_5  g15906(new_n18254_1, new_n18249, new_n18255);
nand_5 g15907(new_n18255, new_n18247, new_n18256);
nand_5 g15908(new_n18256, new_n18246, new_n18257);
nand_5 g15909(new_n18244, new_n12114, new_n18258);
xnor_4 g15910(new_n18258, new_n12110, new_n18259);
xnor_4 g15911(new_n18259, n7569, new_n18260);
xnor_4 g15912(new_n18260, new_n18257, new_n18261);
not_8  g15913(new_n18261, new_n18262);
nor_5  g15914(new_n18262, new_n15417, new_n18263);
not_8  g15915(new_n18263, new_n18264);
xnor_4 g15916(new_n18261, new_n15417, new_n18265);
xnor_4 g15917(new_n18255, new_n18247, new_n18266);
nand_5 g15918(new_n18266, n25751, new_n18267);
xnor_4 g15919(new_n18266, n25751, new_n18268);
not_8  g15920(new_n18268, new_n18269);
xnor_4 g15921(new_n18253, new_n18252, new_n18270);
not_8  g15922(new_n18270, new_n18271);
nor_5  g15923(new_n18271, n26053, new_n18272);
xnor_4 g15924(new_n18270, n26053, new_n18273);
not_8  g15925(new_n18273, new_n18274_1);
nor_5  g15926(new_n17095_1, n7917, new_n18275);
nor_5  g15927(new_n17129, new_n17096, new_n18276);
nor_5  g15928(new_n18276, new_n18275, new_n18277);
nor_5  g15929(new_n18277, new_n18274_1, new_n18278);
nor_5  g15930(new_n18278, new_n18272, new_n18279);
nand_5 g15931(new_n18279, new_n18269, new_n18280);
nand_5 g15932(new_n18280, new_n18267, new_n18281);
nand_5 g15933(new_n18281, new_n18265, new_n18282);
nand_5 g15934(new_n18282, new_n18264, new_n18283);
not_8  g15935(new_n18283, new_n18284);
nor_5  g15936(new_n18258, n4514, new_n18285);
not_8  g15937(new_n18285, new_n18286);
or_5   g15938(new_n18259, new_n12185, new_n18287);
nand_5 g15939(new_n18287, new_n18257, new_n18288_1);
nor_5  g15940(new_n18288_1, new_n18286, new_n18289);
nand_5 g15941(new_n18289, new_n18284, new_n18290_1);
not_8  g15942(new_n18290_1, new_n18291);
and_5  g15943(new_n18259, new_n12185, new_n18292);
xnor_4 g15944(new_n18288_1, new_n18285, new_n18293);
nor_5  g15945(new_n18293, new_n18292, new_n18294);
nand_5 g15946(new_n18294, new_n18283, new_n18295_1);
nor_5  g15947(new_n18295_1, new_n18289, new_n18296);
nor_5  g15948(new_n18296, new_n18291, new_n18297);
nor_5  g15949(new_n18297, new_n18242, new_n18298);
xnor_4 g15950(new_n18294, new_n18283, new_n18299);
not_8  g15951(new_n18299, new_n18300);
xnor_4 g15952(new_n18240, new_n12172, new_n18301_1);
not_8  g15953(new_n18301_1, new_n18302);
nand_5 g15954(new_n18302, new_n18300, new_n18303);
xnor_4 g15955(new_n18302, new_n18299, new_n18304_1);
not_8  g15956(new_n18265, new_n18305);
xnor_4 g15957(new_n18281, new_n18305, new_n18306);
not_8  g15958(new_n18234, new_n18307);
xnor_4 g15959(new_n18238_1, new_n18307, new_n18308);
not_8  g15960(new_n18308, new_n18309);
nand_5 g15961(new_n18309, new_n18306, new_n18310_1);
xnor_4 g15962(new_n18308, new_n18306, new_n18311_1);
xnor_4 g15963(new_n18279, new_n18268, new_n18312);
nand_5 g15964(new_n18312, new_n7216, new_n18313);
xnor_4 g15965(new_n18312, new_n7215, new_n18314);
xnor_4 g15966(new_n18277, new_n18274_1, new_n18315);
nand_5 g15967(new_n18315, new_n7300, new_n18316);
not_8  g15968(new_n17130_1, new_n18317);
nand_5 g15969(new_n18317, new_n7305_1, new_n18318);
nand_5 g15970(new_n17166, new_n17131, new_n18319);
nand_5 g15971(new_n18319, new_n18318, new_n18320);
xnor_4 g15972(new_n18315, new_n7298_1, new_n18321);
nand_5 g15973(new_n18321, new_n18320, new_n18322);
nand_5 g15974(new_n18322, new_n18316, new_n18323_1);
nand_5 g15975(new_n18323_1, new_n18314, new_n18324);
nand_5 g15976(new_n18324, new_n18313, new_n18325);
nand_5 g15977(new_n18325, new_n18311_1, new_n18326);
nand_5 g15978(new_n18326, new_n18310_1, new_n18327);
nand_5 g15979(new_n18327, new_n18304_1, new_n18328);
nand_5 g15980(new_n18328, new_n18303, new_n18329);
nor_5  g15981(new_n18329, new_n18298, new_n18330);
nand_5 g15982(new_n18297, new_n18242, new_n18331);
nand_5 g15983(new_n18331, new_n18290_1, new_n18332_1);
nor_5  g15984(new_n18332_1, new_n18330, n4205);
nor_5  g15985(new_n14047, n22198, new_n18334);
nand_5 g15986(new_n18334, new_n5166, new_n18335);
xnor_4 g15987(new_n18335, new_n5162, new_n18336);
xnor_4 g15988(new_n18336, new_n4998, new_n18337);
xnor_4 g15989(new_n18334, n24327, new_n18338);
not_8  g15990(new_n18338, new_n18339);
nand_5 g15991(new_n18339, new_n8721_1, new_n18340);
xnor_4 g15992(new_n18338, new_n8721_1, new_n18341);
not_8  g15993(new_n14048, new_n18342);
nand_5 g15994(new_n18342, new_n5004, new_n18343_1);
nand_5 g15995(new_n14073, new_n14049, new_n18344);
nand_5 g15996(new_n18344, new_n18343_1, new_n18345_1);
nand_5 g15997(new_n18345_1, new_n18341, new_n18346);
nand_5 g15998(new_n18346, new_n18340, new_n18347);
xnor_4 g15999(new_n18347, new_n18337, new_n18348);
xnor_4 g16000(new_n18348, new_n8202, new_n18349);
xnor_4 g16001(new_n18345_1, new_n18341, new_n18350_1);
not_8  g16002(new_n18350_1, new_n18351);
nor_5  g16003(new_n18351, new_n8207, new_n18352);
xnor_4 g16004(new_n18350_1, new_n8207, new_n18353);
not_8  g16005(new_n18353, new_n18354);
nor_5  g16006(new_n14074, new_n8213, new_n18355);
not_8  g16007(new_n18355, new_n18356);
not_8  g16008(new_n14075, new_n18357);
nand_5 g16009(new_n14106, new_n18357, new_n18358);
nand_5 g16010(new_n18358, new_n18356, new_n18359);
nor_5  g16011(new_n18359, new_n18354, new_n18360);
nor_5  g16012(new_n18360, new_n18352, new_n18361);
xnor_4 g16013(new_n18361, new_n18349, new_n18362_1);
xnor_4 g16014(n21997, n5400, new_n18363);
or_5   g16015(n25119, new_n8795, new_n18364);
xnor_4 g16016(n25119, n23923, new_n18365);
or_5   g16017(n1163, new_n7415, new_n18366);
not_8  g16018(new_n14110, new_n18367);
not_8  g16019(new_n14113, new_n18368);
not_8  g16020(new_n14125, new_n18369);
nand_5 g16021(new_n18369, new_n18368, new_n18370);
nand_5 g16022(new_n18370, new_n14111, new_n18371);
nand_5 g16023(new_n18371, new_n18367, new_n18372);
nand_5 g16024(new_n18372, new_n14109, new_n18373);
nand_5 g16025(new_n18373, new_n18366, new_n18374);
nand_5 g16026(new_n18374, new_n18365, new_n18375);
nand_5 g16027(new_n18375, new_n18364, new_n18376);
xnor_4 g16028(new_n18376, new_n18363, new_n18377_1);
xnor_4 g16029(new_n18377_1, new_n18362_1, new_n18378);
xnor_4 g16030(new_n18374, new_n18365, new_n18379);
xnor_4 g16031(new_n18359, new_n18353, new_n18380);
not_8  g16032(new_n18380, new_n18381);
nor_5  g16033(new_n18381, new_n18379, new_n18382);
not_8  g16034(new_n18382, new_n18383);
xnor_4 g16035(new_n18380, new_n18379, new_n18384);
nor_5  g16036(new_n14129, new_n14108, new_n18385);
nor_5  g16037(new_n14166, new_n14130_1, new_n18386);
nor_5  g16038(new_n18386, new_n18385, new_n18387);
nand_5 g16039(new_n18387, new_n18384, new_n18388);
nand_5 g16040(new_n18388, new_n18383, new_n18389);
xor_4  g16041(new_n18389, new_n18378, n4215);
nand_5 g16042(new_n15206, new_n6312, new_n18391);
xnor_4 g16043(new_n18391, new_n6309, new_n18392);
xnor_4 g16044(new_n18392, new_n5220, new_n18393);
and_5  g16045(new_n15207, n2858, new_n18394);
nor_5  g16046(new_n15207, n2858, new_n18395);
nor_5  g16047(new_n15235, new_n18395, new_n18396);
nor_5  g16048(new_n18396, new_n18394, new_n18397);
xnor_4 g16049(new_n18397, new_n18393, new_n18398);
not_8  g16050(new_n18398, new_n18399);
nand_5 g16051(new_n10263, new_n4504, new_n18400);
xnor_4 g16052(new_n18400, new_n4501, new_n18401);
xnor_4 g16053(new_n18401, new_n7955, new_n18402);
nor_5  g16054(new_n10264, n14440, new_n18403);
not_8  g16055(new_n18403, new_n18404);
xnor_4 g16056(new_n10264, new_n7946, new_n18405_1);
nor_5  g16057(new_n10266, n1654, new_n18406);
not_8  g16058(new_n18406, new_n18407);
not_8  g16059(new_n16799, new_n18408);
not_8  g16060(new_n11308, new_n18409_1);
not_8  g16061(new_n11325_1, new_n18410);
nand_5 g16062(new_n18410, new_n11309, new_n18411);
nand_5 g16063(new_n18411, new_n18409_1, new_n18412);
nand_5 g16064(new_n18412, new_n11307, new_n18413);
nand_5 g16065(new_n18413, new_n18408, new_n18414_1);
nand_5 g16066(new_n18414_1, new_n16798_1, new_n18415);
nand_5 g16067(new_n18415, new_n18407, new_n18416);
nand_5 g16068(new_n18416, new_n18405_1, new_n18417);
nand_5 g16069(new_n18417, new_n18404, new_n18418_1);
xnor_4 g16070(new_n18418_1, new_n18402, new_n18419);
xnor_4 g16071(new_n18419, new_n18399, new_n18420);
not_8  g16072(new_n15236, new_n18421);
xnor_4 g16073(new_n18416, new_n18405_1, new_n18422);
not_8  g16074(new_n18422, new_n18423);
nor_5  g16075(new_n18423, new_n18421, new_n18424);
not_8  g16076(new_n18424, new_n18425);
nand_5 g16077(new_n16803, new_n15238, new_n18426);
not_8  g16078(new_n18426, new_n18427);
xnor_4 g16079(new_n16803, new_n15238, new_n18428);
not_8  g16080(new_n11328, new_n18429);
nor_5  g16081(new_n15241_1, new_n18429, new_n18430);
xnor_4 g16082(new_n15241_1, new_n11328, new_n18431);
not_8  g16083(new_n18431, new_n18432);
nand_5 g16084(new_n15244, new_n11330_1, new_n18433);
not_8  g16085(new_n18433, new_n18434);
xnor_4 g16086(new_n15244, new_n11330_1, new_n18435);
not_8  g16087(new_n11337, new_n18436);
nand_5 g16088(new_n15250, new_n18436, new_n18437_1);
xnor_4 g16089(new_n15250, new_n11337, new_n18438);
nand_5 g16090(new_n10058, new_n15253, new_n18439_1);
nand_5 g16091(new_n10077, new_n10059, new_n18440);
nand_5 g16092(new_n18440, new_n18439_1, new_n18441);
nand_5 g16093(new_n18441, new_n18438, new_n18442);
nand_5 g16094(new_n18442, new_n18437_1, new_n18443);
nor_5  g16095(new_n18443, new_n18435, new_n18444_1);
nor_5  g16096(new_n18444_1, new_n18434, new_n18445_1);
nor_5  g16097(new_n18445_1, new_n18432, new_n18446);
nor_5  g16098(new_n18446, new_n18430, new_n18447);
nor_5  g16099(new_n18447, new_n18428, new_n18448);
nor_5  g16100(new_n18448, new_n18427, new_n18449);
xnor_4 g16101(new_n18423, new_n15236, new_n18450);
nand_5 g16102(new_n18450, new_n18449, new_n18451);
nand_5 g16103(new_n18451, new_n18425, new_n18452_1);
xnor_4 g16104(new_n18452_1, new_n18420, new_n18453);
not_8  g16105(n23166, new_n18454);
nor_5  g16106(new_n15987, n10611, new_n18455);
nand_5 g16107(new_n18455, new_n9683, new_n18456);
nor_5  g16108(new_n18456, n11356, new_n18457);
nand_5 g16109(new_n18457, new_n9678, new_n18458);
nor_5  g16110(new_n18458, n6381, new_n18459);
nand_5 g16111(new_n18459, new_n9672, new_n18460);
xnor_4 g16112(new_n18460, new_n18454, new_n18461);
xnor_4 g16113(new_n18461, new_n8278, new_n18462);
not_8  g16114(new_n18462, new_n18463);
xnor_4 g16115(new_n18459, n10577, new_n18464);
or_5   g16116(new_n18464, n26408, new_n18465);
xnor_4 g16117(new_n18464, new_n8267_1, new_n18466);
xnor_4 g16118(new_n18458, new_n9675, new_n18467_1);
or_5   g16119(new_n18467_1, n18227, new_n18468);
xnor_4 g16120(new_n18467_1, new_n5049, new_n18469);
xnor_4 g16121(new_n18457, n14345, new_n18470);
or_5   g16122(new_n18470, n7377, new_n18471);
xnor_4 g16123(new_n18470, new_n5053, new_n18472);
xnor_4 g16124(new_n18456, new_n11203, new_n18473);
or_5   g16125(new_n18473, n11630, new_n18474);
xnor_4 g16126(new_n18455, n3164, new_n18475);
nor_5  g16127(new_n18475, n13453, new_n18476);
not_8  g16128(new_n18476, new_n18477);
xnor_4 g16129(new_n18475, new_n8268, new_n18478);
not_8  g16130(new_n15988, new_n18479);
nor_5  g16131(new_n18479, new_n8299, new_n18480);
not_8  g16132(new_n15989, new_n18481);
nor_5  g16133(new_n16002, new_n18481, new_n18482_1);
nor_5  g16134(new_n18482_1, new_n18480, new_n18483_1);
nand_5 g16135(new_n18483_1, new_n18478, new_n18484);
nand_5 g16136(new_n18484, new_n18477, new_n18485);
xnor_4 g16137(new_n18473, new_n8290, new_n18486);
nand_5 g16138(new_n18486, new_n18485, new_n18487);
nand_5 g16139(new_n18487, new_n18474, new_n18488);
nand_5 g16140(new_n18488, new_n18472, new_n18489);
nand_5 g16141(new_n18489, new_n18471, new_n18490);
nand_5 g16142(new_n18490, new_n18469, new_n18491);
nand_5 g16143(new_n18491, new_n18468, new_n18492);
nand_5 g16144(new_n18492, new_n18466, new_n18493);
nand_5 g16145(new_n18493, new_n18465, new_n18494);
xnor_4 g16146(new_n18494, new_n18463, new_n18495);
xnor_4 g16147(new_n18495, new_n18453, new_n18496_1);
not_8  g16148(new_n18496_1, new_n18497);
not_8  g16149(new_n18466, new_n18498);
xnor_4 g16150(new_n18492, new_n18498, new_n18499);
xnor_4 g16151(new_n18450, new_n18449, new_n18500);
nand_5 g16152(new_n18500, new_n18499, new_n18501);
not_8  g16153(new_n18500, new_n18502);
xnor_4 g16154(new_n18502, new_n18499, new_n18503);
not_8  g16155(new_n18469, new_n18504);
xnor_4 g16156(new_n18490, new_n18504, new_n18505);
not_8  g16157(new_n18428, new_n18506);
xnor_4 g16158(new_n18447, new_n18506, new_n18507);
nand_5 g16159(new_n18507, new_n18505, new_n18508);
not_8  g16160(new_n18507, new_n18509_1);
xnor_4 g16161(new_n18509_1, new_n18505, new_n18510);
not_8  g16162(new_n18472, new_n18511);
xnor_4 g16163(new_n18488, new_n18511, new_n18512);
xnor_4 g16164(new_n18445_1, new_n18431, new_n18513_1);
nand_5 g16165(new_n18513_1, new_n18512, new_n18514);
not_8  g16166(new_n18513_1, new_n18515_1);
xnor_4 g16167(new_n18515_1, new_n18512, new_n18516);
xnor_4 g16168(new_n18443, new_n18435, new_n18517);
not_8  g16169(new_n18517, new_n18518);
xnor_4 g16170(new_n18486, new_n18485, new_n18519);
not_8  g16171(new_n18519, new_n18520);
nand_5 g16172(new_n18520, new_n18518, new_n18521);
xnor_4 g16173(new_n18520, new_n18517, new_n18522);
xnor_4 g16174(new_n18483_1, new_n18478, new_n18523);
not_8  g16175(new_n18523, new_n18524);
xnor_4 g16176(new_n18441, new_n18438, new_n18525);
nand_5 g16177(new_n18525, new_n18524, new_n18526);
xnor_4 g16178(new_n18525, new_n18523, new_n18527);
nor_5  g16179(new_n16003, new_n10079, new_n18528);
not_8  g16180(new_n18528, new_n18529);
xnor_4 g16181(new_n16003, new_n10078, new_n18530);
nor_5  g16182(new_n16005, new_n10095, new_n18531);
xnor_4 g16183(new_n16005, new_n10095, new_n18532);
not_8  g16184(new_n16010, new_n18533);
nor_5  g16185(new_n18533, new_n10110, new_n18534);
nor_5  g16186(new_n16013_1, new_n10105, new_n18535);
not_8  g16187(new_n18535, new_n18536);
xnor_4 g16188(new_n18533, new_n10110, new_n18537_1);
nor_5  g16189(new_n18537_1, new_n18536, new_n18538);
nor_5  g16190(new_n18538, new_n18534, new_n18539);
nor_5  g16191(new_n18539, new_n18532, new_n18540);
nor_5  g16192(new_n18540, new_n18531, new_n18541);
nand_5 g16193(new_n18541, new_n18530, new_n18542);
nand_5 g16194(new_n18542, new_n18529, new_n18543);
nand_5 g16195(new_n18543, new_n18527, new_n18544);
nand_5 g16196(new_n18544, new_n18526, new_n18545);
nand_5 g16197(new_n18545, new_n18522, new_n18546);
nand_5 g16198(new_n18546, new_n18521, new_n18547);
nand_5 g16199(new_n18547, new_n18516, new_n18548);
nand_5 g16200(new_n18548, new_n18514, new_n18549);
nand_5 g16201(new_n18549, new_n18510, new_n18550);
nand_5 g16202(new_n18550, new_n18508, new_n18551);
nand_5 g16203(new_n18551, new_n18503, new_n18552);
nand_5 g16204(new_n18552, new_n18501, new_n18553);
xnor_4 g16205(new_n18553, new_n18497, n4221);
xnor_4 g16206(new_n11220_1, n18227, new_n18555);
nor_5  g16207(new_n11224, new_n5053, new_n18556);
not_8  g16208(new_n18556, new_n18557);
xnor_4 g16209(new_n11223_1, new_n5053, new_n18558_1);
nand_5 g16210(new_n11228, n11630, new_n18559);
nor_5  g16211(new_n11234_1, new_n8268, new_n18560);
not_8  g16212(new_n13777, new_n18561);
nor_5  g16213(new_n13781_1, new_n18561, new_n18562);
nor_5  g16214(new_n18562, new_n18560, new_n18563);
not_8  g16215(new_n18563, new_n18564);
xnor_4 g16216(new_n11228, new_n8290, new_n18565);
nand_5 g16217(new_n18565, new_n18564, new_n18566);
nand_5 g16218(new_n18566, new_n18559, new_n18567);
nand_5 g16219(new_n18567, new_n18558_1, new_n18568);
nand_5 g16220(new_n18568, new_n18557, new_n18569);
xnor_4 g16221(new_n18569, new_n18555, new_n18570);
xnor_4 g16222(new_n18570, new_n17236_1, new_n18571);
not_8  g16223(new_n9032_1, new_n18572_1);
xnor_4 g16224(new_n18567, new_n18558_1, new_n18573);
nor_5  g16225(new_n18573, new_n18572_1, new_n18574_1);
not_8  g16226(new_n18574_1, new_n18575);
xnor_4 g16227(new_n18573, new_n9032_1, new_n18576_1);
xnor_4 g16228(new_n18565, new_n18563, new_n18577);
nand_5 g16229(new_n18577, new_n9064, new_n18578_1);
xnor_4 g16230(new_n18577, new_n9065, new_n18579);
nand_5 g16231(new_n13782, new_n9071, new_n18580);
xnor_4 g16232(new_n13782, new_n17247, new_n18581);
nor_5  g16233(new_n9078, new_n13798_1, new_n18582_1);
not_8  g16234(new_n18582_1, new_n18583_1);
xnor_4 g16235(new_n9078, new_n6978, new_n18584_1);
nor_5  g16236(new_n9084, new_n7014, new_n18585);
xnor_4 g16237(new_n9082, new_n7014, new_n18586);
not_8  g16238(new_n18586, new_n18587);
nor_5  g16239(new_n9088, new_n7020, new_n18588);
nor_5  g16240(new_n9091, new_n7023, new_n18589);
not_8  g16241(new_n18589, new_n18590);
xnor_4 g16242(new_n9087, new_n7020, new_n18591);
not_8  g16243(new_n18591, new_n18592);
nor_5  g16244(new_n18592, new_n18590, new_n18593);
nor_5  g16245(new_n18593, new_n18588, new_n18594);
nor_5  g16246(new_n18594, new_n18587, new_n18595);
nor_5  g16247(new_n18595, new_n18585, new_n18596);
not_8  g16248(new_n18596, new_n18597);
nand_5 g16249(new_n18597, new_n18584_1, new_n18598);
nand_5 g16250(new_n18598, new_n18583_1, new_n18599);
nand_5 g16251(new_n18599, new_n18581, new_n18600);
nand_5 g16252(new_n18600, new_n18580, new_n18601);
nand_5 g16253(new_n18601, new_n18579, new_n18602);
nand_5 g16254(new_n18602, new_n18578_1, new_n18603);
nand_5 g16255(new_n18603, new_n18576_1, new_n18604);
nand_5 g16256(new_n18604, new_n18575, new_n18605);
xnor_4 g16257(new_n18605, new_n18571, n4224);
xor_4  g16258(new_n11382, new_n11381, n4231);
xnor_4 g16259(new_n15056, new_n13449, new_n18608);
nand_5 g16260(new_n15061, new_n12518, new_n18609);
nand_5 g16261(new_n17867, new_n17860, new_n18610_1);
nand_5 g16262(new_n18610_1, new_n18609, new_n18611);
xnor_4 g16263(new_n18611, new_n18608, new_n18612);
xnor_4 g16264(new_n18612, new_n5042, new_n18613);
nand_5 g16265(new_n17868, n647, new_n18614);
nand_5 g16266(new_n17877_1, new_n17869, new_n18615);
nand_5 g16267(new_n18615, new_n18614, new_n18616);
xnor_4 g16268(new_n18616, new_n18613, new_n18617);
xnor_4 g16269(new_n18617, new_n12637, new_n18618);
nand_5 g16270(new_n17878, new_n12641, new_n18619);
nand_5 g16271(new_n17888, new_n17879, new_n18620);
nand_5 g16272(new_n18620, new_n18619, new_n18621);
xnor_4 g16273(new_n18621, new_n18618, n4266);
xnor_4 g16274(new_n7347, new_n7318, n4340);
xnor_4 g16275(new_n17471, new_n6276_1, new_n18624);
xnor_4 g16276(new_n18624, new_n13897, new_n18625);
nor_5  g16277(new_n17472, new_n13904, new_n18626);
not_8  g16278(new_n18626, new_n18627);
nand_5 g16279(new_n17473, new_n17469, new_n18628);
nand_5 g16280(new_n18628, new_n18627, new_n18629);
xnor_4 g16281(new_n18629, new_n18625, new_n18630);
xnor_4 g16282(new_n18630, new_n5261, new_n18631);
and_5  g16283(new_n17474, new_n17467, new_n18632);
nor_5  g16284(new_n18632, new_n17466_1, new_n18633);
xnor_4 g16285(new_n18633, new_n18631, n4374);
xnor_4 g16286(new_n11900, new_n11847, n4401);
xnor_4 g16287(new_n13842, new_n13841, n4424);
nand_5 g16288(new_n11458, n1881, new_n18637);
not_8  g16289(n1881, new_n18638);
xnor_4 g16290(new_n11458, new_n18638, new_n18639);
nor_5  g16291(new_n11452, n5834, new_n18640);
xnor_4 g16292(new_n11452, n5834, new_n18641);
nand_5 g16293(new_n11445, n13851, new_n18642);
xnor_4 g16294(new_n11446, n13851, new_n18643);
nand_5 g16295(new_n11437, n24937, new_n18644);
nand_5 g16296(new_n17353, new_n17341, new_n18645);
nand_5 g16297(new_n18645, new_n18644, new_n18646);
nand_5 g16298(new_n18646, new_n18643, new_n18647);
nand_5 g16299(new_n18647, new_n18642, new_n18648);
nor_5  g16300(new_n18648, new_n18641, new_n18649_1);
nor_5  g16301(new_n18649_1, new_n18640, new_n18650);
nand_5 g16302(new_n18650, new_n18639, new_n18651);
nand_5 g16303(new_n18651, new_n18637, new_n18652);
nor_5  g16304(n8827, n4306, new_n18653_1);
not_8  g16305(new_n18653_1, new_n18654);
nand_5 g16306(new_n11457, new_n11454, new_n18655);
nand_5 g16307(new_n18655, new_n18654, new_n18656);
xnor_4 g16308(new_n18656, new_n18652, new_n18657);
xnor_4 g16309(new_n18657, new_n10618, new_n18658);
not_8  g16310(new_n10623, new_n18659);
not_8  g16311(new_n18639, new_n18660);
xnor_4 g16312(new_n18650, new_n18660, new_n18661);
nand_5 g16313(new_n18661, new_n18659, new_n18662);
xnor_4 g16314(new_n18661, new_n10623, new_n18663);
not_8  g16315(new_n10628_1, new_n18664);
xnor_4 g16316(new_n18648, new_n18641, new_n18665);
nand_5 g16317(new_n18665, new_n18664, new_n18666);
not_8  g16318(new_n18643, new_n18667);
xnor_4 g16319(new_n18646, new_n18667, new_n18668);
not_8  g16320(new_n18668, new_n18669);
nand_5 g16321(new_n18669, new_n10633, new_n18670);
xnor_4 g16322(new_n18668, new_n10633, new_n18671);
not_8  g16323(new_n17354, new_n18672);
nand_5 g16324(new_n18672, new_n10638, new_n18673);
nand_5 g16325(new_n17365, new_n17355, new_n18674);
nand_5 g16326(new_n18674, new_n18673, new_n18675);
nand_5 g16327(new_n18675, new_n18671, new_n18676);
nand_5 g16328(new_n18676, new_n18670, new_n18677);
not_8  g16329(new_n18677, new_n18678);
xnor_4 g16330(new_n18665, new_n10628_1, new_n18679_1);
nand_5 g16331(new_n18679_1, new_n18678, new_n18680);
nand_5 g16332(new_n18680, new_n18666, new_n18681);
nand_5 g16333(new_n18681, new_n18663, new_n18682);
nand_5 g16334(new_n18682, new_n18662, new_n18683);
xnor_4 g16335(new_n18683, new_n18658, n4432);
xnor_4 g16336(new_n15706, new_n15705, n4441);
nor_5  g16337(n27120, n23065, new_n18686);
nand_5 g16338(new_n18686, new_n9145, new_n18687);
nor_5  g16339(new_n18687, n25370, new_n18688);
nand_5 g16340(new_n18688, new_n9111, new_n18689);
nor_5  g16341(new_n18689, n19042, new_n18690_1);
nand_5 g16342(new_n18690_1, new_n7223, new_n18691);
xnor_4 g16343(new_n18691, new_n7219, new_n18692);
xnor_4 g16344(new_n18692, new_n17934, new_n18693_1);
not_8  g16345(new_n18693_1, new_n18694);
xnor_4 g16346(new_n18690_1, n1293, new_n18695);
nor_5  g16347(new_n18695, new_n17936, new_n18696);
xnor_4 g16348(new_n18695, new_n17936, new_n18697);
xnor_4 g16349(new_n18689, new_n7227, new_n18698);
nor_5  g16350(new_n18698, new_n17941, new_n18699);
xnor_4 g16351(new_n18688, n19472, new_n18700);
nor_5  g16352(new_n18700, new_n9136, new_n18701);
xnor_4 g16353(new_n18700, new_n9136, new_n18702);
not_8  g16354(new_n9139, new_n18703);
xnor_4 g16355(new_n18687, new_n9165, new_n18704);
not_8  g16356(new_n18704, new_n18705);
nor_5  g16357(new_n18705, new_n18703, new_n18706);
not_8  g16358(new_n18706, new_n18707);
xnor_4 g16359(new_n18705, new_n9139, new_n18708_1);
xnor_4 g16360(new_n18686, n24786, new_n18709);
nor_5  g16361(new_n18709, new_n9142, new_n18710);
xnor_4 g16362(new_n18709, new_n9142, new_n18711);
not_8  g16363(new_n9159, new_n18712);
xnor_4 g16364(n27120, new_n9148, new_n18713);
nor_5  g16365(new_n18713, new_n9154, new_n18714);
nor_5  g16366(new_n18714, new_n18712, new_n18715);
nor_5  g16367(new_n18715, new_n18711, new_n18716);
nor_5  g16368(new_n18716, new_n18710, new_n18717);
nand_5 g16369(new_n18717, new_n18708_1, new_n18718);
nand_5 g16370(new_n18718, new_n18707, new_n18719);
nor_5  g16371(new_n18719, new_n18702, new_n18720);
nor_5  g16372(new_n18720, new_n18701, new_n18721_1);
xnor_4 g16373(new_n18698, new_n17941, new_n18722);
nor_5  g16374(new_n18722, new_n18721_1, new_n18723);
nor_5  g16375(new_n18723, new_n18699, new_n18724);
nor_5  g16376(new_n18724, new_n18697, new_n18725_1);
nor_5  g16377(new_n18725_1, new_n18696, new_n18726);
xnor_4 g16378(new_n18726, new_n18694, new_n18727);
nand_5 g16379(new_n12837, new_n9291, new_n18728);
xnor_4 g16380(new_n18728, new_n9349, new_n18729);
xnor_4 g16381(new_n18729, new_n5620, new_n18730);
not_8  g16382(new_n12838, new_n18731);
nand_5 g16383(new_n18731, new_n5627, new_n18732);
nand_5 g16384(new_n12875_1, new_n12839, new_n18733);
nand_5 g16385(new_n18733, new_n18732, new_n18734);
xnor_4 g16386(new_n18734, new_n18730, new_n18735);
xnor_4 g16387(new_n18735, new_n18727, new_n18736);
not_8  g16388(new_n12876, new_n18737_1);
not_8  g16389(new_n18697, new_n18738);
xnor_4 g16390(new_n18724, new_n18738, new_n18739);
nand_5 g16391(new_n18739, new_n18737_1, new_n18740);
xnor_4 g16392(new_n18739, new_n12876, new_n18741);
xnor_4 g16393(new_n18722, new_n18721_1, new_n18742);
not_8  g16394(new_n18742, new_n18743);
nand_5 g16395(new_n18743, new_n12916, new_n18744);
xnor_4 g16396(new_n18742, new_n12916, new_n18745_1);
xnor_4 g16397(new_n18719, new_n18702, new_n18746);
not_8  g16398(new_n18746, new_n18747);
nor_5  g16399(new_n18747, new_n12920, new_n18748);
xnor_4 g16400(new_n18717, new_n18708_1, new_n18749);
nand_5 g16401(new_n18749, new_n12925, new_n18750);
xnor_4 g16402(new_n18749, new_n12926, new_n18751_1);
xnor_4 g16403(new_n18715, new_n18711, new_n18752);
not_8  g16404(new_n18752, new_n18753);
nor_5  g16405(new_n18753, new_n12936, new_n18754);
nor_5  g16406(new_n18752, new_n12931, new_n18755);
not_8  g16407(new_n9160, new_n18756);
xnor_4 g16408(new_n18713, new_n18756, new_n18757);
not_8  g16409(new_n18757, new_n18758);
nor_5  g16410(new_n18758, new_n12940, new_n18759);
not_8  g16411(new_n18759, new_n18760);
nor_5  g16412(new_n12943, new_n9180, new_n18761);
not_8  g16413(new_n18761, new_n18762);
xnor_4 g16414(new_n18757, new_n12940, new_n18763);
nand_5 g16415(new_n18763, new_n18762, new_n18764);
nand_5 g16416(new_n18764, new_n18760, new_n18765);
nor_5  g16417(new_n18765, new_n18755, new_n18766);
nor_5  g16418(new_n18766, new_n18754, new_n18767);
nand_5 g16419(new_n18767, new_n18751_1, new_n18768);
nand_5 g16420(new_n18768, new_n18750, new_n18769);
xnor_4 g16421(new_n18746, new_n12919, new_n18770);
nor_5  g16422(new_n18770, new_n18769, new_n18771);
nor_5  g16423(new_n18771, new_n18748, new_n18772);
nand_5 g16424(new_n18772, new_n18745_1, new_n18773);
nand_5 g16425(new_n18773, new_n18744, new_n18774);
nand_5 g16426(new_n18774, new_n18741, new_n18775);
nand_5 g16427(new_n18775, new_n18740, new_n18776);
xnor_4 g16428(new_n18776, new_n18736, n4451);
xnor_4 g16429(n25494, n6659, new_n18778);
or_5   g16430(new_n17002, n10117, new_n18779);
xnor_4 g16431(n23250, n10117, new_n18780_1);
or_5   g16432(n13460, new_n16920, new_n18781);
xnor_4 g16433(n13460, n11455, new_n18782_1);
or_5   g16434(n6104, new_n16923, new_n18783);
xnor_4 g16435(n6104, n3945, new_n18784);
or_5   g16436(new_n16926, n4119, new_n18785);
nand_5 g16437(new_n5450, new_n5427, new_n18786);
nand_5 g16438(new_n18786, new_n18785, new_n18787);
nand_5 g16439(new_n18787, new_n18784, new_n18788);
nand_5 g16440(new_n18788, new_n18783, new_n18789);
nand_5 g16441(new_n18789, new_n18782_1, new_n18790);
nand_5 g16442(new_n18790, new_n18781, new_n18791);
nand_5 g16443(new_n18791, new_n18780_1, new_n18792);
nand_5 g16444(new_n18792, new_n18779, new_n18793);
xnor_4 g16445(new_n18793, new_n18778, new_n18794);
xnor_4 g16446(new_n18794, new_n14005, new_n18795);
not_8  g16447(new_n18795, new_n18796);
not_8  g16448(new_n18780_1, new_n18797);
xnor_4 g16449(new_n18791, new_n18797, new_n18798);
nor_5  g16450(new_n18798, new_n14010, new_n18799);
xnor_4 g16451(new_n18798, new_n14010, new_n18800);
not_8  g16452(new_n18782_1, new_n18801);
xnor_4 g16453(new_n18789, new_n18801, new_n18802_1);
nor_5  g16454(new_n18802_1, new_n14015, new_n18803);
xnor_4 g16455(new_n18802_1, new_n14015, new_n18804);
not_8  g16456(new_n14021, new_n18805);
xnor_4 g16457(new_n18787, new_n18784, new_n18806);
nor_5  g16458(new_n18806, new_n18805, new_n18807);
not_8  g16459(new_n18807, new_n18808);
xnor_4 g16460(new_n18806, new_n14021, new_n18809);
nor_5  g16461(new_n5451_1, new_n5426, new_n18810);
not_8  g16462(new_n18810, new_n18811);
not_8  g16463(new_n5452, new_n18812);
nand_5 g16464(new_n5485_1, new_n18812, new_n18813);
nand_5 g16465(new_n18813, new_n18811, new_n18814);
nand_5 g16466(new_n18814, new_n18809, new_n18815);
nand_5 g16467(new_n18815, new_n18808, new_n18816);
nor_5  g16468(new_n18816, new_n18804, new_n18817);
nor_5  g16469(new_n18817, new_n18803, new_n18818);
nor_5  g16470(new_n18818, new_n18800, new_n18819);
nor_5  g16471(new_n18819, new_n18799, new_n18820);
xnor_4 g16472(new_n18820, new_n18796, n4476);
nor_5  g16473(new_n4175, n12398, new_n18822);
nand_5 g16474(new_n18822, new_n14812, new_n18823);
nor_5  g16475(new_n18823, n18452, new_n18824);
nand_5 g16476(new_n18824, new_n14804, new_n18825);
nor_5  g16477(new_n18825, n1831, new_n18826);
xnor_4 g16478(new_n18826, new_n6571, new_n18827);
xnor_4 g16479(new_n18825, new_n6478, new_n18828);
not_8  g16480(new_n18828, new_n18829);
nand_5 g16481(new_n18829, new_n6577, new_n18830_1);
not_8  g16482(new_n18830_1, new_n18831_1);
xnor_4 g16483(new_n18824, n13137, new_n18832);
nor_5  g16484(new_n18832, new_n6579, new_n18833);
xnor_4 g16485(new_n18832, new_n6579, new_n18834);
xnor_4 g16486(new_n18823, new_n14808, new_n18835);
nor_5  g16487(new_n18835, new_n6585, new_n18836);
xnor_4 g16488(new_n18835, new_n6585, new_n18837);
xnor_4 g16489(new_n18822, n21317, new_n18838);
not_8  g16490(new_n18838, new_n18839);
nor_5  g16491(new_n18839, new_n6591, new_n18840);
not_8  g16492(new_n18840, new_n18841);
xnor_4 g16493(new_n18838, new_n6591, new_n18842);
not_8  g16494(new_n4176_1, new_n18843_1);
nor_5  g16495(new_n4217, new_n18843_1, new_n18844);
not_8  g16496(new_n18844, new_n18845);
nand_5 g16497(new_n4255, new_n4218, new_n18846);
nand_5 g16498(new_n18846, new_n18845, new_n18847);
nand_5 g16499(new_n18847, new_n18842, new_n18848);
nand_5 g16500(new_n18848, new_n18841, new_n18849);
nor_5  g16501(new_n18849, new_n18837, new_n18850);
nor_5  g16502(new_n18850, new_n18836, new_n18851);
nor_5  g16503(new_n18851, new_n18834, new_n18852);
nor_5  g16504(new_n18852, new_n18833, new_n18853);
xnor_4 g16505(new_n18829, new_n6577, new_n18854);
nor_5  g16506(new_n18854, new_n18853, new_n18855);
nor_5  g16507(new_n18855, new_n18831_1, new_n18856);
xnor_4 g16508(new_n18856, new_n18827, new_n18857);
xnor_4 g16509(new_n18857, new_n12392, new_n18858_1);
not_8  g16510(new_n18854, new_n18859_1);
xnor_4 g16511(new_n18859_1, new_n18853, new_n18860);
nand_5 g16512(new_n18860, new_n12398_1, new_n18861);
xnor_4 g16513(new_n18860, new_n12453, new_n18862);
not_8  g16514(new_n18834, new_n18863);
xnor_4 g16515(new_n18851, new_n18863, new_n18864_1);
nand_5 g16516(new_n18864_1, new_n12402, new_n18865_1);
xnor_4 g16517(new_n18864_1, new_n12401, new_n18866);
not_8  g16518(new_n18849, new_n18867);
xnor_4 g16519(new_n18867, new_n18837, new_n18868);
nand_5 g16520(new_n18868, new_n12407, new_n18869);
xnor_4 g16521(new_n18868, new_n12406, new_n18870);
xnor_4 g16522(new_n18847, new_n18842, new_n18871);
nand_5 g16523(new_n18871, new_n12412, new_n18872);
xnor_4 g16524(new_n18871, new_n12411, new_n18873);
nand_5 g16525(new_n4256_1, new_n12416, new_n18874);
nand_5 g16526(new_n4291, new_n4257, new_n18875);
nand_5 g16527(new_n18875, new_n18874, new_n18876);
nand_5 g16528(new_n18876, new_n18873, new_n18877);
nand_5 g16529(new_n18877, new_n18872, new_n18878);
nand_5 g16530(new_n18878, new_n18870, new_n18879);
nand_5 g16531(new_n18879, new_n18869, new_n18880_1);
nand_5 g16532(new_n18880_1, new_n18866, new_n18881);
nand_5 g16533(new_n18881, new_n18865_1, new_n18882);
nand_5 g16534(new_n18882, new_n18862, new_n18883);
nand_5 g16535(new_n18883, new_n18861, new_n18884);
xnor_4 g16536(new_n18884, new_n18858_1, n4478);
xnor_4 g16537(new_n13284, new_n13246, n4529);
xnor_4 g16538(new_n6471, new_n6422, n4552);
xnor_4 g16539(new_n6467, new_n6434, n4595);
xnor_4 g16540(new_n15187, new_n15144, n4624);
nor_5  g16541(new_n18335, n2659, new_n18890);
xnor_4 g16542(new_n18890, n2858, new_n18891);
not_8  g16543(new_n18891, new_n18892);
nand_5 g16544(new_n18892, new_n4995, new_n18893);
xnor_4 g16545(new_n18891, new_n4995, new_n18894);
not_8  g16546(new_n18336, new_n18895);
nand_5 g16547(new_n18895, new_n4998, new_n18896);
nand_5 g16548(new_n18347, new_n18337, new_n18897);
nand_5 g16549(new_n18897, new_n18896, new_n18898);
nand_5 g16550(new_n18898, new_n18894, new_n18899);
nand_5 g16551(new_n18899, new_n18893, new_n18900);
nand_5 g16552(new_n18890, new_n5158_1, new_n18901_1);
xnor_4 g16553(new_n18901_1, new_n5220, new_n18902);
xnor_4 g16554(new_n18902, new_n4992, new_n18903);
xnor_4 g16555(new_n18903, new_n18900, new_n18904);
not_8  g16556(new_n18904, new_n18905);
nor_5  g16557(new_n18905, new_n8191, new_n18906);
not_8  g16558(new_n18906, new_n18907_1);
xnor_4 g16559(new_n18904, new_n8191, new_n18908);
xnor_4 g16560(new_n18898, new_n18894, new_n18909);
not_8  g16561(new_n18909, new_n18910);
nor_5  g16562(new_n18910, new_n8198, new_n18911);
not_8  g16563(new_n18911, new_n18912);
xnor_4 g16564(new_n18909, new_n8198, new_n18913);
not_8  g16565(new_n18348, new_n18914);
nor_5  g16566(new_n18914, new_n8202, new_n18915);
not_8  g16567(new_n18915, new_n18916);
not_8  g16568(new_n18352, new_n18917);
not_8  g16569(new_n18360, new_n18918);
nand_5 g16570(new_n18918, new_n18917, new_n18919_1);
nand_5 g16571(new_n18919_1, new_n18349, new_n18920);
nand_5 g16572(new_n18920, new_n18916, new_n18921);
nand_5 g16573(new_n18921, new_n18913, new_n18922);
nand_5 g16574(new_n18922, new_n18912, new_n18923);
nand_5 g16575(new_n18923, new_n18908, new_n18924);
nand_5 g16576(new_n18924, new_n18907_1, new_n18925);
nor_5  g16577(new_n18901_1, n3740, new_n18926_1);
not_8  g16578(new_n18926_1, new_n18927);
and_5  g16579(new_n18902, n3506, new_n18928);
nor_5  g16580(new_n18902, n3506, new_n18929);
nor_5  g16581(new_n18929, new_n18900, new_n18930);
nor_5  g16582(new_n18930, new_n18928, new_n18931);
nand_5 g16583(new_n18931, new_n18927, new_n18932);
xnor_4 g16584(new_n18932, new_n18925, new_n18933);
xnor_4 g16585(new_n18933, new_n8139_1, new_n18934);
xnor_4 g16586(new_n18934, new_n14512, new_n18935);
xnor_4 g16587(new_n18923, new_n18908, new_n18936);
nand_5 g16588(new_n18936, new_n8338, new_n18937);
not_8  g16589(new_n18913, new_n18938);
xnor_4 g16590(new_n18921, new_n18938, new_n18939);
not_8  g16591(new_n18939, new_n18940_1);
nand_5 g16592(new_n18940_1, new_n8344, new_n18941);
xnor_4 g16593(new_n18939, new_n8344, new_n18942);
not_8  g16594(new_n18362_1, new_n18943);
nand_5 g16595(new_n18943, new_n8349, new_n18944);
xnor_4 g16596(new_n18362_1, new_n8349, new_n18945_1);
nand_5 g16597(new_n18381, new_n8355, new_n18946);
xnor_4 g16598(new_n18380, new_n8355, new_n18947);
nor_5  g16599(new_n14107_1, new_n8361, new_n18948);
not_8  g16600(new_n14132, new_n18949);
nand_5 g16601(new_n18949, new_n8365, new_n18950);
nand_5 g16602(new_n18191, new_n18174, new_n18951);
nand_5 g16603(new_n18951, new_n18950, new_n18952);
xnor_4 g16604(new_n14107_1, new_n8361, new_n18953);
nor_5  g16605(new_n18953, new_n18952, new_n18954);
nor_5  g16606(new_n18954, new_n18948, new_n18955);
nand_5 g16607(new_n18955, new_n18947, new_n18956);
nand_5 g16608(new_n18956, new_n18946, new_n18957);
nand_5 g16609(new_n18957, new_n18945_1, new_n18958);
nand_5 g16610(new_n18958, new_n18944, new_n18959);
nand_5 g16611(new_n18959, new_n18942, new_n18960);
nand_5 g16612(new_n18960, new_n18941, new_n18961);
xnor_4 g16613(new_n8336, new_n8327, new_n18962_1);
xnor_4 g16614(new_n18936, new_n18962_1, new_n18963);
nand_5 g16615(new_n18963, new_n18961, new_n18964);
nand_5 g16616(new_n18964, new_n18937, new_n18965);
not_8  g16617(new_n18965, new_n18966);
xnor_4 g16618(new_n18966, new_n18935, n4646);
xnor_4 g16619(new_n15196, new_n15123, n4674);
xnor_4 g16620(n7057, n3480, new_n18969);
nor_5  g16621(new_n8110, n8381, new_n18970_1);
nor_5  g16622(n16722, new_n5296, new_n18971);
nor_5  g16623(n20235, new_n6097, new_n18972);
not_8  g16624(new_n18972, new_n18973);
nor_5  g16625(new_n5307, n11486, new_n18974);
not_8  g16626(new_n18974, new_n18975);
nor_5  g16627(new_n8119, n12495, new_n18976);
nand_5 g16628(new_n18976, new_n18975, new_n18977_1);
nand_5 g16629(new_n18977_1, new_n18973, new_n18978);
not_8  g16630(new_n18978, new_n18979);
nor_5  g16631(new_n18979, new_n18971, new_n18980);
nor_5  g16632(new_n18980, new_n18970_1, new_n18981);
xnor_4 g16633(new_n18981, new_n18969, new_n18982_1);
xnor_4 g16634(new_n18982_1, new_n3123, new_n18983);
xnor_4 g16635(n16722, n8381, new_n18984);
xnor_4 g16636(new_n18984, new_n18979, new_n18985);
not_8  g16637(new_n18985, new_n18986);
nor_5  g16638(new_n18986, new_n3130, new_n18987);
not_8  g16639(new_n18987, new_n18988);
xnor_4 g16640(new_n18986, new_n3129, new_n18989);
xnor_4 g16641(n13781, n12495, new_n18990);
nor_5  g16642(new_n18990, new_n3138, new_n18991);
nor_5  g16643(new_n18991, new_n3144, new_n18992);
xnor_4 g16644(new_n18991, new_n3144, new_n18993);
xnor_4 g16645(n20235, n11486, new_n18994);
xnor_4 g16646(new_n18994, new_n18976, new_n18995);
nor_5  g16647(new_n18995, new_n18993, new_n18996);
nor_5  g16648(new_n18996, new_n18992, new_n18997);
not_8  g16649(new_n18997, new_n18998);
nand_5 g16650(new_n18998, new_n18989, new_n18999_1);
nand_5 g16651(new_n18999_1, new_n18988, new_n19000);
xnor_4 g16652(new_n19000, new_n18983, n4693);
xnor_4 g16653(new_n11384, new_n11375_1, n4731);
nand_5 g16654(new_n6355, n8526, new_n19003);
nand_5 g16655(new_n6409, new_n6356_1, new_n19004);
nand_5 g16656(new_n19004, new_n19003, new_n19005_1);
or_5   g16657(n21784, n3582, new_n19006);
nand_5 g16658(new_n6354_1, new_n6310, new_n19007);
nand_5 g16659(new_n19007, new_n19006, new_n19008);
not_8  g16660(new_n19008, new_n19009);
nand_5 g16661(new_n19009, new_n19005_1, new_n19010);
not_8  g16662(new_n19010, new_n19011);
xnor_4 g16663(new_n19011, new_n16363, new_n19012);
xnor_4 g16664(new_n19009, new_n19005_1, new_n19013);
nand_5 g16665(new_n19013, new_n16367_1, new_n19014);
not_8  g16666(new_n19013, new_n19015);
xnor_4 g16667(new_n19015, new_n16367_1, new_n19016);
nand_5 g16668(new_n13708_1, new_n6410, new_n19017);
nand_5 g16669(new_n13751, new_n13709, new_n19018);
nand_5 g16670(new_n19018, new_n19017, new_n19019);
nand_5 g16671(new_n19019, new_n19016, new_n19020);
nand_5 g16672(new_n19020, new_n19014, new_n19021);
xnor_4 g16673(new_n19021, new_n19012, n4745);
xnor_4 g16674(new_n6608, new_n2575, new_n19023);
xnor_4 g16675(new_n19023, new_n10354, n4747);
xnor_4 g16676(new_n6060, new_n6059, n4766);
xnor_4 g16677(new_n14610, new_n14588, n4770);
xnor_4 g16678(new_n17503, new_n16594, n4777);
xnor_4 g16679(n17959, n6861, new_n19028);
nor_5  g16680(new_n3401, n7566, new_n19029);
not_8  g16681(new_n19029, new_n19030);
xnor_4 g16682(n19357, n7566, new_n19031);
nor_5  g16683(n7731, new_n3405, new_n19032);
xnor_4 g16684(n7731, n2328, new_n19033_1);
nor_5  g16685(n15053, new_n5760, new_n19034);
not_8  g16686(n15053, new_n19035);
nor_5  g16687(new_n19035, n12341, new_n19036);
nor_5  g16688(n25471, new_n5763, new_n19037);
not_8  g16689(n25471, new_n19038);
nor_5  g16690(new_n19038, n20986, new_n19039);
nand_5 g16691(new_n3486, n12384, new_n19040);
nor_5  g16692(new_n19040, new_n19039, new_n19041);
nor_5  g16693(new_n19041, new_n19037, new_n19042_1);
nor_5  g16694(new_n19042_1, new_n19036, new_n19043);
nor_5  g16695(new_n19043, new_n19034, new_n19044_1);
and_5  g16696(new_n19044_1, new_n19033_1, new_n19045);
nor_5  g16697(new_n19045, new_n19032, new_n19046);
not_8  g16698(new_n19046, new_n19047);
nand_5 g16699(new_n19047, new_n19031, new_n19048);
nand_5 g16700(new_n19048, new_n19030, new_n19049);
xnor_4 g16701(new_n19049, new_n19028, new_n19050);
nor_5  g16702(n20077, n6794, new_n19051);
nand_5 g16703(new_n19051, new_n2445, new_n19052);
nor_5  g16704(new_n19052, n8745, new_n19053);
nand_5 g16705(new_n19053, new_n2437, new_n19054);
xnor_4 g16706(new_n19054, new_n2433, new_n19055);
xnor_4 g16707(new_n19055, n11580, new_n19056);
xnor_4 g16708(new_n19053, n1777, new_n19057);
not_8  g16709(new_n19057, new_n19058);
nand_5 g16710(new_n19058, n15884, new_n19059);
xnor_4 g16711(new_n19057, n15884, new_n19060);
xnor_4 g16712(new_n19052, new_n2441, new_n19061);
not_8  g16713(new_n19061, new_n19062);
nand_5 g16714(new_n19062, n6356, new_n19063);
xnor_4 g16715(new_n19061, n6356, new_n19064);
xnor_4 g16716(new_n19051, n15636, new_n19065);
not_8  g16717(new_n19065, new_n19066);
nand_5 g16718(new_n19066, n27104, new_n19067);
xnor_4 g16719(new_n19065, n27104, new_n19068);
xnor_4 g16720(n20077, n6794, new_n19069);
nand_5 g16721(new_n19069, n27188, new_n19070);
nor_5  g16722(n6794, new_n9555, new_n19071);
xnor_4 g16723(new_n19069, new_n5882_1, new_n19072);
nand_5 g16724(new_n19072, new_n19071, new_n19073);
nand_5 g16725(new_n19073, new_n19070, new_n19074);
nand_5 g16726(new_n19074, new_n19068, new_n19075);
nand_5 g16727(new_n19075, new_n19067, new_n19076);
nand_5 g16728(new_n19076, new_n19064, new_n19077);
nand_5 g16729(new_n19077, new_n19063, new_n19078);
nand_5 g16730(new_n19078, new_n19060, new_n19079);
nand_5 g16731(new_n19079, new_n19059, new_n19080);
xnor_4 g16732(new_n19080, new_n19056, new_n19081_1);
xnor_4 g16733(new_n19081_1, new_n16899, new_n19082);
not_8  g16734(new_n16247_1, new_n19083);
xnor_4 g16735(new_n19078, new_n19060, new_n19084);
nand_5 g16736(new_n19084, new_n19083, new_n19085);
xnor_4 g16737(new_n19076, new_n19064, new_n19086);
nor_5  g16738(new_n19086, new_n16252, new_n19087);
xnor_4 g16739(new_n19086, new_n16252, new_n19088);
not_8  g16740(new_n5305, new_n19089);
xnor_4 g16741(new_n19074, new_n19068, new_n19090);
nand_5 g16742(new_n19090, new_n19089, new_n19091);
xnor_4 g16743(new_n19090, new_n5305, new_n19092);
xnor_4 g16744(new_n19072, new_n19071, new_n19093);
nand_5 g16745(new_n19093, new_n5342, new_n19094);
xnor_4 g16746(n6794, n6611, new_n19095);
nor_5  g16747(new_n19095, new_n5309, new_n19096);
xnor_4 g16748(new_n19093, new_n5314, new_n19097);
nand_5 g16749(new_n19097, new_n19096, new_n19098);
nand_5 g16750(new_n19098, new_n19094, new_n19099);
nand_5 g16751(new_n19099, new_n19092, new_n19100);
nand_5 g16752(new_n19100, new_n19091, new_n19101);
nor_5  g16753(new_n19101, new_n19088, new_n19102);
nor_5  g16754(new_n19102, new_n19087, new_n19103);
xnor_4 g16755(new_n19084, new_n16247_1, new_n19104);
nand_5 g16756(new_n19104, new_n19103, new_n19105);
nand_5 g16757(new_n19105, new_n19085, new_n19106);
xnor_4 g16758(new_n19106, new_n19082, new_n19107_1);
xnor_4 g16759(new_n19107_1, new_n19050, new_n19108);
xnor_4 g16760(new_n19046, new_n19031, new_n19109);
xnor_4 g16761(new_n19104, new_n19103, new_n19110);
not_8  g16762(new_n19110, new_n19111);
nor_5  g16763(new_n19111, new_n19109, new_n19112);
not_8  g16764(new_n19112, new_n19113);
xnor_4 g16765(new_n19110, new_n19109, new_n19114);
xnor_4 g16766(new_n19101, new_n19088, new_n19115);
xnor_4 g16767(new_n19044_1, new_n19033_1, new_n19116_1);
not_8  g16768(new_n19116_1, new_n19117);
nor_5  g16769(new_n19117, new_n19115, new_n19118);
not_8  g16770(new_n19118, new_n19119);
xnor_4 g16771(new_n19116_1, new_n19115, new_n19120);
xnor_4 g16772(new_n19099, new_n19092, new_n19121);
not_8  g16773(new_n19121, new_n19122);
xnor_4 g16774(n15053, n12341, new_n19123);
xnor_4 g16775(new_n19123, new_n19042_1, new_n19124);
not_8  g16776(new_n19124, new_n19125_1);
nor_5  g16777(new_n19125_1, new_n19122, new_n19126);
not_8  g16778(new_n19126, new_n19127);
xnor_4 g16779(new_n19125_1, new_n19121, new_n19128);
xnor_4 g16780(new_n19095, new_n5308, new_n19129);
not_8  g16781(new_n19129, new_n19130);
xnor_4 g16782(n16502, n12384, new_n19131);
nor_5  g16783(new_n19131, new_n19130, new_n19132);
xnor_4 g16784(n25471, n20986, new_n19133);
xnor_4 g16785(new_n19133, new_n19040, new_n19134);
not_8  g16786(new_n19134, new_n19135);
nor_5  g16787(new_n19135, new_n19132, new_n19136);
xnor_4 g16788(new_n19097, new_n19096, new_n19137);
xnor_4 g16789(new_n19134, new_n19132, new_n19138);
nand_5 g16790(new_n19138, new_n19137, new_n19139);
not_8  g16791(new_n19139, new_n19140);
nor_5  g16792(new_n19140, new_n19136, new_n19141_1);
not_8  g16793(new_n19141_1, new_n19142);
nand_5 g16794(new_n19142, new_n19128, new_n19143);
nand_5 g16795(new_n19143, new_n19127, new_n19144_1);
nand_5 g16796(new_n19144_1, new_n19120, new_n19145);
nand_5 g16797(new_n19145, new_n19119, new_n19146);
nand_5 g16798(new_n19146, new_n19114, new_n19147);
nand_5 g16799(new_n19147, new_n19113, new_n19148);
xor_4  g16800(new_n19148, new_n19108, n4785);
xnor_4 g16801(new_n14946, new_n14912, n4804);
xnor_4 g16802(new_n16604, new_n16584_1, n4810);
or_5   g16803(new_n18454, n18105, new_n19152);
nand_5 g16804(new_n9713, new_n9671, new_n19153);
nand_5 g16805(new_n19153, new_n19152, new_n19154);
not_8  g16806(new_n19154, new_n19155);
nand_5 g16807(new_n11460, new_n16342, new_n19156);
nand_5 g16808(new_n11514, new_n11461, new_n19157);
nand_5 g16809(new_n19157, new_n19156, new_n19158);
nand_5 g16810(new_n11459, new_n11453, new_n19159);
not_8  g16811(new_n18656, new_n19160);
nand_5 g16812(new_n19160, new_n19159, new_n19161);
nor_5  g16813(new_n19159, new_n18654, new_n19162);
not_8  g16814(new_n19162, new_n19163_1);
nand_5 g16815(new_n19163_1, new_n19161, new_n19164_1);
xnor_4 g16816(new_n19164_1, new_n8528, new_n19165);
xnor_4 g16817(new_n19165, new_n19158, new_n19166);
nand_5 g16818(new_n19166, new_n19155, new_n19167);
xnor_4 g16819(new_n19166, new_n19154, new_n19168);
not_8  g16820(new_n9714, new_n19169);
nand_5 g16821(new_n11515_1, new_n19169, new_n19170);
nand_5 g16822(new_n11570, new_n11516, new_n19171);
nand_5 g16823(new_n19171, new_n19170, new_n19172);
nand_5 g16824(new_n19172, new_n19168, new_n19173);
nand_5 g16825(new_n19173, new_n19167, new_n19174_1);
not_8  g16826(new_n19174_1, new_n19175);
not_8  g16827(new_n19158, new_n19176_1);
nand_5 g16828(new_n19164_1, new_n8528, new_n19177);
nand_5 g16829(new_n19177, new_n19176_1, new_n19178);
nor_5  g16830(new_n19164_1, new_n8528, new_n19179);
nor_5  g16831(new_n19179, new_n19162, new_n19180);
nand_5 g16832(new_n19180, new_n19178, new_n19181);
nand_5 g16833(new_n19181, new_n19175, n4814);
xnor_4 g16834(new_n17265, new_n17264, n4850);
xnor_4 g16835(new_n18158, new_n18114, n4891);
xnor_4 g16836(new_n18327, new_n18304_1, n4925);
xnor_4 g16837(new_n17271, new_n17248, n4947);
xnor_4 g16838(new_n10007, new_n10006, n4952);
xnor_4 g16839(n25068, n6790, new_n19188);
nor_5  g16840(n22879, new_n8488, new_n19189);
xnor_4 g16841(n22879, n2331, new_n19190);
not_8  g16842(new_n19190, new_n19191);
nor_5  g16843(new_n8493, n2117, new_n19192);
xnor_4 g16844(n22631, n2117, new_n19193);
not_8  g16845(new_n19193, new_n19194);
nor_5  g16846(n16743, new_n10475, new_n19195);
not_8  g16847(new_n19195, new_n19196_1);
nor_5  g16848(new_n8495, n5882, new_n19197);
not_8  g16849(new_n19197, new_n19198);
nor_5  g16850(n15258, new_n10485, new_n19199);
not_8  g16851(new_n19199, new_n19200);
nor_5  g16852(new_n10482, n4588, new_n19201);
nor_5  g16853(new_n8501, n11775, new_n19202_1);
not_8  g16854(new_n19202_1, new_n19203);
nand_5 g16855(new_n19203, new_n19201, new_n19204);
nand_5 g16856(new_n19204, new_n19200, new_n19205);
nand_5 g16857(new_n19205, new_n19198, new_n19206);
nand_5 g16858(new_n19206, new_n19196_1, new_n19207);
nor_5  g16859(new_n19207, new_n19194, new_n19208);
nor_5  g16860(new_n19208, new_n19192, new_n19209);
nor_5  g16861(new_n19209, new_n19191, new_n19210);
nor_5  g16862(new_n19210, new_n19189, new_n19211);
xnor_4 g16863(new_n19211, new_n19188, new_n19212);
xnor_4 g16864(new_n19212, new_n16193, new_n19213);
xnor_4 g16865(new_n19209, new_n19190, new_n19214);
nor_5  g16866(new_n19214, new_n16199, new_n19215);
xnor_4 g16867(new_n19214, new_n16199, new_n19216);
xnor_4 g16868(new_n19207, new_n19193, new_n19217);
nor_5  g16869(new_n19217, new_n16205, new_n19218);
xnor_4 g16870(new_n19217, new_n16205, new_n19219);
xnor_4 g16871(n16743, n5882, new_n19220_1);
xnor_4 g16872(new_n19220_1, new_n19205, new_n19221_1);
not_8  g16873(new_n19221_1, new_n19222);
nor_5  g16874(new_n19222, new_n16210, new_n19223_1);
not_8  g16875(new_n19223_1, new_n19224_1);
xnor_4 g16876(new_n19221_1, new_n16210, new_n19225);
xnor_4 g16877(n15258, n11775, new_n19226);
xnor_4 g16878(new_n19226, new_n19201, new_n19227);
nand_5 g16879(new_n19227, new_n16214, new_n19228_1);
nor_5  g16880(new_n15983, new_n16216, new_n19229);
not_8  g16881(new_n19228_1, new_n19230);
nor_5  g16882(new_n19227, new_n16214, new_n19231);
nor_5  g16883(new_n19231, new_n19230, new_n19232);
nand_5 g16884(new_n19232, new_n19229, new_n19233_1);
nand_5 g16885(new_n19233_1, new_n19228_1, new_n19234_1);
nand_5 g16886(new_n19234_1, new_n19225, new_n19235);
nand_5 g16887(new_n19235, new_n19224_1, new_n19236);
nor_5  g16888(new_n19236, new_n19219, new_n19237);
nor_5  g16889(new_n19237, new_n19218, new_n19238);
nor_5  g16890(new_n19238, new_n19216, new_n19239);
nor_5  g16891(new_n19239, new_n19215, new_n19240);
xnor_4 g16892(new_n19240, new_n19213, new_n19241);
xnor_4 g16893(new_n19241, new_n16120, new_n19242);
not_8  g16894(new_n16125, new_n19243);
not_8  g16895(new_n19216, new_n19244_1);
xnor_4 g16896(new_n19238, new_n19244_1, new_n19245);
nand_5 g16897(new_n19245, new_n19243, new_n19246);
xnor_4 g16898(new_n19245, new_n16125, new_n19247);
xnor_4 g16899(new_n19236, new_n19219, new_n19248);
not_8  g16900(new_n19248, new_n19249);
nand_5 g16901(new_n19249, new_n16129, new_n19250);
xnor_4 g16902(new_n19248, new_n16129, new_n19251);
xnor_4 g16903(new_n19234_1, new_n19225, new_n19252);
not_8  g16904(new_n19252, new_n19253);
nor_5  g16905(new_n19253, new_n14454, new_n19254);
not_8  g16906(new_n19254, new_n19255);
xnor_4 g16907(new_n19252, new_n14454, new_n19256);
not_8  g16908(new_n15984, new_n19257);
nor_5  g16909(new_n19257, new_n10587, new_n19258);
nor_5  g16910(new_n19258, new_n14464_1, new_n19259);
xnor_4 g16911(new_n19258, new_n14464_1, new_n19260);
xnor_4 g16912(new_n19232, new_n19229, new_n19261);
not_8  g16913(new_n19261, new_n19262);
nor_5  g16914(new_n19262, new_n19260, new_n19263);
nor_5  g16915(new_n19263, new_n19259, new_n19264);
not_8  g16916(new_n19264, new_n19265);
nand_5 g16917(new_n19265, new_n19256, new_n19266);
nand_5 g16918(new_n19266, new_n19255, new_n19267);
nand_5 g16919(new_n19267, new_n19251, new_n19268);
nand_5 g16920(new_n19268, new_n19250, new_n19269);
nand_5 g16921(new_n19269, new_n19247, new_n19270_1);
nand_5 g16922(new_n19270_1, new_n19246, new_n19271);
xnor_4 g16923(new_n19271, new_n19242, n4966);
xnor_4 g16924(new_n18679_1, new_n18678, n4972);
nor_5  g16925(new_n7994, n23895, new_n19274);
xnor_4 g16926(new_n7994, new_n5737, new_n19275);
not_8  g16927(new_n19275, new_n19276);
nand_5 g16928(new_n7999_1, n17351, new_n19277);
xnor_4 g16929(new_n7998, n17351, new_n19278);
nand_5 g16930(new_n8005, n11736, new_n19279);
nand_5 g16931(new_n17967, new_n17955, new_n19280);
nand_5 g16932(new_n19280, new_n19279, new_n19281);
nand_5 g16933(new_n19281, new_n19278, new_n19282_1);
nand_5 g16934(new_n19282_1, new_n19277, new_n19283);
nor_5  g16935(new_n19283, new_n19276, new_n19284);
nor_5  g16936(new_n19284, new_n19274, new_n19285);
nand_5 g16937(new_n19285, new_n7986, new_n19286);
not_8  g16938(new_n19286, new_n19287);
nor_5  g16939(new_n17918, n2289, new_n19288);
nand_5 g16940(new_n19288, new_n7114, new_n19289);
xnor_4 g16941(new_n19289, new_n7886, new_n19290);
xnor_4 g16942(new_n19290, new_n13864, new_n19291);
xnor_4 g16943(new_n19288, n23697, new_n19292);
and_5  g16944(new_n19292, n337, new_n19293);
nor_5  g16945(new_n19292, n337, new_n19294);
not_8  g16946(new_n17919, new_n19295);
nor_5  g16947(new_n19295, new_n3390_1, new_n19296);
nor_5  g16948(new_n17919, n3228, new_n19297);
nor_5  g16949(new_n17933, new_n19297, new_n19298);
nor_5  g16950(new_n19298, new_n19296, new_n19299);
nor_5  g16951(new_n19299, new_n19294, new_n19300);
nor_5  g16952(new_n19300, new_n19293, new_n19301);
xnor_4 g16953(new_n19301, new_n19291, new_n19302);
nor_5  g16954(new_n19302, n25972, new_n19303);
not_8  g16955(new_n19303, new_n19304);
xnor_4 g16956(new_n19302, new_n12752, new_n19305);
xnor_4 g16957(new_n19292, new_n3387, new_n19306);
xnor_4 g16958(new_n19306, new_n19299, new_n19307);
nor_5  g16959(new_n19307, n21915, new_n19308);
not_8  g16960(new_n19308, new_n19309);
nor_5  g16961(new_n17934, n13775, new_n19310);
not_8  g16962(new_n19310, new_n19311);
nand_5 g16963(new_n17953, new_n17935, new_n19312);
nand_5 g16964(new_n19312, new_n19311, new_n19313);
xnor_4 g16965(new_n19307, new_n9196, new_n19314_1);
nand_5 g16966(new_n19314_1, new_n19313, new_n19315_1);
nand_5 g16967(new_n19315_1, new_n19309, new_n19316);
nand_5 g16968(new_n19316, new_n19305, new_n19317);
nand_5 g16969(new_n19317, new_n19304, new_n19318);
nor_5  g16970(new_n19289, n2978, new_n19319);
not_8  g16971(new_n19319, new_n19320);
not_8  g16972(new_n19290, new_n19321);
nor_5  g16973(new_n19321, new_n13864, new_n19322);
nor_5  g16974(new_n19290, n7593, new_n19323_1);
nor_5  g16975(new_n19301, new_n19323_1, new_n19324);
nor_5  g16976(new_n19324, new_n19322, new_n19325);
nand_5 g16977(new_n19325, new_n19320, new_n19326);
nor_5  g16978(new_n19326, new_n19318, new_n19327_1);
xnor_4 g16979(new_n19285, new_n7989, new_n19328);
not_8  g16980(new_n19328, new_n19329);
xnor_4 g16981(new_n19326, new_n19318, new_n19330);
nand_5 g16982(new_n19330, new_n19329, new_n19331);
xnor_4 g16983(new_n19330, new_n19328, new_n19332);
xnor_4 g16984(new_n19283, new_n19275, new_n19333_1);
not_8  g16985(new_n19305, new_n19334);
xnor_4 g16986(new_n19316, new_n19334, new_n19335);
nor_5  g16987(new_n19335, new_n19333_1, new_n19336);
xnor_4 g16988(new_n19335, new_n19333_1, new_n19337);
xnor_4 g16989(new_n19281, new_n19278, new_n19338);
not_8  g16990(new_n19338, new_n19339);
xnor_4 g16991(new_n19314_1, new_n19313, new_n19340);
nand_5 g16992(new_n19340, new_n19339, new_n19341);
not_8  g16993(new_n19341, new_n19342);
not_8  g16994(new_n17954_1, new_n19343);
nand_5 g16995(new_n17968_1, new_n19343, new_n19344);
nand_5 g16996(new_n17994, new_n17969, new_n19345);
nand_5 g16997(new_n19345, new_n19344, new_n19346);
xnor_4 g16998(new_n19340, new_n19339, new_n19347);
nor_5  g16999(new_n19347, new_n19346, new_n19348_1);
nor_5  g17000(new_n19348_1, new_n19342, new_n19349);
nor_5  g17001(new_n19349, new_n19337, new_n19350);
nor_5  g17002(new_n19350, new_n19336, new_n19351);
nand_5 g17003(new_n19351, new_n19332, new_n19352);
nand_5 g17004(new_n19352, new_n19331, new_n19353);
xnor_4 g17005(new_n19353, new_n19327_1, new_n19354_1);
xnor_4 g17006(new_n19354_1, new_n19287, n5011);
or_5   g17007(new_n10741, n2944, new_n19356);
xnor_4 g17008(n11220, n2944, new_n19357_1);
not_8  g17009(n22379, new_n19358);
or_5   g17010(new_n19358, n767, new_n19359);
nand_5 g17011(new_n2939, new_n2899, new_n19360);
nand_5 g17012(new_n19360, new_n19359, new_n19361_1);
nand_5 g17013(new_n19361_1, new_n19357_1, new_n19362);
nand_5 g17014(new_n19362, new_n19356, new_n19363);
not_8  g17015(new_n19363, new_n19364);
or_5   g17016(new_n9530, new_n12514, new_n19365);
not_8  g17017(new_n19365, new_n19366);
nor_5  g17018(n16544, n2160, new_n19367_1);
or_5   g17019(n10763, n6814, new_n19368);
nand_5 g17020(new_n2984, new_n2942, new_n19369);
nand_5 g17021(new_n19369, new_n19368, new_n19370);
nor_5  g17022(new_n19370, new_n19367_1, new_n19371);
nor_5  g17023(new_n19371, new_n19366, new_n19372);
nor_5  g17024(new_n19372, new_n16057, new_n19373);
xnor_4 g17025(new_n19372, new_n16054, new_n19374);
not_8  g17026(new_n19374, new_n19375);
xnor_4 g17027(n16544, new_n12514, new_n19376);
xnor_4 g17028(new_n19376, new_n19370, new_n19377);
not_8  g17029(new_n19377, new_n19378);
nor_5  g17030(new_n19378, new_n16026, new_n19379);
xnor_4 g17031(new_n19377, new_n16026, new_n19380);
not_8  g17032(new_n19380, new_n19381);
not_8  g17033(new_n2985_1, new_n19382);
nor_5  g17034(new_n3032, new_n19382, new_n19383);
not_8  g17035(new_n3033, new_n19384);
nor_5  g17036(new_n3099, new_n19384, new_n19385_1);
nor_5  g17037(new_n19385_1, new_n19383, new_n19386);
nor_5  g17038(new_n19386, new_n19381, new_n19387);
nor_5  g17039(new_n19387, new_n19379, new_n19388);
nor_5  g17040(new_n19388, new_n19375, new_n19389_1);
nor_5  g17041(new_n19389_1, new_n19373, new_n19390);
not_8  g17042(new_n19390, new_n19391);
nand_5 g17043(new_n19391, new_n19364, new_n19392);
xnor_4 g17044(new_n19388, new_n19374, new_n19393);
not_8  g17045(new_n19393, new_n19394);
nand_5 g17046(new_n19394, new_n19363, new_n19395);
nand_5 g17047(new_n19393, new_n19364, new_n19396);
xnor_4 g17048(new_n19361_1, new_n19357_1, new_n19397);
xnor_4 g17049(new_n19386, new_n19380, new_n19398);
not_8  g17050(new_n19398, new_n19399);
nand_5 g17051(new_n19399, new_n19397, new_n19400);
xnor_4 g17052(new_n19398, new_n19397, new_n19401_1);
not_8  g17053(new_n3100, new_n19402);
nand_5 g17054(new_n19402, new_n2940, new_n19403);
nand_5 g17055(new_n3161_1, new_n3101, new_n19404);
nand_5 g17056(new_n19404, new_n19403, new_n19405);
nand_5 g17057(new_n19405, new_n19401_1, new_n19406);
nand_5 g17058(new_n19406, new_n19400, new_n19407);
nand_5 g17059(new_n19407, new_n19396, new_n19408);
nand_5 g17060(new_n19408, new_n19395, new_n19409);
nand_5 g17061(new_n19409, new_n19392, new_n19410);
nand_5 g17062(new_n19390, new_n19363, new_n19411);
nand_5 g17063(new_n19411, new_n19408, new_n19412);
nand_5 g17064(new_n19412, new_n19410, new_n19413);
not_8  g17065(new_n19413, n5020);
nor_5  g17066(n13781, n11486, new_n19415);
nand_5 g17067(new_n19415, new_n8110, new_n19416);
nor_5  g17068(new_n19416, n3480, new_n19417);
xnor_4 g17069(new_n19417, n3018, new_n19418);
xnor_4 g17070(new_n19418, new_n3056, new_n19419);
xnor_4 g17071(new_n19416, new_n2398, new_n19420);
nor_5  g17072(new_n19420, new_n3063, new_n19421);
xnor_4 g17073(new_n19420, new_n3063, new_n19422);
xnor_4 g17074(new_n19415, n16722, new_n19423);
nor_5  g17075(new_n19423, new_n3068, new_n19424_1);
xnor_4 g17076(new_n19423, new_n3068, new_n19425);
xnor_4 g17077(n13781, new_n6097, new_n19426);
nor_5  g17078(new_n19426, new_n3074, new_n19427);
nor_5  g17079(new_n3080, n13781, new_n19428);
not_8  g17080(new_n19428, new_n19429);
xnor_4 g17081(new_n19426, new_n3074, new_n19430);
nor_5  g17082(new_n19430, new_n19429, new_n19431);
nor_5  g17083(new_n19431, new_n19427, new_n19432);
nor_5  g17084(new_n19432, new_n19425, new_n19433);
nor_5  g17085(new_n19433, new_n19424_1, new_n19434);
nor_5  g17086(new_n19434, new_n19422, new_n19435);
nor_5  g17087(new_n19435, new_n19421, new_n19436);
xnor_4 g17088(new_n19436, new_n19419, new_n19437);
xnor_4 g17089(new_n19437, new_n7312, new_n19438);
xnor_4 g17090(new_n19434, new_n19422, new_n19439);
nor_5  g17091(new_n19439, new_n7320, new_n19440);
not_8  g17092(new_n19440, new_n19441);
xnor_4 g17093(new_n19439, new_n7319, new_n19442);
not_8  g17094(new_n19442, new_n19443);
xnor_4 g17095(new_n19432, new_n19425, new_n19444);
nor_5  g17096(new_n19444, new_n7327, new_n19445);
xnor_4 g17097(new_n19430, new_n19428, new_n19446);
not_8  g17098(new_n19446, new_n19447);
nor_5  g17099(new_n19447, new_n7339_1, new_n19448);
xnor_4 g17100(new_n3079, n13781, new_n19449);
nor_5  g17101(new_n19449, new_n7335_1, new_n19450_1);
xnor_4 g17102(new_n19446, new_n7339_1, new_n19451);
not_8  g17103(new_n19451, new_n19452);
nor_5  g17104(new_n19452, new_n19450_1, new_n19453);
nor_5  g17105(new_n19453, new_n19448, new_n19454_1);
xnor_4 g17106(new_n19444, new_n7326, new_n19455);
not_8  g17107(new_n19455, new_n19456);
nor_5  g17108(new_n19456, new_n19454_1, new_n19457);
nor_5  g17109(new_n19457, new_n19445, new_n19458_1);
nor_5  g17110(new_n19458_1, new_n19443, new_n19459);
not_8  g17111(new_n19459, new_n19460);
nand_5 g17112(new_n19460, new_n19441, new_n19461);
xnor_4 g17113(new_n19461, new_n19438, n5024);
xnor_4 g17114(new_n3867, new_n3833, n5046);
xnor_4 g17115(new_n6171_1, new_n3947, n5062);
xnor_4 g17116(new_n13339, new_n13310, n5064);
xnor_4 g17117(n12495, new_n7384, new_n19466);
xnor_4 g17118(new_n19466, new_n2383, new_n19467_1);
xnor_4 g17119(n9251, n7428, new_n19468);
nor_5  g17120(new_n19468, new_n19467_1, new_n19469);
nor_5  g17121(new_n3650, n7428, new_n19470);
xnor_4 g17122(n20138, n10372, new_n19471);
xnor_4 g17123(new_n19471, new_n19470, new_n19472_1);
xnor_4 g17124(new_n19472_1, new_n19469, new_n19473);
nor_5  g17125(new_n19466, new_n2382, new_n19474);
nand_5 g17126(n12495, n11479, new_n19475);
xnor_4 g17127(n20235, n8259, new_n19476);
xnor_4 g17128(new_n19476, new_n19475, new_n19477_1);
xnor_4 g17129(new_n19477_1, new_n2387_1, new_n19478);
xnor_4 g17130(new_n19478, new_n19474, new_n19479);
not_8  g17131(new_n19479, new_n19480);
xnor_4 g17132(new_n19480, new_n19473, n5082);
xnor_4 g17133(new_n14601, new_n14600, n5120);
xnor_4 g17134(new_n15848, new_n15839, n5158);
xnor_4 g17135(new_n17269, new_n17254, n5168);
not_8  g17136(n6659, new_n19485);
xnor_4 g17137(new_n18398, new_n19485, new_n19486);
not_8  g17138(new_n19486, new_n19487);
nand_5 g17139(new_n18421, new_n17002, new_n19488);
xnor_4 g17140(new_n15236, new_n17002, new_n19489);
nand_5 g17141(new_n15238, new_n16920, new_n19490);
xnor_4 g17142(new_n15238, n11455, new_n19491);
not_8  g17143(new_n15241_1, new_n19492);
nand_5 g17144(new_n19492, new_n16923, new_n19493);
xnor_4 g17145(new_n15241_1, new_n16923, new_n19494_1);
nor_5  g17146(new_n15244, new_n16926, new_n19495);
xnor_4 g17147(new_n15244, n5255, new_n19496_1);
not_8  g17148(new_n19496_1, new_n19497);
nor_5  g17149(new_n15249, new_n5428, new_n19498);
not_8  g17150(new_n16265, new_n19499);
nor_5  g17151(new_n16281, new_n19499, new_n19500);
nor_5  g17152(new_n19500, new_n19498, new_n19501);
nor_5  g17153(new_n19501, new_n19497, new_n19502);
nor_5  g17154(new_n19502, new_n19495, new_n19503);
nand_5 g17155(new_n19503, new_n19494_1, new_n19504);
nand_5 g17156(new_n19504, new_n19493, new_n19505);
nand_5 g17157(new_n19505, new_n19491, new_n19506);
nand_5 g17158(new_n19506, new_n19490, new_n19507);
nand_5 g17159(new_n19507, new_n19489, new_n19508);
nand_5 g17160(new_n19508, new_n19488, new_n19509);
xnor_4 g17161(new_n19509, new_n19487, new_n19510);
xnor_4 g17162(new_n19510, new_n16917, new_n19511);
not_8  g17163(new_n19489, new_n19512);
xnor_4 g17164(new_n19507, new_n19512, new_n19513);
nand_5 g17165(new_n19513, new_n17012, new_n19514_1);
xnor_4 g17166(new_n19513, new_n17011, new_n19515_1);
xnor_4 g17167(new_n19505, new_n19491, new_n19516);
not_8  g17168(new_n19516, new_n19517);
nand_5 g17169(new_n19517, new_n17018, new_n19518);
xnor_4 g17170(new_n19516, new_n17018, new_n19519);
xnor_4 g17171(new_n19503, new_n19494_1, new_n19520);
not_8  g17172(new_n19520, new_n19521);
nand_5 g17173(new_n19521, new_n17024, new_n19522);
xnor_4 g17174(new_n19520, new_n17024, new_n19523_1);
xnor_4 g17175(new_n19501, new_n19496_1, new_n19524);
not_8  g17176(new_n19524, new_n19525);
nand_5 g17177(new_n19525, new_n17030, new_n19526);
xnor_4 g17178(new_n19524, new_n17030, new_n19527);
not_8  g17179(new_n16282, new_n19528);
nand_5 g17180(new_n19528, new_n16264, new_n19529);
nand_5 g17181(new_n16306, new_n16283, new_n19530);
nand_5 g17182(new_n19530, new_n19529, new_n19531_1);
nand_5 g17183(new_n19531_1, new_n19527, new_n19532);
nand_5 g17184(new_n19532, new_n19526, new_n19533);
nand_5 g17185(new_n19533, new_n19523_1, new_n19534);
nand_5 g17186(new_n19534, new_n19522, new_n19535);
nand_5 g17187(new_n19535, new_n19519, new_n19536);
nand_5 g17188(new_n19536, new_n19518, new_n19537);
nand_5 g17189(new_n19537, new_n19515_1, new_n19538);
nand_5 g17190(new_n19538, new_n19514_1, new_n19539_1);
xnor_4 g17191(new_n19539_1, new_n19511, n5184);
nor_5  g17192(new_n4732, new_n4610, new_n19541);
nand_5 g17193(new_n4819, new_n19541, new_n19542);
not_8  g17194(new_n4610, new_n19543);
nor_5  g17195(new_n4731_1, new_n19543, new_n19544);
not_8  g17196(new_n4819, new_n19545);
nand_5 g17197(new_n19545, new_n19544, new_n19546);
nand_5 g17198(new_n19546, new_n19542, n5228);
or_5   g17199(n25494, new_n8720, new_n19548);
nand_5 g17200(new_n12010, new_n11994, new_n19549);
nand_5 g17201(new_n19549, new_n19548, new_n19550);
not_8  g17202(new_n19550, new_n19551);
xnor_4 g17203(new_n19551, new_n7631, new_n19552);
nand_5 g17204(new_n12011_1, new_n7542, new_n19553);
xnor_4 g17205(new_n12011_1, new_n7541, new_n19554);
nand_5 g17206(new_n12030, new_n7547, new_n19555);
nand_5 g17207(new_n13341, new_n13308, new_n19556);
nand_5 g17208(new_n19556, new_n19555, new_n19557);
nand_5 g17209(new_n19557, new_n19554, new_n19558);
nand_5 g17210(new_n19558, new_n19553, new_n19559);
xnor_4 g17211(new_n19559, new_n19552, n5256);
xnor_4 g17212(new_n7031, new_n7019, n5265);
xnor_4 g17213(new_n18160, new_n18108, n5273);
xnor_4 g17214(n20946, n2289, new_n19563);
or_5   g17215(new_n2430, n1112, new_n19564);
xnor_4 g17216(n7751, n1112, new_n19565);
or_5   g17217(new_n2434, n20179, new_n19566);
not_8  g17218(new_n17792, new_n19567);
nand_5 g17219(new_n19567, new_n17775, new_n19568);
nand_5 g17220(new_n19568, new_n19566, new_n19569);
nand_5 g17221(new_n19569, new_n19565, new_n19570_1);
nand_5 g17222(new_n19570_1, new_n19564, new_n19571);
xnor_4 g17223(new_n19571, new_n19563, new_n19572);
xnor_4 g17224(new_n19572, new_n7821, new_n19573);
xnor_4 g17225(new_n19569, new_n19565, new_n19574);
nand_5 g17226(new_n19574, new_n7827, new_n19575_1);
xnor_4 g17227(new_n19574, new_n7826, new_n19576);
not_8  g17228(new_n17793, new_n19577);
nand_5 g17229(new_n19577, new_n7833, new_n19578);
nand_5 g17230(new_n17818, new_n17794, new_n19579);
nand_5 g17231(new_n19579, new_n19578, new_n19580);
nand_5 g17232(new_n19580, new_n19576, new_n19581);
nand_5 g17233(new_n19581, new_n19575_1, new_n19582);
xnor_4 g17234(new_n19582, new_n19573, n5274);
nor_5  g17235(n25316, n20385, new_n19584_1);
nand_5 g17236(new_n19584_1, new_n4327, new_n19585);
nor_5  g17237(new_n19585, n3918, new_n19586);
xnor_4 g17238(new_n19586, new_n6659_1, new_n19587);
xnor_4 g17239(new_n19587, new_n11889, new_n19588);
xnor_4 g17240(new_n19585, n3918, new_n19589);
nand_5 g17241(new_n19589, new_n9371_1, new_n19590);
xnor_4 g17242(new_n19584_1, new_n4327, new_n19591);
nand_5 g17243(new_n19591, new_n9379, new_n19592);
xnor_4 g17244(new_n19591, new_n9380_1, new_n19593);
xnor_4 g17245(n25316, n20385, new_n19594);
nor_5  g17246(new_n19594, new_n9385, new_n19595);
nor_5  g17247(new_n9388, new_n4342, new_n19596);
not_8  g17248(new_n19596, new_n19597);
xnor_4 g17249(new_n19594, new_n9385, new_n19598);
nor_5  g17250(new_n19598, new_n19597, new_n19599);
nor_5  g17251(new_n19599, new_n19595, new_n19600);
nand_5 g17252(new_n19600, new_n19593, new_n19601);
nand_5 g17253(new_n19601, new_n19592, new_n19602_1);
xnor_4 g17254(new_n19589, new_n9372_1, new_n19603);
nand_5 g17255(new_n19603, new_n19602_1, new_n19604);
nand_5 g17256(new_n19604, new_n19590, new_n19605);
xnor_4 g17257(new_n19605, new_n19588, new_n19606);
xnor_4 g17258(new_n17558, n19472, new_n19607);
nand_5 g17259(new_n17562, n25370, new_n19608_1);
xnor_4 g17260(new_n17562, new_n9165, new_n19609);
not_8  g17261(new_n4311, new_n19610);
nand_5 g17262(new_n19610, n24786, new_n19611);
xnor_4 g17263(new_n4311, n24786, new_n19612);
nand_5 g17264(new_n4315, n27120, new_n19613);
nor_5  g17265(new_n4319_1, n23065, new_n19614);
not_8  g17266(new_n19614, new_n19615);
xnor_4 g17267(new_n4315, new_n9155, new_n19616);
nand_5 g17268(new_n19616, new_n19615, new_n19617_1);
nand_5 g17269(new_n19617_1, new_n19613, new_n19618_1);
nand_5 g17270(new_n19618_1, new_n19612, new_n19619);
nand_5 g17271(new_n19619, new_n19611, new_n19620);
nand_5 g17272(new_n19620, new_n19609, new_n19621);
nand_5 g17273(new_n19621, new_n19608_1, new_n19622);
xnor_4 g17274(new_n19622, new_n19607, new_n19623_1);
xnor_4 g17275(new_n19623_1, new_n19606, new_n19624);
xnor_4 g17276(new_n19620, new_n19609, new_n19625);
xnor_4 g17277(new_n19603, new_n19602_1, new_n19626);
not_8  g17278(new_n19626, new_n19627);
nand_5 g17279(new_n19627, new_n19625, new_n19628);
xnor_4 g17280(new_n19626, new_n19625, new_n19629);
xnor_4 g17281(new_n19618_1, new_n19612, new_n19630);
xnor_4 g17282(new_n19600, new_n19593, new_n19631);
not_8  g17283(new_n19631, new_n19632);
nand_5 g17284(new_n19632, new_n19630, new_n19633);
xnor_4 g17285(new_n19631, new_n19630, new_n19634);
xnor_4 g17286(new_n19598, new_n19596, new_n19635);
xnor_4 g17287(new_n19616, new_n19614, new_n19636);
nor_5  g17288(new_n19636, new_n19635, new_n19637);
not_8  g17289(new_n19637, new_n19638);
not_8  g17290(new_n9481, new_n19639);
xnor_4 g17291(new_n4319_1, new_n9148, new_n19640);
nor_5  g17292(new_n19640, new_n19639, new_n19641_1);
not_8  g17293(new_n19641_1, new_n19642);
not_8  g17294(new_n19636, new_n19643);
xnor_4 g17295(new_n19643, new_n19635, new_n19644);
nand_5 g17296(new_n19644, new_n19642, new_n19645);
nand_5 g17297(new_n19645, new_n19638, new_n19646);
nand_5 g17298(new_n19646, new_n19634, new_n19647);
nand_5 g17299(new_n19647, new_n19633, new_n19648_1);
nand_5 g17300(new_n19648_1, new_n19629, new_n19649);
nand_5 g17301(new_n19649, new_n19628, new_n19650);
xnor_4 g17302(new_n19650, new_n19624, n5300);
nor_5  g17303(new_n13965, new_n7620, new_n19652_1);
nor_5  g17304(new_n7630_1, new_n7626, new_n19653);
nor_5  g17305(new_n19653, new_n19652_1, new_n19654);
nor_5  g17306(new_n19654, new_n19551, new_n19655);
xnor_4 g17307(new_n19654, new_n19550, new_n19656);
not_8  g17308(new_n19656, new_n19657);
nand_5 g17309(new_n19550, new_n7631, new_n19658);
nand_5 g17310(new_n19559, new_n19552, new_n19659);
nand_5 g17311(new_n19659, new_n19658, new_n19660);
nor_5  g17312(new_n19660, new_n19657, new_n19661);
nor_5  g17313(new_n19661, new_n19655, n5325);
xnor_4 g17314(n25120, new_n11675, new_n19663);
not_8  g17315(new_n19663, new_n19664_1);
or_5   g17316(n8363, n1222, new_n19665);
xnor_4 g17317(n8363, new_n11678, new_n19666);
or_5   g17318(n25240, n14680, new_n19667);
xnor_4 g17319(n25240, new_n14989_1, new_n19668);
or_5   g17320(n17250, n10125, new_n19669);
xnor_4 g17321(n17250, new_n7647_1, new_n19670);
or_5   g17322(new_n11283, new_n7650, new_n19671);
not_8  g17323(new_n19671, new_n19672);
nor_5  g17324(n23160, n8067, new_n19673);
nor_5  g17325(n20923, n16524, new_n19674);
not_8  g17326(new_n13783_1, new_n19675);
nor_5  g17327(new_n13787, new_n19675, new_n19676);
nor_5  g17328(new_n19676, new_n19674, new_n19677);
not_8  g17329(new_n19677, new_n19678);
nor_5  g17330(new_n19678, new_n19673, new_n19679);
nor_5  g17331(new_n19679, new_n19672, new_n19680_1);
nand_5 g17332(new_n19680_1, new_n19670, new_n19681);
nand_5 g17333(new_n19681, new_n19669, new_n19682);
nand_5 g17334(new_n19682, new_n19668, new_n19683);
nand_5 g17335(new_n19683, new_n19667, new_n19684);
nand_5 g17336(new_n19684, new_n19666, new_n19685);
nand_5 g17337(new_n19685, new_n19665, new_n19686);
xnor_4 g17338(new_n19686, new_n19664_1, new_n19687);
nand_5 g17339(new_n19687, new_n4548, new_n19688);
xnor_4 g17340(new_n19687, n23272, new_n19689);
not_8  g17341(new_n19666, new_n19690);
xnor_4 g17342(new_n19684, new_n19690, new_n19691);
nand_5 g17343(new_n19691, new_n4552_1, new_n19692);
xnor_4 g17344(new_n19691, n11481, new_n19693);
not_8  g17345(new_n19668, new_n19694);
xnor_4 g17346(new_n19682, new_n19694, new_n19695);
nand_5 g17347(new_n19695, new_n4556, new_n19696);
xnor_4 g17348(new_n19695, n16439, new_n19697);
xnor_4 g17349(new_n19680_1, new_n19670, new_n19698);
not_8  g17350(new_n19698, new_n19699);
nand_5 g17351(new_n19699, new_n4560, new_n19700);
xnor_4 g17352(new_n19698, new_n4560, new_n19701_1);
xnor_4 g17353(n23160, new_n7650, new_n19702);
xnor_4 g17354(new_n19702, new_n19678, new_n19703);
not_8  g17355(new_n19703, new_n19704);
nand_5 g17356(new_n19704, new_n4564, new_n19705);
xnor_4 g17357(new_n19703, new_n4564, new_n19706);
nand_5 g17358(new_n13788, new_n4568, new_n19707);
not_8  g17359(new_n13794, new_n19708);
nand_5 g17360(new_n19708, new_n13789, new_n19709);
nand_5 g17361(new_n19709, new_n19707, new_n19710);
nand_5 g17362(new_n19710, new_n19706, new_n19711);
nand_5 g17363(new_n19711, new_n19705, new_n19712);
nand_5 g17364(new_n19712, new_n19701_1, new_n19713);
nand_5 g17365(new_n19713, new_n19700, new_n19714);
nand_5 g17366(new_n19714, new_n19697, new_n19715);
nand_5 g17367(new_n19715, new_n19696, new_n19716);
nand_5 g17368(new_n19716, new_n19693, new_n19717);
nand_5 g17369(new_n19717, new_n19692, new_n19718);
nand_5 g17370(new_n19718, new_n19689, new_n19719);
nand_5 g17371(new_n19719, new_n19688, new_n19720);
or_5   g17372(n25120, n17458, new_n19721);
nand_5 g17373(new_n19686, new_n19663, new_n19722);
nand_5 g17374(new_n19722, new_n19721, new_n19723);
nor_5  g17375(new_n19723, new_n19720, new_n19724);
xnor_4 g17376(n12702, new_n9274, new_n19725);
nor_5  g17377(n26797, n15077, new_n19726);
xnor_4 g17378(n26797, new_n9341, new_n19727);
not_8  g17379(new_n19727, new_n19728);
nor_5  g17380(n23913, n3710, new_n19729);
xnor_4 g17381(n23913, new_n9349, new_n19730);
not_8  g17382(new_n19730, new_n19731);
nor_5  g17383(n26318, n22554, new_n19732);
xnor_4 g17384(n26318, new_n5836, new_n19733);
not_8  g17385(new_n19733, new_n19734);
nor_5  g17386(n26054, n20429, new_n19735);
xnor_4 g17387(n26054, new_n5862, new_n19736_1);
not_8  g17388(new_n19736_1, new_n19737);
nor_5  g17389(n19081, n3909, new_n19738);
xnor_4 g17390(n19081, new_n5837, new_n19739);
not_8  g17391(new_n19739, new_n19740);
nor_5  g17392(n23974, n8309, new_n19741);
xnor_4 g17393(n23974, new_n9306, new_n19742);
nand_5 g17394(n19144, n2146, new_n19743);
not_8  g17395(new_n19743, new_n19744);
nor_5  g17396(n19144, n2146, new_n19745);
nor_5  g17397(n22173, n12593, new_n19746);
not_8  g17398(new_n17767, new_n19747);
nor_5  g17399(new_n17768, new_n19747, new_n19748);
nor_5  g17400(new_n19748, new_n19746, new_n19749_1);
not_8  g17401(new_n19749_1, new_n19750);
nor_5  g17402(new_n19750, new_n19745, new_n19751);
nor_5  g17403(new_n19751, new_n19744, new_n19752);
nand_5 g17404(new_n19752, new_n19742, new_n19753);
not_8  g17405(new_n19753, new_n19754);
nor_5  g17406(new_n19754, new_n19741, new_n19755);
nor_5  g17407(new_n19755, new_n19740, new_n19756_1);
nor_5  g17408(new_n19756_1, new_n19738, new_n19757);
nor_5  g17409(new_n19757, new_n19737, new_n19758);
nor_5  g17410(new_n19758, new_n19735, new_n19759);
nor_5  g17411(new_n19759, new_n19734, new_n19760);
nor_5  g17412(new_n19760, new_n19732, new_n19761);
nor_5  g17413(new_n19761, new_n19731, new_n19762);
nor_5  g17414(new_n19762, new_n19729, new_n19763);
nor_5  g17415(new_n19763, new_n19728, new_n19764);
nor_5  g17416(new_n19764, new_n19726, new_n19765);
xnor_4 g17417(new_n19765, new_n19725, new_n19766);
nand_5 g17418(new_n19766, new_n5904_1, new_n19767_1);
xnor_4 g17419(new_n19766, n12650, new_n19768);
xnor_4 g17420(new_n19763, new_n19727, new_n19769);
nand_5 g17421(new_n19769, new_n5835, new_n19770_1);
xnor_4 g17422(new_n19769, n10201, new_n19771);
xnor_4 g17423(new_n19761, new_n19730, new_n19772);
nand_5 g17424(new_n19772, new_n5850_1, new_n19773);
xnor_4 g17425(new_n19772, n10593, new_n19774);
xnor_4 g17426(new_n19759, new_n19733, new_n19775);
nand_5 g17427(new_n19775, new_n5856, new_n19776);
xnor_4 g17428(new_n19757, new_n19736_1, new_n19777);
nand_5 g17429(new_n19777, new_n5861, new_n19778);
xnor_4 g17430(new_n19777, n11580, new_n19779);
xnor_4 g17431(new_n19755, new_n19739, new_n19780_1);
nand_5 g17432(new_n19780_1, new_n5867, new_n19781);
xnor_4 g17433(new_n19780_1, n15884, new_n19782);
xnor_4 g17434(new_n19752, new_n19742, new_n19783);
nor_5  g17435(new_n19783, n6356, new_n19784);
xnor_4 g17436(n19144, n2146, new_n19785);
xnor_4 g17437(new_n19785, new_n19749_1, new_n19786);
nand_5 g17438(new_n19786, n27104, new_n19787);
xnor_4 g17439(new_n19786, new_n5877, new_n19788);
and_5  g17440(new_n17769, new_n5882_1, new_n19789_1);
nor_5  g17441(new_n17770, new_n17766, new_n19790);
nor_5  g17442(new_n19790, new_n19789_1, new_n19791);
nand_5 g17443(new_n19791, new_n19788, new_n19792_1);
nand_5 g17444(new_n19792_1, new_n19787, new_n19793);
xnor_4 g17445(new_n19783, new_n5872, new_n19794);
not_8  g17446(new_n19794, new_n19795);
nor_5  g17447(new_n19795, new_n19793, new_n19796);
nor_5  g17448(new_n19796, new_n19784, new_n19797);
not_8  g17449(new_n19797, new_n19798_1);
nand_5 g17450(new_n19798_1, new_n19782, new_n19799);
nand_5 g17451(new_n19799, new_n19781, new_n19800);
nand_5 g17452(new_n19800, new_n19779, new_n19801);
nand_5 g17453(new_n19801, new_n19778, new_n19802);
xnor_4 g17454(new_n19775, n18290, new_n19803_1);
nand_5 g17455(new_n19803_1, new_n19802, new_n19804);
nand_5 g17456(new_n19804, new_n19776, new_n19805);
nand_5 g17457(new_n19805, new_n19774, new_n19806);
nand_5 g17458(new_n19806, new_n19773, new_n19807);
nand_5 g17459(new_n19807, new_n19771, new_n19808);
nand_5 g17460(new_n19808, new_n19770_1, new_n19809);
nand_5 g17461(new_n19809, new_n19768, new_n19810);
nand_5 g17462(new_n19810, new_n19767_1, new_n19811);
or_5   g17463(n12702, n12507, new_n19812);
not_8  g17464(new_n19765, new_n19813);
nand_5 g17465(new_n19813, new_n19725, new_n19814);
nand_5 g17466(new_n19814, new_n19812, new_n19815);
nor_5  g17467(new_n19815, new_n19811, new_n19816);
xnor_4 g17468(new_n19816, new_n19724, new_n19817);
xnor_4 g17469(new_n19723, new_n19720, new_n19818);
not_8  g17470(new_n19818, new_n19819);
xnor_4 g17471(new_n19815, new_n19811, new_n19820);
nand_5 g17472(new_n19820, new_n19819, new_n19821);
xnor_4 g17473(new_n19820, new_n19818, new_n19822);
xnor_4 g17474(new_n19718, new_n19689, new_n19823);
xnor_4 g17475(new_n19809, new_n19768, new_n19824);
not_8  g17476(new_n19824, new_n19825);
nand_5 g17477(new_n19825, new_n19823, new_n19826);
xnor_4 g17478(new_n19824, new_n19823, new_n19827);
xnor_4 g17479(new_n19716, new_n19693, new_n19828);
not_8  g17480(new_n19771, new_n19829);
xnor_4 g17481(new_n19807, new_n19829, new_n19830);
nand_5 g17482(new_n19830, new_n19828, new_n19831);
not_8  g17483(new_n19828, new_n19832);
xnor_4 g17484(new_n19830, new_n19832, new_n19833);
xnor_4 g17485(new_n19714, new_n19697, new_n19834);
not_8  g17486(new_n19774, new_n19835);
xnor_4 g17487(new_n19805, new_n19835, new_n19836);
nand_5 g17488(new_n19836, new_n19834, new_n19837);
not_8  g17489(new_n19834, new_n19838);
xnor_4 g17490(new_n19836, new_n19838, new_n19839);
not_8  g17491(new_n19701_1, new_n19840);
xnor_4 g17492(new_n19712, new_n19840, new_n19841);
not_8  g17493(new_n19841, new_n19842);
not_8  g17494(new_n19803_1, new_n19843);
xnor_4 g17495(new_n19843, new_n19802, new_n19844);
nand_5 g17496(new_n19844, new_n19842, new_n19845);
xnor_4 g17497(new_n19844, new_n19841, new_n19846);
not_8  g17498(new_n19779, new_n19847);
xnor_4 g17499(new_n19800, new_n19847, new_n19848);
xnor_4 g17500(new_n19710, new_n19706, new_n19849);
nand_5 g17501(new_n19849, new_n19848, new_n19850);
not_8  g17502(new_n19849, new_n19851);
xnor_4 g17503(new_n19851, new_n19848, new_n19852);
xnor_4 g17504(new_n19797, new_n19782, new_n19853);
nand_5 g17505(new_n19853, new_n13796, new_n19854);
xnor_4 g17506(new_n19853, new_n13795, new_n19855);
xnor_4 g17507(new_n19794, new_n19793, new_n19856);
not_8  g17508(new_n19856, new_n19857);
nor_5  g17509(new_n19857, new_n7011, new_n19858);
xnor_4 g17510(new_n19791, new_n19788, new_n19859);
not_8  g17511(new_n19859, new_n19860);
nor_5  g17512(new_n19860, new_n7016, new_n19861);
xnor_4 g17513(new_n19859, new_n7016, new_n19862);
not_8  g17514(new_n19862, new_n19863);
nor_5  g17515(new_n17772, new_n17765, new_n19864);
nor_5  g17516(new_n17773, new_n7021, new_n19865);
nor_5  g17517(new_n19865, new_n19864, new_n19866);
not_8  g17518(new_n19866, new_n19867);
nor_5  g17519(new_n19867, new_n19863, new_n19868);
nor_5  g17520(new_n19868, new_n19861, new_n19869);
xnor_4 g17521(new_n19856, new_n7011, new_n19870);
not_8  g17522(new_n19870, new_n19871);
nor_5  g17523(new_n19871, new_n19869, new_n19872);
nor_5  g17524(new_n19872, new_n19858, new_n19873_1);
not_8  g17525(new_n19873_1, new_n19874);
nand_5 g17526(new_n19874, new_n19855, new_n19875);
nand_5 g17527(new_n19875, new_n19854, new_n19876);
nand_5 g17528(new_n19876, new_n19852, new_n19877);
nand_5 g17529(new_n19877, new_n19850, new_n19878);
nand_5 g17530(new_n19878, new_n19846, new_n19879);
nand_5 g17531(new_n19879, new_n19845, new_n19880);
nand_5 g17532(new_n19880, new_n19839, new_n19881);
nand_5 g17533(new_n19881, new_n19837, new_n19882);
nand_5 g17534(new_n19882, new_n19833, new_n19883);
nand_5 g17535(new_n19883, new_n19831, new_n19884);
nand_5 g17536(new_n19884, new_n19827, new_n19885);
nand_5 g17537(new_n19885, new_n19826, new_n19886);
nand_5 g17538(new_n19886, new_n19822, new_n19887);
nand_5 g17539(new_n19887, new_n19821, new_n19888);
xnor_4 g17540(new_n19888, new_n19817, n5351);
nand_5 g17541(new_n17458_1, new_n17449, new_n19890);
not_8  g17542(new_n19890, n5353);
nor_5  g17543(new_n12558, n2160, new_n19892);
not_8  g17544(new_n12559, new_n19893);
nor_5  g17545(new_n12611, new_n19893, new_n19894);
nor_5  g17546(new_n19894, new_n19892, new_n19895);
or_5   g17547(n9934, n2272, new_n19896);
nand_5 g17548(new_n12557, new_n12515_1, new_n19897);
nand_5 g17549(new_n19897, new_n19896, new_n19898);
nand_5 g17550(new_n19898, new_n19895, new_n19899);
nor_5  g17551(new_n12618, n21784, new_n19900);
not_8  g17552(new_n19900, new_n19901);
nand_5 g17553(new_n19901, new_n7704, new_n19902);
not_8  g17554(new_n19902, new_n19903);
not_8  g17555(new_n12619, new_n19904);
nand_5 g17556(new_n19904, new_n7707, new_n19905_1);
nand_5 g17557(new_n12636, new_n12620_1, new_n19906);
nand_5 g17558(new_n19906, new_n19905_1, new_n19907);
nand_5 g17559(new_n19907, new_n19903, new_n19908);
not_8  g17560(new_n19908, new_n19909_1);
xnor_4 g17561(new_n19909_1, new_n19899, new_n19910);
xnor_4 g17562(new_n19898, new_n19895, new_n19911_1);
not_8  g17563(new_n19911_1, new_n19912);
xnor_4 g17564(new_n19900, new_n7704, new_n19913);
xnor_4 g17565(new_n19913, new_n19907, new_n19914);
nand_5 g17566(new_n19914, new_n19912, new_n19915);
xnor_4 g17567(new_n19914, new_n19911_1, new_n19916_1);
not_8  g17568(new_n12637, new_n19917);
nand_5 g17569(new_n19917, new_n12613, new_n19918);
nand_5 g17570(new_n12692, new_n12638, new_n19919);
nand_5 g17571(new_n19919, new_n19918, new_n19920);
nand_5 g17572(new_n19920, new_n19916_1, new_n19921);
nand_5 g17573(new_n19921, new_n19915, new_n19922_1);
xnor_4 g17574(new_n19922_1, new_n19910, n5399);
nand_5 g17575(new_n18612, n2979, new_n19924);
nand_5 g17576(new_n18616, new_n18613, new_n19925);
nand_5 g17577(new_n19925, new_n19924, new_n19926);
nand_5 g17578(new_n15056, n9934, new_n19927);
nor_5  g17579(new_n15056, n9934, new_n19928);
nor_5  g17580(new_n18611, new_n19928, new_n19929);
nor_5  g17581(new_n19929, new_n15109, new_n19930_1);
and_5  g17582(new_n19930_1, new_n19927, new_n19931);
nand_5 g17583(new_n19931, new_n19926, new_n19932);
xnor_4 g17584(new_n19932, new_n19909_1, new_n19933);
not_8  g17585(new_n19926, new_n19934);
xnor_4 g17586(new_n19931, new_n19934, new_n19935);
not_8  g17587(new_n19935, new_n19936);
nand_5 g17588(new_n19936, new_n19914, new_n19937);
nand_5 g17589(new_n18617, new_n19917, new_n19938);
nand_5 g17590(new_n18621, new_n18618, new_n19939);
nand_5 g17591(new_n19939, new_n19938, new_n19940);
xnor_4 g17592(new_n19935, new_n19914, new_n19941_1);
nand_5 g17593(new_n19941_1, new_n19940, new_n19942);
nand_5 g17594(new_n19942, new_n19937, new_n19943);
xnor_4 g17595(new_n19943, new_n19933, n5403);
xnor_4 g17596(new_n16608_1, new_n16573, n5430);
not_8  g17597(new_n15517, new_n19946);
nor_5  g17598(new_n15523, new_n19946, new_n19947);
not_8  g17599(new_n15512, new_n19948);
nand_5 g17600(new_n19948, new_n11089, new_n19949);
nand_5 g17601(new_n15512, new_n11093, new_n19950);
nand_5 g17602(new_n15524, new_n19950, new_n19951);
nand_5 g17603(new_n19951, new_n19949, new_n19952);
nor_5  g17604(new_n19952, new_n10941, new_n19953);
not_8  g17605(new_n19953, new_n19954);
nor_5  g17606(new_n19954, new_n19947, n5439);
xnor_4 g17607(new_n13048_1, new_n13027, n5472);
xnor_4 g17608(new_n8909_1, new_n8867, n5485);
xnor_4 g17609(new_n19351, new_n19332, n5524);
nand_5 g17610(new_n17471, new_n6276_1, new_n19959);
nor_5  g17611(new_n19959, new_n14315, new_n19960);
nand_5 g17612(new_n19960, new_n6263, new_n19961);
nor_5  g17613(new_n19961, new_n6259, new_n19962);
nand_5 g17614(new_n19962, new_n6252, new_n19963);
nor_5  g17615(new_n19963, new_n6247, new_n19964);
not_8  g17616(new_n19964, new_n19965);
nor_5  g17617(new_n19965, new_n6240, new_n19966);
xnor_4 g17618(new_n19966, new_n6236, new_n19967);
not_8  g17619(new_n19967, new_n19968_1);
nand_5 g17620(new_n19968_1, new_n14646, new_n19969);
xnor_4 g17621(new_n19967, new_n14646, new_n19970);
not_8  g17622(new_n14651, new_n19971);
xnor_4 g17623(new_n19964, new_n6240, new_n19972);
not_8  g17624(new_n19972, new_n19973);
nand_5 g17625(new_n19973, new_n19971, new_n19974);
xnor_4 g17626(new_n19972, new_n19971, new_n19975);
not_8  g17627(new_n14655, new_n19976);
xnor_4 g17628(new_n19963, new_n6247, new_n19977);
nand_5 g17629(new_n19977, new_n19976, new_n19978);
xnor_4 g17630(new_n19977, new_n14655, new_n19979);
xnor_4 g17631(new_n19962, new_n6252, new_n19980);
nand_5 g17632(new_n19980, new_n14659, new_n19981);
xnor_4 g17633(new_n19980, new_n14660, new_n19982);
xnor_4 g17634(new_n19961, new_n6259, new_n19983);
nand_5 g17635(new_n19983, new_n14663, new_n19984);
xnor_4 g17636(new_n19983, new_n14664, new_n19985);
xnor_4 g17637(new_n19960, new_n14310_1, new_n19986);
not_8  g17638(new_n19986, new_n19987);
nand_5 g17639(new_n19987, new_n14667, new_n19988_1);
xnor_4 g17640(new_n19986, new_n14667, new_n19989);
xnor_4 g17641(new_n19959, new_n6269, new_n19990);
not_8  g17642(new_n19990, new_n19991);
not_8  g17643(new_n13897, new_n19992);
nand_5 g17644(new_n18624, new_n19992, new_n19993);
nand_5 g17645(new_n18629, new_n18625, new_n19994);
nand_5 g17646(new_n19994, new_n19993, new_n19995);
nand_5 g17647(new_n19995, new_n19991, new_n19996);
xnor_4 g17648(new_n19995, new_n19990, new_n19997);
nand_5 g17649(new_n19997, new_n13894, new_n19998);
nand_5 g17650(new_n19998, new_n19996, new_n19999);
nand_5 g17651(new_n19999, new_n19989, new_n20000);
nand_5 g17652(new_n20000, new_n19988_1, new_n20001);
nand_5 g17653(new_n20001, new_n19985, new_n20002);
nand_5 g17654(new_n20002, new_n19984, new_n20003);
nand_5 g17655(new_n20003, new_n19982, new_n20004_1);
nand_5 g17656(new_n20004_1, new_n19981, new_n20005);
nand_5 g17657(new_n20005, new_n19979, new_n20006);
nand_5 g17658(new_n20006, new_n19978, new_n20007);
nand_5 g17659(new_n20007, new_n19975, new_n20008);
nand_5 g17660(new_n20008, new_n19974, new_n20009);
nand_5 g17661(new_n20009, new_n19970, new_n20010);
nand_5 g17662(new_n20010, new_n19969, new_n20011);
not_8  g17663(new_n19966, new_n20012);
nor_5  g17664(new_n20012, new_n6236, new_n20013_1);
nor_5  g17665(new_n20013_1, new_n14286, new_n20014);
nand_5 g17666(new_n20013_1, new_n14283, new_n20015);
not_8  g17667(new_n20015, new_n20016);
nor_5  g17668(new_n20016, new_n20014, new_n20017_1);
xnor_4 g17669(new_n20017_1, new_n14695, new_n20018);
xnor_4 g17670(new_n20018, new_n20011, new_n20019);
nand_5 g17671(new_n20019, new_n5040, new_n20020);
xnor_4 g17672(new_n20019, new_n5041, new_n20021);
xnor_4 g17673(new_n20009, new_n19970, new_n20022);
not_8  g17674(new_n20022, new_n20023);
nand_5 g17675(new_n20023, new_n5219, new_n20024);
xnor_4 g17676(new_n20022, new_n5219, new_n20025);
xnor_4 g17677(new_n20007, new_n19975, new_n20026);
not_8  g17678(new_n20026, new_n20027);
nand_5 g17679(new_n20027, new_n5226_1, new_n20028);
xnor_4 g17680(new_n20026, new_n5226_1, new_n20029);
xnor_4 g17681(new_n20005, new_n19979, new_n20030);
not_8  g17682(new_n20030, new_n20031);
nand_5 g17683(new_n20031, new_n5230, new_n20032);
xnor_4 g17684(new_n20030, new_n5230, new_n20033_1);
xnor_4 g17685(new_n20003, new_n19982, new_n20034);
not_8  g17686(new_n20034, new_n20035);
nand_5 g17687(new_n20035, new_n5235, new_n20036_1);
xnor_4 g17688(new_n20034, new_n5235, new_n20037);
xnor_4 g17689(new_n20001, new_n19985, new_n20038);
not_8  g17690(new_n20038, new_n20039);
nand_5 g17691(new_n20039, new_n5241, new_n20040_1);
xnor_4 g17692(new_n20038, new_n5241, new_n20041);
xnor_4 g17693(new_n19999, new_n19989, new_n20042);
not_8  g17694(new_n20042, new_n20043);
nand_5 g17695(new_n20043, new_n5247, new_n20044);
xnor_4 g17696(new_n20042, new_n5247, new_n20045);
xnor_4 g17697(new_n19997, new_n13894, new_n20046);
not_8  g17698(new_n20046, new_n20047);
nand_5 g17699(new_n20047, new_n5252, new_n20048);
xnor_4 g17700(new_n20046, new_n5252, new_n20049);
and_5  g17701(new_n18630, new_n5263, new_n20050);
not_8  g17702(new_n18631, new_n20051);
nor_5  g17703(new_n18633, new_n20051, new_n20052);
nor_5  g17704(new_n20052, new_n20050, new_n20053);
nand_5 g17705(new_n20053, new_n20049, new_n20054);
nand_5 g17706(new_n20054, new_n20048, new_n20055);
nand_5 g17707(new_n20055, new_n20045, new_n20056);
nand_5 g17708(new_n20056, new_n20044, new_n20057);
nand_5 g17709(new_n20057, new_n20041, new_n20058);
nand_5 g17710(new_n20058, new_n20040_1, new_n20059);
nand_5 g17711(new_n20059, new_n20037, new_n20060);
nand_5 g17712(new_n20060, new_n20036_1, new_n20061_1);
nand_5 g17713(new_n20061_1, new_n20033_1, new_n20062);
nand_5 g17714(new_n20062, new_n20032, new_n20063);
nand_5 g17715(new_n20063, new_n20029, new_n20064);
nand_5 g17716(new_n20064, new_n20028, new_n20065);
nand_5 g17717(new_n20065, new_n20025, new_n20066);
nand_5 g17718(new_n20066, new_n20024, new_n20067);
nand_5 g17719(new_n20067, new_n20021, new_n20068);
nand_5 g17720(new_n20068, new_n20020, new_n20069_1);
not_8  g17721(new_n20017_1, new_n20070);
nand_5 g17722(new_n20070, new_n14696, new_n20071);
nand_5 g17723(new_n20017_1, new_n14695, new_n20072);
nand_5 g17724(new_n20072, new_n20011, new_n20073);
nand_5 g17725(new_n20073, new_n20071, new_n20074);
nand_5 g17726(new_n20074, new_n20015, new_n20075);
not_8  g17727(new_n20075, new_n20076);
xnor_4 g17728(new_n20076, new_n20069_1, n5564);
xnor_4 g17729(new_n7343, new_n7330_1, n5593);
xnor_4 g17730(new_n18669, new_n15135, new_n20079);
nand_5 g17731(new_n17354, new_n15142, new_n20080);
xnor_4 g17732(new_n18672, new_n15142, new_n20081);
nand_5 g17733(new_n17356, new_n15147, new_n20082);
xnor_4 g17734(new_n17356, new_n15149, new_n20083);
nand_5 g17735(new_n16324, new_n15153, new_n20084);
xnor_4 g17736(new_n17360, new_n15153, new_n20085);
nor_5  g17737(new_n16327_1, new_n15158, new_n20086_1);
not_8  g17738(new_n18194, new_n20087);
not_8  g17739(new_n18207, new_n20088);
nor_5  g17740(new_n20088, new_n20087, new_n20089);
nor_5  g17741(new_n20089, new_n20086_1, new_n20090);
not_8  g17742(new_n20090, new_n20091);
nand_5 g17743(new_n20091, new_n20085, new_n20092);
nand_5 g17744(new_n20092, new_n20084, new_n20093);
nand_5 g17745(new_n20093, new_n20083, new_n20094);
nand_5 g17746(new_n20094, new_n20082, new_n20095);
nand_5 g17747(new_n20095, new_n20081, new_n20096_1);
nand_5 g17748(new_n20096_1, new_n20080, new_n20097);
xnor_4 g17749(new_n20097, new_n20079, n5603);
xnor_4 g17750(n17911, n14440, new_n20099);
not_8  g17751(new_n20099, new_n20100);
nor_5  g17752(new_n16889, n1654, new_n20101);
xnor_4 g17753(n21997, n1654, new_n20102);
not_8  g17754(new_n20102, new_n20103_1);
nor_5  g17755(new_n16894, n13783, new_n20104);
xnor_4 g17756(n25119, n13783, new_n20105);
not_8  g17757(new_n20105, new_n20106);
nor_5  g17758(n26660, new_n9035, new_n20107);
xnor_4 g17759(n26660, n1163, new_n20108);
not_8  g17760(new_n20108, new_n20109);
nor_5  g17761(new_n16237, n3018, new_n20110);
nor_5  g17762(n18537, new_n11311, new_n20111);
nor_5  g17763(n7057, new_n2398, new_n20112);
not_8  g17764(new_n18969, new_n20113);
nor_5  g17765(new_n18981, new_n20113, new_n20114);
nor_5  g17766(new_n20114, new_n20112, new_n20115);
not_8  g17767(new_n20115, new_n20116);
nor_5  g17768(new_n20116, new_n20111, new_n20117);
nor_5  g17769(new_n20117, new_n20110, new_n20118);
nor_5  g17770(new_n20118, new_n20109, new_n20119);
nor_5  g17771(new_n20119, new_n20107, new_n20120);
nor_5  g17772(new_n20120, new_n20106, new_n20121);
nor_5  g17773(new_n20121, new_n20104, new_n20122);
nor_5  g17774(new_n20122, new_n20103_1, new_n20123);
nor_5  g17775(new_n20123, new_n20101, new_n20124);
xnor_4 g17776(new_n20124, new_n20100, new_n20125);
xnor_4 g17777(new_n20125, new_n3100, new_n20126_1);
not_8  g17778(new_n20126_1, new_n20127);
xnor_4 g17779(new_n20122, new_n20102, new_n20128);
nor_5  g17780(new_n20128, new_n3103, new_n20129);
xnor_4 g17781(new_n20128, new_n3104, new_n20130);
not_8  g17782(new_n20130, new_n20131);
xnor_4 g17783(new_n20120, new_n20105, new_n20132);
nor_5  g17784(new_n20132, new_n3108, new_n20133);
xnor_4 g17785(new_n20132, new_n3109, new_n20134);
not_8  g17786(new_n20134, new_n20135);
xnor_4 g17787(new_n20118, new_n20108, new_n20136);
not_8  g17788(new_n20136, new_n20137);
nand_5 g17789(new_n20137, new_n3114, new_n20138_1);
xnor_4 g17790(new_n20136, new_n3114, new_n20139);
xnor_4 g17791(n18537, n3018, new_n20140);
xnor_4 g17792(new_n20140, new_n20115, new_n20141);
nor_5  g17793(new_n20141, new_n3118, new_n20142);
not_8  g17794(new_n20142, new_n20143);
nor_5  g17795(new_n18982_1, new_n3122, new_n20144);
not_8  g17796(new_n20144, new_n20145);
not_8  g17797(new_n19000, new_n20146);
nand_5 g17798(new_n20146, new_n18983, new_n20147);
nand_5 g17799(new_n20147, new_n20145, new_n20148);
xnor_4 g17800(new_n20141, new_n3120, new_n20149_1);
nand_5 g17801(new_n20149_1, new_n20148, new_n20150);
nand_5 g17802(new_n20150, new_n20143, new_n20151_1);
not_8  g17803(new_n20151_1, new_n20152);
nand_5 g17804(new_n20152, new_n20139, new_n20153);
nand_5 g17805(new_n20153, new_n20138_1, new_n20154);
not_8  g17806(new_n20154, new_n20155);
nor_5  g17807(new_n20155, new_n20135, new_n20156);
nor_5  g17808(new_n20156, new_n20133, new_n20157);
nor_5  g17809(new_n20157, new_n20131, new_n20158);
nor_5  g17810(new_n20158, new_n20129, new_n20159);
xnor_4 g17811(new_n20159, new_n20127, n5609);
xnor_4 g17812(new_n14220, new_n14199, n5634);
not_8  g17813(new_n7766, new_n20162);
or_5   g17814(new_n3294, n2978, new_n20163);
xnor_4 g17815(n3425, n2978, new_n20164);
or_5   g17816(n23697, new_n3295, new_n20165);
xnor_4 g17817(n23697, n9967, new_n20166);
or_5   g17818(new_n3317, n2289, new_n20167);
nand_5 g17819(new_n19571, new_n19563, new_n20168);
nand_5 g17820(new_n20168, new_n20167, new_n20169_1);
nand_5 g17821(new_n20169_1, new_n20166, new_n20170);
nand_5 g17822(new_n20170, new_n20165, new_n20171);
nand_5 g17823(new_n20171, new_n20164, new_n20172);
nand_5 g17824(new_n20172, new_n20163, new_n20173);
nand_5 g17825(new_n20173, new_n20162, new_n20174);
not_8  g17826(new_n20173, new_n20175);
nand_5 g17827(new_n20175, new_n7766, new_n20176);
xnor_4 g17828(new_n20171, new_n20164, new_n20177);
nand_5 g17829(new_n20177, new_n7811_1, new_n20178);
xnor_4 g17830(new_n20177, new_n7813, new_n20179_1);
xnor_4 g17831(new_n20169_1, new_n20166, new_n20180);
nand_5 g17832(new_n20180, new_n7817, new_n20181);
xnor_4 g17833(new_n20180, new_n7816, new_n20182);
nand_5 g17834(new_n19572, new_n7822, new_n20183);
nand_5 g17835(new_n19582, new_n19573, new_n20184);
nand_5 g17836(new_n20184, new_n20183, new_n20185);
nand_5 g17837(new_n20185, new_n20182, new_n20186);
nand_5 g17838(new_n20186, new_n20181, new_n20187_1);
nand_5 g17839(new_n20187_1, new_n20179_1, new_n20188);
nand_5 g17840(new_n20188, new_n20178, new_n20189);
nand_5 g17841(new_n20189, new_n20176, new_n20190);
nand_5 g17842(new_n20190, new_n20174, new_n20191);
nor_5  g17843(new_n7704, new_n7684, new_n20192);
not_8  g17844(new_n20192, new_n20193);
nand_5 g17845(new_n7765, new_n7705, new_n20194);
nand_5 g17846(new_n20194, new_n20193, new_n20195);
xnor_4 g17847(new_n20195, new_n20173, new_n20196);
xnor_4 g17848(new_n20196, new_n20191, n5643);
xnor_4 g17849(n18035, n5834, new_n20198);
not_8  g17850(new_n20198, new_n20199);
nor_5  g17851(n13851, new_n11194, new_n20200);
nor_5  g17852(new_n16408, new_n16390, new_n20201);
nor_5  g17853(new_n20201, new_n20200, new_n20202);
xnor_4 g17854(new_n20202, new_n20199, new_n20203);
xnor_4 g17855(new_n20203, new_n15914, new_n20204);
nand_5 g17856(new_n16409, new_n15944, new_n20205);
xnor_4 g17857(new_n16408, new_n16389, new_n20206);
xnor_4 g17858(new_n20206, new_n15944, new_n20207);
nand_5 g17859(new_n16412, new_n15949, new_n20208);
xnor_4 g17860(new_n16411, new_n15949, new_n20209);
nand_5 g17861(new_n16416, new_n15954, new_n20210);
xnor_4 g17862(new_n16415, new_n15954, new_n20211);
nand_5 g17863(new_n16419_1, new_n15956_1, new_n20212);
nand_5 g17864(new_n14761, new_n14483, new_n20213_1);
xnor_4 g17865(new_n14761, new_n16422, new_n20214);
nand_5 g17866(new_n14778, new_n14488, new_n20215);
xnor_4 g17867(new_n14778, new_n14489, new_n20216);
nor_5  g17868(new_n14786, new_n14491, new_n20217);
nor_5  g17869(new_n20217, new_n14498, new_n20218);
xnor_4 g17870(new_n20217, new_n14497, new_n20219);
not_8  g17871(new_n20219, new_n20220);
nor_5  g17872(new_n20220, new_n14792, new_n20221);
nor_5  g17873(new_n20221, new_n20218, new_n20222);
not_8  g17874(new_n20222, new_n20223);
nand_5 g17875(new_n20223, new_n20216, new_n20224);
nand_5 g17876(new_n20224, new_n20215, new_n20225);
nand_5 g17877(new_n20225, new_n20214, new_n20226);
nand_5 g17878(new_n20226, new_n20213_1, new_n20227);
xnor_4 g17879(new_n16419_1, new_n15960, new_n20228);
nand_5 g17880(new_n20228, new_n20227, new_n20229);
nand_5 g17881(new_n20229, new_n20212, new_n20230);
nand_5 g17882(new_n20230, new_n20211, new_n20231);
nand_5 g17883(new_n20231, new_n20210, new_n20232);
nand_5 g17884(new_n20232, new_n20209, new_n20233);
nand_5 g17885(new_n20233, new_n20208, new_n20234);
nand_5 g17886(new_n20234, new_n20207, new_n20235_1);
nand_5 g17887(new_n20235_1, new_n20205, new_n20236);
xor_4  g17888(new_n20236, new_n20204, n5680);
xnor_4 g17889(new_n15621, new_n15619, n5687);
xnor_4 g17890(new_n16750, new_n16741, n5700);
not_8  g17891(new_n11101_1, new_n20240);
xnor_4 g17892(new_n11167, new_n20240, n5732);
xnor_4 g17893(n23775, new_n5296, new_n20242);
nor_5  g17894(n20235, n8259, new_n20243);
not_8  g17895(new_n19475, new_n20244);
nor_5  g17896(new_n19476, new_n20244, new_n20245);
nor_5  g17897(new_n20245, new_n20243, new_n20246);
xnor_4 g17898(new_n20246, new_n20242, new_n20247);
xnor_4 g17899(new_n20247, new_n2395, new_n20248);
nor_5  g17900(new_n19477_1, new_n2387_1, new_n20249);
nor_5  g17901(new_n19478, new_n19474, new_n20250_1);
nor_5  g17902(new_n20250_1, new_n20249, new_n20251);
xnor_4 g17903(new_n20251, new_n20248, new_n20252);
xnor_4 g17904(n8869, n6385, new_n20253);
nand_5 g17905(n20138, new_n7431, new_n20254);
nand_5 g17906(new_n19471, new_n19470, new_n20255);
nand_5 g17907(new_n20255, new_n20254, new_n20256);
xnor_4 g17908(new_n20256, new_n20253, new_n20257);
not_8  g17909(new_n20257, new_n20258);
xnor_4 g17910(new_n20258, new_n20252, new_n20259_1);
not_8  g17911(new_n20259_1, new_n20260);
nand_5 g17912(new_n19472_1, new_n19469, new_n20261);
nor_5  g17913(new_n19479, new_n19473, new_n20262);
not_8  g17914(new_n20262, new_n20263);
nand_5 g17915(new_n20263, new_n20261, new_n20264);
xnor_4 g17916(new_n20264, new_n20260, n5742);
xnor_4 g17917(new_n14507, new_n14505, n5765);
xnor_4 g17918(new_n13286, new_n13240, n5776);
xnor_4 g17919(new_n2891, new_n2848, n5782);
xnor_4 g17920(n18901, new_n9035, new_n20269);
nor_5  g17921(n18537, n4376, new_n20270);
xnor_4 g17922(n18537, new_n7371, new_n20271);
not_8  g17923(new_n20271, new_n20272);
nor_5  g17924(n14570, n7057, new_n20273);
xnor_4 g17925(new_n7375, n7057, new_n20274);
not_8  g17926(new_n20274, new_n20275);
nor_5  g17927(n23775, n8381, new_n20276);
not_8  g17928(new_n20242, new_n20277);
nor_5  g17929(new_n20246, new_n20277, new_n20278);
nor_5  g17930(new_n20278, new_n20276, new_n20279_1);
nor_5  g17931(new_n20279_1, new_n20275, new_n20280);
nor_5  g17932(new_n20280, new_n20273, new_n20281);
nor_5  g17933(new_n20281, new_n20272, new_n20282);
nor_5  g17934(new_n20282, new_n20270, new_n20283);
xnor_4 g17935(new_n20283, new_n20269, new_n20284);
xnor_4 g17936(new_n20284, new_n2420_1, new_n20285);
xnor_4 g17937(new_n20281, new_n20271, new_n20286);
not_8  g17938(new_n20286, new_n20287_1);
nor_5  g17939(new_n20287_1, new_n2472, new_n20288);
xnor_4 g17940(new_n20279_1, new_n20274, new_n20289);
nand_5 g17941(new_n20247, new_n2396, new_n20290);
nand_5 g17942(new_n20251, new_n20248, new_n20291);
nand_5 g17943(new_n20291, new_n20290, new_n20292);
nand_5 g17944(new_n20292, new_n20289, new_n20293);
not_8  g17945(new_n20293, new_n20294);
xnor_4 g17946(new_n20292, new_n20289, new_n20295);
nor_5  g17947(new_n20295, new_n2404, new_n20296);
nor_5  g17948(new_n20296, new_n20294, new_n20297);
xnor_4 g17949(new_n20287_1, new_n2413, new_n20298);
not_8  g17950(new_n20298, new_n20299);
nor_5  g17951(new_n20299, new_n20297, new_n20300);
nor_5  g17952(new_n20300, new_n20288, new_n20301_1);
xnor_4 g17953(new_n20301_1, new_n20285, new_n20302);
not_8  g17954(new_n20302, new_n20303);
xnor_4 g17955(n23068, n7099, new_n20304);
nor_5  g17956(n19514, new_n12575, new_n20305);
xnor_4 g17957(n19514, n12811, new_n20306);
not_8  g17958(new_n20306, new_n20307);
nor_5  g17959(n10053, new_n2959, new_n20308);
xnor_4 g17960(n10053, n1118, new_n20309);
nor_5  g17961(n25974, new_n3009, new_n20310);
nor_5  g17962(new_n12584, n8399, new_n20311);
nor_5  g17963(new_n3975, n1630, new_n20312);
nor_5  g17964(n9507, new_n12586, new_n20313);
nand_5 g17965(n26979, new_n12671, new_n20314);
nor_5  g17966(new_n20314, new_n20313, new_n20315);
nor_5  g17967(new_n20315, new_n20312, new_n20316);
nor_5  g17968(new_n20316, new_n20311, new_n20317);
nor_5  g17969(new_n20317, new_n20310, new_n20318);
and_5  g17970(new_n20318, new_n20309, new_n20319);
nor_5  g17971(new_n20319, new_n20308, new_n20320);
nor_5  g17972(new_n20320, new_n20307, new_n20321);
nor_5  g17973(new_n20321, new_n20305, new_n20322);
xnor_4 g17974(new_n20322, new_n20304, new_n20323);
xnor_4 g17975(new_n20323, new_n20303, new_n20324);
xnor_4 g17976(new_n20320, new_n20307, new_n20325);
xnor_4 g17977(new_n20298, new_n20297, new_n20326);
nor_5  g17978(new_n20326, new_n20325, new_n20327);
not_8  g17979(new_n20327, new_n20328);
xnor_4 g17980(new_n20295, new_n2404, new_n20329);
xnor_4 g17981(new_n20318, new_n20309, new_n20330_1);
not_8  g17982(new_n20330_1, new_n20331);
nor_5  g17983(new_n20331, new_n20329, new_n20332);
xnor_4 g17984(new_n20331, new_n20329, new_n20333_1);
xnor_4 g17985(n25974, n8399, new_n20334);
xnor_4 g17986(new_n20334, new_n20316, new_n20335);
not_8  g17987(new_n20335, new_n20336);
nor_5  g17988(new_n20336, new_n20252, new_n20337);
xnor_4 g17989(new_n20335, new_n20252, new_n20338);
not_8  g17990(new_n20338, new_n20339);
xnor_4 g17991(n26979, n1451, new_n20340);
nor_5  g17992(new_n20340, new_n19467_1, new_n20341);
xnor_4 g17993(n9507, n1630, new_n20342);
xnor_4 g17994(new_n20342, new_n20314, new_n20343);
not_8  g17995(new_n20343, new_n20344);
nor_5  g17996(new_n20344, new_n20341, new_n20345);
xnor_4 g17997(new_n20343, new_n20341, new_n20346);
not_8  g17998(new_n20346, new_n20347);
nor_5  g17999(new_n20347, new_n19480, new_n20348);
nor_5  g18000(new_n20348, new_n20345, new_n20349_1);
nor_5  g18001(new_n20349_1, new_n20339, new_n20350);
nor_5  g18002(new_n20350, new_n20337, new_n20351);
nor_5  g18003(new_n20351, new_n20333_1, new_n20352);
nor_5  g18004(new_n20352, new_n20332, new_n20353);
not_8  g18005(new_n20326, new_n20354);
xnor_4 g18006(new_n20354, new_n20325, new_n20355_1);
nand_5 g18007(new_n20355_1, new_n20353, new_n20356);
nand_5 g18008(new_n20356, new_n20328, new_n20357);
xnor_4 g18009(new_n20357, new_n20324, n5833);
xnor_4 g18010(new_n13282, new_n13252, n5840);
xor_4  g18011(new_n20149_1, new_n20148, n5841);
xnor_4 g18012(new_n13766, new_n13764_1, n5850);
xnor_4 g18013(new_n20225, new_n20214, n5903);
xnor_4 g18014(new_n17554, new_n7227, new_n20363);
not_8  g18015(new_n20363, new_n20364);
nand_5 g18016(new_n17559, n19472, new_n20365);
nand_5 g18017(new_n19622, new_n19607, new_n20366_1);
nand_5 g18018(new_n20366_1, new_n20365, new_n20367);
xnor_4 g18019(new_n20367, new_n20364, new_n20368);
nand_5 g18020(new_n19586, new_n6659_1, new_n20369);
xnor_4 g18021(new_n20369, n26752, new_n20370);
xnor_4 g18022(new_n20370, new_n9360, new_n20371);
nand_5 g18023(new_n19587, new_n9366, new_n20372);
nand_5 g18024(new_n19605, new_n19588, new_n20373);
nand_5 g18025(new_n20373, new_n20372, new_n20374);
xnor_4 g18026(new_n20374, new_n20371, new_n20375);
xnor_4 g18027(new_n20375, new_n20368, new_n20376);
not_8  g18028(new_n19606, new_n20377);
nand_5 g18029(new_n19623_1, new_n20377, new_n20378);
nand_5 g18030(new_n19650, new_n19624, new_n20379);
nand_5 g18031(new_n20379, new_n20378, new_n20380);
xnor_4 g18032(new_n20380, new_n20376, n5904);
xnor_4 g18033(n27089, n6814, new_n20382);
or_5   g18034(new_n9535, n11841, new_n20383);
xnor_4 g18035(n19701, n11841, new_n20384);
or_5   g18036(new_n9538, n10710, new_n20385_1);
xnor_4 g18037(n23529, n10710, new_n20386);
or_5   g18038(new_n9541, n20929, new_n20387);
xnor_4 g18039(n24620, n20929, new_n20388_1);
nor_5  g18040(n8006, new_n2955, new_n20389);
xnor_4 g18041(n8006, n5211, new_n20390);
nor_5  g18042(n25074, new_n9546, new_n20391);
not_8  g18043(new_n20391, new_n20392);
xnor_4 g18044(n25074, n12956, new_n20393);
nor_5  g18045(n18295, new_n4521, new_n20394);
nor_5  g18046(new_n2963, n16396, new_n20395);
nor_5  g18047(new_n4525, n6502, new_n20396);
nor_5  g18048(n9399, new_n9553, new_n20397);
nor_5  g18049(n15780, new_n3078, new_n20398);
not_8  g18050(new_n20398, new_n20399);
nor_5  g18051(new_n20399, new_n20397, new_n20400);
nor_5  g18052(new_n20400, new_n20396, new_n20401);
nor_5  g18053(new_n20401, new_n20395, new_n20402_1);
nor_5  g18054(new_n20402_1, new_n20394, new_n20403_1);
nand_5 g18055(new_n20403_1, new_n20393, new_n20404);
nand_5 g18056(new_n20404, new_n20392, new_n20405);
and_5  g18057(new_n20405, new_n20390, new_n20406);
nor_5  g18058(new_n20406, new_n20389, new_n20407);
not_8  g18059(new_n20407, new_n20408);
nand_5 g18060(new_n20408, new_n20388_1, new_n20409_1);
nand_5 g18061(new_n20409_1, new_n20387, new_n20410);
nand_5 g18062(new_n20410, new_n20386, new_n20411_1);
nand_5 g18063(new_n20411_1, new_n20385_1, new_n20412);
nand_5 g18064(new_n20412, new_n20384, new_n20413);
nand_5 g18065(new_n20413, new_n20383, new_n20414);
xnor_4 g18066(new_n20414, new_n20382, new_n20415);
xnor_4 g18067(new_n20415, new_n10830, new_n20416);
xnor_4 g18068(new_n20412, new_n20384, new_n20417);
nand_5 g18069(new_n20417, new_n10833, new_n20418);
xnor_4 g18070(new_n20417, new_n10835, new_n20419);
xnor_4 g18071(new_n20410, new_n20386, new_n20420);
nand_5 g18072(new_n20420, new_n10838, new_n20421);
xnor_4 g18073(new_n20420, new_n10840, new_n20422);
xnor_4 g18074(new_n20408, new_n20388_1, new_n20423);
nand_5 g18075(new_n20423, new_n10843, new_n20424_1);
not_8  g18076(new_n20390, new_n20425);
xnor_4 g18077(new_n20405, new_n20425, new_n20426);
not_8  g18078(new_n20426, new_n20427);
nand_5 g18079(new_n20427, new_n10848, new_n20428);
xnor_4 g18080(new_n20426, new_n10848, new_n20429_1);
xnor_4 g18081(new_n20403_1, new_n20393, new_n20430);
not_8  g18082(new_n20430, new_n20431);
nor_5  g18083(new_n20431, new_n10852, new_n20432);
not_8  g18084(new_n20432, new_n20433);
xnor_4 g18085(n18295, n16396, new_n20434);
xnor_4 g18086(new_n20434, new_n20401, new_n20435);
not_8  g18087(new_n20435, new_n20436_1);
nor_5  g18088(new_n20436_1, new_n10858, new_n20437);
not_8  g18089(new_n20437, new_n20438);
xnor_4 g18090(new_n20436_1, new_n10857, new_n20439);
xnor_4 g18091(n15780, n2088, new_n20440);
nor_5  g18092(new_n20440, new_n10865, new_n20441_1);
xnor_4 g18093(n9399, n6502, new_n20442);
xnor_4 g18094(new_n20442, new_n20399, new_n20443);
not_8  g18095(new_n20443, new_n20444);
and_5  g18096(new_n20444, new_n20441_1, new_n20445_1);
xnor_4 g18097(new_n20443, new_n20441_1, new_n20446);
and_5  g18098(new_n20446, new_n10872, new_n20447);
nor_5  g18099(new_n20447, new_n20445_1, new_n20448);
nand_5 g18100(new_n20448, new_n20439, new_n20449);
nand_5 g18101(new_n20449, new_n20438, new_n20450_1);
xnor_4 g18102(new_n20431, new_n10851_1, new_n20451);
nand_5 g18103(new_n20451, new_n20450_1, new_n20452);
nand_5 g18104(new_n20452, new_n20433, new_n20453);
nand_5 g18105(new_n20453, new_n20429_1, new_n20454);
nand_5 g18106(new_n20454, new_n20428, new_n20455_1);
xnor_4 g18107(new_n20423, new_n10883, new_n20456);
nand_5 g18108(new_n20456, new_n20455_1, new_n20457);
nand_5 g18109(new_n20457, new_n20424_1, new_n20458);
nand_5 g18110(new_n20458, new_n20422, new_n20459);
nand_5 g18111(new_n20459, new_n20421, new_n20460);
nand_5 g18112(new_n20460, new_n20419, new_n20461);
nand_5 g18113(new_n20461, new_n20418, new_n20462);
xnor_4 g18114(new_n20462, new_n20416, n5911);
xnor_4 g18115(new_n12672, new_n4080, n5936);
xnor_4 g18116(new_n10686, new_n10640, n5943);
xnor_4 g18117(new_n15185, new_n15150, n5964);
not_8  g18118(new_n16966, new_n20467);
nor_5  g18119(new_n16977, n11184, new_n20468);
not_8  g18120(new_n20468, new_n20469);
nor_5  g18121(new_n5322, n23146, new_n20470_1);
not_8  g18122(new_n20470_1, new_n20471);
nor_5  g18123(new_n5326, n17968, new_n20472);
nand_5 g18124(new_n20472, new_n5340, new_n20473);
nand_5 g18125(new_n20473, new_n20471, new_n20474);
nand_5 g18126(new_n20474, new_n5337_1, new_n20475);
nand_5 g18127(new_n20475, new_n20469, new_n20476);
nor_5  g18128(new_n20476, new_n16972, new_n20477);
not_8  g18129(new_n20477, new_n20478_1);
nand_5 g18130(new_n20476, new_n16983, new_n20479);
nand_5 g18131(new_n20479, n8255, new_n20480);
nand_5 g18132(new_n20480, new_n20478_1, new_n20481);
nand_5 g18133(new_n20481, new_n20467, new_n20482);
not_8  g18134(new_n20482, new_n20483);
nor_5  g18135(new_n20481, new_n16969, new_n20484);
nor_5  g18136(new_n20484, new_n16968_1, new_n20485);
nor_5  g18137(new_n20485, new_n20483, new_n20486);
nor_5  g18138(new_n20486, new_n16961, new_n20487);
not_8  g18139(new_n20487, new_n20488);
nand_5 g18140(new_n20486, new_n16965, new_n20489_1);
nand_5 g18141(new_n20489_1, n12380, new_n20490_1);
nand_5 g18142(new_n20490_1, new_n20488, new_n20491);
nand_5 g18143(new_n20491, new_n16958, new_n20492);
not_8  g18144(new_n20492, new_n20493);
not_8  g18145(n8694, new_n20494);
nor_5  g18146(new_n20491, new_n16991, new_n20495_1);
nor_5  g18147(new_n20495_1, new_n20494, new_n20496);
nor_5  g18148(new_n20496, new_n20493, new_n20497);
not_8  g18149(new_n20497, new_n20498);
nand_5 g18150(new_n20498, new_n16955, new_n20499);
nand_5 g18151(new_n20497, new_n16995, new_n20500);
nand_5 g18152(new_n20500, n15602, new_n20501);
nand_5 g18153(new_n20501, new_n20499, new_n20502);
xnor_4 g18154(new_n20502, new_n16954_1, new_n20503);
xnor_4 g18155(new_n20503, new_n3313, new_n20504);
xnor_4 g18156(new_n20498, new_n16995, new_n20505);
not_8  g18157(new_n20505, new_n20506);
nor_5  g18158(new_n20506, new_n3319, new_n20507);
not_8  g18159(new_n20507, new_n20508);
xnor_4 g18160(new_n20505, new_n3319, new_n20509);
xnor_4 g18161(new_n20491, new_n16991, new_n20510);
nor_5  g18162(new_n20510, new_n3324_1, new_n20511);
not_8  g18163(new_n20511, new_n20512);
xnor_4 g18164(new_n20510, new_n3324_1, new_n20513);
not_8  g18165(new_n20513, new_n20514);
xnor_4 g18166(new_n20486, new_n16964, new_n20515_1);
not_8  g18167(new_n20515_1, new_n20516);
nor_5  g18168(new_n20516, new_n3329, new_n20517);
not_8  g18169(new_n20517, new_n20518);
xnor_4 g18170(new_n20515_1, new_n3329, new_n20519);
xnor_4 g18171(new_n20481, new_n16970, new_n20520);
not_8  g18172(new_n20520, new_n20521);
nor_5  g18173(new_n20521, new_n3334, new_n20522);
xnor_4 g18174(new_n20520, new_n3334, new_n20523);
not_8  g18175(new_n20523, new_n20524);
xnor_4 g18176(new_n20476, new_n16984, new_n20525);
not_8  g18177(new_n20525, new_n20526);
nor_5  g18178(new_n20526, new_n3339, new_n20527);
xnor_4 g18179(new_n20525, new_n3339, new_n20528);
not_8  g18180(new_n20528, new_n20529);
xnor_4 g18181(new_n20474, new_n16980, new_n20530);
not_8  g18182(new_n20530, new_n20531);
nor_5  g18183(new_n20531, new_n3344, new_n20532);
xnor_4 g18184(new_n20530, new_n3344, new_n20533_1);
not_8  g18185(new_n20533_1, new_n20534);
xnor_4 g18186(new_n20472, new_n5328, new_n20535);
and_5  g18187(new_n20535, new_n3355, new_n20536);
nor_5  g18188(new_n5349, new_n3351, new_n20537);
xnor_4 g18189(new_n20535, new_n3495, new_n20538);
not_8  g18190(new_n20538, new_n20539);
nor_5  g18191(new_n20539, new_n20537, new_n20540);
nor_5  g18192(new_n20540, new_n20536, new_n20541);
nor_5  g18193(new_n20541, new_n20534, new_n20542);
nor_5  g18194(new_n20542, new_n20532, new_n20543);
nor_5  g18195(new_n20543, new_n20529, new_n20544);
nor_5  g18196(new_n20544, new_n20527, new_n20545);
nor_5  g18197(new_n20545, new_n20524, new_n20546);
nor_5  g18198(new_n20546, new_n20522, new_n20547);
not_8  g18199(new_n20547, new_n20548);
nand_5 g18200(new_n20548, new_n20519, new_n20549);
nand_5 g18201(new_n20549, new_n20518, new_n20550);
nand_5 g18202(new_n20550, new_n20514, new_n20551);
nand_5 g18203(new_n20551, new_n20512, new_n20552);
nand_5 g18204(new_n20552, new_n20509, new_n20553);
nand_5 g18205(new_n20553, new_n20508, new_n20554);
xnor_4 g18206(new_n20554, new_n20504, n5980);
xnor_4 g18207(new_n11967, new_n11941, n6012);
nand_5 g18208(new_n10764, new_n9530, new_n20557);
xnor_4 g18209(new_n10763_1, new_n9530, new_n20558);
not_8  g18210(new_n10767, new_n20559);
nand_5 g18211(new_n20559, new_n2941, new_n20560);
xnor_4 g18212(new_n10767, new_n2941, new_n20561);
nand_5 g18213(new_n10771, new_n9535, new_n20562);
xnor_4 g18214(new_n10771, n19701, new_n20563);
nand_5 g18215(new_n9868, new_n9538, new_n20564);
nand_5 g18216(new_n9907, new_n9869, new_n20565);
nand_5 g18217(new_n20565, new_n20564, new_n20566);
nand_5 g18218(new_n20566, new_n20563, new_n20567);
nand_5 g18219(new_n20567, new_n20562, new_n20568);
nand_5 g18220(new_n20568, new_n20561, new_n20569);
nand_5 g18221(new_n20569, new_n20560, new_n20570);
nand_5 g18222(new_n20570, new_n20558, new_n20571);
nand_5 g18223(new_n20571, new_n20557, new_n20572);
nor_5  g18224(new_n20572, new_n10757, new_n20573);
not_8  g18225(new_n20573, new_n20574);
nor_5  g18226(new_n15000, n3582, new_n20575);
xnor_4 g18227(new_n15000, n3582, new_n20576);
not_8  g18228(new_n15005, new_n20577);
nor_5  g18229(new_n20577, n2145, new_n20578);
xnor_4 g18230(new_n15005, new_n6312, new_n20579);
nor_5  g18231(new_n15008, n5031, new_n20580);
xnor_4 g18232(new_n15008, n5031, new_n20581);
nor_5  g18233(new_n9938_1, new_n8147, new_n20582_1);
nor_5  g18234(new_n9975, new_n9940, new_n20583);
nor_5  g18235(new_n20583, new_n20582_1, new_n20584);
not_8  g18236(new_n20584, new_n20585);
nor_5  g18237(new_n20585, new_n20581, new_n20586);
nor_5  g18238(new_n20586, new_n20580, new_n20587);
nor_5  g18239(new_n20587, new_n20579, new_n20588);
nor_5  g18240(new_n20588, new_n20578, new_n20589);
nor_5  g18241(new_n20589, new_n20576, new_n20590_1);
nor_5  g18242(new_n20590_1, new_n20575, new_n20591);
nand_5 g18243(new_n20591, new_n15051, new_n20592);
xnor_4 g18244(new_n20592, new_n20574, new_n20593);
not_8  g18245(new_n10757, new_n20594);
xnor_4 g18246(new_n20572, new_n20594, new_n20595);
not_8  g18247(new_n20595, new_n20596);
xnor_4 g18248(new_n20591, new_n15051, new_n20597);
not_8  g18249(new_n20597, new_n20598);
nand_5 g18250(new_n20598, new_n20596, new_n20599);
xnor_4 g18251(new_n20597, new_n20596, new_n20600);
not_8  g18252(new_n20558, new_n20601);
xnor_4 g18253(new_n20570, new_n20601, new_n20602_1);
not_8  g18254(new_n20576, new_n20603);
xnor_4 g18255(new_n20589, new_n20603, new_n20604_1);
not_8  g18256(new_n20604_1, new_n20605);
nand_5 g18257(new_n20605, new_n20602_1, new_n20606);
xnor_4 g18258(new_n20604_1, new_n20602_1, new_n20607);
not_8  g18259(new_n20561, new_n20608);
xnor_4 g18260(new_n20568, new_n20608, new_n20609_1);
not_8  g18261(new_n20579, new_n20610);
xnor_4 g18262(new_n20587, new_n20610, new_n20611);
not_8  g18263(new_n20611, new_n20612);
nand_5 g18264(new_n20612, new_n20609_1, new_n20613);
xnor_4 g18265(new_n20611, new_n20609_1, new_n20614);
not_8  g18266(new_n20563, new_n20615);
xnor_4 g18267(new_n20566, new_n20615, new_n20616);
xnor_4 g18268(new_n20584, new_n20581, new_n20617);
not_8  g18269(new_n20617, new_n20618);
nand_5 g18270(new_n20618, new_n20616, new_n20619);
xnor_4 g18271(new_n20617, new_n20616, new_n20620);
not_8  g18272(new_n9976, new_n20621);
nand_5 g18273(new_n20621, new_n9908, new_n20622);
nand_5 g18274(new_n10023, new_n9977, new_n20623_1);
nand_5 g18275(new_n20623_1, new_n20622, new_n20624);
nand_5 g18276(new_n20624, new_n20620, new_n20625);
nand_5 g18277(new_n20625, new_n20619, new_n20626);
nand_5 g18278(new_n20626, new_n20614, new_n20627);
nand_5 g18279(new_n20627, new_n20613, new_n20628);
nand_5 g18280(new_n20628, new_n20607, new_n20629_1);
nand_5 g18281(new_n20629_1, new_n20606, new_n20630);
nand_5 g18282(new_n20630, new_n20600, new_n20631);
nand_5 g18283(new_n20631, new_n20599, new_n20632);
xnor_4 g18284(new_n20632, new_n20593, n6022);
xnor_4 g18285(new_n20230, new_n20211, n6031);
nand_5 g18286(new_n17630, new_n11678, new_n20635);
xnor_4 g18287(new_n20635, new_n11675, new_n20636);
xnor_4 g18288(new_n20636, new_n9274, new_n20637);
not_8  g18289(new_n17631, new_n20638);
nand_5 g18290(new_n20638, new_n9341, new_n20639);
nand_5 g18291(new_n17673, new_n17632, new_n20640);
nand_5 g18292(new_n20640, new_n20639, new_n20641);
xnor_4 g18293(new_n20641, new_n20637, new_n20642);
xnor_4 g18294(new_n20642, new_n5905, new_n20643);
nor_5  g18295(new_n17674, n26797, new_n20644);
not_8  g18296(new_n17675, new_n20645);
nor_5  g18297(new_n17714, new_n20645, new_n20646);
nor_5  g18298(new_n20646, new_n20644, new_n20647);
xnor_4 g18299(new_n20647, new_n20643, new_n20648);
xnor_4 g18300(new_n20648, new_n8641, new_n20649);
nand_5 g18301(new_n17715, new_n8648, new_n20650);
nand_5 g18302(new_n17760, new_n17716, new_n20651);
nand_5 g18303(new_n20651, new_n20650, new_n20652);
xnor_4 g18304(new_n20652, new_n20649, n6044);
nor_5  g18305(new_n9714, new_n9670, new_n20654);
nor_5  g18306(new_n9785, new_n9715, new_n20655);
nor_5  g18307(new_n20655, new_n20654, new_n20656);
or_5   g18308(new_n9668, n4306, new_n20657);
xnor_4 g18309(new_n19155, new_n20657, new_n20658_1);
not_8  g18310(new_n20658_1, new_n20659);
xnor_4 g18311(new_n20659, new_n20656, new_n20660);
nor_5  g18312(new_n20660, new_n4735, new_n20661_1);
not_8  g18313(new_n20661_1, new_n20662);
xnor_4 g18314(new_n20660, new_n4739, new_n20663);
nor_5  g18315(new_n9786, new_n4744, new_n20664);
not_8  g18316(new_n20664, new_n20665);
nand_5 g18317(new_n9836, new_n9787, new_n20666);
nand_5 g18318(new_n20666, new_n20665, new_n20667);
nand_5 g18319(new_n20667, new_n20663, new_n20668);
nand_5 g18320(new_n20668, new_n20662, new_n20669);
nand_5 g18321(new_n19154, new_n20657, new_n20670);
not_8  g18322(new_n20670, new_n20671);
nand_5 g18323(new_n20671, new_n20656, new_n20672);
nor_5  g18324(new_n20672, new_n4610, new_n20673_1);
nand_5 g18325(new_n20673_1, new_n20669, new_n20674);
not_8  g18326(new_n20669, new_n20675);
and_5  g18327(new_n20672, new_n4610, new_n20676);
nand_5 g18328(new_n20676, new_n20675, new_n20677);
nand_5 g18329(new_n20677, new_n20674, n6046);
xnor_4 g18330(n17077, n7437, new_n20679);
not_8  g18331(new_n20679, new_n20680_1);
or_5   g18332(n26510, new_n2947, new_n20681);
xnor_4 g18333(n26510, n20700, new_n20682);
or_5   g18334(n23068, new_n2951, new_n20683);
not_8  g18335(new_n20322, new_n20684);
nand_5 g18336(new_n20684, new_n20304, new_n20685_1);
nand_5 g18337(new_n20685_1, new_n20683, new_n20686);
nand_5 g18338(new_n20686, new_n20682, new_n20687);
nand_5 g18339(new_n20687, new_n20681, new_n20688);
xnor_4 g18340(new_n20688, new_n20680_1, new_n20689);
xnor_4 g18341(n21997, new_n7362, new_n20690);
not_8  g18342(new_n20690, new_n20691_1);
or_5   g18343(new_n16894, new_n7365, new_n20692);
not_8  g18344(new_n20692, new_n20693);
nor_5  g18345(n25119, n21934, new_n20694);
nor_5  g18346(n18901, n1163, new_n20695);
not_8  g18347(new_n20269, new_n20696_1);
nor_5  g18348(new_n20283, new_n20696_1, new_n20697);
nor_5  g18349(new_n20697, new_n20695, new_n20698);
not_8  g18350(new_n20698, new_n20699);
nor_5  g18351(new_n20699, new_n20694, new_n20700_1);
nor_5  g18352(new_n20700_1, new_n20693, new_n20701);
xnor_4 g18353(new_n20701, new_n20691_1, new_n20702);
xnor_4 g18354(new_n20702, new_n7943_1, new_n20703);
xnor_4 g18355(n25119, new_n7365, new_n20704_1);
xnor_4 g18356(new_n20704_1, new_n20699, new_n20705_1);
nor_5  g18357(new_n20705_1, new_n2428, new_n20706);
not_8  g18358(new_n20706, new_n20707);
nor_5  g18359(new_n20284, new_n2466, new_n20708);
nand_5 g18360(new_n20301_1, new_n20285, new_n20709_1);
not_8  g18361(new_n20709_1, new_n20710);
nor_5  g18362(new_n20710, new_n20708, new_n20711);
xnor_4 g18363(new_n20705_1, new_n7933, new_n20712);
nand_5 g18364(new_n20712, new_n20711, new_n20713_1);
nand_5 g18365(new_n20713_1, new_n20707, new_n20714);
xnor_4 g18366(new_n20714, new_n20703, new_n20715);
xnor_4 g18367(new_n20715, new_n20689, new_n20716);
xnor_4 g18368(new_n20686, new_n20682, new_n20717);
xnor_4 g18369(new_n20712, new_n20711, new_n20718);
not_8  g18370(new_n20718, new_n20719);
nor_5  g18371(new_n20719, new_n20717, new_n20720);
not_8  g18372(new_n20720, new_n20721);
nor_5  g18373(new_n20323, new_n20303, new_n20722_1);
nor_5  g18374(new_n20357, new_n20324, new_n20723_1);
nor_5  g18375(new_n20723_1, new_n20722_1, new_n20724);
xnor_4 g18376(new_n20718, new_n20717, new_n20725);
nand_5 g18377(new_n20725, new_n20724, new_n20726);
nand_5 g18378(new_n20726, new_n20721, new_n20727);
xnor_4 g18379(new_n20727, new_n20716, n6084);
not_8  g18380(new_n10872, new_n20729);
xnor_4 g18381(new_n20446, new_n20729, n6160);
xnor_4 g18382(new_n20451, new_n20450_1, n6171);
or_5   g18383(n22359, new_n8422, new_n20732);
nand_5 g18384(new_n16112, new_n10546, new_n20733);
nand_5 g18385(new_n20733, new_n20732, new_n20734);
xnor_4 g18386(new_n20734, new_n10551, new_n20735);
xnor_4 g18387(n26264, n21905, new_n20736);
or_5   g18388(n22918, new_n8470, new_n20737);
xnor_4 g18389(n22918, n7841, new_n20738);
or_5   g18390(n25923, new_n8475, new_n20739);
xnor_4 g18391(n25923, n16812, new_n20740);
nand_5 g18392(n25068, new_n10461, new_n20741);
not_8  g18393(new_n19211, new_n20742);
nand_5 g18394(new_n20742, new_n19188, new_n20743);
nand_5 g18395(new_n20743, new_n20741, new_n20744);
nand_5 g18396(new_n20744, new_n20740, new_n20745);
nand_5 g18397(new_n20745, new_n20739, new_n20746);
nand_5 g18398(new_n20746, new_n20738, new_n20747);
nand_5 g18399(new_n20747, new_n20737, new_n20748_1);
xnor_4 g18400(new_n20748_1, new_n20736, new_n20749);
xnor_4 g18401(new_n20749, new_n16460_1, new_n20750);
not_8  g18402(new_n20738, new_n20751);
xnor_4 g18403(new_n20746, new_n20751, new_n20752);
nor_5  g18404(new_n20752, new_n16185_1, new_n20753);
xnor_4 g18405(new_n20752, new_n16185_1, new_n20754);
xnor_4 g18406(new_n20744, new_n20740, new_n20755);
nor_5  g18407(new_n20755, new_n16188, new_n20756);
not_8  g18408(new_n20756, new_n20757);
xnor_4 g18409(new_n20755, new_n16187, new_n20758);
nand_5 g18410(new_n19212, new_n16197, new_n20759);
nand_5 g18411(new_n19240, new_n19213, new_n20760);
nand_5 g18412(new_n20760, new_n20759, new_n20761_1);
nand_5 g18413(new_n20761_1, new_n20758, new_n20762);
nand_5 g18414(new_n20762, new_n20757, new_n20763);
nor_5  g18415(new_n20763, new_n20754, new_n20764);
nor_5  g18416(new_n20764, new_n20753, new_n20765);
xnor_4 g18417(new_n20765, new_n20750, new_n20766);
xnor_4 g18418(new_n20766, new_n20735, new_n20767);
not_8  g18419(new_n16113, new_n20768);
xnor_4 g18420(new_n20763, new_n20754, new_n20769);
not_8  g18421(new_n20769, new_n20770);
nand_5 g18422(new_n20770, new_n20768, new_n20771);
xnor_4 g18423(new_n20769, new_n20768, new_n20772);
not_8  g18424(new_n20758, new_n20773);
xnor_4 g18425(new_n20761_1, new_n20773, new_n20774_1);
not_8  g18426(new_n20774_1, new_n20775);
nand_5 g18427(new_n20775, new_n16117, new_n20776);
xnor_4 g18428(new_n20774_1, new_n16117, new_n20777);
nand_5 g18429(new_n19241, new_n16123, new_n20778);
nand_5 g18430(new_n19271, new_n19242, new_n20779);
nand_5 g18431(new_n20779, new_n20778, new_n20780);
nand_5 g18432(new_n20780, new_n20777, new_n20781);
nand_5 g18433(new_n20781, new_n20776, new_n20782);
nand_5 g18434(new_n20782, new_n20772, new_n20783);
nand_5 g18435(new_n20783, new_n20771, new_n20784);
xnor_4 g18436(new_n20784, new_n20767, n6183);
xnor_4 g18437(n14702, n14345, new_n20786);
not_8  g18438(new_n20786, new_n20787);
nor_5  g18439(new_n11203, n2999, new_n20788_1);
xnor_4 g18440(n11356, n2999, new_n20789);
not_8  g18441(new_n20789, new_n20790);
nor_5  g18442(new_n9683, n2547, new_n20791);
xnor_4 g18443(n3164, n2547, new_n20792);
nor_5  g18444(n10611, new_n11408, new_n20793);
not_8  g18445(new_n14952, new_n20794_1);
nor_5  g18446(new_n14961, new_n20794_1, new_n20795_1);
nor_5  g18447(new_n20795_1, new_n20793, new_n20796);
and_5  g18448(new_n20796, new_n20792, new_n20797);
nor_5  g18449(new_n20797, new_n20791, new_n20798);
nor_5  g18450(new_n20798, new_n20790, new_n20799);
nor_5  g18451(new_n20799, new_n20788_1, new_n20800);
xnor_4 g18452(new_n20800, new_n20787, new_n20801);
xnor_4 g18453(new_n20801, new_n9596, new_n20802);
xnor_4 g18454(new_n20798, new_n20789, new_n20803_1);
nor_5  g18455(new_n20803_1, new_n9602, new_n20804);
not_8  g18456(new_n20804, new_n20805);
xnor_4 g18457(new_n20803_1, new_n9603, new_n20806);
xnor_4 g18458(new_n20796, new_n20792, new_n20807);
not_8  g18459(new_n20807, new_n20808);
nor_5  g18460(new_n20808, new_n9609, new_n20809);
not_8  g18461(new_n20809, new_n20810);
xnor_4 g18462(new_n20807, new_n9609, new_n20811);
nand_5 g18463(new_n14962, new_n9614, new_n20812);
nand_5 g18464(new_n14983, new_n14963, new_n20813);
nand_5 g18465(new_n20813, new_n20812, new_n20814);
nand_5 g18466(new_n20814, new_n20811, new_n20815);
nand_5 g18467(new_n20815, new_n20810, new_n20816);
nand_5 g18468(new_n20816, new_n20806, new_n20817);
nand_5 g18469(new_n20817, new_n20805, new_n20818);
xor_4  g18470(new_n20818, new_n20802, n6189);
xnor_4 g18471(n20036, n15167, new_n20820);
nor_5  g18472(new_n6836, n11192, new_n20821);
nor_5  g18473(n21095, new_n4305, new_n20822);
nor_5  g18474(n9380, new_n15544, new_n20823);
not_8  g18475(new_n20823, new_n20824);
nor_5  g18476(new_n20824, new_n20822, new_n20825);
nor_5  g18477(new_n20825, new_n20821, new_n20826_1);
xnor_4 g18478(new_n20826_1, new_n20820, new_n20827);
xnor_4 g18479(new_n20827, new_n19253, new_n20828);
xnor_4 g18480(n9380, n8656, new_n20829);
nor_5  g18481(new_n20829, new_n19257, new_n20830);
xnor_4 g18482(n21095, n11192, new_n20831);
xnor_4 g18483(new_n20831, new_n20824, new_n20832);
not_8  g18484(new_n20832, new_n20833);
nor_5  g18485(new_n20833, new_n20830, new_n20834);
not_8  g18486(new_n20834, new_n20835);
xnor_4 g18487(new_n20832, new_n20830, new_n20836);
nand_5 g18488(new_n20836, new_n19261, new_n20837);
nand_5 g18489(new_n20837, new_n20835, new_n20838);
xnor_4 g18490(new_n20838, new_n20828, n6223);
xnor_4 g18491(new_n14980, new_n14970, n6233);
xnor_4 g18492(new_n19920, new_n19916_1, n6245);
xnor_4 g18493(new_n10875, new_n10864, n6248);
xnor_4 g18494(n21839, n16544, new_n20843);
or_5   g18495(n27089, new_n2941, new_n20844);
nand_5 g18496(new_n20414, new_n20382, new_n20845);
nand_5 g18497(new_n20845, new_n20844, new_n20846);
xnor_4 g18498(new_n20846, new_n20843, new_n20847);
xnor_4 g18499(new_n20847, new_n10823, new_n20848);
nand_5 g18500(new_n20415, new_n10828, new_n20849);
nand_5 g18501(new_n20462, new_n20416, new_n20850);
nand_5 g18502(new_n20850, new_n20849, new_n20851);
xnor_4 g18503(new_n20851, new_n20848, n6256);
xnor_4 g18504(new_n15850, new_n15834, n6271);
or_5   g18505(new_n8417_1, n13549, new_n20854);
not_8  g18506(n23493, new_n20855);
or_5   g18507(new_n20855, n8405, new_n20856);
nand_5 g18508(new_n20734, new_n10550, new_n20857);
nand_5 g18509(new_n20857, new_n20856, new_n20858);
nand_5 g18510(new_n20858, new_n10554, new_n20859);
nand_5 g18511(new_n20859, new_n20854, new_n20860);
not_8  g18512(new_n20860, new_n20861);
nor_5  g18513(n13951, new_n2717, new_n20862);
xnor_4 g18514(n13951, n2944, new_n20863);
not_8  g18515(new_n20863, new_n20864);
nor_5  g18516(n22793, new_n2720, new_n20865);
nor_5  g18517(new_n15883, new_n15859_1, new_n20866);
nor_5  g18518(new_n20866, new_n20865, new_n20867);
nor_5  g18519(new_n20867, new_n20864, new_n20868);
nor_5  g18520(new_n20868, new_n20862, new_n20869_1);
nand_5 g18521(new_n20869_1, new_n20861, new_n20870);
xnor_4 g18522(new_n20867, new_n20864, new_n20871);
xnor_4 g18523(new_n20858, new_n10610, new_n20872);
not_8  g18524(new_n20872, new_n20873);
nand_5 g18525(new_n20873, new_n20871, new_n20874);
xnor_4 g18526(new_n20872, new_n20871, new_n20875);
not_8  g18527(new_n20735, new_n20876);
nor_5  g18528(new_n20876, new_n15884_1, new_n20877);
xnor_4 g18529(new_n20876, new_n15884_1, new_n20878);
not_8  g18530(new_n15886, new_n20879_1);
nand_5 g18531(new_n20768, new_n20879_1, new_n20880);
not_8  g18532(new_n16114, new_n20881);
nand_5 g18533(new_n16139, new_n20881, new_n20882);
nand_5 g18534(new_n20882, new_n20880, new_n20883);
nor_5  g18535(new_n20883, new_n20878, new_n20884);
nor_5  g18536(new_n20884, new_n20877, new_n20885);
nand_5 g18537(new_n20885, new_n20875, new_n20886);
nand_5 g18538(new_n20886, new_n20874, new_n20887);
xnor_4 g18539(new_n20869_1, new_n20860, new_n20888);
nand_5 g18540(new_n20888, new_n20887, new_n20889);
nand_5 g18541(new_n20889, new_n20870, new_n20890);
nor_5  g18542(new_n13680, n1881, new_n20891);
xnor_4 g18543(n8827, n1881, new_n20892);
not_8  g18544(new_n20892, new_n20893);
nor_5  g18545(new_n13699, n5834, new_n20894);
nor_5  g18546(new_n20202, new_n20199, new_n20895);
nor_5  g18547(new_n20895, new_n20894, new_n20896);
nor_5  g18548(new_n20896, new_n20893, new_n20897);
nor_5  g18549(new_n20897, new_n20891, new_n20898);
not_8  g18550(new_n20898, new_n20899);
xnor_4 g18551(new_n20899, new_n20890, new_n20900);
not_8  g18552(new_n20888, new_n20901);
xnor_4 g18553(new_n20901, new_n20887, new_n20902);
nand_5 g18554(new_n20902, new_n20899, new_n20903);
xnor_4 g18555(new_n20902, new_n20898, new_n20904);
xnor_4 g18556(new_n20896, new_n20893, new_n20905);
not_8  g18557(new_n20875, new_n20906);
xnor_4 g18558(new_n20885, new_n20906, new_n20907);
nor_5  g18559(new_n20907, new_n20905, new_n20908);
xnor_4 g18560(new_n20883, new_n20878, new_n20909);
nand_5 g18561(new_n20909, new_n20203, new_n20910);
xnor_4 g18562(new_n20202, new_n20198, new_n20911);
xnor_4 g18563(new_n20909, new_n20911, new_n20912);
nor_5  g18564(new_n16409, new_n16140, new_n20913);
nor_5  g18565(new_n16432, new_n16410, new_n20914);
nor_5  g18566(new_n20914, new_n20913, new_n20915_1);
nand_5 g18567(new_n20915_1, new_n20912, new_n20916);
nand_5 g18568(new_n20916, new_n20910, new_n20917);
xnor_4 g18569(new_n20907, new_n20905, new_n20918);
nor_5  g18570(new_n20918, new_n20917, new_n20919);
nor_5  g18571(new_n20919, new_n20908, new_n20920);
nand_5 g18572(new_n20920, new_n20904, new_n20921);
nand_5 g18573(new_n20921, new_n20903, new_n20922);
xnor_4 g18574(new_n20922, new_n20900, n6276);
xnor_4 g18575(new_n19871, new_n19869, n6308);
xnor_4 g18576(new_n17856, new_n17842, n6311);
xnor_4 g18577(new_n17612, new_n17596, n6323);
nor_5  g18578(new_n6236, new_n6186, new_n20927);
not_8  g18579(new_n6237, new_n20928);
nor_5  g18580(new_n6306, new_n20928, new_n20929_1);
nor_5  g18581(new_n20929_1, new_n20927, new_n20930);
not_8  g18582(new_n20930, new_n20931);
nand_5 g18583(new_n14286, new_n14691, new_n20932);
not_8  g18584(new_n20932, new_n20933);
nand_5 g18585(new_n20933, new_n20931, new_n20934);
nor_5  g18586(new_n14286, new_n14691, new_n20935_1);
nand_5 g18587(new_n20935_1, new_n20930, new_n20936_1);
nand_5 g18588(new_n20936_1, new_n20934, new_n20937);
nand_5 g18589(new_n20937, new_n19010, new_n20938);
xnor_4 g18590(new_n20937, new_n19011, new_n20939);
xnor_4 g18591(new_n14287, new_n14691, new_n20940);
xnor_4 g18592(new_n20940, new_n20931, new_n20941);
not_8  g18593(new_n20941, new_n20942);
nand_5 g18594(new_n20942, new_n19013, new_n20943);
xnor_4 g18595(new_n20941, new_n19013, new_n20944);
not_8  g18596(new_n6307, new_n20945);
nand_5 g18597(new_n6410, new_n20945, new_n20946_1);
nand_5 g18598(new_n6475, new_n6411, new_n20947);
nand_5 g18599(new_n20947, new_n20946_1, new_n20948);
nand_5 g18600(new_n20948, new_n20944, new_n20949);
nand_5 g18601(new_n20949, new_n20943, new_n20950);
nand_5 g18602(new_n20950, new_n20939, new_n20951);
nand_5 g18603(new_n20951, new_n20938, new_n20952);
nand_5 g18604(new_n20952, new_n20934, new_n20953);
not_8  g18605(new_n20953, n6330);
xnor_4 g18606(new_n9106, new_n9068, n6339);
xnor_4 g18607(new_n14944_1, new_n14917, n6354);
nor_5  g18608(new_n3304, n7335, new_n20957);
or_5   g18609(new_n3312, n5696, new_n20958);
xnor_4 g18610(new_n3312, new_n3168, new_n20959);
or_5   g18611(new_n3318, n13367, new_n20960);
xnor_4 g18612(new_n3321, n13367, new_n20961);
or_5   g18613(new_n3323, n932, new_n20962);
xnor_4 g18614(new_n3323, new_n3175, new_n20963);
or_5   g18615(new_n3328, n6691, new_n20964);
xnor_4 g18616(new_n3328, new_n3179, new_n20965);
nand_5 g18617(new_n3336, new_n3183, new_n20966);
xnor_4 g18618(new_n3333, new_n3183, new_n20967);
nand_5 g18619(new_n3341, new_n3187, new_n20968);
nand_5 g18620(new_n3346, new_n3191, new_n20969);
xnor_4 g18621(new_n3343_1, new_n3191, new_n20970);
not_8  g18622(n11121, new_n20971);
not_8  g18623(new_n3356, new_n20972);
nand_5 g18624(new_n20972, new_n20971, new_n20973);
not_8  g18625(new_n20973, new_n20974);
nand_5 g18626(n16217, n12315, new_n20975);
xnor_4 g18627(new_n3356, new_n20971, new_n20976);
and_5  g18628(new_n20976, new_n20975, new_n20977);
nor_5  g18629(new_n20977, new_n20974, new_n20978);
not_8  g18630(new_n20978, new_n20979);
nand_5 g18631(new_n20979, new_n20970, new_n20980);
nand_5 g18632(new_n20980, new_n20969, new_n20981);
xnor_4 g18633(new_n3338, new_n3187, new_n20982);
nand_5 g18634(new_n20982, new_n20981, new_n20983);
nand_5 g18635(new_n20983, new_n20968, new_n20984);
nand_5 g18636(new_n20984, new_n20967, new_n20985);
nand_5 g18637(new_n20985, new_n20966, new_n20986_1);
nand_5 g18638(new_n20986_1, new_n20965, new_n20987);
nand_5 g18639(new_n20987, new_n20964, new_n20988);
nand_5 g18640(new_n20988, new_n20963, new_n20989);
nand_5 g18641(new_n20989, new_n20962, new_n20990);
nand_5 g18642(new_n20990, new_n20961, new_n20991);
nand_5 g18643(new_n20991, new_n20960, new_n20992);
nand_5 g18644(new_n20992, new_n20959, new_n20993);
nand_5 g18645(new_n20993, new_n20958, new_n20994);
nor_5  g18646(new_n20994, new_n20957, new_n20995);
not_8  g18647(n7335, new_n20996);
nor_5  g18648(new_n3305, new_n20996, new_n20997);
nor_5  g18649(new_n20997, new_n3309, new_n20998);
not_8  g18650(new_n20998, new_n20999);
nor_5  g18651(new_n20999, new_n20995, new_n21000);
nand_5 g18652(new_n21000, new_n18041, new_n21001);
not_8  g18653(new_n21000, new_n21002);
nand_5 g18654(new_n21002, new_n18087, new_n21003);
xnor_4 g18655(new_n21000, new_n18087, new_n21004);
xnor_4 g18656(new_n3304, new_n20996, new_n21005);
xnor_4 g18657(new_n21005, new_n20994, new_n21006);
not_8  g18658(new_n21006, new_n21007);
nand_5 g18659(new_n21007, new_n18091, new_n21008_1);
xnor_4 g18660(new_n21006, new_n18091, new_n21009);
xnor_4 g18661(new_n20992, new_n20959, new_n21010);
not_8  g18662(new_n21010, new_n21011);
nand_5 g18663(new_n21011, new_n18100, new_n21012);
xnor_4 g18664(new_n21010, new_n18100, new_n21013);
xnor_4 g18665(new_n20990, new_n20961, new_n21014);
not_8  g18666(new_n21014, new_n21015);
nand_5 g18667(new_n21015, new_n18106, new_n21016);
xnor_4 g18668(new_n21014, new_n18106, new_n21017_1);
xnor_4 g18669(new_n20988, new_n20963, new_n21018);
not_8  g18670(new_n21018, new_n21019);
nand_5 g18671(new_n21019, new_n18112, new_n21020);
xnor_4 g18672(new_n21018, new_n18112, new_n21021);
xnor_4 g18673(new_n20986_1, new_n20965, new_n21022);
not_8  g18674(new_n21022, new_n21023);
nand_5 g18675(new_n21023, new_n18118, new_n21024);
xnor_4 g18676(new_n21022, new_n18118, new_n21025);
not_8  g18677(new_n20967, new_n21026);
xnor_4 g18678(new_n20984, new_n21026, new_n21027);
nand_5 g18679(new_n21027, new_n18124, new_n21028);
xnor_4 g18680(new_n21027, new_n18123, new_n21029);
xnor_4 g18681(new_n20982, new_n20981, new_n21030);
nor_5  g18682(new_n21030, new_n18128, new_n21031);
not_8  g18683(new_n21031, new_n21032);
xnor_4 g18684(new_n21030, new_n18127, new_n21033);
xnor_4 g18685(new_n20978, new_n20970, new_n21034_1);
nor_5  g18686(new_n21034_1, new_n18135, new_n21035);
xnor_4 g18687(new_n21034_1, new_n18135, new_n21036);
nor_5  g18688(new_n20976, new_n18139, new_n21037);
not_8  g18689(new_n21037, new_n21038);
nor_5  g18690(new_n20976, new_n20975, new_n21039);
nor_5  g18691(new_n21039, new_n20977, new_n21040);
nor_5  g18692(new_n21040, new_n18138, new_n21041);
not_8  g18693(new_n21041, new_n21042);
xnor_4 g18694(n16217, new_n3349_1, new_n21043);
and_5  g18695(new_n21043, new_n18146, new_n21044);
not_8  g18696(new_n21044, new_n21045);
nand_5 g18697(new_n21045, new_n21042, new_n21046_1);
nand_5 g18698(new_n21046_1, new_n21038, new_n21047);
nor_5  g18699(new_n21047, new_n21036, new_n21048);
nor_5  g18700(new_n21048, new_n21035, new_n21049);
nand_5 g18701(new_n21049, new_n21033, new_n21050);
nand_5 g18702(new_n21050, new_n21032, new_n21051);
nand_5 g18703(new_n21051, new_n21029, new_n21052);
nand_5 g18704(new_n21052, new_n21028, new_n21053);
nand_5 g18705(new_n21053, new_n21025, new_n21054);
nand_5 g18706(new_n21054, new_n21024, new_n21055);
nand_5 g18707(new_n21055, new_n21021, new_n21056);
nand_5 g18708(new_n21056, new_n21020, new_n21057);
nand_5 g18709(new_n21057, new_n21017_1, new_n21058);
nand_5 g18710(new_n21058, new_n21016, new_n21059);
nand_5 g18711(new_n21059, new_n21013, new_n21060);
nand_5 g18712(new_n21060, new_n21012, new_n21061);
nand_5 g18713(new_n21061, new_n21009, new_n21062_1);
nand_5 g18714(new_n21062_1, new_n21008_1, new_n21063);
nand_5 g18715(new_n21063, new_n21004, new_n21064);
nand_5 g18716(new_n21064, new_n21003, new_n21065);
nand_5 g18717(new_n21065, new_n21001, new_n21066);
nand_5 g18718(new_n21002, new_n18040, new_n21067);
nand_5 g18719(new_n21067, new_n21064, new_n21068);
nand_5 g18720(new_n21068, new_n21066, new_n21069);
not_8  g18721(new_n21069, n6375);
xnor_4 g18722(new_n20057, new_n20041, n6383);
xnor_4 g18723(new_n15367, new_n15324, n6407);
xnor_4 g18724(new_n9096, new_n9094, n6431);
xnor_4 g18725(new_n17441, new_n17436_1, n6437);
xnor_4 g18726(new_n4348, new_n4346, n6457);
xnor_4 g18727(new_n13054_1, new_n13021, n6465);
and_5  g18728(new_n18392, n3740, new_n21077);
nor_5  g18729(new_n18391, n3582, new_n21078_1);
nor_5  g18730(new_n18392, n3740, new_n21079);
nor_5  g18731(new_n18397, new_n21079, new_n21080);
nor_5  g18732(new_n21080, new_n21078_1, new_n21081);
not_8  g18733(new_n21081, new_n21082);
nor_5  g18734(new_n21082, new_n21077, new_n21083);
xnor_4 g18735(new_n21083, new_n8854, new_n21084);
nor_5  g18736(new_n18399, new_n8845, new_n21085);
not_8  g18737(new_n21085, new_n21086);
xnor_4 g18738(new_n18398, new_n8845, new_n21087);
nor_5  g18739(new_n15236, new_n3610, new_n21088);
nor_5  g18740(new_n15277, new_n15237, new_n21089);
nor_5  g18741(new_n21089, new_n21088, new_n21090);
nand_5 g18742(new_n21090, new_n21087, new_n21091);
nand_5 g18743(new_n21091, new_n21086, new_n21092);
xnor_4 g18744(new_n21092, new_n21084, new_n21093_1);
nor_5  g18745(new_n3736, n2743, new_n21094_1);
nor_5  g18746(new_n3742, new_n3675, new_n21095_1);
nor_5  g18747(new_n3741, n7026, new_n21096);
nor_5  g18748(new_n15312, new_n21096, new_n21097);
nor_5  g18749(new_n21097, new_n21095_1, new_n21098);
nor_5  g18750(new_n21098, new_n21094_1, new_n21099);
nor_5  g18751(new_n3735, n9259, new_n21100);
not_8  g18752(new_n3736, new_n21101);
nor_5  g18753(new_n21101, new_n14355, new_n21102);
nor_5  g18754(new_n21102, new_n21100, new_n21103);
not_8  g18755(new_n21103, new_n21104);
nor_5  g18756(new_n21104, new_n21099, new_n21105);
not_8  g18757(new_n21105, new_n21106);
xnor_4 g18758(new_n21106, new_n21093_1, new_n21107);
xnor_4 g18759(new_n21090, new_n21087, new_n21108);
not_8  g18760(new_n21108, new_n21109);
xnor_4 g18761(new_n3736, new_n14355, new_n21110);
xnor_4 g18762(new_n21110, new_n21098, new_n21111);
nor_5  g18763(new_n21111, new_n21109, new_n21112);
xnor_4 g18764(new_n21111, new_n21109, new_n21113);
nor_5  g18765(new_n15313, new_n15278, new_n21114);
nor_5  g18766(new_n15371, new_n15314, new_n21115);
nor_5  g18767(new_n21115, new_n21114, new_n21116);
nor_5  g18768(new_n21116, new_n21113, new_n21117);
nor_5  g18769(new_n21117, new_n21112, new_n21118);
xnor_4 g18770(new_n21118, new_n21107, n6470);
xnor_4 g18771(new_n12266, new_n12240, n6476);
xnor_4 g18772(new_n19533, new_n19523_1, n6506);
not_8  g18773(new_n17674, new_n21122);
not_8  g18774(new_n9938_1, new_n21123_1);
not_8  g18775(new_n9954, new_n21124);
nor_5  g18776(new_n9960, new_n9957, new_n21125);
not_8  g18777(new_n21125, new_n21126);
nor_5  g18778(new_n21126, new_n21124, new_n21127);
nand_5 g18779(new_n21127, new_n9950, new_n21128);
nor_5  g18780(new_n21128, new_n9945, new_n21129);
nand_5 g18781(new_n21129, new_n9941, new_n21130);
nor_5  g18782(new_n21130, new_n21123_1, new_n21131);
not_8  g18783(new_n21131, new_n21132);
nor_5  g18784(new_n21132, new_n15008, new_n21133);
xnor_4 g18785(new_n21133, new_n15005, new_n21134_1);
xnor_4 g18786(new_n21134_1, new_n10767, new_n21135);
not_8  g18787(new_n21135, new_n21136);
xnor_4 g18788(new_n21132, new_n15008, new_n21137);
nand_5 g18789(new_n21137, new_n10771, new_n21138_1);
xnor_4 g18790(new_n21137, new_n10772, new_n21139);
xnor_4 g18791(new_n21130, new_n21123_1, new_n21140);
nand_5 g18792(new_n21140, new_n9868, new_n21141);
xnor_4 g18793(new_n21140, new_n10776, new_n21142);
xnor_4 g18794(new_n21129, new_n9941, new_n21143);
nand_5 g18795(new_n21143, new_n9871, new_n21144);
xnor_4 g18796(new_n21143, new_n10778, new_n21145);
xnor_4 g18797(new_n21128, new_n9946_1, new_n21146);
not_8  g18798(new_n21146, new_n21147);
nand_5 g18799(new_n21147, new_n9874, new_n21148);
xnor_4 g18800(new_n21146, new_n9874, new_n21149);
xnor_4 g18801(new_n21127, new_n9950, new_n21150);
nand_5 g18802(new_n21150, new_n9877, new_n21151);
xnor_4 g18803(new_n21125, new_n9954, new_n21152);
nand_5 g18804(new_n21152, new_n9882, new_n21153);
xnor_4 g18805(new_n21152, new_n9882, new_n21154_1);
not_8  g18806(new_n21154_1, new_n21155);
nor_5  g18807(new_n9961, new_n9891, new_n21156);
nor_5  g18808(new_n21156, new_n10791, new_n21157_1);
nor_5  g18809(new_n9961, new_n9927, new_n21158);
nor_5  g18810(new_n21158, new_n21125, new_n21159);
not_8  g18811(new_n21156, new_n21160);
nor_5  g18812(new_n21160, new_n9857, new_n21161);
nor_5  g18813(new_n21161, new_n21157_1, new_n21162);
not_8  g18814(new_n21162, new_n21163);
nor_5  g18815(new_n21163, new_n21159, new_n21164);
nor_5  g18816(new_n21164, new_n21157_1, new_n21165);
not_8  g18817(new_n21165, new_n21166);
nand_5 g18818(new_n21166, new_n21155, new_n21167);
nand_5 g18819(new_n21167, new_n21153, new_n21168_1);
xnor_4 g18820(new_n21150, new_n9878, new_n21169);
nand_5 g18821(new_n21169, new_n21168_1, new_n21170);
nand_5 g18822(new_n21170, new_n21151, new_n21171);
nand_5 g18823(new_n21171, new_n21149, new_n21172);
nand_5 g18824(new_n21172, new_n21148, new_n21173_1);
nand_5 g18825(new_n21173_1, new_n21145, new_n21174);
nand_5 g18826(new_n21174, new_n21144, new_n21175);
nand_5 g18827(new_n21175, new_n21142, new_n21176_1);
nand_5 g18828(new_n21176_1, new_n21141, new_n21177);
nand_5 g18829(new_n21177, new_n21139, new_n21178);
nand_5 g18830(new_n21178, new_n21138_1, new_n21179);
xnor_4 g18831(new_n21179, new_n21136, new_n21180);
xnor_4 g18832(new_n21180, new_n21122, new_n21181);
not_8  g18833(new_n21139, new_n21182_1);
xnor_4 g18834(new_n21177, new_n21182_1, new_n21183);
not_8  g18835(new_n21183, new_n21184);
nor_5  g18836(new_n21184, new_n17676, new_n21185);
xnor_4 g18837(new_n21183, new_n17676, new_n21186);
not_8  g18838(new_n21186, new_n21187);
not_8  g18839(new_n21142, new_n21188);
xnor_4 g18840(new_n21175, new_n21188, new_n21189);
not_8  g18841(new_n21189, new_n21190);
nor_5  g18842(new_n21190, new_n17680, new_n21191);
xnor_4 g18843(new_n21189, new_n17680, new_n21192);
not_8  g18844(new_n21192, new_n21193_1);
xnor_4 g18845(new_n21173_1, new_n21145, new_n21194);
nor_5  g18846(new_n21194, new_n17683, new_n21195);
xnor_4 g18847(new_n21194, new_n17683, new_n21196);
not_8  g18848(new_n17686, new_n21197);
not_8  g18849(new_n21149, new_n21198);
xnor_4 g18850(new_n21171, new_n21198, new_n21199);
nor_5  g18851(new_n21199, new_n21197, new_n21200);
not_8  g18852(new_n21200, new_n21201);
xnor_4 g18853(new_n21169, new_n21168_1, new_n21202);
nand_5 g18854(new_n21202, new_n17689, new_n21203_1);
not_8  g18855(new_n21203_1, new_n21204);
xnor_4 g18856(new_n21202, new_n17689, new_n21205);
xnor_4 g18857(new_n21165, new_n21154_1, new_n21206);
nand_5 g18858(new_n21206, new_n17692, new_n21207);
not_8  g18859(new_n21207, new_n21208);
xnor_4 g18860(new_n21206, new_n17692, new_n21209);
not_8  g18861(new_n17695, new_n21210);
xnor_4 g18862(new_n21162, new_n21159, new_n21211);
nor_5  g18863(new_n21211, new_n21210, new_n21212);
xnor_4 g18864(new_n9960, new_n9891, new_n21213);
and_5  g18865(new_n21213, new_n17697, new_n21214);
xnor_4 g18866(new_n21211, new_n17695, new_n21215);
nand_5 g18867(new_n21215, new_n21214, new_n21216);
not_8  g18868(new_n21216, new_n21217);
nor_5  g18869(new_n21217, new_n21212, new_n21218);
nor_5  g18870(new_n21218, new_n21209, new_n21219);
nor_5  g18871(new_n21219, new_n21208, new_n21220);
nor_5  g18872(new_n21220, new_n21205, new_n21221);
nor_5  g18873(new_n21221, new_n21204, new_n21222_1);
not_8  g18874(new_n21222_1, new_n21223);
xnor_4 g18875(new_n21199, new_n17686, new_n21224);
nand_5 g18876(new_n21224, new_n21223, new_n21225_1);
nand_5 g18877(new_n21225_1, new_n21201, new_n21226_1);
nor_5  g18878(new_n21226_1, new_n21196, new_n21227);
nor_5  g18879(new_n21227, new_n21195, new_n21228);
nor_5  g18880(new_n21228, new_n21193_1, new_n21229);
nor_5  g18881(new_n21229, new_n21191, new_n21230);
nor_5  g18882(new_n21230, new_n21187, new_n21231);
nor_5  g18883(new_n21231, new_n21185, new_n21232);
xnor_4 g18884(new_n21232, new_n21181, n6514);
not_8  g18885(new_n12131_1, new_n21234);
nand_5 g18886(new_n12227, new_n21234, new_n21235);
nand_5 g18887(new_n12270, new_n12228_1, new_n21236);
nand_5 g18888(new_n21236, new_n21235, new_n21237);
not_8  g18889(new_n12226, new_n21238_1);
xnor_4 g18890(new_n12182, new_n12761, new_n21239);
not_8  g18891(new_n21239, new_n21240);
nor_5  g18892(new_n21240, new_n21238_1, new_n21241);
nor_5  g18893(new_n12182, new_n16062_1, new_n21242);
not_8  g18894(new_n21242, new_n21243);
nand_5 g18895(new_n21238_1, new_n21243, new_n21244);
nor_5  g18896(new_n21244, new_n21239, new_n21245);
nor_5  g18897(new_n21245, new_n21241, new_n21246);
xnor_4 g18898(new_n21246, new_n21237, n6542);
xnor_4 g18899(new_n16304, new_n16288, n6558);
xnor_4 g18900(new_n18995, new_n18993, n6560);
xnor_4 g18901(new_n6598, n10405, new_n21250);
nor_5  g18902(new_n6601, new_n4199, new_n21251);
xnor_4 g18903(new_n6601, n11302, new_n21252);
nor_5  g18904(new_n6606, n17090, new_n21253);
nor_5  g18905(new_n6609, new_n2575, new_n21254_1);
xnor_4 g18906(new_n6605, n17090, new_n21255);
not_8  g18907(new_n21255, new_n21256);
nor_5  g18908(new_n21256, new_n21254_1, new_n21257);
nor_5  g18909(new_n21257, new_n21253, new_n21258);
nand_5 g18910(new_n21258, new_n21252, new_n21259);
not_8  g18911(new_n21259, new_n21260);
nor_5  g18912(new_n21260, new_n21251, new_n21261);
xnor_4 g18913(new_n21261, new_n21250, new_n21262);
xnor_4 g18914(new_n21262, new_n10341, new_n21263);
not_8  g18915(new_n21263, new_n21264);
xnor_4 g18916(new_n21258, new_n21252, new_n21265);
and_5  g18917(new_n21265, new_n10344, new_n21266);
xnor_4 g18918(new_n21265, new_n10345_1, new_n21267);
not_8  g18919(new_n21267, new_n21268);
xnor_4 g18920(new_n21255, new_n21254_1, new_n21269);
and_5  g18921(new_n21269, new_n10351, new_n21270);
nor_5  g18922(new_n19023, new_n10354, new_n21271);
not_8  g18923(new_n21271, new_n21272);
xnor_4 g18924(new_n21269, new_n10350, new_n21273);
not_8  g18925(new_n21273, new_n21274);
nor_5  g18926(new_n21274, new_n21272, new_n21275);
nor_5  g18927(new_n21275, new_n21270, new_n21276_1);
nor_5  g18928(new_n21276_1, new_n21268, new_n21277);
nor_5  g18929(new_n21277, new_n21266, new_n21278);
xnor_4 g18930(new_n21278, new_n21264, n6567);
nor_5  g18931(new_n14525, n8324, new_n21280);
nand_5 g18932(new_n21280, new_n8585, new_n21281);
nor_5  g18933(new_n21281, n9445, new_n21282);
nand_5 g18934(new_n21282, new_n8577, new_n21283);
xnor_4 g18935(new_n21283, new_n8573, new_n21284);
not_8  g18936(new_n21284, new_n21285);
xnor_4 g18937(new_n21285, new_n4663, new_n21286);
not_8  g18938(new_n21286, new_n21287_1);
xnor_4 g18939(new_n21282, new_n8577, new_n21288);
nand_5 g18940(new_n21288, new_n4672, new_n21289);
xnor_4 g18941(new_n21288, new_n4671, new_n21290);
xnor_4 g18942(new_n21281, n9445, new_n21291);
nand_5 g18943(new_n21291, new_n4677, new_n21292);
xnor_4 g18944(new_n21291, new_n4676, new_n21293);
xnor_4 g18945(new_n21280, n1279, new_n21294);
not_8  g18946(new_n21294, new_n21295);
nand_5 g18947(new_n21295, new_n4683, new_n21296);
xnor_4 g18948(new_n21295, new_n4682, new_n21297);
nand_5 g18949(new_n14527, new_n4686, new_n21298_1);
nand_5 g18950(new_n14553, new_n14528, new_n21299);
nand_5 g18951(new_n21299, new_n21298_1, new_n21300);
nand_5 g18952(new_n21300, new_n21297, new_n21301);
nand_5 g18953(new_n21301, new_n21296, new_n21302_1);
nand_5 g18954(new_n21302_1, new_n21293, new_n21303);
nand_5 g18955(new_n21303, new_n21292, new_n21304);
nand_5 g18956(new_n21304, new_n21290, new_n21305);
nand_5 g18957(new_n21305, new_n21289, new_n21306);
xnor_4 g18958(new_n21306, new_n21287_1, new_n21307);
xnor_4 g18959(new_n8574, n23272, new_n21308);
nand_5 g18960(new_n8578, new_n4552_1, new_n21309);
xnor_4 g18961(new_n8578, n11481, new_n21310);
nand_5 g18962(new_n8582, new_n4556, new_n21311);
xnor_4 g18963(new_n8582, n16439, new_n21312);
nand_5 g18964(new_n8586, new_n4560, new_n21313);
nor_5  g18965(new_n8590, new_n4564, new_n21314);
nor_5  g18966(new_n14574, new_n14555, new_n21315);
nor_5  g18967(new_n21315, new_n21314, new_n21316);
xnor_4 g18968(new_n8586, n15241, new_n21317_1);
nand_5 g18969(new_n21317_1, new_n21316, new_n21318);
nand_5 g18970(new_n21318, new_n21313, new_n21319);
nand_5 g18971(new_n21319, new_n21312, new_n21320);
nand_5 g18972(new_n21320, new_n21311, new_n21321);
nand_5 g18973(new_n21321, new_n21310, new_n21322);
nand_5 g18974(new_n21322, new_n21309, new_n21323);
xnor_4 g18975(new_n21323, new_n21308, new_n21324);
xnor_4 g18976(new_n21324, new_n21307, new_n21325);
not_8  g18977(new_n21290, new_n21326);
xnor_4 g18978(new_n21304, new_n21326, new_n21327);
xnor_4 g18979(new_n21321, new_n21310, new_n21328);
not_8  g18980(new_n21328, new_n21329);
nand_5 g18981(new_n21329, new_n21327, new_n21330);
xnor_4 g18982(new_n21328, new_n21327, new_n21331);
not_8  g18983(new_n21293, new_n21332);
xnor_4 g18984(new_n21302_1, new_n21332, new_n21333);
xnor_4 g18985(new_n21319, new_n21312, new_n21334);
not_8  g18986(new_n21334, new_n21335);
nand_5 g18987(new_n21335, new_n21333, new_n21336);
xnor_4 g18988(new_n21334, new_n21333, new_n21337);
not_8  g18989(new_n21297, new_n21338);
xnor_4 g18990(new_n21300, new_n21338, new_n21339);
xnor_4 g18991(new_n21317_1, new_n21316, new_n21340);
not_8  g18992(new_n21340, new_n21341);
nand_5 g18993(new_n21341, new_n21339, new_n21342);
xnor_4 g18994(new_n21340, new_n21339, new_n21343);
not_8  g18995(new_n14554, new_n21344);
nand_5 g18996(new_n14575_1, new_n21344, new_n21345);
nand_5 g18997(new_n14614, new_n14576_1, new_n21346);
nand_5 g18998(new_n21346, new_n21345, new_n21347);
nand_5 g18999(new_n21347, new_n21343, new_n21348);
nand_5 g19000(new_n21348, new_n21342, new_n21349_1);
nand_5 g19001(new_n21349_1, new_n21337, new_n21350);
nand_5 g19002(new_n21350, new_n21336, new_n21351);
nand_5 g19003(new_n21351, new_n21331, new_n21352);
nand_5 g19004(new_n21352, new_n21330, new_n21353);
xnor_4 g19005(new_n21353, new_n21325, n6576);
xnor_4 g19006(new_n21040, new_n18138, new_n21355);
xnor_4 g19007(new_n21355, new_n21044, n6587);
xnor_4 g19008(new_n19884, new_n19827, n6612);
not_8  g19009(new_n18461, new_n21358);
nand_5 g19010(new_n21358, new_n11458, new_n21359);
xnor_4 g19011(new_n18461, new_n11458, new_n21360);
not_8  g19012(new_n18464, new_n21361);
nand_5 g19013(new_n21361, new_n11452, new_n21362);
xnor_4 g19014(new_n18464, new_n11452, new_n21363);
not_8  g19015(new_n18467_1, new_n21364);
nand_5 g19016(new_n21364, new_n11445, new_n21365_1);
xnor_4 g19017(new_n18467_1, new_n11445, new_n21366);
not_8  g19018(new_n18470, new_n21367_1);
nand_5 g19019(new_n21367_1, new_n11437, new_n21368);
xnor_4 g19020(new_n18470, new_n11437, new_n21369);
not_8  g19021(new_n18473, new_n21370);
nand_5 g19022(new_n21370, new_n17343, new_n21371);
xnor_4 g19023(new_n21370, new_n11429, new_n21372);
nor_5  g19024(new_n18475, new_n11421, new_n21373);
not_8  g19025(new_n21373, new_n21374);
xnor_4 g19026(new_n18475, new_n11421, new_n21375);
not_8  g19027(new_n21375, new_n21376);
nor_5  g19028(new_n15988, new_n11414, new_n21377);
not_8  g19029(new_n21377, new_n21378);
xnor_4 g19030(new_n18479, new_n11414, new_n21379);
nor_5  g19031(new_n15991, new_n11406, new_n21380);
nor_5  g19032(new_n11489, n18, new_n21381);
nand_5 g19033(new_n21381, new_n9693, new_n21382);
not_8  g19034(new_n21382, new_n21383);
nor_5  g19035(new_n21381, new_n15995, new_n21384);
nor_5  g19036(new_n21384, new_n21383, new_n21385);
nand_5 g19037(new_n21385, new_n11397, new_n21386);
nand_5 g19038(new_n21386, new_n21382, new_n21387);
xnor_4 g19039(new_n15991, new_n11405, new_n21388);
not_8  g19040(new_n21388, new_n21389);
nor_5  g19041(new_n21389, new_n21387, new_n21390);
nor_5  g19042(new_n21390, new_n21380, new_n21391);
nand_5 g19043(new_n21391, new_n21379, new_n21392);
nand_5 g19044(new_n21392, new_n21378, new_n21393);
nand_5 g19045(new_n21393, new_n21376, new_n21394);
nand_5 g19046(new_n21394, new_n21374, new_n21395);
nand_5 g19047(new_n21395, new_n21372, new_n21396_1);
nand_5 g19048(new_n21396_1, new_n21371, new_n21397);
nand_5 g19049(new_n21397, new_n21369, new_n21398_1);
nand_5 g19050(new_n21398_1, new_n21368, new_n21399_1);
nand_5 g19051(new_n21399_1, new_n21366, new_n21400);
nand_5 g19052(new_n21400, new_n21365_1, new_n21401);
nand_5 g19053(new_n21401, new_n21363, new_n21402);
nand_5 g19054(new_n21402, new_n21362, new_n21403);
nand_5 g19055(new_n21403, new_n21360, new_n21404_1);
nand_5 g19056(new_n21404_1, new_n21359, new_n21405);
nor_5  g19057(new_n18460, n23166, new_n21406);
nand_5 g19058(new_n18656, new_n21406, new_n21407);
nor_5  g19059(new_n21407, new_n21405, new_n21408);
nor_5  g19060(new_n18656, new_n21406, new_n21409);
nand_5 g19061(new_n21409, new_n21405, new_n21410);
not_8  g19062(new_n21410, new_n21411);
nor_5  g19063(new_n21411, new_n21408, new_n21412);
xnor_4 g19064(new_n19160, new_n21406, new_n21413);
not_8  g19065(new_n21413, new_n21414);
xnor_4 g19066(new_n21414, new_n21405, new_n21415);
not_8  g19067(new_n21415, new_n21416);
nand_5 g19068(new_n21416, new_n20597, new_n21417);
xnor_4 g19069(new_n21415, new_n20597, new_n21418);
xnor_4 g19070(new_n21403, new_n21360, new_n21419);
not_8  g19071(new_n21419, new_n21420);
nand_5 g19072(new_n21420, new_n20604_1, new_n21421);
xnor_4 g19073(new_n21419, new_n20604_1, new_n21422);
xnor_4 g19074(new_n21401, new_n21363, new_n21423);
not_8  g19075(new_n21423, new_n21424);
nand_5 g19076(new_n21424, new_n20611, new_n21425);
xnor_4 g19077(new_n21423, new_n20611, new_n21426);
xnor_4 g19078(new_n21399_1, new_n21366, new_n21427);
not_8  g19079(new_n21427, new_n21428);
nand_5 g19080(new_n21428, new_n20617, new_n21429);
xnor_4 g19081(new_n21427, new_n20617, new_n21430);
xnor_4 g19082(new_n21397, new_n21369, new_n21431);
not_8  g19083(new_n21431, new_n21432);
nand_5 g19084(new_n21432, new_n9976, new_n21433);
xnor_4 g19085(new_n21431, new_n9976, new_n21434);
not_8  g19086(new_n21372, new_n21435);
xnor_4 g19087(new_n21395, new_n21435, new_n21436);
nand_5 g19088(new_n21436, new_n9982, new_n21437);
xnor_4 g19089(new_n21436, new_n9980, new_n21438);
xnor_4 g19090(new_n21393, new_n21376, new_n21439);
not_8  g19091(new_n21439, new_n21440);
nand_5 g19092(new_n21440, new_n9987, new_n21441);
xnor_4 g19093(new_n21439, new_n9987, new_n21442);
not_8  g19094(new_n21379, new_n21443);
xnor_4 g19095(new_n21391, new_n21443, new_n21444);
nand_5 g19096(new_n21444, new_n9993, new_n21445);
xnor_4 g19097(new_n21444, new_n9991, new_n21446_1);
xnor_4 g19098(new_n21388, new_n21387, new_n21447);
nor_5  g19099(new_n21447, new_n9999, new_n21448);
not_8  g19100(new_n21448, new_n21449);
xnor_4 g19101(new_n21447, new_n9997, new_n21450);
xnor_4 g19102(new_n21385, new_n11396, new_n21451);
not_8  g19103(new_n21451, new_n21452);
nor_5  g19104(new_n21452, new_n10010_1, new_n21453);
not_8  g19105(new_n21453, new_n21454);
xnor_4 g19106(new_n11393, n18, new_n21455);
nor_5  g19107(new_n21455, new_n10006, new_n21456);
not_8  g19108(new_n21456, new_n21457);
xnor_4 g19109(new_n21451, new_n10010_1, new_n21458);
nand_5 g19110(new_n21458, new_n21457, new_n21459);
nand_5 g19111(new_n21459, new_n21454, new_n21460);
nand_5 g19112(new_n21460, new_n21450, new_n21461);
nand_5 g19113(new_n21461, new_n21449, new_n21462);
nand_5 g19114(new_n21462, new_n21446_1, new_n21463);
nand_5 g19115(new_n21463, new_n21445, new_n21464);
nand_5 g19116(new_n21464, new_n21442, new_n21465);
nand_5 g19117(new_n21465, new_n21441, new_n21466);
nand_5 g19118(new_n21466, new_n21438, new_n21467);
nand_5 g19119(new_n21467, new_n21437, new_n21468);
nand_5 g19120(new_n21468, new_n21434, new_n21469);
nand_5 g19121(new_n21469, new_n21433, new_n21470);
nand_5 g19122(new_n21470, new_n21430, new_n21471_1);
nand_5 g19123(new_n21471_1, new_n21429, new_n21472_1);
nand_5 g19124(new_n21472_1, new_n21426, new_n21473);
nand_5 g19125(new_n21473, new_n21425, new_n21474);
nand_5 g19126(new_n21474, new_n21422, new_n21475);
nand_5 g19127(new_n21475, new_n21421, new_n21476);
nand_5 g19128(new_n21476, new_n21418, new_n21477);
nand_5 g19129(new_n21477, new_n21417, new_n21478);
xnor_4 g19130(new_n21478, new_n20592, new_n21479);
xnor_4 g19131(new_n21479, new_n21412, n6628);
xnor_4 g19132(new_n2885, new_n2865, n6630);
xnor_4 g19133(n25331, new_n16884, new_n21482);
not_8  g19134(new_n21482, new_n21483);
or_5   g19135(n21997, n18483, new_n21484);
nand_5 g19136(new_n20701, new_n20690, new_n21485);
nand_5 g19137(new_n21485, new_n21484, new_n21486);
xnor_4 g19138(new_n21486, new_n21483, new_n21487);
xnor_4 g19139(new_n21487, new_n7952, new_n21488);
not_8  g19140(new_n21488, new_n21489_1);
not_8  g19141(new_n7943_1, new_n21490);
nor_5  g19142(new_n20702, new_n21490, new_n21491);
not_8  g19143(new_n21491, new_n21492);
not_8  g19144(new_n20714, new_n21493);
nand_5 g19145(new_n21493, new_n20703, new_n21494);
nand_5 g19146(new_n21494, new_n21492, new_n21495);
xnor_4 g19147(new_n21495, new_n21489_1, new_n21496);
xnor_4 g19148(n14130, n468, new_n21497);
not_8  g19149(new_n21497, new_n21498);
nor_5  g19150(n16482, new_n7408_1, new_n21499);
xnor_4 g19151(n16482, n5400, new_n21500);
not_8  g19152(new_n21500, new_n21501);
nor_5  g19153(new_n8795, n9942, new_n21502);
nor_5  g19154(n25643, new_n7415, new_n21503);
xnor_4 g19155(n25643, n329, new_n21504);
not_8  g19156(new_n21504, new_n21505);
nor_5  g19157(new_n8803_1, n9557, new_n21506);
xnor_4 g19158(n24170, n9557, new_n21507);
not_8  g19159(new_n21507, new_n21508);
or_5   g19160(new_n3576, n2409, new_n21509);
xnor_4 g19161(n3136, n2409, new_n21510);
nand_5 g19162(new_n8807, n6385, new_n21511);
nand_5 g19163(new_n20256, new_n20253, new_n21512);
nand_5 g19164(new_n21512, new_n21511, new_n21513);
nand_5 g19165(new_n21513, new_n21510, new_n21514);
nand_5 g19166(new_n21514, new_n21509, new_n21515);
nor_5  g19167(new_n21515, new_n21508, new_n21516);
nor_5  g19168(new_n21516, new_n21506, new_n21517);
nor_5  g19169(new_n21517, new_n21505, new_n21518);
nor_5  g19170(new_n21518, new_n21503, new_n21519);
xnor_4 g19171(n23923, n9942, new_n21520);
not_8  g19172(new_n21520, new_n21521);
nor_5  g19173(new_n21521, new_n21519, new_n21522);
nor_5  g19174(new_n21522, new_n21502, new_n21523);
nor_5  g19175(new_n21523, new_n21501, new_n21524);
nor_5  g19176(new_n21524, new_n21499, new_n21525_1);
xnor_4 g19177(new_n21525_1, new_n21498, new_n21526);
xnor_4 g19178(new_n21526, new_n21496, new_n21527);
xnor_4 g19179(new_n21523, new_n21500, new_n21528);
nor_5  g19180(new_n21528, new_n20715, new_n21529);
xnor_4 g19181(new_n21528, new_n20715, new_n21530);
xnor_4 g19182(new_n21521, new_n21519, new_n21531);
nor_5  g19183(new_n21531, new_n20719, new_n21532);
not_8  g19184(new_n21532, new_n21533);
xnor_4 g19185(new_n21517, new_n21504, new_n21534);
nor_5  g19186(new_n21534, new_n20303, new_n21535);
xnor_4 g19187(new_n21534, new_n20302, new_n21536);
not_8  g19188(new_n21536, new_n21537);
xnor_4 g19189(new_n21515, new_n21507, new_n21538_1);
nor_5  g19190(new_n21538_1, new_n20354, new_n21539);
xnor_4 g19191(new_n21538_1, new_n20326, new_n21540);
not_8  g19192(new_n21540, new_n21541);
xnor_4 g19193(new_n21513, new_n21510, new_n21542);
nor_5  g19194(new_n21542, new_n20329, new_n21543);
xnor_4 g19195(new_n21542, new_n20329, new_n21544);
nor_5  g19196(new_n20257, new_n20252, new_n21545);
nor_5  g19197(new_n20264, new_n20260, new_n21546);
nor_5  g19198(new_n21546, new_n21545, new_n21547);
nor_5  g19199(new_n21547, new_n21544, new_n21548);
nor_5  g19200(new_n21548, new_n21543, new_n21549_1);
nor_5  g19201(new_n21549_1, new_n21541, new_n21550);
nor_5  g19202(new_n21550, new_n21539, new_n21551);
nor_5  g19203(new_n21551, new_n21537, new_n21552);
nor_5  g19204(new_n21552, new_n21535, new_n21553);
xnor_4 g19205(new_n21531, new_n20718, new_n21554);
nand_5 g19206(new_n21554, new_n21553, new_n21555);
nand_5 g19207(new_n21555, new_n21533, new_n21556);
nor_5  g19208(new_n21556, new_n21530, new_n21557);
nor_5  g19209(new_n21557, new_n21529, new_n21558);
nand_5 g19210(new_n21558, new_n21527, new_n21559);
not_8  g19211(new_n21559, new_n21560);
nor_5  g19212(new_n21558, new_n21527, new_n21561);
nor_5  g19213(new_n21561, new_n21560, n6634);
xnor_4 g19214(new_n6932, new_n6915, n6652);
xnor_4 g19215(new_n13332, new_n13316, n6655);
xnor_4 g19216(new_n12815, new_n12790, n6669);
xnor_4 g19217(new_n10016, new_n9995, n6671);
xnor_4 g19218(new_n14410, new_n14388, n6673);
nand_5 g19219(new_n21246, new_n21237, new_n21568);
nor_5  g19220(new_n12182, new_n12696, new_n21569);
not_8  g19221(new_n21244, new_n21570);
nand_5 g19222(new_n21570, new_n21569, new_n21571);
nand_5 g19223(new_n21571, new_n21568, n6674);
xnor_4 g19224(new_n17610, new_n17600, n6684);
xnor_4 g19225(new_n13062, new_n13013, n6706);
xnor_4 g19226(n12702, new_n6526, new_n21575);
nor_5  g19227(n26797, n15182, new_n21576);
xnor_4 g19228(n26797, new_n6542_1, new_n21577);
not_8  g19229(new_n21577, new_n21578);
nor_5  g19230(n27037, n23913, new_n21579);
xnor_4 g19231(n27037, new_n5851, new_n21580);
not_8  g19232(new_n21580, new_n21581);
nor_5  g19233(n22554, n8964, new_n21582);
xnor_4 g19234(n22554, new_n6551, new_n21583);
not_8  g19235(new_n21583, new_n21584);
nor_5  g19236(n20429, n20151, new_n21585);
xnor_4 g19237(n20429, new_n6557, new_n21586);
not_8  g19238(new_n21586, new_n21587);
nor_5  g19239(n7693, n3909, new_n21588);
xnor_4 g19240(n7693, new_n5837, new_n21589);
not_8  g19241(new_n21589, new_n21590);
nor_5  g19242(n23974, n10405, new_n21591);
xnor_4 g19243(n23974, new_n4189, new_n21592);
not_8  g19244(new_n21592, new_n21593);
nand_5 g19245(n11302, n2146, new_n21594);
nor_5  g19246(n11302, n2146, new_n21595);
not_8  g19247(new_n21595, new_n21596);
nor_5  g19248(n22173, n17090, new_n21597);
not_8  g19249(new_n16644, new_n21598);
nor_5  g19250(new_n21598, new_n16643, new_n21599_1);
nor_5  g19251(new_n21599_1, new_n21597, new_n21600);
nand_5 g19252(new_n21600, new_n21596, new_n21601);
nand_5 g19253(new_n21601, new_n21594, new_n21602);
nor_5  g19254(new_n21602, new_n21593, new_n21603);
nor_5  g19255(new_n21603, new_n21591, new_n21604);
nor_5  g19256(new_n21604, new_n21590, new_n21605);
nor_5  g19257(new_n21605, new_n21588, new_n21606);
nor_5  g19258(new_n21606, new_n21587, new_n21607);
nor_5  g19259(new_n21607, new_n21585, new_n21608);
nor_5  g19260(new_n21608, new_n21584, new_n21609);
nor_5  g19261(new_n21609, new_n21582, new_n21610);
nor_5  g19262(new_n21610, new_n21581, new_n21611);
nor_5  g19263(new_n21611, new_n21579, new_n21612);
nor_5  g19264(new_n21612, new_n21578, new_n21613);
nor_5  g19265(new_n21613, new_n21576, new_n21614);
xnor_4 g19266(new_n21614, new_n21575, new_n21615_1);
nand_5 g19267(new_n21615_1, n1831, new_n21616);
xnor_4 g19268(new_n21615_1, new_n6478, new_n21617);
xnor_4 g19269(new_n21612, new_n21577, new_n21618);
nand_5 g19270(new_n21618, n13137, new_n21619);
xnor_4 g19271(new_n21618, new_n14804, new_n21620);
xnor_4 g19272(new_n21610, new_n21580, new_n21621);
nand_5 g19273(new_n21621, n18452, new_n21622);
xnor_4 g19274(new_n21621, new_n14808, new_n21623);
xnor_4 g19275(new_n21608, new_n21583, new_n21624);
nand_5 g19276(new_n21624, n21317, new_n21625);
xnor_4 g19277(new_n21624, new_n14812, new_n21626);
xnor_4 g19278(new_n21606, new_n21586, new_n21627);
nand_5 g19279(new_n21627, n12398, new_n21628_1);
xnor_4 g19280(new_n21627, new_n4169, new_n21629);
xnor_4 g19281(new_n21604, new_n21589, new_n21630);
nand_5 g19282(new_n21630, n19789, new_n21631);
xnor_4 g19283(new_n21630, new_n4170, new_n21632);
xnor_4 g19284(new_n21602, new_n21592, new_n21633);
nand_5 g19285(new_n21633, n20169, new_n21634);
xnor_4 g19286(new_n21633, new_n4227, new_n21635);
xnor_4 g19287(n11302, new_n5838, new_n21636);
xnor_4 g19288(new_n21636, new_n21600, new_n21637_1);
nand_5 g19289(new_n21637_1, n8285, new_n21638);
xnor_4 g19290(new_n21637_1, new_n4171, new_n21639);
not_8  g19291(new_n16640_1, new_n21640);
not_8  g19292(new_n16645, new_n21641);
nor_5  g19293(new_n21641, new_n16641, new_n21642);
nor_5  g19294(new_n21642, new_n21640, new_n21643);
not_8  g19295(new_n21643, new_n21644);
nand_5 g19296(new_n21644, new_n21639, new_n21645_1);
nand_5 g19297(new_n21645_1, new_n21638, new_n21646);
nand_5 g19298(new_n21646, new_n21635, new_n21647);
nand_5 g19299(new_n21647, new_n21634, new_n21648);
nand_5 g19300(new_n21648, new_n21632, new_n21649_1);
nand_5 g19301(new_n21649_1, new_n21631, new_n21650);
nand_5 g19302(new_n21650, new_n21629, new_n21651);
nand_5 g19303(new_n21651, new_n21628_1, new_n21652);
nand_5 g19304(new_n21652, new_n21626, new_n21653);
nand_5 g19305(new_n21653, new_n21625, new_n21654_1);
nand_5 g19306(new_n21654_1, new_n21623, new_n21655);
nand_5 g19307(new_n21655, new_n21622, new_n21656);
nand_5 g19308(new_n21656, new_n21620, new_n21657);
nand_5 g19309(new_n21657, new_n21619, new_n21658);
nand_5 g19310(new_n21658, new_n21617, new_n21659);
nand_5 g19311(new_n21659, new_n21616, new_n21660);
or_5   g19312(n12702, n8614, new_n21661);
not_8  g19313(new_n21614, new_n21662);
nand_5 g19314(new_n21662, new_n21575, new_n21663);
nand_5 g19315(new_n21663, new_n21661, new_n21664);
xnor_4 g19316(new_n21664, new_n21660, new_n21665_1);
nor_5  g19317(new_n21285, new_n4664, new_n21666);
nor_5  g19318(new_n21306, new_n21287_1, new_n21667);
nor_5  g19319(new_n21667, new_n21666, new_n21668);
nor_5  g19320(new_n21283, n1536, new_n21669);
xnor_4 g19321(new_n21669, new_n4645, new_n21670);
xnor_4 g19322(new_n21670, new_n21668, new_n21671);
xnor_4 g19323(new_n21671, new_n21665_1, new_n21672);
xnor_4 g19324(new_n21658, new_n21617, new_n21673);
not_8  g19325(new_n21673, new_n21674_1);
nand_5 g19326(new_n21674_1, new_n21307, new_n21675);
xnor_4 g19327(new_n21673, new_n21307, new_n21676);
xnor_4 g19328(new_n21656, new_n21620, new_n21677);
not_8  g19329(new_n21677, new_n21678);
nand_5 g19330(new_n21678, new_n21327, new_n21679);
xnor_4 g19331(new_n21677, new_n21327, new_n21680_1);
xnor_4 g19332(new_n21654_1, new_n21623, new_n21681);
not_8  g19333(new_n21681, new_n21682);
nand_5 g19334(new_n21682, new_n21333, new_n21683);
xnor_4 g19335(new_n21681, new_n21333, new_n21684);
xnor_4 g19336(new_n21652, new_n21626, new_n21685_1);
not_8  g19337(new_n21685_1, new_n21686);
nand_5 g19338(new_n21686, new_n21339, new_n21687_1);
xnor_4 g19339(new_n21685_1, new_n21339, new_n21688);
xnor_4 g19340(new_n21650, new_n21629, new_n21689);
not_8  g19341(new_n21689, new_n21690);
nand_5 g19342(new_n21690, new_n21344, new_n21691);
xnor_4 g19343(new_n21690, new_n14554, new_n21692);
xnor_4 g19344(new_n21648, new_n21632, new_n21693);
not_8  g19345(new_n21693, new_n21694);
nand_5 g19346(new_n21694, new_n14580, new_n21695);
xnor_4 g19347(new_n21693, new_n14580, new_n21696);
not_8  g19348(new_n21635, new_n21697);
xnor_4 g19349(new_n21646, new_n21697, new_n21698);
nand_5 g19350(new_n21698, new_n14584, new_n21699);
xnor_4 g19351(new_n21698, new_n14583, new_n21700);
xnor_4 g19352(new_n21643, new_n21639, new_n21701);
nor_5  g19353(new_n21701, new_n14589, new_n21702);
not_8  g19354(new_n16646, new_n21703);
nor_5  g19355(new_n21703, new_n14594, new_n21704);
not_8  g19356(new_n21704, new_n21705);
nand_5 g19357(new_n16647, new_n16635, new_n21706);
nand_5 g19358(new_n21706, new_n21705, new_n21707);
xnor_4 g19359(new_n21701, new_n14589, new_n21708);
nor_5  g19360(new_n21708, new_n21707, new_n21709);
nor_5  g19361(new_n21709, new_n21702, new_n21710);
nand_5 g19362(new_n21710, new_n21700, new_n21711);
nand_5 g19363(new_n21711, new_n21699, new_n21712);
nand_5 g19364(new_n21712, new_n21696, new_n21713);
nand_5 g19365(new_n21713, new_n21695, new_n21714);
nand_5 g19366(new_n21714, new_n21692, new_n21715);
nand_5 g19367(new_n21715, new_n21691, new_n21716);
nand_5 g19368(new_n21716, new_n21688, new_n21717_1);
nand_5 g19369(new_n21717_1, new_n21687_1, new_n21718);
nand_5 g19370(new_n21718, new_n21684, new_n21719_1);
nand_5 g19371(new_n21719_1, new_n21683, new_n21720);
nand_5 g19372(new_n21720, new_n21680_1, new_n21721);
nand_5 g19373(new_n21721, new_n21679, new_n21722);
nand_5 g19374(new_n21722, new_n21676, new_n21723);
nand_5 g19375(new_n21723, new_n21675, new_n21724);
xnor_4 g19376(new_n21724, new_n21672, n6707);
xnor_4 g19377(new_n13921, new_n13651, n6736);
xnor_4 g19378(n23895, n5101, new_n21727);
nand_5 g19379(new_n5740, n16507, new_n21728);
xnor_4 g19380(n17351, n16507, new_n21729);
nand_5 g19381(n22470, new_n5743, new_n21730);
xnor_4 g19382(n22470, n11736, new_n21731);
nand_5 g19383(new_n5746, n19116, new_n21732);
or_5   g19384(n17959, new_n3397, new_n21733);
nand_5 g19385(new_n19049, new_n19028, new_n21734);
nand_5 g19386(new_n21734, new_n21733, new_n21735_1);
xnor_4 g19387(n23200, n19116, new_n21736);
nand_5 g19388(new_n21736, new_n21735_1, new_n21737);
nand_5 g19389(new_n21737, new_n21732, new_n21738);
nand_5 g19390(new_n21738, new_n21731, new_n21739);
nand_5 g19391(new_n21739, new_n21730, new_n21740);
nand_5 g19392(new_n21740, new_n21729, new_n21741);
nand_5 g19393(new_n21741, new_n21728, new_n21742);
xnor_4 g19394(new_n21742, new_n21727, new_n21743);
nor_5  g19395(new_n19054, n22660, new_n21744);
nand_5 g19396(new_n21744, new_n5796, new_n21745);
nor_5  g19397(new_n21745, n9655, new_n21746);
nand_5 g19398(new_n21746, new_n5790, new_n21747);
xnor_4 g19399(new_n21747, new_n5787, new_n21748);
xnor_4 g19400(new_n21748, n12650, new_n21749_1);
xnor_4 g19401(new_n21746, n25345, new_n21750_1);
not_8  g19402(new_n21750_1, new_n21751);
nand_5 g19403(new_n21751, n10201, new_n21752);
xnor_4 g19404(new_n21750_1, n10201, new_n21753_1);
xnor_4 g19405(new_n21745, new_n5793, new_n21754);
not_8  g19406(new_n21754, new_n21755);
nand_5 g19407(new_n21755, n10593, new_n21756);
xnor_4 g19408(new_n21754, n10593, new_n21757);
xnor_4 g19409(new_n21744, n13490, new_n21758);
not_8  g19410(new_n21758, new_n21759);
nand_5 g19411(new_n21759, n18290, new_n21760);
xnor_4 g19412(new_n21758, n18290, new_n21761);
not_8  g19413(new_n19055, new_n21762);
nand_5 g19414(new_n21762, n11580, new_n21763);
nand_5 g19415(new_n19080, new_n19056, new_n21764);
nand_5 g19416(new_n21764, new_n21763, new_n21765_1);
nand_5 g19417(new_n21765_1, new_n21761, new_n21766);
nand_5 g19418(new_n21766, new_n21760, new_n21767);
nand_5 g19419(new_n21767, new_n21757, new_n21768);
nand_5 g19420(new_n21768, new_n21756, new_n21769);
nand_5 g19421(new_n21769, new_n21753_1, new_n21770);
nand_5 g19422(new_n21770, new_n21752, new_n21771);
xnor_4 g19423(new_n21771, new_n21749_1, new_n21772);
xnor_4 g19424(new_n21772, new_n16882, new_n21773);
xnor_4 g19425(new_n21769, new_n21753_1, new_n21774);
nand_5 g19426(new_n21774, new_n16886, new_n21775);
xnor_4 g19427(new_n21767, new_n21757, new_n21776);
nor_5  g19428(new_n21776, new_n16891, new_n21777);
xnor_4 g19429(new_n21776, new_n16891, new_n21778);
xnor_4 g19430(new_n21765_1, new_n21761, new_n21779_1);
nand_5 g19431(new_n21779_1, new_n16896, new_n21780);
xnor_4 g19432(new_n21779_1, new_n16895, new_n21781);
nand_5 g19433(new_n19081_1, new_n16900, new_n21782);
nand_5 g19434(new_n19106, new_n19082, new_n21783);
nand_5 g19435(new_n21783, new_n21782, new_n21784_1);
nand_5 g19436(new_n21784_1, new_n21781, new_n21785);
nand_5 g19437(new_n21785, new_n21780, new_n21786);
nor_5  g19438(new_n21786, new_n21778, new_n21787);
nor_5  g19439(new_n21787, new_n21777, new_n21788);
xnor_4 g19440(new_n21774, new_n16885_1, new_n21789);
nand_5 g19441(new_n21789, new_n21788, new_n21790);
nand_5 g19442(new_n21790, new_n21775, new_n21791);
xnor_4 g19443(new_n21791, new_n21773, new_n21792);
xnor_4 g19444(new_n21792, new_n21743, new_n21793);
not_8  g19445(new_n21729, new_n21794);
xnor_4 g19446(new_n21740, new_n21794, new_n21795);
not_8  g19447(new_n21795, new_n21796);
xnor_4 g19448(new_n21789, new_n21788, new_n21797);
nand_5 g19449(new_n21797, new_n21796, new_n21798);
not_8  g19450(new_n21798, new_n21799);
xnor_4 g19451(new_n21797, new_n21795, new_n21800_1);
not_8  g19452(new_n21800_1, new_n21801);
xnor_4 g19453(new_n21738, new_n21731, new_n21802);
xnor_4 g19454(new_n21786, new_n21778, new_n21803);
not_8  g19455(new_n21803, new_n21804);
nand_5 g19456(new_n21804, new_n21802, new_n21805);
not_8  g19457(new_n21805, new_n21806);
xnor_4 g19458(new_n21803, new_n21802, new_n21807);
not_8  g19459(new_n21807, new_n21808);
xnor_4 g19460(new_n21736, new_n21735_1, new_n21809);
xnor_4 g19461(new_n21784_1, new_n21781, new_n21810);
nor_5  g19462(new_n21810, new_n21809, new_n21811);
xnor_4 g19463(new_n21810, new_n21809, new_n21812);
nor_5  g19464(new_n19107_1, new_n19050, new_n21813);
nor_5  g19465(new_n19148, new_n19108, new_n21814);
nor_5  g19466(new_n21814, new_n21813, new_n21815);
nor_5  g19467(new_n21815, new_n21812, new_n21816);
nor_5  g19468(new_n21816, new_n21811, new_n21817);
not_8  g19469(new_n21817, new_n21818);
nor_5  g19470(new_n21818, new_n21808, new_n21819);
nor_5  g19471(new_n21819, new_n21806, new_n21820_1);
nor_5  g19472(new_n21820_1, new_n21801, new_n21821);
nor_5  g19473(new_n21821, new_n21799, new_n21822);
xnor_4 g19474(new_n21822, new_n21793, n6791);
xnor_4 g19475(new_n3861, new_n3850_1, n6802);
xnor_4 g19476(new_n17273, new_n17244, n6826);
xnor_4 g19477(new_n10681, new_n10650_1, n6835);
not_8  g19478(new_n19372, new_n21827);
nand_5 g19479(new_n19377, n11220, new_n21828);
xnor_4 g19480(new_n19377, new_n10741, new_n21829);
nand_5 g19481(new_n2985_1, n22379, new_n21830);
xnor_4 g19482(new_n2985_1, new_n19358, new_n21831);
not_8  g19483(new_n3034, new_n21832_1);
nand_5 g19484(new_n21832_1, n1662, new_n21833);
xnor_4 g19485(new_n3034, n1662, new_n21834);
nand_5 g19486(new_n3041, n12875, new_n21835);
xnor_4 g19487(new_n3040, n12875, new_n21836);
nor_5  g19488(new_n3047, new_n2906, new_n21837);
nor_5  g19489(new_n3055, n5213, new_n21838);
xnor_4 g19490(new_n3054, n5213, new_n21839_1);
not_8  g19491(new_n21839_1, new_n21840);
nor_5  g19492(new_n3062, n4665, new_n21841);
xnor_4 g19493(new_n3061, n4665, new_n21842);
nor_5  g19494(new_n3067_1, new_n2917, new_n21843);
xnor_4 g19495(new_n3067_1, new_n2917, new_n21844);
nor_5  g19496(new_n3076_1, new_n9889, new_n21845);
nor_5  g19497(new_n21845, n4326, new_n21846);
xnor_4 g19498(new_n21845, n4326, new_n21847);
nor_5  g19499(new_n21847, new_n3073, new_n21848);
nor_5  g19500(new_n21848, new_n21846, new_n21849);
not_8  g19501(new_n21849, new_n21850);
nor_5  g19502(new_n21850, new_n21844, new_n21851);
nor_5  g19503(new_n21851, new_n21843, new_n21852);
nand_5 g19504(new_n21852, new_n21842, new_n21853);
not_8  g19505(new_n21853, new_n21854);
nor_5  g19506(new_n21854, new_n21841, new_n21855);
nor_5  g19507(new_n21855, new_n21840, new_n21856);
nor_5  g19508(new_n21856, new_n21838, new_n21857);
xnor_4 g19509(new_n3047, n2035, new_n21858);
nand_5 g19510(new_n21858, new_n21857, new_n21859);
not_8  g19511(new_n21859, new_n21860);
nor_5  g19512(new_n21860, new_n21837, new_n21861);
not_8  g19513(new_n21861, new_n21862);
nand_5 g19514(new_n21862, new_n21836, new_n21863);
nand_5 g19515(new_n21863, new_n21835, new_n21864);
nand_5 g19516(new_n21864, new_n21834, new_n21865);
nand_5 g19517(new_n21865, new_n21833, new_n21866);
nand_5 g19518(new_n21866, new_n21831, new_n21867);
nand_5 g19519(new_n21867, new_n21830, new_n21868);
nand_5 g19520(new_n21868, new_n21829, new_n21869);
nand_5 g19521(new_n21869, new_n21828, new_n21870);
nand_5 g19522(new_n21870, new_n21827, new_n21871);
xnor_4 g19523(new_n21871, new_n19010, new_n21872);
xnor_4 g19524(new_n21870, new_n21827, new_n21873);
nand_5 g19525(new_n21873, new_n19015, new_n21874_1);
xnor_4 g19526(new_n21873, new_n19013, new_n21875);
xnor_4 g19527(new_n21868, new_n21829, new_n21876);
nand_5 g19528(new_n21876, new_n13679, new_n21877);
xnor_4 g19529(new_n21876, new_n6410, new_n21878);
not_8  g19530(new_n6412, new_n21879);
xnor_4 g19531(new_n21866, new_n21831, new_n21880);
nand_5 g19532(new_n21880, new_n21879, new_n21881);
xnor_4 g19533(new_n21880, new_n6412, new_n21882);
xnor_4 g19534(new_n21864, new_n21834, new_n21883);
nand_5 g19535(new_n21883, new_n13715, new_n21884);
xnor_4 g19536(new_n21883, new_n6420, new_n21885);
not_8  g19537(new_n6425, new_n21886);
xnor_4 g19538(new_n21862, new_n21836, new_n21887);
nand_5 g19539(new_n21887, new_n21886, new_n21888);
xnor_4 g19540(new_n21887, new_n6425, new_n21889);
xnor_4 g19541(new_n21858, new_n21857, new_n21890);
nand_5 g19542(new_n21890, new_n6431_1, new_n21891);
xnor_4 g19543(new_n21890, new_n6432, new_n21892);
xnor_4 g19544(new_n21855, new_n21839_1, new_n21893);
not_8  g19545(new_n21893, new_n21894);
nor_5  g19546(new_n21894, new_n6437_1, new_n21895);
not_8  g19547(new_n21895, new_n21896);
xnor_4 g19548(new_n21893, new_n6437_1, new_n21897);
not_8  g19549(new_n21897, new_n21898_1);
xnor_4 g19550(new_n21852, new_n21842, new_n21899);
nor_5  g19551(new_n21899, new_n6444, new_n21900);
xnor_4 g19552(new_n21899, new_n6441, new_n21901);
not_8  g19553(new_n21901, new_n21902);
xnor_4 g19554(new_n21849, new_n21844, new_n21903);
nor_5  g19555(new_n21903, new_n6447, new_n21904);
xnor_4 g19556(new_n21903, new_n6448, new_n21905_1);
not_8  g19557(new_n21905_1, new_n21906);
xnor_4 g19558(new_n21847, new_n3082, new_n21907);
and_5  g19559(new_n21907, new_n13729, new_n21908);
nor_5  g19560(new_n6111, new_n6110, new_n21909);
not_8  g19561(new_n21909, new_n21910);
xnor_4 g19562(new_n21907, new_n6452, new_n21911);
not_8  g19563(new_n21911, new_n21912);
nor_5  g19564(new_n21912, new_n21910, new_n21913);
nor_5  g19565(new_n21913, new_n21908, new_n21914);
nor_5  g19566(new_n21914, new_n21906, new_n21915_1);
nor_5  g19567(new_n21915_1, new_n21904, new_n21916);
nor_5  g19568(new_n21916, new_n21902, new_n21917);
nor_5  g19569(new_n21917, new_n21900, new_n21918);
nor_5  g19570(new_n21918, new_n21898_1, new_n21919);
not_8  g19571(new_n21919, new_n21920);
nand_5 g19572(new_n21920, new_n21896, new_n21921);
nand_5 g19573(new_n21921, new_n21892, new_n21922);
nand_5 g19574(new_n21922, new_n21891, new_n21923);
nand_5 g19575(new_n21923, new_n21889, new_n21924);
nand_5 g19576(new_n21924, new_n21888, new_n21925);
nand_5 g19577(new_n21925, new_n21885, new_n21926);
nand_5 g19578(new_n21926, new_n21884, new_n21927);
nand_5 g19579(new_n21927, new_n21882, new_n21928);
nand_5 g19580(new_n21928, new_n21881, new_n21929);
nand_5 g19581(new_n21929, new_n21878, new_n21930);
nand_5 g19582(new_n21930, new_n21877, new_n21931);
nand_5 g19583(new_n21931, new_n21875, new_n21932);
nand_5 g19584(new_n21932, new_n21874_1, new_n21933);
xnor_4 g19585(new_n21933, new_n21872, n6853);
xnor_4 g19586(new_n15836, new_n11856, new_n21935);
nor_5  g19587(new_n15841, new_n11861, new_n21936);
xnor_4 g19588(new_n15841, new_n11861, new_n21937);
nor_5  g19589(new_n11864, new_n4383, new_n21938);
not_8  g19590(new_n21938, new_n21939);
nand_5 g19591(new_n13773, new_n13757, new_n21940);
nand_5 g19592(new_n21940, new_n21939, new_n21941);
nor_5  g19593(new_n21941, new_n21937, new_n21942);
nor_5  g19594(new_n21942, new_n21936, new_n21943_1);
xor_4  g19595(new_n21943_1, new_n21935, n6862);
or_5   g19596(new_n7526, n8305, new_n21945);
nand_5 g19597(new_n16830, new_n16815, new_n21946);
nand_5 g19598(new_n21946, new_n21945, new_n21947);
not_8  g19599(new_n21947, new_n21948);
not_8  g19600(n25296, new_n21949);
or_5   g19601(new_n21949, n23717, new_n21950);
nand_5 g19602(new_n12026, new_n12012, new_n21951);
nand_5 g19603(new_n21951, new_n21950, new_n21952);
nand_5 g19604(new_n21952, new_n19550, new_n21953);
not_8  g19605(new_n12011_1, new_n21954);
nand_5 g19606(new_n12028, new_n21954, new_n21955);
nand_5 g19607(new_n12054, new_n12029, new_n21956);
nand_5 g19608(new_n21956, new_n21955, new_n21957_1);
not_8  g19609(new_n21952, new_n21958);
xnor_4 g19610(new_n21958, new_n19550, new_n21959);
nand_5 g19611(new_n21959, new_n21957_1, new_n21960_1);
nand_5 g19612(new_n21960_1, new_n21953, new_n21961);
not_8  g19613(new_n21961, new_n21962);
nand_5 g19614(new_n21962, new_n21948, new_n21963);
nor_5  g19615(new_n16831, new_n12055, new_n21964);
nor_5  g19616(new_n16854, new_n16832, new_n21965);
nor_5  g19617(new_n21965, new_n21964, new_n21966);
not_8  g19618(new_n21966, new_n21967);
nand_5 g19619(new_n21967, new_n21961, new_n21968);
nand_5 g19620(new_n21968, new_n21963, new_n21969);
not_8  g19621(new_n21959, new_n21970);
xnor_4 g19622(new_n21970, new_n21957_1, new_n21971);
not_8  g19623(new_n21971, new_n21972);
nand_5 g19624(new_n21972, new_n21947, new_n21973);
nand_5 g19625(new_n21971, new_n21966, new_n21974);
nand_5 g19626(new_n21974, new_n21973, new_n21975);
nor_5  g19627(new_n21975, new_n21969, n6863);
xnor_4 g19628(new_n6473, new_n6417, n6867);
xnor_4 g19629(new_n18955, new_n18947, n6965);
xnor_4 g19630(new_n7876_1, new_n7829, n6967);
xor_4  g19631(new_n15369, new_n15320, n6975);
xor_4  g19632(new_n21215, new_n21214, n6983);
not_8  g19633(new_n15815_1, new_n21982);
xnor_4 g19634(new_n21982, new_n11842_1, new_n21983);
nand_5 g19635(new_n15821, new_n11845, new_n21984);
xnor_4 g19636(new_n15820, new_n11845, new_n21985);
nor_5  g19637(new_n15824, new_n11848, new_n21986_1);
not_8  g19638(new_n21986_1, new_n21987);
xnor_4 g19639(new_n15824, new_n11849, new_n21988);
nor_5  g19640(new_n15831_1, new_n11853, new_n21989);
nor_5  g19641(new_n15837, new_n11857, new_n21990);
nor_5  g19642(new_n21943_1, new_n21935, new_n21991);
nor_5  g19643(new_n21991, new_n21990, new_n21992);
xnor_4 g19644(new_n15830, new_n11852, new_n21993_1);
nor_5  g19645(new_n21993_1, new_n21992, new_n21994);
nor_5  g19646(new_n21994, new_n21989, new_n21995);
nand_5 g19647(new_n21995, new_n21988, new_n21996);
nand_5 g19648(new_n21996, new_n21987, new_n21997_1);
nand_5 g19649(new_n21997_1, new_n21985, new_n21998);
nand_5 g19650(new_n21998, new_n21984, new_n21999);
xnor_4 g19651(new_n21999, new_n21983, n6985);
xnor_4 g19652(new_n15637, new_n15592, n6998);
xnor_4 g19653(new_n11807, new_n9453, n7032);
xnor_4 g19654(new_n21057, new_n21017_1, n7038);
xnor_4 g19655(new_n18763, new_n18762, n7079);
xnor_4 g19656(new_n7863, new_n17809, n7190);
xnor_4 g19657(new_n16785, new_n16781, n7229);
xnor_4 g19658(new_n9099, new_n9086, n7230);
xnor_4 g19659(new_n20228, new_n20227, n7233);
xnor_4 g19660(new_n14032, new_n14024, n7236);
xnor_4 g19661(new_n17152, new_n7334, n7253);
or_5   g19662(new_n20635, n17458, new_n22011);
or_5   g19663(new_n20636, n12507, new_n22012);
nand_5 g19664(new_n20636, n12507, new_n22013);
nand_5 g19665(new_n20641, new_n22013, new_n22014);
nand_5 g19666(new_n22014, new_n22012, new_n22015);
nand_5 g19667(new_n22015, new_n22011, new_n22016_1);
nand_5 g19668(new_n21133, new_n15005, new_n22017);
xnor_4 g19669(new_n22017, new_n15000, new_n22018);
nand_5 g19670(new_n22018, new_n10764, new_n22019);
xnor_4 g19671(new_n22018, new_n10763_1, new_n22020);
nand_5 g19672(new_n21134_1, new_n20559, new_n22021);
nand_5 g19673(new_n21179, new_n21135, new_n22022);
nand_5 g19674(new_n22022, new_n22021, new_n22023);
nand_5 g19675(new_n22023, new_n22020, new_n22024);
nand_5 g19676(new_n22024, new_n22019, new_n22025);
not_8  g19677(new_n22025, new_n22026);
nor_5  g19678(new_n22017, new_n15000, new_n22027_1);
nor_5  g19679(new_n22027_1, new_n15050, new_n22028);
nand_5 g19680(new_n22027_1, new_n15047, new_n22029);
not_8  g19681(new_n22029, new_n22030);
nor_5  g19682(new_n22030, new_n22028, new_n22031);
xnor_4 g19683(new_n22031, new_n10757, new_n22032);
xnor_4 g19684(new_n22032, new_n22026, new_n22033);
nand_5 g19685(new_n22033, new_n22016_1, new_n22034);
not_8  g19686(new_n22034, new_n22035);
xnor_4 g19687(new_n22033, new_n22016_1, new_n22036);
not_8  g19688(new_n20642, new_n22037);
not_8  g19689(new_n22020, new_n22038);
xnor_4 g19690(new_n22023, new_n22038, new_n22039);
nor_5  g19691(new_n22039, new_n22037, new_n22040);
not_8  g19692(new_n22040, new_n22041);
nor_5  g19693(new_n21180, new_n21122, new_n22042);
not_8  g19694(new_n22042, new_n22043_1);
not_8  g19695(new_n21181, new_n22044);
nand_5 g19696(new_n21232, new_n22044, new_n22045);
nand_5 g19697(new_n22045, new_n22043_1, new_n22046);
xnor_4 g19698(new_n22039, new_n22037, new_n22047);
not_8  g19699(new_n22047, new_n22048);
nand_5 g19700(new_n22048, new_n22046, new_n22049);
nand_5 g19701(new_n22049, new_n22041, new_n22050_1);
nor_5  g19702(new_n22050_1, new_n22036, new_n22051);
nor_5  g19703(new_n22051, new_n22035, new_n22052);
and_5  g19704(new_n22031, new_n20594, new_n22053);
nor_5  g19705(new_n22031, new_n20594, new_n22054);
nor_5  g19706(new_n22054, new_n22025, new_n22055);
nor_5  g19707(new_n22055, new_n22030, new_n22056);
not_8  g19708(new_n22056, new_n22057);
nor_5  g19709(new_n22057, new_n22053, new_n22058);
not_8  g19710(new_n22058, new_n22059);
xnor_4 g19711(new_n22059, new_n22052, n7256);
or_5   g19712(new_n8416, n2416, new_n22061);
xnor_4 g19713(n22764, n2416, new_n22062);
or_5   g19714(new_n8466, n21905, new_n22063_1);
nand_5 g19715(new_n20748_1, new_n20736, new_n22064);
nand_5 g19716(new_n22064, new_n22063_1, new_n22065);
nand_5 g19717(new_n22065, new_n22062, new_n22066);
nand_5 g19718(new_n22066, new_n22061, new_n22067);
not_8  g19719(new_n22067, new_n22068_1);
xnor_4 g19720(new_n22065, new_n22062, new_n22069);
nor_5  g19721(new_n22069, new_n16457, new_n22070);
not_8  g19722(new_n22070, new_n22071);
xnor_4 g19723(new_n22069, new_n16456, new_n22072_1);
not_8  g19724(new_n16460_1, new_n22073);
nor_5  g19725(new_n20749, new_n22073, new_n22074);
not_8  g19726(new_n22074, new_n22075);
nand_5 g19727(new_n20765, new_n20750, new_n22076_1);
nand_5 g19728(new_n22076_1, new_n22075, new_n22077);
nand_5 g19729(new_n22077, new_n22072_1, new_n22078);
nand_5 g19730(new_n22078, new_n22071, new_n22079);
xnor_4 g19731(new_n22079, new_n22068_1, new_n22080);
xnor_4 g19732(new_n22080, new_n16453, new_n22081);
xnor_4 g19733(new_n22081, new_n20860, new_n22082);
xnor_4 g19734(new_n22077, new_n22072_1, new_n22083);
nand_5 g19735(new_n22083, new_n20873, new_n22084);
xnor_4 g19736(new_n22083, new_n20872, new_n22085);
nand_5 g19737(new_n20766, new_n20876, new_n22086);
nand_5 g19738(new_n20784, new_n20767, new_n22087);
nand_5 g19739(new_n22087, new_n22086, new_n22088);
nand_5 g19740(new_n22088, new_n22085, new_n22089);
nand_5 g19741(new_n22089, new_n22084, new_n22090_1);
xnor_4 g19742(new_n22090_1, new_n22082, n7268);
nand_5 g19743(new_n11582, new_n12314, new_n22092);
nor_5  g19744(new_n22092, n2175, new_n22093);
nand_5 g19745(new_n22093, new_n12272, new_n22094);
nor_5  g19746(new_n22094, n23912, new_n22095);
not_8  g19747(new_n22095, new_n22096);
not_8  g19748(n10514, new_n22097);
not_8  g19749(n23912, new_n22098);
xnor_4 g19750(new_n22094, new_n22098, new_n22099);
or_5   g19751(new_n22099, new_n22097, new_n22100);
xnor_4 g19752(new_n22099, n10514, new_n22101);
xnor_4 g19753(new_n22093, n13026, new_n22102);
not_8  g19754(new_n22102, new_n22103);
nand_5 g19755(new_n22103, n18649, new_n22104);
xnor_4 g19756(new_n22102, n18649, new_n22105);
xnor_4 g19757(new_n22092, new_n12310, new_n22106);
not_8  g19758(new_n22106, new_n22107_1);
nand_5 g19759(new_n22107_1, n6218, new_n22108);
xnor_4 g19760(new_n22106, n6218, new_n22109);
nand_5 g19761(new_n11584, n20470, new_n22110);
xnor_4 g19762(new_n11583, n20470, new_n22111);
nand_5 g19763(new_n11588, n21222, new_n22112);
xnor_4 g19764(new_n11587, n21222, new_n22113_1);
nand_5 g19765(new_n11592, n9832, new_n22114);
xnor_4 g19766(new_n11591_1, n9832, new_n22115);
nand_5 g19767(new_n11597, n1558, new_n22116);
xnor_4 g19768(new_n11596, n1558, new_n22117);
nand_5 g19769(new_n11600, n21749, new_n22118);
xnor_4 g19770(new_n11599, n21749, new_n22119);
nand_5 g19771(new_n11604, n7769, new_n22120);
nor_5  g19772(new_n9482, n15506, new_n22121);
xnor_4 g19773(new_n11604, new_n10133, new_n22122);
nand_5 g19774(new_n22122, new_n22121, new_n22123);
nand_5 g19775(new_n22123, new_n22120, new_n22124_1);
nand_5 g19776(new_n22124_1, new_n22119, new_n22125);
nand_5 g19777(new_n22125, new_n22118, new_n22126_1);
nand_5 g19778(new_n22126_1, new_n22117, new_n22127);
nand_5 g19779(new_n22127, new_n22116, new_n22128);
nand_5 g19780(new_n22128, new_n22115, new_n22129);
nand_5 g19781(new_n22129, new_n22114, new_n22130_1);
nand_5 g19782(new_n22130_1, new_n22113_1, new_n22131);
nand_5 g19783(new_n22131, new_n22112, new_n22132);
nand_5 g19784(new_n22132, new_n22111, new_n22133);
nand_5 g19785(new_n22133, new_n22110, new_n22134);
nand_5 g19786(new_n22134, new_n22109, new_n22135);
nand_5 g19787(new_n22135, new_n22108, new_n22136);
nand_5 g19788(new_n22136, new_n22105, new_n22137);
nand_5 g19789(new_n22137, new_n22104, new_n22138);
nand_5 g19790(new_n22138, new_n22101, new_n22139);
nand_5 g19791(new_n22139, new_n22100, new_n22140);
nor_5  g19792(new_n22140, new_n22096, new_n22141);
not_8  g19793(n9872, new_n22142);
xnor_4 g19794(new_n22138, new_n22101, new_n22143);
nand_5 g19795(new_n22143, new_n22142, new_n22144_1);
xnor_4 g19796(new_n22143, n9872, new_n22145);
not_8  g19797(n5842, new_n22146);
xnor_4 g19798(new_n22136, new_n22105, new_n22147);
nand_5 g19799(new_n22147, new_n22146, new_n22148);
xnor_4 g19800(new_n22147, n5842, new_n22149);
not_8  g19801(n6379, new_n22150_1);
xnor_4 g19802(new_n22134, new_n22109, new_n22151);
nand_5 g19803(new_n22151, new_n22150_1, new_n22152);
xnor_4 g19804(new_n22151, n6379, new_n22153);
not_8  g19805(n2102, new_n22154);
xnor_4 g19806(new_n22132, new_n22111, new_n22155);
nand_5 g19807(new_n22155, new_n22154, new_n22156);
xnor_4 g19808(new_n22155, n2102, new_n22157_1);
not_8  g19809(n17954, new_n22158);
xnor_4 g19810(new_n22130_1, new_n22113_1, new_n22159);
nand_5 g19811(new_n22159, new_n22158, new_n22160);
not_8  g19812(n8256, new_n22161);
xnor_4 g19813(new_n22128, new_n22115, new_n22162);
nand_5 g19814(new_n22162, new_n22161, new_n22163);
xnor_4 g19815(new_n22162, n8256, new_n22164);
not_8  g19816(n24150, new_n22165);
xnor_4 g19817(new_n22126_1, new_n22117, new_n22166);
nand_5 g19818(new_n22166, new_n22165, new_n22167);
xnor_4 g19819(new_n22166, n24150, new_n22168);
xnor_4 g19820(new_n22124_1, new_n22119, new_n22169);
nand_5 g19821(new_n22169, new_n17478, new_n22170);
xnor_4 g19822(new_n22169, n19584, new_n22171);
xnor_4 g19823(new_n22122, new_n22121, new_n22172);
nor_5  g19824(new_n22172, new_n17488, new_n22173_1);
not_8  g19825(new_n22172, new_n22174);
nor_5  g19826(new_n22174, n5060, new_n22175);
xnor_4 g19827(n21138, n15506, new_n22176);
nand_5 g19828(new_n22176, n15332, new_n22177);
nor_5  g19829(new_n22177, new_n22175, new_n22178);
nor_5  g19830(new_n22178, new_n22173_1, new_n22179);
nand_5 g19831(new_n22179, new_n22171, new_n22180);
nand_5 g19832(new_n22180, new_n22170, new_n22181);
nand_5 g19833(new_n22181, new_n22168, new_n22182);
nand_5 g19834(new_n22182, new_n22167, new_n22183);
nand_5 g19835(new_n22183, new_n22164, new_n22184);
nand_5 g19836(new_n22184, new_n22163, new_n22185);
xnor_4 g19837(new_n22159, n17954, new_n22186);
nand_5 g19838(new_n22186, new_n22185, new_n22187);
nand_5 g19839(new_n22187, new_n22160, new_n22188);
nand_5 g19840(new_n22188, new_n22157_1, new_n22189);
nand_5 g19841(new_n22189, new_n22156, new_n22190);
nand_5 g19842(new_n22190, new_n22153, new_n22191);
nand_5 g19843(new_n22191, new_n22152, new_n22192);
nand_5 g19844(new_n22192, new_n22149, new_n22193);
nand_5 g19845(new_n22193, new_n22148, new_n22194);
nand_5 g19846(new_n22194, new_n22145, new_n22195);
nand_5 g19847(new_n22195, new_n22144_1, new_n22196);
nand_5 g19848(new_n22196, new_n22141, new_n22197);
not_8  g19849(new_n22196, new_n22198_1);
nand_5 g19850(new_n22140, new_n22096, new_n22199);
not_8  g19851(new_n22199, new_n22200);
nand_5 g19852(new_n22200, new_n22198_1, new_n22201_1);
nand_5 g19853(new_n22201_1, new_n22197, new_n22202);
xnor_4 g19854(new_n22202, new_n15579, new_n22203);
xnor_4 g19855(new_n22140, new_n22095, new_n22204);
xnor_4 g19856(new_n22204, new_n22198_1, new_n22205);
nand_5 g19857(new_n22205, new_n15583, new_n22206);
xnor_4 g19858(new_n22205, new_n15584, new_n22207);
xnor_4 g19859(new_n22194, new_n22145, new_n22208);
nand_5 g19860(new_n22208, new_n2702, new_n22209);
xnor_4 g19861(new_n22208, new_n2701, new_n22210);
xnor_4 g19862(new_n22192, new_n22149, new_n22211);
nand_5 g19863(new_n22211, new_n2832, new_n22212);
xnor_4 g19864(new_n22190, new_n22153, new_n22213_1);
nand_5 g19865(new_n22213_1, new_n2837, new_n22214);
xnor_4 g19866(new_n22213_1, new_n2838, new_n22215);
xnor_4 g19867(new_n22188, new_n22157_1, new_n22216);
nand_5 g19868(new_n22216, new_n2847, new_n22217);
xnor_4 g19869(new_n22216, new_n2843, new_n22218);
xnor_4 g19870(new_n22186, new_n22185, new_n22219);
nand_5 g19871(new_n22219, new_n2850, new_n22220);
xnor_4 g19872(new_n22219, new_n15599, new_n22221);
xnor_4 g19873(new_n22183, new_n22164, new_n22222);
nand_5 g19874(new_n22222, new_n2858_1, new_n22223);
xnor_4 g19875(new_n22222, new_n2854, new_n22224);
xnor_4 g19876(new_n22181, new_n22168, new_n22225);
nand_5 g19877(new_n22225, new_n2864, new_n22226);
xnor_4 g19878(new_n22225, new_n2861, new_n22227);
not_8  g19879(new_n22171, new_n22228);
xnor_4 g19880(new_n22179, new_n22228, new_n22229);
not_8  g19881(new_n22229, new_n22230);
nand_5 g19882(new_n22230, new_n2869, new_n22231);
xnor_4 g19883(new_n22229, new_n2869, new_n22232);
xnor_4 g19884(new_n22172, n5060, new_n22233);
xnor_4 g19885(new_n22233, new_n22177, new_n22234);
nand_5 g19886(new_n22234, new_n2873, new_n22235);
xnor_4 g19887(new_n22176, new_n17502, new_n22236);
nor_5  g19888(new_n22236, new_n2876, new_n22237);
not_8  g19889(new_n22237, new_n22238);
xnor_4 g19890(new_n22234, new_n2880, new_n22239);
nand_5 g19891(new_n22239, new_n22238, new_n22240);
nand_5 g19892(new_n22240, new_n22235, new_n22241);
nand_5 g19893(new_n22241, new_n22232, new_n22242);
nand_5 g19894(new_n22242, new_n22231, new_n22243);
nand_5 g19895(new_n22243, new_n22227, new_n22244);
nand_5 g19896(new_n22244, new_n22226, new_n22245);
nand_5 g19897(new_n22245, new_n22224, new_n22246);
nand_5 g19898(new_n22246, new_n22223, new_n22247);
nand_5 g19899(new_n22247, new_n22221, new_n22248);
nand_5 g19900(new_n22248, new_n22220, new_n22249);
nand_5 g19901(new_n22249, new_n22218, new_n22250);
nand_5 g19902(new_n22250, new_n22217, new_n22251);
nand_5 g19903(new_n22251, new_n22215, new_n22252);
nand_5 g19904(new_n22252, new_n22214, new_n22253_1);
xnor_4 g19905(new_n22211, new_n2831, new_n22254);
nand_5 g19906(new_n22254, new_n22253_1, new_n22255);
nand_5 g19907(new_n22255, new_n22212, new_n22256);
nand_5 g19908(new_n22256, new_n22210, new_n22257);
nand_5 g19909(new_n22257, new_n22209, new_n22258);
nand_5 g19910(new_n22258, new_n22207, new_n22259);
nand_5 g19911(new_n22259, new_n22206, new_n22260);
xnor_4 g19912(new_n22260, new_n22203, n7277);
xnor_4 g19913(new_n14214, new_n14206, n7280);
xnor_4 g19914(new_n6066, new_n6037, n7298);
xnor_4 g19915(new_n20626, new_n20614, n7308);
xnor_4 g19916(new_n20869_1, new_n7684, new_n22265);
not_8  g19917(new_n7706, new_n22266);
not_8  g19918(new_n20871, new_n22267);
nand_5 g19919(new_n22267, new_n22266, new_n22268);
xnor_4 g19920(new_n20871, new_n7706, new_n22269);
not_8  g19921(new_n22269, new_n22270_1);
not_8  g19922(new_n15884_1, new_n22271);
nand_5 g19923(new_n22271, new_n7713, new_n22272);
nand_5 g19924(new_n15913, new_n15885_1, new_n22273);
nand_5 g19925(new_n22273, new_n22272, new_n22274_1);
nand_5 g19926(new_n22274_1, new_n22270_1, new_n22275);
nand_5 g19927(new_n22275, new_n22268, new_n22276);
xnor_4 g19928(new_n22276, new_n22265, new_n22277);
xnor_4 g19929(new_n22277, new_n20898, new_n22278);
xnor_4 g19930(new_n22274_1, new_n22269, new_n22279);
not_8  g19931(new_n22279, new_n22280);
nand_5 g19932(new_n22280, new_n20905, new_n22281);
nor_5  g19933(new_n20203, new_n15914, new_n22282);
nor_5  g19934(new_n20236, new_n20204, new_n22283_1);
nor_5  g19935(new_n22283_1, new_n22282, new_n22284);
xnor_4 g19936(new_n22279, new_n20905, new_n22285);
nand_5 g19937(new_n22285, new_n22284, new_n22286);
nand_5 g19938(new_n22286, new_n22281, new_n22287);
xnor_4 g19939(new_n22287, new_n22278, n7313);
xnor_4 g19940(new_n3865, new_n3839, n7346);
xnor_4 g19941(new_n21952, new_n14900, new_n22290_1);
nand_5 g19942(new_n21952, new_n14903, new_n22291);
xnor_4 g19943(new_n21958, new_n14903, new_n22292);
nand_5 g19944(new_n14911, new_n12027, new_n22293);
xnor_4 g19945(new_n14908, new_n12027, new_n22294);
nand_5 g19946(new_n14915, new_n12032, new_n22295);
xnor_4 g19947(new_n14914, new_n12032, new_n22296);
nand_5 g19948(new_n14920, new_n12038, new_n22297);
nor_5  g19949(new_n6902, new_n6769, new_n22298);
not_8  g19950(new_n6903, new_n22299);
nor_5  g19951(new_n6938, new_n22299, new_n22300);
nor_5  g19952(new_n22300, new_n22298, new_n22301);
xnor_4 g19953(new_n14920, new_n12039, new_n22302);
nand_5 g19954(new_n22302, new_n22301, new_n22303);
nand_5 g19955(new_n22303, new_n22297, new_n22304);
nand_5 g19956(new_n22304, new_n22296, new_n22305);
nand_5 g19957(new_n22305, new_n22295, new_n22306);
nand_5 g19958(new_n22306, new_n22294, new_n22307);
nand_5 g19959(new_n22307, new_n22293, new_n22308);
nand_5 g19960(new_n22308, new_n22292, new_n22309_1);
nand_5 g19961(new_n22309_1, new_n22291, new_n22310);
xnor_4 g19962(new_n22310, new_n22290_1, n7349);
xnor_4 g19963(new_n22256, new_n22210, n7363);
or_5   g19964(n21839, new_n9530, new_n22313);
nand_5 g19965(new_n20846, new_n20843, new_n22314);
nand_5 g19966(new_n22314, new_n22313, new_n22315);
not_8  g19967(new_n22315, new_n22316);
xnor_4 g19968(new_n22316, new_n10820, new_n22317_1);
nand_5 g19969(new_n20847, new_n10824, new_n22318);
nand_5 g19970(new_n20851, new_n20848, new_n22319);
nand_5 g19971(new_n22319, new_n22318, new_n22320);
xnor_4 g19972(new_n22320, new_n22317_1, n7390);
xnor_4 g19973(new_n9640, new_n9639, n7403);
xnor_4 g19974(new_n9834, new_n9791, n7408);
xnor_4 g19975(new_n21226_1, new_n21196, n7432);
nand_5 g19976(new_n19010, new_n16363, new_n22325);
nand_5 g19977(new_n19021, new_n19012, new_n22326);
nand_5 g19978(new_n22326, new_n22325, n7475);
xnor_4 g19979(new_n5476, new_n5475, n7477);
xnor_4 g19980(new_n9468, new_n9440, n7507);
nand_5 g19981(new_n12703, n23895, new_n22330);
xnor_4 g19982(new_n12702_1, n23895, new_n22331);
nand_5 g19983(new_n12706, n17351, new_n22332_1);
nand_5 g19984(new_n7293, new_n7251, new_n22333);
nand_5 g19985(new_n22333, new_n22332_1, new_n22334);
nand_5 g19986(new_n22334, new_n22331, new_n22335_1);
nand_5 g19987(new_n22335_1, new_n22330, new_n22336);
xnor_4 g19988(new_n22336, new_n12757, new_n22337);
xnor_4 g19989(new_n22337, new_n18301_1, new_n22338);
xnor_4 g19990(new_n22334, new_n22331, new_n22339);
nand_5 g19991(new_n22339, new_n18308, new_n22340);
xnor_4 g19992(new_n22339, new_n18309, new_n22341_1);
nand_5 g19993(new_n7294, new_n7215, new_n22342);
nand_5 g19994(new_n7356, new_n7295, new_n22343);
nand_5 g19995(new_n22343, new_n22342, new_n22344);
nand_5 g19996(new_n22344, new_n22341_1, new_n22345);
nand_5 g19997(new_n22345, new_n22340, new_n22346);
xnor_4 g19998(new_n22346, new_n22338, n7514);
xnor_4 g19999(new_n11562, new_n11534, n7558);
xnor_4 g20000(new_n12808, new_n12806, n7572);
xnor_4 g20001(new_n6597, n7693, new_n22350);
nor_5  g20002(new_n6598, new_n4189, new_n22351);
not_8  g20003(new_n21250, new_n22352);
nor_5  g20004(new_n21261, new_n22352, new_n22353_1);
nor_5  g20005(new_n22353_1, new_n22351, new_n22354);
xnor_4 g20006(new_n22354, new_n22350, new_n22355);
xnor_4 g20007(new_n22355, new_n10331, new_n22356);
not_8  g20008(new_n22356, new_n22357);
nor_5  g20009(new_n21262, new_n10338, new_n22358_1);
nor_5  g20010(new_n21278, new_n21264, new_n22359_1);
nor_5  g20011(new_n22359_1, new_n22358_1, new_n22360);
xnor_4 g20012(new_n22360, new_n22357, n7575);
xnor_4 g20013(new_n22102, new_n10258, new_n22362);
nor_5  g20014(new_n22107_1, new_n10313, new_n22363);
xnor_4 g20015(new_n22107_1, new_n10313, new_n22364);
nor_5  g20016(new_n11584, new_n10319, new_n22365);
nor_5  g20017(new_n11619, new_n11585, new_n22366);
nor_5  g20018(new_n22366, new_n22365, new_n22367);
nor_5  g20019(new_n22367, new_n22364, new_n22368);
nor_5  g20020(new_n22368, new_n22363, new_n22369);
xnor_4 g20021(new_n22369, new_n22362, new_n22370);
xnor_4 g20022(new_n22370, new_n12237, new_n22371);
xnor_4 g20023(new_n22367, new_n22364, new_n22372);
nor_5  g20024(new_n22372, new_n12244, new_n22373);
xnor_4 g20025(new_n22372, new_n12244, new_n22374);
nand_5 g20026(new_n12250, new_n11620, new_n22375);
nand_5 g20027(new_n11673, new_n11635, new_n22376);
nand_5 g20028(new_n22376, new_n22375, new_n22377);
nor_5  g20029(new_n22377, new_n22374, new_n22378);
nor_5  g20030(new_n22378, new_n22373, new_n22379_1);
nor_5  g20031(new_n22379_1, new_n22371, new_n22380);
and_5  g20032(new_n22379_1, new_n22371, new_n22381);
nor_5  g20033(new_n22381, new_n22380, n7585);
xnor_4 g20034(new_n21792, new_n8193, new_n22383);
nand_5 g20035(new_n21797, new_n8197, new_n22384);
xnor_4 g20036(new_n21797, new_n8196, new_n22385);
nand_5 g20037(new_n21804, new_n8201, new_n22386);
xnor_4 g20038(new_n21803, new_n8201, new_n22387);
nand_5 g20039(new_n21810, new_n8206, new_n22388);
xnor_4 g20040(new_n21810, new_n8209, new_n22389);
nand_5 g20041(new_n19107_1, new_n8212, new_n22390);
xnor_4 g20042(new_n19107_1, new_n8211, new_n22391);
nand_5 g20043(new_n19110, new_n8218, new_n22392);
xnor_4 g20044(new_n19110, new_n8217, new_n22393);
not_8  g20045(new_n19115, new_n22394);
nand_5 g20046(new_n22394, new_n8223, new_n22395);
xnor_4 g20047(new_n19115, new_n8223, new_n22396);
nor_5  g20048(new_n19122, new_n8234, new_n22397);
xnor_4 g20049(new_n19121, new_n8234, new_n22398);
not_8  g20050(new_n22398, new_n22399);
nor_5  g20051(new_n19130, new_n8242, new_n22400);
nor_5  g20052(new_n22400, new_n8238, new_n22401);
not_8  g20053(new_n22401, new_n22402);
xnor_4 g20054(new_n22400, new_n8237, new_n22403);
nand_5 g20055(new_n22403, new_n19137, new_n22404);
nand_5 g20056(new_n22404, new_n22402, new_n22405);
not_8  g20057(new_n22405, new_n22406);
nor_5  g20058(new_n22406, new_n22399, new_n22407);
nor_5  g20059(new_n22407, new_n22397, new_n22408);
not_8  g20060(new_n22408, new_n22409);
nand_5 g20061(new_n22409, new_n22396, new_n22410);
nand_5 g20062(new_n22410, new_n22395, new_n22411);
nand_5 g20063(new_n22411, new_n22393, new_n22412);
nand_5 g20064(new_n22412, new_n22392, new_n22413);
nand_5 g20065(new_n22413, new_n22391, new_n22414);
nand_5 g20066(new_n22414, new_n22390, new_n22415);
nand_5 g20067(new_n22415, new_n22389, new_n22416);
nand_5 g20068(new_n22416, new_n22388, new_n22417);
nand_5 g20069(new_n22417, new_n22387, new_n22418);
nand_5 g20070(new_n22418, new_n22386, new_n22419);
nand_5 g20071(new_n22419, new_n22385, new_n22420);
nand_5 g20072(new_n22420, new_n22384, new_n22421);
xnor_4 g20073(new_n22421, new_n22383, n7588);
not_8  g20074(new_n15278, new_n22423);
nand_5 g20075(new_n7038_1, new_n2353, new_n22424);
nor_5  g20076(new_n22424, n21753, new_n22425);
nand_5 g20077(new_n22425, new_n11911, new_n22426);
nor_5  g20078(new_n22426, n13074, new_n22427);
xnor_4 g20079(new_n22427, n23463, new_n22428);
xnor_4 g20080(new_n22428, new_n17002, new_n22429);
xnor_4 g20081(new_n22426, new_n3171, new_n22430);
or_5   g20082(new_n22430, n11455, new_n22431);
xnor_4 g20083(new_n22430, new_n16920, new_n22432);
xnor_4 g20084(new_n22425, n10739, new_n22433_1);
or_5   g20085(new_n22433_1, n3945, new_n22434);
xnor_4 g20086(new_n22433_1, new_n16923, new_n22435);
xnor_4 g20087(new_n22424, new_n2350, new_n22436);
or_5   g20088(new_n22436, n5255, new_n22437);
xnor_4 g20089(new_n22436, new_n16926, new_n22438);
not_8  g20090(new_n7039, new_n22439);
nand_5 g20091(new_n22439, new_n5428, new_n22440);
xnor_4 g20092(new_n7039, new_n5428, new_n22441);
not_8  g20093(new_n7058, new_n22442_1);
nand_5 g20094(new_n22442_1, new_n5432, new_n22443);
nand_5 g20095(new_n7080, new_n5436, new_n22444_1);
xnor_4 g20096(new_n7076, new_n5436, new_n22445);
not_8  g20097(new_n7071, new_n22446);
nand_5 g20098(new_n22446, new_n5332, new_n22447);
nand_5 g20099(n21654, n2387, new_n22448);
xnor_4 g20100(new_n7071, new_n5332, new_n22449);
nand_5 g20101(new_n22449, new_n22448, new_n22450);
nand_5 g20102(new_n22450, new_n22447, new_n22451);
nand_5 g20103(new_n22451, new_n22445, new_n22452);
nand_5 g20104(new_n22452, new_n22444_1, new_n22453);
xnor_4 g20105(new_n7058, new_n5432, new_n22454);
nand_5 g20106(new_n22454, new_n22453, new_n22455);
nand_5 g20107(new_n22455, new_n22443, new_n22456);
nand_5 g20108(new_n22456, new_n22441, new_n22457);
nand_5 g20109(new_n22457, new_n22440, new_n22458);
nand_5 g20110(new_n22458, new_n22438, new_n22459);
nand_5 g20111(new_n22459, new_n22437, new_n22460);
nand_5 g20112(new_n22460, new_n22435, new_n22461);
nand_5 g20113(new_n22461, new_n22434, new_n22462);
nand_5 g20114(new_n22462, new_n22432, new_n22463);
nand_5 g20115(new_n22463, new_n22431, new_n22464);
xnor_4 g20116(new_n22464, new_n22429, new_n22465);
xnor_4 g20117(new_n22465, new_n22423, new_n22466);
not_8  g20118(new_n22466, new_n22467_1);
xnor_4 g20119(new_n22462, new_n22432, new_n22468);
nor_5  g20120(new_n22468, new_n15316, new_n22469);
xnor_4 g20121(new_n22468, new_n15316, new_n22470_1);
xnor_4 g20122(new_n22460, new_n22435, new_n22471);
nand_5 g20123(new_n22471, new_n15322, new_n22472);
not_8  g20124(new_n15322, new_n22473);
xnor_4 g20125(new_n22471, new_n22473, new_n22474);
xnor_4 g20126(new_n22458, new_n22438, new_n22475);
nand_5 g20127(new_n22475, new_n15327_1, new_n22476);
xnor_4 g20128(new_n22456, new_n22441, new_n22477);
nand_5 g20129(new_n22477, new_n15332_1, new_n22478);
not_8  g20130(new_n15338, new_n22479);
xnor_4 g20131(new_n22454, new_n22453, new_n22480);
nand_5 g20132(new_n22480, new_n22479, new_n22481);
xnor_4 g20133(new_n22480, new_n15338, new_n22482);
not_8  g20134(new_n15343, new_n22483);
xnor_4 g20135(new_n22451, new_n22445, new_n22484_1);
nand_5 g20136(new_n22484_1, new_n22483, new_n22485);
xnor_4 g20137(new_n22484_1, new_n15343, new_n22486);
nor_5  g20138(new_n22449, new_n15349, new_n22487);
not_8  g20139(new_n22448, new_n22488);
xnor_4 g20140(new_n22449, new_n22488, new_n22489_1);
nor_5  g20141(new_n22489_1, new_n15348, new_n22490);
xnor_4 g20142(n21654, new_n2368, new_n22491);
and_5  g20143(new_n22491, new_n15354, new_n22492_1);
nor_5  g20144(new_n22492_1, new_n22490, new_n22493);
nor_5  g20145(new_n22493, new_n22487, new_n22494_1);
nand_5 g20146(new_n22494_1, new_n22486, new_n22495);
nand_5 g20147(new_n22495, new_n22485, new_n22496);
nand_5 g20148(new_n22496, new_n22482, new_n22497);
nand_5 g20149(new_n22497, new_n22481, new_n22498);
xnor_4 g20150(new_n22477, new_n15333, new_n22499);
nand_5 g20151(new_n22499, new_n22498, new_n22500);
nand_5 g20152(new_n22500, new_n22478, new_n22501);
xnor_4 g20153(new_n22475, new_n15326, new_n22502);
nand_5 g20154(new_n22502, new_n22501, new_n22503);
nand_5 g20155(new_n22503, new_n22476, new_n22504);
nand_5 g20156(new_n22504, new_n22474, new_n22505);
nand_5 g20157(new_n22505, new_n22472, new_n22506);
nor_5  g20158(new_n22506, new_n22470_1, new_n22507);
nor_5  g20159(new_n22507, new_n22469, new_n22508);
xnor_4 g20160(new_n22508, new_n22467_1, n7598);
xnor_4 g20161(new_n19019, new_n19016, n7607);
xnor_4 g20162(new_n5282, new_n5251, n7610);
xnor_4 g20163(new_n3503, new_n3485, n7616);
xnor_4 g20164(n10514, new_n6641, new_n22513);
nor_5  g20165(n18649, n3795, new_n22514);
xnor_4 g20166(n18649, new_n6645, new_n22515);
not_8  g20167(new_n22515, new_n22516);
nor_5  g20168(n25464, n6218, new_n22517);
xnor_4 g20169(n25464, new_n12116, new_n22518);
not_8  g20170(new_n22518, new_n22519);
nor_5  g20171(n20470, n4590, new_n22520);
xnor_4 g20172(n20470, new_n6652_1, new_n22521);
not_8  g20173(new_n22521, new_n22522);
nor_5  g20174(n26752, n21222, new_n22523);
xnor_4 g20175(n26752, new_n11623, new_n22524);
not_8  g20176(new_n22524, new_n22525);
nor_5  g20177(n9832, n6513, new_n22526);
xnor_4 g20178(n9832, new_n6659_1, new_n22527);
not_8  g20179(new_n22527, new_n22528);
nand_5 g20180(n3918, n1558, new_n22529);
nor_5  g20181(n3918, n1558, new_n22530);
not_8  g20182(new_n22530, new_n22531);
nor_5  g20183(n21749, n919, new_n22532);
not_8  g20184(new_n17479, new_n22533_1);
nor_5  g20185(new_n17485, new_n22533_1, new_n22534);
nor_5  g20186(new_n22534, new_n22532, new_n22535);
nand_5 g20187(new_n22535, new_n22531, new_n22536);
nand_5 g20188(new_n22536, new_n22529, new_n22537);
nor_5  g20189(new_n22537, new_n22528, new_n22538);
nor_5  g20190(new_n22538, new_n22526, new_n22539);
nor_5  g20191(new_n22539, new_n22525, new_n22540);
nor_5  g20192(new_n22540, new_n22523, new_n22541);
nor_5  g20193(new_n22541, new_n22522, new_n22542);
nor_5  g20194(new_n22542, new_n22520, new_n22543);
nor_5  g20195(new_n22543, new_n22519, new_n22544);
nor_5  g20196(new_n22544, new_n22517, new_n22545);
nor_5  g20197(new_n22545, new_n22516, new_n22546);
nor_5  g20198(new_n22546, new_n22514, new_n22547);
xnor_4 g20199(new_n22547, new_n22513, new_n22548);
nand_5 g20200(new_n22548, n9872, new_n22549);
xnor_4 g20201(new_n22548, new_n22142, new_n22550);
xnor_4 g20202(new_n22545, new_n22515, new_n22551);
nand_5 g20203(new_n22551, n5842, new_n22552);
xnor_4 g20204(new_n22551, new_n22146, new_n22553);
xnor_4 g20205(new_n22543, new_n22518, new_n22554_1);
nand_5 g20206(new_n22554_1, n6379, new_n22555);
xnor_4 g20207(new_n22554_1, new_n22150_1, new_n22556);
xnor_4 g20208(new_n22541, new_n22521, new_n22557);
nand_5 g20209(new_n22557, n2102, new_n22558);
xnor_4 g20210(new_n22557, new_n22154, new_n22559);
xnor_4 g20211(new_n22539, new_n22524, new_n22560);
nand_5 g20212(new_n22560, n17954, new_n22561);
xnor_4 g20213(new_n22560, new_n22158, new_n22562);
xnor_4 g20214(new_n22537, new_n22527, new_n22563);
nand_5 g20215(new_n22563, n8256, new_n22564);
xnor_4 g20216(new_n22563, new_n22161, new_n22565);
xnor_4 g20217(n3918, new_n10124, new_n22566);
xnor_4 g20218(new_n22566, new_n22535, new_n22567);
nand_5 g20219(new_n22567, n24150, new_n22568);
xnor_4 g20220(new_n22567, new_n22165, new_n22569);
nand_5 g20221(new_n17486, n19584, new_n22570);
nand_5 g20222(new_n17497, new_n17487, new_n22571);
nand_5 g20223(new_n22571, new_n22570, new_n22572);
nand_5 g20224(new_n22572, new_n22569, new_n22573);
nand_5 g20225(new_n22573, new_n22568, new_n22574);
nand_5 g20226(new_n22574, new_n22565, new_n22575);
nand_5 g20227(new_n22575, new_n22564, new_n22576);
nand_5 g20228(new_n22576, new_n22562, new_n22577);
nand_5 g20229(new_n22577, new_n22561, new_n22578);
nand_5 g20230(new_n22578, new_n22559, new_n22579);
nand_5 g20231(new_n22579, new_n22558, new_n22580);
nand_5 g20232(new_n22580, new_n22556, new_n22581);
nand_5 g20233(new_n22581, new_n22555, new_n22582);
nand_5 g20234(new_n22582, new_n22553, new_n22583);
nand_5 g20235(new_n22583, new_n22552, new_n22584_1);
nand_5 g20236(new_n22584_1, new_n22550, new_n22585);
nand_5 g20237(new_n22585, new_n22549, new_n22586);
or_5   g20238(n10514, n6105, new_n22587);
not_8  g20239(new_n22547, new_n22588_1);
nand_5 g20240(new_n22588_1, new_n22513, new_n22589_1);
nand_5 g20241(new_n22589_1, new_n22587, new_n22590);
nand_5 g20242(new_n22590, new_n22586, new_n22591_1);
xnor_4 g20243(new_n22591_1, new_n16624, new_n22592);
xnor_4 g20244(new_n22590, new_n22586, new_n22593);
nor_5  g20245(new_n22593, new_n16502_1, new_n22594);
xnor_4 g20246(new_n22593, new_n16502_1, new_n22595);
xnor_4 g20247(new_n22584_1, new_n22550, new_n22596);
not_8  g20248(new_n22596, new_n22597_1);
nand_5 g20249(new_n22597_1, new_n16551, new_n22598);
xnor_4 g20250(new_n22596, new_n16551, new_n22599);
xnor_4 g20251(new_n22582, new_n22553, new_n22600);
not_8  g20252(new_n22600, new_n22601);
nand_5 g20253(new_n22601, new_n16556, new_n22602);
xnor_4 g20254(new_n22600, new_n16556, new_n22603);
xnor_4 g20255(new_n22580, new_n22556, new_n22604);
not_8  g20256(new_n22604, new_n22605);
nand_5 g20257(new_n22605, new_n16561, new_n22606);
xnor_4 g20258(new_n22604, new_n16561, new_n22607);
xnor_4 g20259(new_n22578, new_n22559, new_n22608);
not_8  g20260(new_n22608, new_n22609);
nand_5 g20261(new_n22609, new_n16566, new_n22610);
xnor_4 g20262(new_n22608, new_n16566, new_n22611);
xnor_4 g20263(new_n22576, new_n22562, new_n22612);
not_8  g20264(new_n22612, new_n22613);
nand_5 g20265(new_n22613, new_n16571, new_n22614);
xnor_4 g20266(new_n22612, new_n16571, new_n22615);
xnor_4 g20267(new_n22574, new_n22565, new_n22616);
not_8  g20268(new_n22616, new_n22617);
nand_5 g20269(new_n22617, new_n16576, new_n22618);
xnor_4 g20270(new_n22616, new_n16576, new_n22619_1);
not_8  g20271(new_n22569, new_n22620_1);
xnor_4 g20272(new_n22572, new_n22620_1, new_n22621);
nand_5 g20273(new_n22621, new_n16581, new_n22622);
xnor_4 g20274(new_n22621, new_n16583_1, new_n22623_1);
not_8  g20275(new_n17498, new_n22624);
nand_5 g20276(new_n22624, new_n16587, new_n22625);
nand_5 g20277(new_n17508, new_n17499, new_n22626_1);
nand_5 g20278(new_n22626_1, new_n22625, new_n22627);
nand_5 g20279(new_n22627, new_n22623_1, new_n22628);
nand_5 g20280(new_n22628, new_n22622, new_n22629);
nand_5 g20281(new_n22629, new_n22619_1, new_n22630);
nand_5 g20282(new_n22630, new_n22618, new_n22631_1);
nand_5 g20283(new_n22631_1, new_n22615, new_n22632);
nand_5 g20284(new_n22632, new_n22614, new_n22633);
nand_5 g20285(new_n22633, new_n22611, new_n22634);
nand_5 g20286(new_n22634, new_n22610, new_n22635);
nand_5 g20287(new_n22635, new_n22607, new_n22636);
nand_5 g20288(new_n22636, new_n22606, new_n22637);
nand_5 g20289(new_n22637, new_n22603, new_n22638);
nand_5 g20290(new_n22638, new_n22602, new_n22639);
nand_5 g20291(new_n22639, new_n22599, new_n22640);
nand_5 g20292(new_n22640, new_n22598, new_n22641);
not_8  g20293(new_n22641, new_n22642);
nor_5  g20294(new_n22642, new_n22595, new_n22643);
nor_5  g20295(new_n22643, new_n22594, new_n22644);
xnor_4 g20296(new_n22644, new_n22592, n7630);
nand_5 g20297(new_n19932, new_n19908, new_n22646);
nand_5 g20298(new_n19943, new_n19933, new_n22647);
nand_5 g20299(new_n22647, new_n22646, new_n22648);
not_8  g20300(new_n22648, n7643);
xnor_4 g20301(new_n12955, new_n12924, n7647);
xnor_4 g20302(new_n10684, new_n10646, n7679);
xnor_4 g20303(new_n21466, new_n21438, n7686);
xnor_4 g20304(new_n19390, new_n19363, new_n22653);
xnor_4 g20305(new_n22653, new_n19409, n7698);
xnor_4 g20306(new_n20628, new_n20607, n7708);
xnor_4 g20307(new_n19377, new_n16856, new_n22656);
not_8  g20308(new_n22656, new_n22657);
nor_5  g20309(new_n19382, new_n16884, new_n22658);
xnor_4 g20310(new_n2985_1, new_n16884, new_n22659);
not_8  g20311(new_n22659, new_n22660_1);
nor_5  g20312(new_n21832_1, n21997, new_n22661);
not_8  g20313(new_n22661, new_n22662);
xnor_4 g20314(new_n3034, n21997, new_n22663);
nor_5  g20315(new_n3041, n25119, new_n22664);
not_8  g20316(new_n22664, new_n22665);
nand_5 g20317(new_n9061, new_n9033, new_n22666);
nand_5 g20318(new_n22666, new_n22665, new_n22667);
nand_5 g20319(new_n22667, new_n22663, new_n22668);
nand_5 g20320(new_n22668, new_n22662, new_n22669);
nor_5  g20321(new_n22669, new_n22660_1, new_n22670);
nor_5  g20322(new_n22670, new_n22658, new_n22671);
xnor_4 g20323(new_n22671, new_n22657, new_n22672);
xnor_4 g20324(new_n6355, new_n5220, new_n22673);
nor_5  g20325(new_n6357, n2858, new_n22674);
nor_5  g20326(new_n17229, new_n17222, new_n22675);
nor_5  g20327(new_n22675, new_n22674, new_n22676);
xnor_4 g20328(new_n22676, new_n22673, new_n22677);
xnor_4 g20329(new_n22677, new_n22672, new_n22678);
xnor_4 g20330(new_n22669, new_n22660_1, new_n22679);
nand_5 g20331(new_n22679, new_n17230, new_n22680);
xnor_4 g20332(new_n22679, new_n17231, new_n22681);
not_8  g20333(new_n22663, new_n22682);
xnor_4 g20334(new_n22667, new_n22682, new_n22683);
nand_5 g20335(new_n22683, new_n17236_1, new_n22684);
xnor_4 g20336(new_n22683, new_n17233, new_n22685);
nand_5 g20337(new_n9062, new_n18572_1, new_n22686);
nand_5 g20338(new_n9108, new_n9063, new_n22687);
nand_5 g20339(new_n22687, new_n22686, new_n22688);
nand_5 g20340(new_n22688, new_n22685, new_n22689);
nand_5 g20341(new_n22689, new_n22684, new_n22690);
nand_5 g20342(new_n22690, new_n22681, new_n22691);
nand_5 g20343(new_n22691, new_n22680, new_n22692);
xnor_4 g20344(new_n22692, new_n22678, n7780);
not_8  g20345(new_n15578, new_n22694);
nor_5  g20346(new_n2634, new_n4661, new_n22695);
xnor_4 g20347(new_n2634, new_n4661, new_n22696);
nor_5  g20348(new_n2638, new_n4618, new_n22697_1);
xnor_4 g20349(new_n2638, new_n4618, new_n22698);
nor_5  g20350(new_n10257, new_n22698, new_n22699);
nor_5  g20351(new_n22699, new_n22697_1, new_n22700);
nor_5  g20352(new_n22700, new_n22696, new_n22701);
nor_5  g20353(new_n22701, new_n22695, new_n22702);
xnor_4 g20354(new_n22702, new_n22694, new_n22703);
not_8  g20355(new_n22703, new_n22704);
not_8  g20356(new_n18401, new_n22705);
nor_5  g20357(new_n22705, new_n2766, new_n22706);
xnor_4 g20358(new_n18401, new_n2766, new_n22707);
not_8  g20359(new_n22707, new_n22708);
not_8  g20360(new_n10264, new_n22709);
nor_5  g20361(new_n22709, new_n2771, new_n22710);
not_8  g20362(new_n10265, new_n22711);
nor_5  g20363(new_n10310, new_n22711, new_n22712);
nor_5  g20364(new_n22712, new_n22710, new_n22713);
nor_5  g20365(new_n22713, new_n22708, new_n22714_1);
nor_5  g20366(new_n22714_1, new_n22706, new_n22715);
nor_5  g20367(new_n18400, n21839, new_n22716);
xnor_4 g20368(new_n22716, new_n16776, new_n22717);
xnor_4 g20369(new_n22717, new_n22715, new_n22718);
xnor_4 g20370(new_n22718, new_n22704, new_n22719);
xnor_4 g20371(new_n22700, new_n22696, new_n22720);
not_8  g20372(new_n22720, new_n22721);
xnor_4 g20373(new_n22713, new_n22707, new_n22722);
nor_5  g20374(new_n22722, new_n22721, new_n22723);
xnor_4 g20375(new_n22722, new_n22721, new_n22724);
nor_5  g20376(new_n10311, new_n10258, new_n22725);
nor_5  g20377(new_n10372_1, new_n10312, new_n22726);
nor_5  g20378(new_n22726, new_n22725, new_n22727);
nor_5  g20379(new_n22727, new_n22724, new_n22728);
nor_5  g20380(new_n22728, new_n22723, new_n22729);
xnor_4 g20381(new_n22729, new_n22719, n7794);
xnor_4 g20382(new_n18594, new_n18587, n7811);
xor_4  g20383(new_n18539, new_n18532, n7830);
xnor_4 g20384(new_n22417, new_n22387, n7834);
xnor_4 g20385(new_n11667_1, new_n11652, n7884);
xnor_4 g20386(new_n3146, new_n3144, n7937);
xnor_4 g20387(new_n3159, new_n3106, n7943);
xor_4  g20388(new_n10366, new_n10330_1, n7950);
xnor_4 g20389(new_n20902, new_n16452, new_n22738);
not_8  g20390(new_n22738, new_n22739);
nand_5 g20391(new_n20907, new_n16457, new_n22740);
nand_5 g20392(new_n20909, new_n22073, new_n22741);
xnor_4 g20393(new_n20909, new_n16460_1, new_n22742);
not_8  g20394(new_n16185_1, new_n22743);
nand_5 g20395(new_n22743, new_n16140, new_n22744);
nand_5 g20396(new_n16234, new_n16186, new_n22745);
nand_5 g20397(new_n22745, new_n22744, new_n22746);
nand_5 g20398(new_n22746, new_n22742, new_n22747);
nand_5 g20399(new_n22747, new_n22741, new_n22748);
xnor_4 g20400(new_n20907, new_n16456, new_n22749);
nand_5 g20401(new_n22749, new_n22748, new_n22750);
nand_5 g20402(new_n22750, new_n22740, new_n22751);
xnor_4 g20403(new_n22751, new_n22739, n7959);
xnor_4 g20404(new_n18599, new_n18581, n7968);
xnor_4 g20405(new_n19644, new_n19642, n7992);
xnor_4 g20406(new_n13693, new_n8278, new_n22755);
not_8  g20407(new_n22755, new_n22756);
nand_5 g20408(new_n13696, n26408, new_n22757);
xnor_4 g20409(new_n13696, new_n8267_1, new_n22758);
nor_5  g20410(new_n11220_1, n18227, new_n22759);
nor_5  g20411(new_n18569, new_n18555, new_n22760);
nor_5  g20412(new_n22760, new_n22759, new_n22761_1);
nand_5 g20413(new_n22761_1, new_n22758, new_n22762);
nand_5 g20414(new_n22762, new_n22757, new_n22763);
xnor_4 g20415(new_n22763, new_n22756, new_n22764_1);
xnor_4 g20416(new_n22764_1, new_n19823, new_n22765);
not_8  g20417(new_n22758, new_n22766);
xnor_4 g20418(new_n22761_1, new_n22766, new_n22767);
nand_5 g20419(new_n22767, new_n19832, new_n22768);
xnor_4 g20420(new_n22767, new_n19828, new_n22769);
nand_5 g20421(new_n19838, new_n18570, new_n22770);
xnor_4 g20422(new_n19834, new_n18570, new_n22771);
not_8  g20423(new_n18573, new_n22772);
nand_5 g20424(new_n19841, new_n22772, new_n22773);
xnor_4 g20425(new_n19841, new_n18573, new_n22774);
nand_5 g20426(new_n19851, new_n18577, new_n22775);
xnor_4 g20427(new_n19849, new_n18577, new_n22776);
not_8  g20428(new_n13782, new_n22777);
nor_5  g20429(new_n13796, new_n22777, new_n22778);
not_8  g20430(new_n22778, new_n22779_1);
nand_5 g20431(new_n13802, new_n13797, new_n22780);
nand_5 g20432(new_n22780, new_n22779_1, new_n22781);
nand_5 g20433(new_n22781, new_n22776, new_n22782);
nand_5 g20434(new_n22782, new_n22775, new_n22783);
nand_5 g20435(new_n22783, new_n22774, new_n22784);
nand_5 g20436(new_n22784, new_n22773, new_n22785);
nand_5 g20437(new_n22785, new_n22771, new_n22786);
nand_5 g20438(new_n22786, new_n22770, new_n22787_1);
nand_5 g20439(new_n22787_1, new_n22769, new_n22788);
nand_5 g20440(new_n22788, new_n22768, new_n22789);
xnor_4 g20441(new_n22789, new_n22765, n7999);
xnor_4 g20442(new_n19267, new_n19251, n8027);
nor_5  g20443(new_n22702, new_n15578, new_n22792);
nor_5  g20444(new_n6575, new_n6526, new_n22793_1);
xnor_4 g20445(new_n6574, new_n6526, new_n22794);
not_8  g20446(new_n22794, new_n22795);
nor_5  g20447(new_n6582, new_n6542_1, new_n22796);
nor_5  g20448(new_n13170, n27037, new_n22797);
not_8  g20449(new_n22797, new_n22798);
xnor_4 g20450(new_n6587_1, n27037, new_n22799);
nor_5  g20451(new_n13206, n8964, new_n22800);
not_8  g20452(new_n22800, new_n22801);
xnor_4 g20453(new_n6590_1, n8964, new_n22802);
nor_5  g20454(new_n6593, new_n6557, new_n22803);
nor_5  g20455(new_n6597, new_n4185, new_n22804);
not_8  g20456(new_n22350, new_n22805);
nor_5  g20457(new_n22354, new_n22805, new_n22806);
nor_5  g20458(new_n22806, new_n22804, new_n22807);
xnor_4 g20459(new_n6593, n20151, new_n22808);
not_8  g20460(new_n22808, new_n22809);
nor_5  g20461(new_n22809, new_n22807, new_n22810);
nor_5  g20462(new_n22810, new_n22803, new_n22811);
nand_5 g20463(new_n22811, new_n22802, new_n22812);
nand_5 g20464(new_n22812, new_n22801, new_n22813);
nand_5 g20465(new_n22813, new_n22799, new_n22814);
nand_5 g20466(new_n22814, new_n22798, new_n22815);
xnor_4 g20467(new_n6581, new_n6542_1, new_n22816);
not_8  g20468(new_n22816, new_n22817);
nor_5  g20469(new_n22817, new_n22815, new_n22818);
nor_5  g20470(new_n22818, new_n22796, new_n22819_1);
nor_5  g20471(new_n22819_1, new_n22795, new_n22820);
nor_5  g20472(new_n22820, new_n22793_1, new_n22821);
nor_5  g20473(new_n22821, new_n6525, new_n22822);
not_8  g20474(new_n22822, new_n22823);
nand_5 g20475(new_n22823, new_n22792, new_n22824);
not_8  g20476(new_n22792, new_n22825);
nand_5 g20477(new_n22822, new_n22825, new_n22826);
xnor_4 g20478(new_n22821, new_n13111, new_n22827);
not_8  g20479(new_n22827, new_n22828);
nand_5 g20480(new_n22828, new_n22703, new_n22829);
xnor_4 g20481(new_n22827, new_n22703, new_n22830);
xnor_4 g20482(new_n22819_1, new_n22795, new_n22831);
nand_5 g20483(new_n22831, new_n22721, new_n22832);
xnor_4 g20484(new_n22831, new_n22720, new_n22833);
xnor_4 g20485(new_n22816, new_n22815, new_n22834);
not_8  g20486(new_n22834, new_n22835);
nand_5 g20487(new_n22835, new_n10258, new_n22836);
xnor_4 g20488(new_n22834, new_n10258, new_n22837);
not_8  g20489(new_n10313, new_n22838);
not_8  g20490(new_n22799, new_n22839);
xnor_4 g20491(new_n22813, new_n22839, new_n22840);
nand_5 g20492(new_n22840, new_n22838, new_n22841);
xnor_4 g20493(new_n22840, new_n10313, new_n22842);
not_8  g20494(new_n22802, new_n22843_1);
xnor_4 g20495(new_n22811, new_n22843_1, new_n22844);
nand_5 g20496(new_n22844, new_n10320, new_n22845);
xnor_4 g20497(new_n22844, new_n10319, new_n22846);
not_8  g20498(new_n10325, new_n22847);
xnor_4 g20499(new_n22809, new_n22807, new_n22848);
nand_5 g20500(new_n22848, new_n22847, new_n22849);
xnor_4 g20501(new_n22848, new_n10325, new_n22850);
nor_5  g20502(new_n22355, new_n10332, new_n22851);
nor_5  g20503(new_n22360, new_n22357, new_n22852);
nor_5  g20504(new_n22852, new_n22851, new_n22853);
not_8  g20505(new_n22853, new_n22854);
nand_5 g20506(new_n22854, new_n22850, new_n22855);
nand_5 g20507(new_n22855, new_n22849, new_n22856);
nand_5 g20508(new_n22856, new_n22846, new_n22857);
nand_5 g20509(new_n22857, new_n22845, new_n22858_1);
nand_5 g20510(new_n22858_1, new_n22842, new_n22859);
nand_5 g20511(new_n22859, new_n22841, new_n22860);
nand_5 g20512(new_n22860, new_n22837, new_n22861);
nand_5 g20513(new_n22861, new_n22836, new_n22862);
nand_5 g20514(new_n22862, new_n22833, new_n22863);
nand_5 g20515(new_n22863, new_n22832, new_n22864);
nand_5 g20516(new_n22864, new_n22830, new_n22865);
nand_5 g20517(new_n22865, new_n22829, new_n22866);
nand_5 g20518(new_n22866, new_n22826, new_n22867);
nand_5 g20519(new_n22867, new_n22824, n8031);
not_8  g20520(new_n21083, new_n22869);
nor_5  g20521(new_n22705, new_n7955, new_n22870_1);
not_8  g20522(new_n22870_1, new_n22871_1);
nor_5  g20523(new_n18401, n22626, new_n22872);
nor_5  g20524(new_n18418_1, new_n22872, new_n22873);
nor_5  g20525(new_n22873, new_n22716, new_n22874);
nand_5 g20526(new_n22874, new_n22871_1, new_n22875);
nor_5  g20527(new_n22875, new_n22869, new_n22876);
xnor_4 g20528(new_n22875, new_n21083, new_n22877);
not_8  g20529(new_n22877, new_n22878);
nor_5  g20530(new_n18419, new_n18398, new_n22879_1);
not_8  g20531(new_n18420, new_n22880);
nor_5  g20532(new_n18452_1, new_n22880, new_n22881);
nor_5  g20533(new_n22881, new_n22879_1, new_n22882);
nor_5  g20534(new_n22882, new_n22878, new_n22883);
nor_5  g20535(new_n22883, new_n22876, new_n22884);
not_8  g20536(new_n22884, new_n22885);
nor_5  g20537(new_n18461, n9554, new_n22886);
nor_5  g20538(new_n18494, new_n22886, new_n22887);
nor_5  g20539(new_n21358, new_n8278, new_n22888);
nor_5  g20540(new_n22888, new_n21406, new_n22889);
not_8  g20541(new_n22889, new_n22890);
nor_5  g20542(new_n22890, new_n22887, new_n22891_1);
nor_5  g20543(new_n22891_1, new_n22885, new_n22892);
xnor_4 g20544(new_n22891_1, new_n22884, new_n22893);
not_8  g20545(new_n22893, new_n22894);
not_8  g20546(new_n22891_1, new_n22895);
xnor_4 g20547(new_n22882, new_n22878, new_n22896);
not_8  g20548(new_n22896, new_n22897_1);
nor_5  g20549(new_n22897_1, new_n22895, new_n22898);
xnor_4 g20550(new_n22896, new_n22891_1, new_n22899);
nor_5  g20551(new_n18495, new_n18453, new_n22900);
nor_5  g20552(new_n18553, new_n18496_1, new_n22901);
nor_5  g20553(new_n22901, new_n22900, new_n22902);
nor_5  g20554(new_n22902, new_n22899, new_n22903_1);
nor_5  g20555(new_n22903_1, new_n22898, new_n22904);
nor_5  g20556(new_n22904, new_n22894, new_n22905);
nor_5  g20557(new_n22905, new_n22892, n8042);
not_8  g20558(new_n10510, new_n22907_1);
nand_5 g20559(new_n10614_1, new_n22907_1, new_n22908);
nand_5 g20560(new_n10696, new_n10615, new_n22909);
nand_5 g20561(new_n22909, new_n22908, n8095);
nor_5  g20562(new_n18454, n4306, new_n22911);
xnor_4 g20563(n23166, n4306, new_n22912);
not_8  g20564(new_n22912, new_n22913);
nor_5  g20565(new_n9672, n3279, new_n22914_1);
xnor_4 g20566(n10577, n3279, new_n22915);
not_8  g20567(new_n22915, new_n22916);
nor_5  g20568(n13914, new_n9675, new_n22917);
xnor_4 g20569(n13914, n6381, new_n22918_1);
not_8  g20570(new_n22918_1, new_n22919);
nor_5  g20571(n14702, new_n9678, new_n22920);
nor_5  g20572(new_n20800, new_n20787, new_n22921);
nor_5  g20573(new_n22921, new_n22920, new_n22922);
nor_5  g20574(new_n22922, new_n22919, new_n22923);
nor_5  g20575(new_n22923, new_n22917, new_n22924);
nor_5  g20576(new_n22924, new_n22916, new_n22925);
nor_5  g20577(new_n22925, new_n22914_1, new_n22926);
nor_5  g20578(new_n22926, new_n22913, new_n22927);
nor_5  g20579(new_n22927, new_n22911, new_n22928);
xnor_4 g20580(new_n22928, new_n9529, new_n22929);
xnor_4 g20581(new_n22926, new_n22913, new_n22930);
nand_5 g20582(new_n22930, new_n9582, new_n22931);
xnor_4 g20583(new_n22930, new_n9581, new_n22932);
xnor_4 g20584(new_n22924, new_n22916, new_n22933);
nand_5 g20585(new_n22933, new_n9587, new_n22934);
xnor_4 g20586(new_n22933, new_n9586, new_n22935);
xnor_4 g20587(new_n22922, new_n22918_1, new_n22936);
not_8  g20588(new_n22936, new_n22937);
nand_5 g20589(new_n22937, new_n9591, new_n22938);
xnor_4 g20590(new_n22936, new_n9591, new_n22939_1);
nor_5  g20591(new_n20801, new_n9596, new_n22940);
nor_5  g20592(new_n20818, new_n20802, new_n22941);
nor_5  g20593(new_n22941, new_n22940, new_n22942);
nand_5 g20594(new_n22942, new_n22939_1, new_n22943);
nand_5 g20595(new_n22943, new_n22938, new_n22944);
nand_5 g20596(new_n22944, new_n22935, new_n22945);
nand_5 g20597(new_n22945, new_n22934, new_n22946);
nand_5 g20598(new_n22946, new_n22932, new_n22947);
nand_5 g20599(new_n22947, new_n22931, new_n22948);
xnor_4 g20600(new_n22948, new_n22929, n8103);
xnor_4 g20601(new_n20095, new_n20081, n8109);
not_8  g20602(new_n20592, new_n22951);
nand_5 g20603(new_n22951, new_n20574, new_n22952);
nand_5 g20604(new_n20632, new_n20593, new_n22953);
nand_5 g20605(new_n22953, new_n22952, n8127);
xnor_4 g20606(new_n17886, new_n17883, n8130);
or_5   g20607(n8856, new_n3164_1, new_n22956);
xnor_4 g20608(n8856, n4319, new_n22957);
or_5   g20609(new_n12485, n14130, new_n22958);
xnor_4 g20610(n23463, n14130, new_n22959);
or_5   g20611(n16482, new_n3171, new_n22960);
xnor_4 g20612(n16482, n13074, new_n22961);
or_5   g20613(new_n11911, n9942, new_n22962);
nand_5 g20614(new_n2380, new_n2349, new_n22963);
nand_5 g20615(new_n22963, new_n22962, new_n22964);
nand_5 g20616(new_n22964, new_n22961, new_n22965);
nand_5 g20617(new_n22965, new_n22960, new_n22966);
nand_5 g20618(new_n22966, new_n22959, new_n22967);
nand_5 g20619(new_n22967, new_n22958, new_n22968);
nand_5 g20620(new_n22968, new_n22957, new_n22969);
nand_5 g20621(new_n22969, new_n22956, new_n22970);
not_8  g20622(new_n22970, new_n22971);
xnor_4 g20623(new_n22971, new_n8020, new_n22972);
nand_5 g20624(new_n22970, new_n8023, new_n22973);
xnor_4 g20625(new_n22971, new_n8023, new_n22974);
xnor_4 g20626(new_n22968, new_n22957, new_n22975);
nand_5 g20627(new_n22975, new_n8028, new_n22976);
xnor_4 g20628(new_n22975, new_n8027_1, new_n22977);
xnor_4 g20629(new_n22966, new_n22959, new_n22978);
nand_5 g20630(new_n22978, new_n8033, new_n22979);
xnor_4 g20631(new_n22978, new_n8032, new_n22980);
xnor_4 g20632(new_n22964, new_n22961, new_n22981);
nor_5  g20633(new_n22981, new_n8038, new_n22982);
xnor_4 g20634(new_n22981, new_n8038, new_n22983);
nor_5  g20635(new_n2518, new_n2381, new_n22984);
nor_5  g20636(new_n2566, new_n2519, new_n22985);
nor_5  g20637(new_n22985, new_n22984, new_n22986);
nor_5  g20638(new_n22986, new_n22983, new_n22987);
nor_5  g20639(new_n22987, new_n22982, new_n22988);
nand_5 g20640(new_n22988, new_n22980, new_n22989);
nand_5 g20641(new_n22989, new_n22979, new_n22990);
nand_5 g20642(new_n22990, new_n22977, new_n22991);
nand_5 g20643(new_n22991, new_n22976, new_n22992);
nand_5 g20644(new_n22992, new_n22974, new_n22993);
nand_5 g20645(new_n22993, new_n22973, new_n22994);
xnor_4 g20646(new_n22994, new_n22972, n8135);
xnor_4 g20647(new_n8071, new_n2555_1, n8139);
nand_5 g20648(new_n19417, new_n11311, new_n22997);
nor_5  g20649(new_n22997, n26660, new_n22998_1);
xnor_4 g20650(new_n22998_1, n13783, new_n22999);
xnor_4 g20651(new_n22999, new_n3042, new_n23000);
xnor_4 g20652(new_n22997, new_n8101, new_n23001);
nand_5 g20653(new_n23001, new_n3050, new_n23002);
xnor_4 g20654(new_n23001, new_n3049, new_n23003);
nand_5 g20655(new_n19418, new_n3057, new_n23004);
nand_5 g20656(new_n19436, new_n19419, new_n23005);
nand_5 g20657(new_n23005, new_n23004, new_n23006_1);
nand_5 g20658(new_n23006_1, new_n23003, new_n23007_1);
nand_5 g20659(new_n23007_1, new_n23002, new_n23008);
xnor_4 g20660(new_n23008, new_n23000, new_n23009_1);
xnor_4 g20661(new_n23009_1, new_n7303, new_n23010);
xnor_4 g20662(new_n23006_1, new_n23003, new_n23011);
nand_5 g20663(new_n23011, new_n7310, new_n23012);
xnor_4 g20664(new_n23011, new_n7308_1, new_n23013);
nand_5 g20665(new_n19437, new_n7313_1, new_n23014_1);
nand_5 g20666(new_n19461, new_n19438, new_n23015);
nand_5 g20667(new_n23015, new_n23014_1, new_n23016);
nand_5 g20668(new_n23016, new_n23013, new_n23017);
nand_5 g20669(new_n23017, new_n23012, new_n23018);
xnor_4 g20670(new_n23018, new_n23010, n8148);
xor_4  g20671(new_n18770, new_n18769, n8149);
xnor_4 g20672(new_n4087, new_n4069, n8159);
xnor_4 g20673(new_n12431, new_n2582_1, n8179);
xnor_4 g20674(new_n15846_1, new_n15843, n8215);
xnor_4 g20675(new_n20093, new_n20083, n8267);
xnor_4 g20676(new_n21273, new_n21271, n8276);
nand_5 g20677(new_n22998_1, new_n2422, new_n23026);
nor_5  g20678(new_n23026, n1654, new_n23027);
and_5  g20679(new_n23027, new_n7946, new_n23028);
xnor_4 g20680(new_n23028, n22626, new_n23029);
not_8  g20681(new_n23029, new_n23030);
nand_5 g20682(new_n23030, new_n16026, new_n23031);
not_8  g20683(new_n23031, new_n23032);
xnor_4 g20684(new_n23030, new_n16026, new_n23033);
xnor_4 g20685(new_n23027, n14440, new_n23034);
nor_5  g20686(new_n23034, new_n3031, new_n23035_1);
xnor_4 g20687(new_n23034, new_n3031, new_n23036);
xnor_4 g20688(new_n23026, new_n7935, new_n23037);
nand_5 g20689(new_n23037, new_n3037, new_n23038);
nand_5 g20690(new_n22999, new_n3043, new_n23039_1);
nand_5 g20691(new_n23008, new_n23000, new_n23040);
nand_5 g20692(new_n23040, new_n23039_1, new_n23041);
xnor_4 g20693(new_n23037, new_n3035, new_n23042);
nand_5 g20694(new_n23042, new_n23041, new_n23043);
nand_5 g20695(new_n23043, new_n23038, new_n23044);
nor_5  g20696(new_n23044, new_n23036, new_n23045);
nor_5  g20697(new_n23045, new_n23035_1, new_n23046);
nor_5  g20698(new_n23046, new_n23033, new_n23047_1);
nor_5  g20699(new_n23047_1, new_n23032, new_n23048);
and_5  g20700(new_n23028, new_n7955, new_n23049);
xnor_4 g20701(new_n23049, new_n16054, new_n23050);
xnor_4 g20702(new_n23050, new_n23048, new_n23051);
nand_5 g20703(new_n23051, new_n18302, new_n23052);
xnor_4 g20704(new_n23051, new_n18301_1, new_n23053);
not_8  g20705(new_n23033, new_n23054);
xnor_4 g20706(new_n23046, new_n23054, new_n23055);
nand_5 g20707(new_n23055, new_n18309, new_n23056);
xnor_4 g20708(new_n23055, new_n18308, new_n23057);
not_8  g20709(new_n23036, new_n23058_1);
xnor_4 g20710(new_n23044, new_n23058_1, new_n23059);
nand_5 g20711(new_n23059, new_n7216, new_n23060);
xnor_4 g20712(new_n23042, new_n23041, new_n23061);
nand_5 g20713(new_n23061, new_n7300, new_n23062);
xnor_4 g20714(new_n23061, new_n7298_1, new_n23063);
nand_5 g20715(new_n23009_1, new_n7305_1, new_n23064);
nand_5 g20716(new_n23018, new_n23010, new_n23065_1);
nand_5 g20717(new_n23065_1, new_n23064, new_n23066_1);
nand_5 g20718(new_n23066_1, new_n23063, new_n23067_1);
nand_5 g20719(new_n23067_1, new_n23062, new_n23068_1);
xnor_4 g20720(new_n23059, new_n7215, new_n23069);
nand_5 g20721(new_n23069, new_n23068_1, new_n23070);
nand_5 g20722(new_n23070, new_n23060, new_n23071);
nand_5 g20723(new_n23071, new_n23057, new_n23072);
nand_5 g20724(new_n23072, new_n23056, new_n23073);
nand_5 g20725(new_n23073, new_n23053, new_n23074);
nand_5 g20726(new_n23074, new_n23052, new_n23075);
nor_5  g20727(new_n23075, new_n18241_1, new_n23076);
not_8  g20728(new_n23048, new_n23077);
nor_5  g20729(new_n23049, new_n16054, new_n23078);
and_5  g20730(new_n23078, new_n23077, new_n23079);
nand_5 g20731(new_n23075, new_n18241_1, new_n23080);
nand_5 g20732(new_n23049, new_n16054, new_n23081);
nor_5  g20733(new_n23081, new_n23077, new_n23082);
nor_5  g20734(new_n23082, new_n23080, new_n23083);
nor_5  g20735(new_n23083, new_n23079, new_n23084);
nor_5  g20736(new_n23084, new_n23076, n8288);
xnor_4 g20737(new_n11971, new_n7855, n8306);
xor_4  g20738(new_n8408_1, new_n8351, n8320);
xnor_4 g20739(new_n13280, new_n13258, n8321);
xnor_4 g20740(new_n17445, new_n17428, n8339);
xnor_4 g20741(new_n9648_1, new_n9594, n8376);
xor_4  g20742(new_n20440, new_n10865, n8408);
not_8  g20743(new_n15354, new_n23092);
xnor_4 g20744(new_n23092, new_n15353_1, n8417);
xnor_4 g20745(new_n13741, new_n13722_1, n8432);
nor_5  g20746(new_n16776, new_n10757, new_n23095);
nor_5  g20747(new_n10819, new_n10762, new_n23096);
nor_5  g20748(new_n23096, new_n23095, new_n23097);
not_8  g20749(new_n23097, new_n23098);
nand_5 g20750(new_n23098, new_n10739_1, new_n23099);
nand_5 g20751(new_n10820, new_n10738, new_n23100);
nand_5 g20752(new_n10894, new_n10821, new_n23101);
nand_5 g20753(new_n23101, new_n23100, new_n23102);
nand_5 g20754(new_n23102, new_n23099, new_n23103);
nand_5 g20755(new_n23097, new_n10738, new_n23104);
nand_5 g20756(new_n23104, new_n23101, new_n23105);
nand_5 g20757(new_n23105, new_n23103, new_n23106);
not_8  g20758(new_n23106, n8453);
xnor_4 g20759(new_n16633, new_n14601, n8480);
xnor_4 g20760(new_n17614, new_n17593, n8489);
xnor_4 g20761(new_n22990, new_n22977, n8505);
xnor_4 g20762(new_n20920, new_n20904, n8510);
xnor_4 g20763(new_n12943, new_n9179, n8519);
xnor_4 g20764(new_n10358, new_n10356_1, n8535);
xnor_4 g20765(new_n20624, new_n20620, n8550);
xnor_4 g20766(new_n21914, new_n21906, n8563);
xnor_4 g20767(new_n14212, new_n14210, n8594);
xnor_4 g20768(new_n7345, new_n7324, n8608);
not_8  g20769(new_n4795, new_n23118);
xnor_4 g20770(new_n23118, new_n4794, n8620);
xnor_4 g20771(new_n7880, new_n7819, n8637);
xnor_4 g20772(new_n18321, new_n18320, n8662);
xnor_4 g20773(new_n20152, new_n20139, n8716);
xnor_4 g20774(new_n8355, new_n8352, new_n23123);
xnor_4 g20775(new_n23123, new_n8406, n8744);
nand_5 g20776(new_n13693, n9554, new_n23125);
nand_5 g20777(new_n22763, new_n22755, new_n23126);
nand_5 g20778(new_n23126, new_n23125, new_n23127);
xnor_4 g20779(new_n23127, new_n16361, new_n23128);
nand_5 g20780(new_n6355, n3740, new_n23129);
nand_5 g20781(new_n22676, new_n22673, new_n23130);
nand_5 g20782(new_n23130, new_n23129, new_n23131);
xnor_4 g20783(new_n23131, new_n19008, new_n23132);
not_8  g20784(new_n23132, new_n23133);
xnor_4 g20785(new_n23133, new_n23128, new_n23134);
nand_5 g20786(new_n22764_1, new_n22677, new_n23135);
not_8  g20787(new_n22677, new_n23136);
xnor_4 g20788(new_n22764_1, new_n23136, new_n23137);
nor_5  g20789(new_n22767, new_n17231, new_n23138);
xnor_4 g20790(new_n22767, new_n17231, new_n23139);
nand_5 g20791(new_n18570, new_n17233, new_n23140);
nand_5 g20792(new_n18605, new_n18571, new_n23141);
nand_5 g20793(new_n23141, new_n23140, new_n23142);
nor_5  g20794(new_n23142, new_n23139, new_n23143);
nor_5  g20795(new_n23143, new_n23138, new_n23144);
nand_5 g20796(new_n23144, new_n23137, new_n23145);
nand_5 g20797(new_n23145, new_n23135, new_n23146_1);
xnor_4 g20798(new_n23146_1, new_n23134, n8803);
nor_5  g20799(new_n21747, n13494, new_n23148);
not_8  g20800(new_n21748, new_n23149);
nand_5 g20801(new_n23149, n12650, new_n23150);
nand_5 g20802(new_n21771, new_n21749_1, new_n23151);
nand_5 g20803(new_n23151, new_n23150, new_n23152);
not_8  g20804(new_n23152, new_n23153);
xnor_4 g20805(new_n23153, new_n23148, new_n23154);
or_5   g20806(n16544, n4319, new_n23155);
not_8  g20807(new_n16881, new_n23156);
nand_5 g20808(new_n23156, new_n16857, new_n23157);
nand_5 g20809(new_n23157, new_n23155, new_n23158);
not_8  g20810(new_n23158, new_n23159);
xnor_4 g20811(new_n23159, new_n23154, new_n23160_1);
not_8  g20812(new_n16882, new_n23161);
nand_5 g20813(new_n21772, new_n23161, new_n23162);
nand_5 g20814(new_n21791, new_n21773, new_n23163);
nand_5 g20815(new_n23163, new_n23162, new_n23164);
xnor_4 g20816(new_n23164, new_n23160_1, new_n23165);
xnor_4 g20817(new_n23165, new_n12479, new_n23166_1);
nand_5 g20818(new_n21792, new_n8190, new_n23167);
nand_5 g20819(new_n22421, new_n22383, new_n23168);
nand_5 g20820(new_n23168, new_n23167, new_n23169);
xnor_4 g20821(new_n23169, new_n23166_1, n8809);
nand_5 g20822(new_n23131, new_n19009, new_n23171);
not_8  g20823(new_n23171, new_n23172);
nor_5  g20824(new_n19377, n3324, new_n23173);
not_8  g20825(new_n23173, new_n23174);
nand_5 g20826(new_n22671, new_n22656, new_n23175);
nand_5 g20827(new_n23175, new_n23174, new_n23176);
nor_5  g20828(new_n23176, new_n19372, new_n23177);
xnor_4 g20829(new_n23177, new_n23172, new_n23178);
xnor_4 g20830(new_n23176, new_n19372, new_n23179);
nand_5 g20831(new_n23179, new_n23132, new_n23180);
xnor_4 g20832(new_n23179, new_n23133, new_n23181);
nand_5 g20833(new_n23136, new_n22672, new_n23182);
nand_5 g20834(new_n22692, new_n22678, new_n23183);
nand_5 g20835(new_n23183, new_n23182, new_n23184);
nand_5 g20836(new_n23184, new_n23181, new_n23185);
nand_5 g20837(new_n23185, new_n23180, new_n23186);
xnor_4 g20838(new_n23186, new_n23178, n8821);
xnor_4 g20839(new_n16602, new_n16601, n8824);
xor_4  g20840(new_n18953, new_n18952, n8849);
xnor_4 g20841(new_n14733, new_n14725, n8861);
xnor_4 g20842(n22442, n8856, new_n23191);
nor_5  g20843(n14130, new_n7404, new_n23192);
nor_5  g20844(new_n21525_1, new_n21498, new_n23193);
nor_5  g20845(new_n23193, new_n23192, new_n23194);
xnor_4 g20846(new_n23194, new_n23191, new_n23195);
xnor_4 g20847(n3324, new_n7613, new_n23196);
not_8  g20848(new_n23196, new_n23197);
or_5   g20849(n25331, n17911, new_n23198);
nand_5 g20850(new_n21486, new_n21482, new_n23199);
nand_5 g20851(new_n23199, new_n23198, new_n23200_1);
xnor_4 g20852(new_n23200_1, new_n23197, new_n23201);
xnor_4 g20853(new_n23201, new_n7961, new_n23202);
not_8  g20854(new_n7952, new_n23203);
nor_5  g20855(new_n21487, new_n23203, new_n23204);
not_8  g20856(new_n23204, new_n23205);
nand_5 g20857(new_n21495, new_n21488, new_n23206);
nand_5 g20858(new_n23206, new_n23205, new_n23207);
xnor_4 g20859(new_n23207, new_n23202, new_n23208);
not_8  g20860(new_n23208, new_n23209);
xnor_4 g20861(new_n23209, new_n23195, new_n23210);
not_8  g20862(new_n21496, new_n23211);
nor_5  g20863(new_n21526, new_n23211, new_n23212);
not_8  g20864(new_n23212, new_n23213);
nand_5 g20865(new_n21559, new_n23213, new_n23214);
xnor_4 g20866(new_n23214, new_n23210, n8862);
xor_4  g20867(new_n14608, new_n14607, n8884);
xor_4  g20868(new_n20340, new_n19467_1, n8909);
xnor_4 g20869(new_n12450, new_n12405, n8911);
xnor_4 g20870(new_n11904, new_n11902, n8971);
xnor_4 g20871(new_n22862, new_n22833, n8982);
xnor_4 g20872(new_n5722, new_n5702, n8993);
xor_4  g20873(new_n15363, new_n15362, n9012);
nand_5 g20874(new_n21664, new_n21660, new_n23223);
not_8  g20875(new_n21668, new_n23224);
not_8  g20876(new_n21669, new_n23225);
nand_5 g20877(new_n23225, new_n4645, new_n23226);
nor_5  g20878(new_n23226, new_n23224, new_n23227);
xnor_4 g20879(new_n23227, new_n23223, new_n23228);
not_8  g20880(new_n21665_1, new_n23229);
nand_5 g20881(new_n21671, new_n23229, new_n23230);
nand_5 g20882(new_n21724, new_n21672, new_n23231);
nand_5 g20883(new_n23231, new_n23230, new_n23232);
xnor_4 g20884(new_n23232, new_n23228, n9032);
xnor_4 g20885(new_n17155, new_n17154, n9042);
xnor_4 g20886(new_n18547, new_n18516, n9046);
xnor_4 g20887(new_n8711, new_n8646, n9047);
xnor_4 g20888(new_n16298, new_n16297, n9104);
nand_5 g20889(new_n22079, new_n22067, new_n23238_1);
nand_5 g20890(new_n23238_1, new_n16453, new_n23239);
not_8  g20891(new_n23239, new_n23240);
nor_5  g20892(new_n22079, new_n22067, new_n23241);
nor_5  g20893(new_n23241, new_n16453, new_n23242);
nor_5  g20894(new_n23242, new_n23240, new_n23243);
xnor_4 g20895(new_n23243, new_n20860, new_n23244);
not_8  g20896(new_n22081, new_n23245);
nand_5 g20897(new_n23245, new_n20860, new_n23246);
nand_5 g20898(new_n22090_1, new_n22082, new_n23247_1);
nand_5 g20899(new_n23247_1, new_n23246, new_n23248_1);
xnor_4 g20900(new_n23248_1, new_n23244, n9129);
xnor_4 g20901(new_n20552, new_n20509, n9146);
xnor_4 g20902(new_n9179, new_n7069, n9164);
xnor_4 g20903(new_n13654, new_n13653, n9166);
xnor_4 g20904(new_n19393, new_n19363, new_n23253);
xnor_4 g20905(new_n23253, new_n19407, n9182);
xnor_4 g20906(new_n7602, new_n7565, n9191);
xnor_4 g20907(new_n12456, new_n12396, n9217);
xor_4  g20908(new_n17332, new_n17331, n9220);
xnor_4 g20909(new_n20541, new_n20534, n9261);
xnor_4 g20910(n22626, n3324, new_n23259);
not_8  g20911(new_n23259, new_n23260);
nor_5  g20912(new_n16884, n14440, new_n23261);
nor_5  g20913(new_n20124, new_n20100, new_n23262);
nor_5  g20914(new_n23262, new_n23261, new_n23263);
xnor_4 g20915(new_n23263, new_n23260, new_n23264);
nor_5  g20916(new_n23264, new_n19399, new_n23265);
not_8  g20917(new_n23265, new_n23266);
xnor_4 g20918(new_n23264, new_n19398, new_n23267);
nor_5  g20919(new_n20125, new_n19402, new_n23268);
not_8  g20920(new_n23268, new_n23269);
nand_5 g20921(new_n20159, new_n20126_1, new_n23270_1);
nand_5 g20922(new_n23270_1, new_n23269, new_n23271);
nand_5 g20923(new_n23271, new_n23267, new_n23272_1);
nand_5 g20924(new_n23272_1, new_n23266, new_n23273);
nor_5  g20925(n22626, new_n16856, new_n23274);
nor_5  g20926(new_n23263, new_n23260, new_n23275);
nor_5  g20927(new_n23275, new_n23274, new_n23276);
xnor_4 g20928(new_n23276, new_n19393, new_n23277);
xnor_4 g20929(new_n23277, new_n23273, n9287);
xor_4  g20930(new_n15179, new_n15166, n9308);
xnor_4 g20931(new_n5286, new_n5240, n9344);
xnor_4 g20932(new_n3863, new_n3845, n9364);
not_8  g20933(new_n23273, new_n23282);
nor_5  g20934(new_n23276, new_n19394, new_n23283);
not_8  g20935(new_n23283, new_n23284);
nor_5  g20936(new_n23284, new_n23282, new_n23285);
nand_5 g20937(new_n23285, new_n19390, new_n23286);
not_8  g20938(new_n23276, new_n23287);
nor_5  g20939(new_n23287, new_n19393, new_n23288);
not_8  g20940(new_n23288, new_n23289_1);
nor_5  g20941(new_n23289_1, new_n23273, new_n23290);
nand_5 g20942(new_n23290, new_n19391, new_n23291);
nand_5 g20943(new_n23291, new_n23286, n9371);
xor_4  g20944(new_n10866, new_n10865, n9382);
xnor_4 g20945(new_n22904, new_n22893, n9403);
xnor_4 g20946(new_n13661, new_n13633, n9419);
xnor_4 g20947(new_n22635, new_n22607, n9423);
xnor_4 g20948(new_n20154, new_n20134, n9430);
xnor_4 g20949(n25120, n23272, new_n23298);
not_8  g20950(new_n23298, new_n23299);
and_5  g20951(new_n4552_1, n8363, new_n23300);
xnor_4 g20952(n11481, n8363, new_n23301);
not_8  g20953(new_n23301, new_n23302);
nor_5  g20954(n16439, new_n14989_1, new_n23303);
nor_5  g20955(new_n16796, new_n16793, new_n23304_1);
nor_5  g20956(new_n23304_1, new_n23303, new_n23305_1);
nor_5  g20957(new_n23305_1, new_n23302, new_n23306);
nor_5  g20958(new_n23306, new_n23300, new_n23307);
xnor_4 g20959(new_n23307, new_n23299, new_n23308);
xnor_4 g20960(new_n23308, new_n18419, new_n23309);
xnor_4 g20961(new_n23305_1, new_n23302, new_n23310);
not_8  g20962(new_n23310, new_n23311);
nand_5 g20963(new_n23311, new_n18422, new_n23312);
xnor_4 g20964(new_n23310, new_n18422, new_n23313);
nor_5  g20965(new_n16803, new_n16797, new_n23314);
nor_5  g20966(new_n16807, new_n16804, new_n23315);
nor_5  g20967(new_n23315, new_n23314, new_n23316);
not_8  g20968(new_n23316, new_n23317);
nand_5 g20969(new_n23317, new_n23313, new_n23318);
nand_5 g20970(new_n23318, new_n23312, new_n23319);
xnor_4 g20971(new_n23319, new_n23309, new_n23320);
xnor_4 g20972(new_n23320, new_n18495, new_n23321);
not_8  g20973(new_n23321, new_n23322);
xnor_4 g20974(new_n23316, new_n23313, new_n23323);
not_8  g20975(new_n23323, new_n23324);
nand_5 g20976(new_n23324, new_n18499, new_n23325);
xnor_4 g20977(new_n23323, new_n18499, new_n23326);
nand_5 g20978(new_n18505, new_n16808, new_n23327);
xnor_4 g20979(new_n18490, new_n18469, new_n23328);
xnor_4 g20980(new_n23328, new_n16808, new_n23329);
nand_5 g20981(new_n18512, new_n11362, new_n23330);
xnor_4 g20982(new_n18488, new_n18472, new_n23331);
xnor_4 g20983(new_n23331, new_n11362, new_n23332);
nor_5  g20984(new_n18519, new_n11365, new_n23333_1);
not_8  g20985(new_n23333_1, new_n23334);
xnor_4 g20986(new_n18520, new_n11365, new_n23335);
nor_5  g20987(new_n18524, new_n11370, new_n23336);
not_8  g20988(new_n11372, new_n23337);
not_8  g20989(new_n16003, new_n23338);
nor_5  g20990(new_n23338, new_n23337, new_n23339);
nor_5  g20991(new_n16019, new_n16004, new_n23340);
nor_5  g20992(new_n23340, new_n23339, new_n23341_1);
xnor_4 g20993(new_n18524, new_n11370, new_n23342_1);
nor_5  g20994(new_n23342_1, new_n23341_1, new_n23343);
nor_5  g20995(new_n23343, new_n23336, new_n23344);
nand_5 g20996(new_n23344, new_n23335, new_n23345);
nand_5 g20997(new_n23345, new_n23334, new_n23346);
nand_5 g20998(new_n23346, new_n23332, new_n23347);
nand_5 g20999(new_n23347, new_n23330, new_n23348);
nand_5 g21000(new_n23348, new_n23329, new_n23349);
nand_5 g21001(new_n23349, new_n23327, new_n23350);
nand_5 g21002(new_n23350, new_n23326, new_n23351);
nand_5 g21003(new_n23351, new_n23325, new_n23352);
xnor_4 g21004(new_n23352, new_n23322, n9435);
xnor_4 g21005(new_n17275, new_n17241, n9451);
xnor_4 g21006(n12657, n10763, new_n23355_1);
not_8  g21007(new_n23355_1, new_n23356);
or_5   g21008(n17077, new_n2944_1, new_n23357);
nand_5 g21009(new_n20688, new_n20679, new_n23358);
nand_5 g21010(new_n23358, new_n23357, new_n23359);
xnor_4 g21011(new_n23359, new_n23356, new_n23360);
xnor_4 g21012(new_n23360, new_n21496, new_n23361);
nor_5  g21013(new_n20715, new_n20689, new_n23362);
nor_5  g21014(new_n20727, new_n20716, new_n23363);
nor_5  g21015(new_n23363, new_n23362, new_n23364);
xnor_4 g21016(new_n23364, new_n23361, n9458);
nor_5  g21017(n12507, new_n10741, new_n23366);
xnor_4 g21018(n12507, n11220, new_n23367);
not_8  g21019(new_n23367, new_n23368);
nor_5  g21020(new_n19358, n15077, new_n23369_1);
not_8  g21021(new_n15915, new_n23370);
nor_5  g21022(new_n15939, new_n23370, new_n23371_1);
nor_5  g21023(new_n23371_1, new_n23369_1, new_n23372);
nor_5  g21024(new_n23372, new_n23368, new_n23373);
nor_5  g21025(new_n23373, new_n23366, new_n23374);
xnor_4 g21026(new_n23374, new_n22277, new_n23375);
xnor_4 g21027(new_n23372, new_n23368, new_n23376);
nand_5 g21028(new_n23376, new_n22280, new_n23377);
xnor_4 g21029(new_n23376, new_n22279, new_n23378);
not_8  g21030(new_n15940, new_n23379);
nand_5 g21031(new_n23379, new_n15914, new_n23380);
nand_5 g21032(new_n15973, new_n15941, new_n23381);
nand_5 g21033(new_n23381, new_n23380, new_n23382);
nand_5 g21034(new_n23382, new_n23378, new_n23383);
nand_5 g21035(new_n23383, new_n23377, new_n23384);
xnor_4 g21036(new_n23384, new_n23375, n9459);
xnor_4 g21037(new_n16232, new_n16231, n9508);
xnor_4 g21038(new_n13665, new_n13621, n9552);
xnor_4 g21039(new_n4798, new_n4797, n9556);
xnor_4 g21040(new_n11875, new_n9388, n9558);
xnor_4 g21041(new_n22491, new_n23092, n9616);
xnor_4 g21042(new_n9103, new_n9074, n9622);
xnor_4 g21043(new_n17816, new_n17798, n9626);
xnor_4 g21044(new_n4803, new_n4783, n9633);
and_5  g21045(n25120, new_n4548, new_n23394);
nor_5  g21046(new_n23307, new_n23299, new_n23395);
nor_5  g21047(new_n23395, new_n23394, new_n23396);
not_8  g21048(new_n23396, new_n23397);
nor_5  g21049(new_n23397, new_n22875, new_n23398);
xnor_4 g21050(new_n23397, new_n22875, new_n23399);
not_8  g21051(new_n23308, new_n23400);
nand_5 g21052(new_n23400, new_n18419, new_n23401_1);
nand_5 g21053(new_n23319, new_n23309, new_n23402);
nand_5 g21054(new_n23402, new_n23401_1, new_n23403);
nor_5  g21055(new_n23403, new_n23399, new_n23404);
nor_5  g21056(new_n23404, new_n23398, new_n23405);
not_8  g21057(new_n23405, new_n23406);
nor_5  g21058(new_n23406, new_n5833_1, new_n23407);
xnor_4 g21059(new_n23405, new_n5833_1, new_n23408);
not_8  g21060(new_n23408, new_n23409);
xnor_4 g21061(new_n23403, new_n23399, new_n23410);
not_8  g21062(new_n23410, new_n23411);
nor_5  g21063(new_n23411, new_n5832, new_n23412);
xnor_4 g21064(new_n23410, new_n5832, new_n23413);
not_8  g21065(new_n23413, new_n23414_1);
nand_5 g21066(new_n23320, new_n5834_1, new_n23415);
nor_5  g21067(new_n23324, new_n5914, new_n23416);
xnor_4 g21068(new_n23324, new_n5914, new_n23417);
nor_5  g21069(new_n16808, new_n5919, new_n23418);
nor_5  g21070(new_n16812_1, new_n16809, new_n23419);
nor_5  g21071(new_n23419, new_n23418, new_n23420);
nor_5  g21072(new_n23420, new_n23417, new_n23421);
nor_5  g21073(new_n23421, new_n23416, new_n23422);
xnor_4 g21074(new_n23320, new_n5834_1, new_n23423);
not_8  g21075(new_n23423, new_n23424);
nand_5 g21076(new_n23424, new_n23422, new_n23425);
nand_5 g21077(new_n23425, new_n23415, new_n23426);
nor_5  g21078(new_n23426, new_n23414_1, new_n23427);
nor_5  g21079(new_n23427, new_n23412, new_n23428);
nor_5  g21080(new_n23428, new_n23409, new_n23429_1);
nor_5  g21081(new_n23429_1, new_n23407, n9635);
xnor_4 g21082(new_n20948, new_n20944, n9648);
xnor_4 g21083(new_n5266, new_n5265_1, n9689);
xnor_4 g21084(new_n11560, new_n11538_1, n9695);
xnor_4 g21085(new_n8085, new_n8035, n9699);
xnor_4 g21086(new_n17901, new_n17281, new_n23435);
nand_5 g21087(new_n17294, new_n15744, new_n23436);
nand_5 g21088(new_n17338, new_n17295, new_n23437);
nand_5 g21089(new_n23437, new_n23436, new_n23438);
xnor_4 g21090(new_n23438, new_n23435, n9726);
xnor_4 g21091(new_n14227, new_n10670, n9753);
xnor_4 g21092(new_n3505, new_n3480_1, n9761);
xnor_4 g21093(new_n10688, new_n10635, n9763);
xnor_4 g21094(new_n14605, new_n14604, n9767);
xnor_4 g21095(new_n14785, new_n14491, n9771);
xor_4  g21096(new_n22986, new_n22983, n9778);
xnor_4 g21097(new_n17046, new_n17035_1, n9783);
xnor_4 g21098(new_n7104, new_n7100, n9803);
nand_5 g21099(new_n22427, new_n12485, new_n23448);
nor_5  g21100(new_n23448, n4319, new_n23449);
not_8  g21101(new_n23449, new_n23450_1);
not_8  g21102(new_n19333_1, new_n23451);
xnor_4 g21103(new_n23448, new_n3164_1, new_n23452);
nand_5 g21104(new_n23452, new_n23451, new_n23453);
not_8  g21105(new_n23452, new_n23454);
nand_5 g21106(new_n23454, new_n19333_1, new_n23455);
nand_5 g21107(new_n22428, new_n19339, new_n23456);
not_8  g21108(new_n22428, new_n23457);
nand_5 g21109(new_n23457, new_n19338, new_n23458);
not_8  g21110(new_n17968_1, new_n23459);
nand_5 g21111(new_n22430, new_n23459, new_n23460);
not_8  g21112(new_n22430, new_n23461);
nand_5 g21113(new_n23461, new_n17968_1, new_n23462);
nor_5  g21114(new_n22433_1, new_n17979, new_n23463_1);
not_8  g21115(new_n17983, new_n23464);
nand_5 g21116(new_n22436, new_n23464, new_n23465);
xnor_4 g21117(new_n22436, new_n17983, new_n23466);
nand_5 g21118(new_n9110, new_n7039, new_n23467);
nand_5 g21119(new_n7085, new_n7056, new_n23468);
nand_5 g21120(new_n23468, new_n23467, new_n23469);
nand_5 g21121(new_n23469, new_n23466, new_n23470);
nand_5 g21122(new_n23470, new_n23465, new_n23471_1);
xnor_4 g21123(new_n22433_1, new_n17979, new_n23472);
nor_5  g21124(new_n23472, new_n23471_1, new_n23473);
nor_5  g21125(new_n23473, new_n23463_1, new_n23474);
nand_5 g21126(new_n23474, new_n23462, new_n23475);
nand_5 g21127(new_n23475, new_n23460, new_n23476);
nand_5 g21128(new_n23476, new_n23458, new_n23477);
nand_5 g21129(new_n23477, new_n23456, new_n23478);
nand_5 g21130(new_n23478, new_n23455, new_n23479);
nand_5 g21131(new_n23479, new_n23453, new_n23480_1);
xnor_4 g21132(new_n23480_1, new_n19328, new_n23481);
xnor_4 g21133(new_n23481, new_n23450_1, new_n23482);
not_8  g21134(new_n23482, new_n23483);
nand_5 g21135(new_n23483, new_n3436, new_n23484);
xnor_4 g21136(new_n23482, new_n3436, new_n23485);
xnor_4 g21137(new_n23452, new_n19333_1, new_n23486);
xnor_4 g21138(new_n23486, new_n23478, new_n23487);
nand_5 g21139(new_n23487, new_n3446, new_n23488);
xnor_4 g21140(new_n23487, new_n3445, new_n23489);
xnor_4 g21141(new_n23457, new_n19338, new_n23490);
xnor_4 g21142(new_n23490, new_n23476, new_n23491);
not_8  g21143(new_n23491, new_n23492);
nand_5 g21144(new_n23492, new_n3451_1, new_n23493_1);
xnor_4 g21145(new_n23491, new_n3451_1, new_n23494);
xnor_4 g21146(new_n22430, new_n17968_1, new_n23495);
xnor_4 g21147(new_n23495, new_n23474, new_n23496);
nand_5 g21148(new_n23496, new_n3455, new_n23497);
xnor_4 g21149(new_n23496, new_n3457, new_n23498);
not_8  g21150(new_n23472, new_n23499);
xnor_4 g21151(new_n23499, new_n23471_1, new_n23500);
nand_5 g21152(new_n23500, new_n3460_1, new_n23501);
xnor_4 g21153(new_n23500, new_n3462, new_n23502);
xnor_4 g21154(new_n23469, new_n23466, new_n23503);
nand_5 g21155(new_n23503, new_n3467, new_n23504);
not_8  g21156(new_n3467, new_n23505);
xnor_4 g21157(new_n23503, new_n23505, new_n23506);
not_8  g21158(new_n7086, new_n23507);
nand_5 g21159(new_n23507, new_n3471, new_n23508);
nand_5 g21160(new_n7112, new_n7087, new_n23509);
nand_5 g21161(new_n23509, new_n23508, new_n23510);
nand_5 g21162(new_n23510, new_n23506, new_n23511);
nand_5 g21163(new_n23511, new_n23504, new_n23512);
nand_5 g21164(new_n23512, new_n23502, new_n23513_1);
nand_5 g21165(new_n23513_1, new_n23501, new_n23514);
nand_5 g21166(new_n23514, new_n23498, new_n23515);
nand_5 g21167(new_n23515, new_n23497, new_n23516);
nand_5 g21168(new_n23516, new_n23494, new_n23517);
nand_5 g21169(new_n23517, new_n23493_1, new_n23518);
nand_5 g21170(new_n23518, new_n23489, new_n23519);
nand_5 g21171(new_n23519, new_n23488, new_n23520);
nand_5 g21172(new_n23520, new_n23485, new_n23521);
nand_5 g21173(new_n23521, new_n23484, new_n23522);
nor_5  g21174(new_n23480_1, new_n19328, new_n23523);
xnor_4 g21175(new_n23450_1, new_n19286, new_n23524);
nand_5 g21176(new_n23524, new_n23523, new_n23525);
not_8  g21177(new_n23524, new_n23526);
nand_5 g21178(new_n23526, new_n23480_1, new_n23527);
nand_5 g21179(new_n23527, new_n23525, new_n23528);
nor_5  g21180(new_n23528, new_n23522, new_n23529_1);
not_8  g21181(new_n23480_1, new_n23530);
nor_5  g21182(new_n23449, new_n19286, new_n23531);
nand_5 g21183(new_n23531, new_n23530, new_n23532);
xnor_4 g21184(new_n23532, new_n23529_1, n9833);
nor_5  g21185(new_n18691, n13775, new_n23534);
nand_5 g21186(new_n23534, new_n9196, new_n23535);
or_5   g21187(new_n23535, n25972, new_n23536);
nand_5 g21188(new_n23536, new_n19326, new_n23537);
xnor_4 g21189(new_n23535, new_n12752, new_n23538);
nand_5 g21190(new_n23538, new_n19302, new_n23539);
not_8  g21191(new_n23538, new_n23540);
xnor_4 g21192(new_n23540, new_n19302, new_n23541_1);
xnor_4 g21193(new_n23534, n21915, new_n23542);
nand_5 g21194(new_n23542, new_n19307, new_n23543);
xnor_4 g21195(new_n23534, new_n9196, new_n23544);
xnor_4 g21196(new_n23544, new_n19307, new_n23545);
nand_5 g21197(new_n18692, new_n17934, new_n23546_1);
nand_5 g21198(new_n18726, new_n18694, new_n23547);
nand_5 g21199(new_n23547, new_n23546_1, new_n23548);
nand_5 g21200(new_n23548, new_n23545, new_n23549);
nand_5 g21201(new_n23549, new_n23543, new_n23550_1);
nand_5 g21202(new_n23550_1, new_n23541_1, new_n23551);
nand_5 g21203(new_n23551, new_n23539, new_n23552);
nor_5  g21204(new_n23552, new_n23537, new_n23553);
nor_5  g21205(new_n18728, n3710, new_n23554);
and_5  g21206(new_n23554, new_n9341, new_n23555);
not_8  g21207(new_n23555, new_n23556);
nor_5  g21208(new_n23556, n12507, new_n23557);
xnor_4 g21209(new_n23557, new_n17284, new_n23558);
not_8  g21210(new_n13856, new_n23559);
xnor_4 g21211(new_n23555, n12507, new_n23560);
not_8  g21212(new_n23560, new_n23561);
nand_5 g21213(new_n23561, new_n23559, new_n23562);
not_8  g21214(new_n5580, new_n23563);
xnor_4 g21215(new_n23554, n15077, new_n23564);
not_8  g21216(new_n23564, new_n23565);
nand_5 g21217(new_n23565, new_n23563, new_n23566);
xnor_4 g21218(new_n23565, new_n5580, new_n23567);
not_8  g21219(new_n18729, new_n23568);
nor_5  g21220(new_n23568, new_n5620, new_n23569);
not_8  g21221(new_n18730, new_n23570);
nor_5  g21222(new_n18734, new_n23570, new_n23571);
nor_5  g21223(new_n23571, new_n23569, new_n23572);
nand_5 g21224(new_n23572, new_n23567, new_n23573);
nand_5 g21225(new_n23573, new_n23566, new_n23574);
xnor_4 g21226(new_n23561, new_n13856, new_n23575);
nand_5 g21227(new_n23575, new_n23574, new_n23576);
nand_5 g21228(new_n23576, new_n23562, new_n23577);
xnor_4 g21229(new_n23577, new_n23558, new_n23578);
xnor_4 g21230(new_n23536, new_n19326, new_n23579);
xnor_4 g21231(new_n23579, new_n23552, new_n23580);
nand_5 g21232(new_n23580, new_n23578, new_n23581);
not_8  g21233(new_n23578, new_n23582);
xnor_4 g21234(new_n23580, new_n23582, new_n23583);
xnor_4 g21235(new_n23550_1, new_n23541_1, new_n23584);
xnor_4 g21236(new_n23575, new_n23574, new_n23585_1);
not_8  g21237(new_n23585_1, new_n23586_1);
nand_5 g21238(new_n23586_1, new_n23584, new_n23587);
xnor_4 g21239(new_n23585_1, new_n23584, new_n23588_1);
xnor_4 g21240(new_n23572, new_n23567, new_n23589);
not_8  g21241(new_n23589, new_n23590);
xnor_4 g21242(new_n23548, new_n23545, new_n23591);
nand_5 g21243(new_n23591, new_n23590, new_n23592);
xnor_4 g21244(new_n23591, new_n23589, new_n23593);
not_8  g21245(new_n18735, new_n23594);
nand_5 g21246(new_n23594, new_n18727, new_n23595);
nand_5 g21247(new_n18776, new_n18736, new_n23596);
nand_5 g21248(new_n23596, new_n23595, new_n23597);
nand_5 g21249(new_n23597, new_n23593, new_n23598);
nand_5 g21250(new_n23598, new_n23592, new_n23599);
nand_5 g21251(new_n23599, new_n23588_1, new_n23600);
nand_5 g21252(new_n23600, new_n23587, new_n23601);
nand_5 g21253(new_n23601, new_n23583, new_n23602);
nand_5 g21254(new_n23602, new_n23581, new_n23603);
nand_5 g21255(new_n23603, new_n23553, new_n23604);
xnor_4 g21256(new_n23603, new_n23553, new_n23605);
not_8  g21257(new_n23557, new_n23606);
nand_5 g21258(new_n23606, new_n17284, new_n23607);
not_8  g21259(new_n23607, new_n23608);
nand_5 g21260(new_n23577, new_n23608, new_n23609);
not_8  g21261(new_n23609, new_n23610);
nand_5 g21262(new_n23610, new_n23605, new_n23611);
nand_5 g21263(new_n23611, new_n23604, n9838);
xnor_4 g21264(new_n21116, new_n21113, n9867);
not_8  g21265(new_n8530, new_n23614);
not_8  g21266(new_n22016_1, new_n23615);
nand_5 g21267(new_n20642, n12702, new_n23616);
nand_5 g21268(new_n20647, new_n20643, new_n23617);
nand_5 g21269(new_n23617, new_n23616, new_n23618);
nand_5 g21270(new_n23618, new_n23615, new_n23619_1);
xnor_4 g21271(new_n23618, new_n22016_1, new_n23620);
not_8  g21272(new_n23620, new_n23621);
nand_5 g21273(new_n23621, new_n8635, new_n23622);
nand_5 g21274(new_n20648, new_n8642, new_n23623);
nand_5 g21275(new_n20652, new_n20649, new_n23624_1);
nand_5 g21276(new_n23624_1, new_n23623, new_n23625);
xnor_4 g21277(new_n23620, new_n8635, new_n23626);
nand_5 g21278(new_n23626, new_n23625, new_n23627);
nand_5 g21279(new_n23627, new_n23622, new_n23628_1);
nand_5 g21280(new_n23628_1, new_n23619_1, new_n23629);
nand_5 g21281(new_n23629, new_n23614, new_n23630);
not_8  g21282(new_n23630, n9890);
and_5  g21283(new_n19349, new_n19337, new_n23632);
nor_5  g21284(new_n23632, new_n19350, n9917);
xnor_4 g21285(new_n22304, new_n22296, n9919);
xnor_4 g21286(new_n19535, new_n19519, n9938);
xnor_4 g21287(new_n19138, new_n19137, n9946);
not_8  g21288(new_n18612, new_n23637_1);
xnor_4 g21289(n21784, new_n5220, new_n23638);
not_8  g21290(new_n23638, new_n23639);
or_5   g21291(n5521, n2858, new_n23640);
xnor_4 g21292(n5521, new_n5158_1, new_n23641);
or_5   g21293(n11926, n2659, new_n23642);
xnor_4 g21294(n11926, new_n5162, new_n23643);
or_5   g21295(n24327, n4325, new_n23644);
xnor_4 g21296(n24327, new_n6318, new_n23645);
or_5   g21297(new_n5170, new_n4003, new_n23646);
not_8  g21298(new_n23646, new_n23647);
nor_5  g21299(n22198, n5337, new_n23648);
nor_5  g21300(n20826, n626, new_n23649);
not_8  g21301(new_n13823, new_n23650);
nor_5  g21302(new_n13827, new_n23650, new_n23651);
nor_5  g21303(new_n23651, new_n23649, new_n23652);
not_8  g21304(new_n23652, new_n23653);
nor_5  g21305(new_n23653, new_n23648, new_n23654);
nor_5  g21306(new_n23654, new_n23647, new_n23655);
nand_5 g21307(new_n23655, new_n23645, new_n23656);
nand_5 g21308(new_n23656, new_n23644, new_n23657_1);
nand_5 g21309(new_n23657_1, new_n23643, new_n23658);
nand_5 g21310(new_n23658, new_n23642, new_n23659);
nand_5 g21311(new_n23659, new_n23641, new_n23660);
nand_5 g21312(new_n23660, new_n23640, new_n23661);
xnor_4 g21313(new_n23661, new_n23639, new_n23662);
xnor_4 g21314(new_n23662, new_n5089, new_n23663_1);
not_8  g21315(new_n23641, new_n23664);
xnor_4 g21316(new_n23659, new_n23664, new_n23665);
nand_5 g21317(new_n23665, new_n5094, new_n23666);
xnor_4 g21318(new_n23665, new_n5093, new_n23667);
xnor_4 g21319(new_n23657_1, new_n23643, new_n23668);
not_8  g21320(new_n23668, new_n23669_1);
nand_5 g21321(new_n23669_1, new_n5097, new_n23670);
xnor_4 g21322(new_n23655, new_n23645, new_n23671);
not_8  g21323(new_n23671, new_n23672);
nand_5 g21324(new_n23672, new_n5102, new_n23673);
xnor_4 g21325(new_n23671, new_n5102, new_n23674);
xnor_4 g21326(n22198, new_n4003, new_n23675);
xnor_4 g21327(new_n23675, new_n23653, new_n23676);
nor_5  g21328(new_n23676, new_n5106, new_n23677);
nor_5  g21329(new_n13828, new_n13822, new_n23678);
not_8  g21330(new_n23678, new_n23679);
nand_5 g21331(new_n13830, new_n13807, new_n23680);
nand_5 g21332(new_n23680, new_n23679, new_n23681);
xnor_4 g21333(new_n23676, new_n5107, new_n23682);
not_8  g21334(new_n23682, new_n23683);
nor_5  g21335(new_n23683, new_n23681, new_n23684_1);
nor_5  g21336(new_n23684_1, new_n23677, new_n23685);
not_8  g21337(new_n23685, new_n23686);
nand_5 g21338(new_n23686, new_n23674, new_n23687);
nand_5 g21339(new_n23687, new_n23673, new_n23688);
xnor_4 g21340(new_n23668, new_n5097, new_n23689);
nand_5 g21341(new_n23689, new_n23688, new_n23690_1);
nand_5 g21342(new_n23690_1, new_n23670, new_n23691);
nand_5 g21343(new_n23691, new_n23667, new_n23692);
nand_5 g21344(new_n23692, new_n23666, new_n23693);
xnor_4 g21345(new_n23693, new_n23663_1, new_n23694);
xnor_4 g21346(new_n23694, new_n23637_1, new_n23695);
not_8  g21347(new_n17868, new_n23696);
xnor_4 g21348(new_n23691, new_n23667, new_n23697_1);
not_8  g21349(new_n23697_1, new_n23698);
nand_5 g21350(new_n23698, new_n23696, new_n23699);
not_8  g21351(new_n23699, new_n23700);
xnor_4 g21352(new_n23697_1, new_n23696, new_n23701);
not_8  g21353(new_n23701, new_n23702);
not_8  g21354(new_n17870, new_n23703);
xnor_4 g21355(new_n23689, new_n23688, new_n23704);
not_8  g21356(new_n23704, new_n23705);
nand_5 g21357(new_n23705, new_n23703, new_n23706);
not_8  g21358(new_n23706, new_n23707);
xnor_4 g21359(new_n23704, new_n23703, new_n23708);
not_8  g21360(new_n23708, new_n23709);
not_8  g21361(new_n3925_1, new_n23710);
xnor_4 g21362(new_n23686, new_n23674, new_n23711);
not_8  g21363(new_n23711, new_n23712);
nand_5 g21364(new_n23712, new_n23710, new_n23713);
not_8  g21365(new_n23713, new_n23714_1);
xnor_4 g21366(new_n23711, new_n3925_1, new_n23715);
not_8  g21367(new_n3927, new_n23716);
xnor_4 g21368(new_n23682, new_n23681, new_n23717_1);
nor_5  g21369(new_n23717_1, new_n23716, new_n23718);
nor_5  g21370(new_n13831, new_n13806, new_n23719_1);
nor_5  g21371(new_n13845, new_n13832, new_n23720);
nor_5  g21372(new_n23720, new_n23719_1, new_n23721);
xnor_4 g21373(new_n23717_1, new_n3927, new_n23722);
not_8  g21374(new_n23722, new_n23723);
nor_5  g21375(new_n23723, new_n23721, new_n23724);
nor_5  g21376(new_n23724, new_n23718, new_n23725);
not_8  g21377(new_n23725, new_n23726);
nor_5  g21378(new_n23726, new_n23715, new_n23727);
nor_5  g21379(new_n23727, new_n23714_1, new_n23728);
nor_5  g21380(new_n23728, new_n23709, new_n23729);
nor_5  g21381(new_n23729, new_n23707, new_n23730);
nor_5  g21382(new_n23730, new_n23702, new_n23731);
nor_5  g21383(new_n23731, new_n23700, new_n23732);
xnor_4 g21384(new_n23732, new_n23695, n9968);
nand_5 g21385(new_n21961, new_n14841, new_n23734);
not_8  g21386(new_n23734, new_n23735);
xnor_4 g21387(new_n21961, new_n14842, new_n23736);
not_8  g21388(new_n23736, new_n23737);
nand_5 g21389(new_n21972, new_n14841, new_n23738);
xnor_4 g21390(new_n21971, new_n14841, new_n23739);
nor_5  g21391(new_n12055, new_n11993, new_n23740);
nor_5  g21392(new_n12103, new_n12056, new_n23741);
nor_5  g21393(new_n23741, new_n23740, new_n23742);
nand_5 g21394(new_n23742, new_n23739, new_n23743);
nand_5 g21395(new_n23743, new_n23738, new_n23744);
nor_5  g21396(new_n23744, new_n23737, new_n23745);
nor_5  g21397(new_n23745, new_n23735, n10009);
xnor_4 g21398(new_n22727, new_n22724, n10010);
and_5  g21399(new_n17281, new_n11765, new_n23748_1);
not_8  g21400(new_n15745, new_n23749);
nor_5  g21401(new_n15777, new_n23749, new_n23750);
nor_5  g21402(new_n23750, new_n23748_1, new_n23751);
not_8  g21403(new_n23751, new_n23752);
nor_5  g21404(new_n23752, new_n21982, new_n23753);
xnor_4 g21405(new_n23751, new_n21982, new_n23754);
not_8  g21406(new_n23754, new_n23755_1);
nor_5  g21407(new_n15815_1, new_n15778, new_n23756);
nor_5  g21408(new_n15856, new_n15816_1, new_n23757);
nor_5  g21409(new_n23757, new_n23756, new_n23758);
nor_5  g21410(new_n23758, new_n23755_1, new_n23759);
nor_5  g21411(new_n23759, new_n23753, n10019);
xnor_4 g21412(new_n15641, new_n15586, n10021);
xor_4  g21413(new_n10219, new_n10209, n10055);
xnor_4 g21414(new_n11389, new_n11368, n10101);
xnor_4 g21415(new_n4811, new_n4759, n10111);
nor_5  g21416(n16544, new_n16856, new_n23765);
xnor_4 g21417(n16544, n3324, new_n23766);
not_8  g21418(new_n23766, new_n23767);
nor_5  g21419(new_n16884, n6814, new_n23768);
xnor_4 g21420(n17911, n6814, new_n23769);
not_8  g21421(new_n23769, new_n23770);
nor_5  g21422(new_n16889, n19701, new_n23771);
xnor_4 g21423(n21997, n19701, new_n23772);
not_8  g21424(new_n23772, new_n23773);
nor_5  g21425(new_n16894, n23529, new_n23774);
xnor_4 g21426(n25119, n23529, new_n23775_1);
not_8  g21427(new_n23775_1, new_n23776);
nor_5  g21428(n24620, new_n9035, new_n23777);
xnor_4 g21429(n24620, n1163, new_n23778);
not_8  g21430(new_n23778, new_n23779);
nor_5  g21431(new_n16237, n5211, new_n23780);
nor_5  g21432(n18537, new_n2955, new_n23781);
nor_5  g21433(new_n9546, n7057, new_n23782);
not_8  g21434(new_n10080, new_n23783);
nor_5  g21435(new_n10092, new_n23783, new_n23784);
nor_5  g21436(new_n23784, new_n23782, new_n23785);
not_8  g21437(new_n23785, new_n23786);
nor_5  g21438(new_n23786, new_n23781, new_n23787);
nor_5  g21439(new_n23787, new_n23780, new_n23788);
nor_5  g21440(new_n23788, new_n23779, new_n23789);
nor_5  g21441(new_n23789, new_n23777, new_n23790);
nor_5  g21442(new_n23790, new_n23776, new_n23791);
nor_5  g21443(new_n23791, new_n23774, new_n23792);
nor_5  g21444(new_n23792, new_n23773, new_n23793);
nor_5  g21445(new_n23793, new_n23771, new_n23794);
nor_5  g21446(new_n23794, new_n23770, new_n23795);
nor_5  g21447(new_n23795, new_n23768, new_n23796);
nor_5  g21448(new_n23796, new_n23767, new_n23797);
nor_5  g21449(new_n23797, new_n23765, new_n23798);
xnor_4 g21450(new_n23798, new_n22884, new_n23799);
not_8  g21451(new_n23798, new_n23800);
nor_5  g21452(new_n23800, new_n22897_1, new_n23801);
nor_5  g21453(new_n23798, new_n22896, new_n23802);
xnor_4 g21454(new_n23796, new_n23766, new_n23803);
not_8  g21455(new_n23803, new_n23804);
nand_5 g21456(new_n23804, new_n18453, new_n23805);
xnor_4 g21457(new_n23803, new_n18453, new_n23806);
xnor_4 g21458(new_n23794, new_n23769, new_n23807);
nor_5  g21459(new_n23807, new_n18502, new_n23808);
not_8  g21460(new_n23808, new_n23809);
xnor_4 g21461(new_n23807, new_n18500, new_n23810);
xnor_4 g21462(new_n23792, new_n23772, new_n23811);
nor_5  g21463(new_n23811, new_n18509_1, new_n23812);
not_8  g21464(new_n23812, new_n23813);
xnor_4 g21465(new_n23811, new_n18507, new_n23814);
not_8  g21466(new_n23814, new_n23815);
xnor_4 g21467(new_n23790, new_n23775_1, new_n23816);
nor_5  g21468(new_n23816, new_n18515_1, new_n23817);
xnor_4 g21469(new_n23816, new_n18513_1, new_n23818);
not_8  g21470(new_n23818, new_n23819);
xnor_4 g21471(new_n23788, new_n23778, new_n23820);
nor_5  g21472(new_n23820, new_n18517, new_n23821);
xnor_4 g21473(n18537, n5211, new_n23822);
xnor_4 g21474(new_n23822, new_n23785, new_n23823);
nor_5  g21475(new_n23823, new_n18525, new_n23824);
not_8  g21476(new_n23824, new_n23825);
xnor_4 g21477(new_n23823, new_n18525, new_n23826);
not_8  g21478(new_n23826, new_n23827);
nor_5  g21479(new_n10093, new_n10078, new_n23828);
not_8  g21480(new_n23828, new_n23829);
not_8  g21481(new_n10118, new_n23830);
nand_5 g21482(new_n23830, new_n10094, new_n23831_1);
nand_5 g21483(new_n23831_1, new_n23829, new_n23832);
nand_5 g21484(new_n23832, new_n23827, new_n23833);
nand_5 g21485(new_n23833, new_n23825, new_n23834);
not_8  g21486(new_n23834, new_n23835);
xnor_4 g21487(new_n23820, new_n18518, new_n23836);
nand_5 g21488(new_n23836, new_n23835, new_n23837);
not_8  g21489(new_n23837, new_n23838);
nor_5  g21490(new_n23838, new_n23821, new_n23839);
nor_5  g21491(new_n23839, new_n23819, new_n23840);
nor_5  g21492(new_n23840, new_n23817, new_n23841);
nor_5  g21493(new_n23841, new_n23815, new_n23842_1);
not_8  g21494(new_n23842_1, new_n23843);
nand_5 g21495(new_n23843, new_n23813, new_n23844);
nand_5 g21496(new_n23844, new_n23810, new_n23845);
nand_5 g21497(new_n23845, new_n23809, new_n23846);
nand_5 g21498(new_n23846, new_n23806, new_n23847);
nand_5 g21499(new_n23847, new_n23805, new_n23848);
nor_5  g21500(new_n23848, new_n23802, new_n23849_1);
nor_5  g21501(new_n23849_1, new_n23801, new_n23850);
xnor_4 g21502(new_n23850, new_n23799, n10165);
xnor_4 g21503(new_n13924, new_n13922_1, n10236);
xnor_4 g21504(new_n15502, new_n15476, n10239);
xnor_4 g21505(new_n6752, new_n6705, n10244);
xnor_4 g21506(new_n19458_1, new_n19443, n10261);
xnor_4 g21507(new_n16852, new_n16837_1, n10262);
not_8  g21508(new_n18146, new_n23857);
xnor_4 g21509(new_n23857, new_n18145_1, n10287);
nand_5 g21510(new_n23127, new_n16361, new_n23859);
xnor_4 g21511(new_n23171, new_n23859, new_n23860);
not_8  g21512(new_n23128, new_n23861);
nand_5 g21513(new_n23133, new_n23861, new_n23862);
nand_5 g21514(new_n23146_1, new_n23134, new_n23863);
nand_5 g21515(new_n23863, new_n23862, new_n23864);
xnor_4 g21516(new_n23864, new_n23860, n10295);
xnor_4 g21517(new_n15964, new_n15961, n10321);
xnor_4 g21518(new_n15504, new_n15473, n10326);
xnor_4 g21519(new_n2883, new_n2870, n10327);
xnor_4 g21520(new_n21971, new_n21947, new_n23869);
xnor_4 g21521(new_n23869, new_n21966, n10330);
xnor_4 g21522(new_n22639, new_n22599, n10340);
xnor_4 g21523(new_n18142, new_n18138, new_n23872);
xnor_4 g21524(new_n23872, new_n18147, n10345);
nand_5 g21525(new_n15119, new_n5148, new_n23874);
and_5  g21526(new_n22951, new_n23874, new_n23875);
nand_5 g21527(new_n20597, new_n5152, new_n23876);
xnor_4 g21528(new_n20598, new_n5152, new_n23877);
not_8  g21529(new_n5153, new_n23878);
nand_5 g21530(new_n20604_1, new_n23878, new_n23879);
xnor_4 g21531(new_n20604_1, new_n5153, new_n23880);
not_8  g21532(new_n5156, new_n23881);
nand_5 g21533(new_n20611, new_n23881, new_n23882);
xnor_4 g21534(new_n20611, new_n5156, new_n23883_1);
not_8  g21535(new_n5160, new_n23884);
nand_5 g21536(new_n20617, new_n23884, new_n23885);
xnor_4 g21537(new_n20617, new_n5160, new_n23886);
not_8  g21538(new_n5164, new_n23887);
nand_5 g21539(new_n9976, new_n23887, new_n23888_1);
xnor_4 g21540(new_n9976, new_n5164, new_n23889);
not_8  g21541(new_n5168_1, new_n23890);
nand_5 g21542(new_n9982, new_n23890, new_n23891);
xnor_4 g21543(new_n9980, new_n23890, new_n23892);
not_8  g21544(new_n5172, new_n23893);
nand_5 g21545(new_n9987, new_n23893, new_n23894);
xnor_4 g21546(new_n9985, new_n23893, new_n23895_1);
nor_5  g21547(new_n9991, new_n5177, new_n23896);
xnor_4 g21548(new_n9991, new_n5178, new_n23897);
not_8  g21549(new_n23897, new_n23898);
and_5  g21550(new_n9997, new_n5183, new_n23899_1);
xnor_4 g21551(new_n9999, new_n5183, new_n23900);
not_8  g21552(new_n23900, new_n23901);
nor_5  g21553(new_n10005, new_n5192, new_n23902);
not_8  g21554(new_n23902, new_n23903_1);
nor_5  g21555(new_n23903_1, new_n10010_1, new_n23904);
not_8  g21556(new_n5188, new_n23905);
xnor_4 g21557(new_n23903_1, new_n10002, new_n23906);
not_8  g21558(new_n23906, new_n23907);
nor_5  g21559(new_n23907, new_n23905, new_n23908);
nor_5  g21560(new_n23908, new_n23904, new_n23909);
nor_5  g21561(new_n23909, new_n23901, new_n23910);
nor_5  g21562(new_n23910, new_n23899_1, new_n23911);
nor_5  g21563(new_n23911, new_n23898, new_n23912_1);
nor_5  g21564(new_n23912_1, new_n23896, new_n23913_1);
not_8  g21565(new_n23913_1, new_n23914);
nand_5 g21566(new_n23914, new_n23895_1, new_n23915);
nand_5 g21567(new_n23915, new_n23894, new_n23916);
nand_5 g21568(new_n23916, new_n23892, new_n23917);
nand_5 g21569(new_n23917, new_n23891, new_n23918);
nand_5 g21570(new_n23918, new_n23889, new_n23919);
nand_5 g21571(new_n23919, new_n23888_1, new_n23920);
nand_5 g21572(new_n23920, new_n23886, new_n23921);
nand_5 g21573(new_n23921, new_n23885, new_n23922);
nand_5 g21574(new_n23922, new_n23883_1, new_n23923_1);
nand_5 g21575(new_n23923_1, new_n23882, new_n23924_1);
nand_5 g21576(new_n23924_1, new_n23880, new_n23925);
nand_5 g21577(new_n23925, new_n23879, new_n23926);
nand_5 g21578(new_n23926, new_n23877, new_n23927);
nand_5 g21579(new_n23927, new_n23876, new_n23928);
xnor_4 g21580(new_n20592, new_n23874, new_n23929);
not_8  g21581(new_n23929, new_n23930);
nor_5  g21582(new_n23930, new_n23928, new_n23931);
nor_5  g21583(new_n23931, new_n23875, n10356);
xnor_4 g21584(new_n21224, new_n21222_1, n10385);
nand_5 g21585(new_n21478, new_n20592, new_n23934);
not_8  g21586(new_n23934, new_n23935_1);
nor_5  g21587(new_n21478, new_n20592, new_n23936);
nor_5  g21588(new_n23936, new_n21410, new_n23937);
nor_5  g21589(new_n23937, new_n23935_1, new_n23938);
nor_5  g21590(new_n23938, new_n21408, n10387);
xnor_4 g21591(new_n21712, new_n21696, n10388);
xnor_4 g21592(new_n16612, new_n16563, n10390);
xnor_4 g21593(new_n10104, new_n10103, n10404);
xnor_4 g21594(new_n17044, new_n17040, n10409);
xnor_4 g21595(new_n17263_1, new_n9092, n10420);
xnor_4 g21596(new_n19449, new_n7334, n10432);
not_8  g21597(new_n22099, new_n23946);
xnor_4 g21598(new_n22720, new_n23946, new_n23947);
not_8  g21599(new_n10258, new_n23948);
nor_5  g21600(new_n22103, new_n23948, new_n23949);
nor_5  g21601(new_n22369, new_n22362, new_n23950);
nor_5  g21602(new_n23950, new_n23949, new_n23951);
xnor_4 g21603(new_n23951, new_n23947, new_n23952);
xnor_4 g21604(new_n23952, new_n12231, new_n23953);
not_8  g21605(new_n23953, new_n23954_1);
nor_5  g21606(new_n22370, new_n12237, new_n23955);
nor_5  g21607(new_n22380, new_n23955, new_n23956);
xnor_4 g21608(new_n23956, new_n23954_1, n10484);
xnor_4 g21609(new_n12092, new_n12076, n10489);
xnor_4 g21610(new_n14399, new_n3785_1, n10525);
xnor_4 g21611(new_n18752, new_n12936, new_n23960);
xnor_4 g21612(new_n23960, new_n18765, n10540);
xnor_4 g21613(new_n17164, new_n17134, n10561);
xnor_4 g21614(new_n16616, new_n16553, n10564);
xnor_4 g21615(new_n10670, new_n10668, n10588);
xnor_4 g21616(new_n10674, new_n10671, n10595);
xor_4  g21617(new_n22496, new_n22482, n10617);
xnor_4 g21618(new_n13292, new_n13224, n10628);
xnor_4 g21619(new_n11334, new_n6035, new_n23968);
nand_5 g21620(new_n11343, new_n6039, new_n23969);
xnor_4 g21621(new_n11343, new_n6038, new_n23970);
not_8  g21622(new_n11346, new_n23971);
nor_5  g21623(new_n23971, new_n6043, new_n23972);
xnor_4 g21624(new_n11346, new_n6043, new_n23973);
not_8  g21625(new_n23973, new_n23974_1);
nor_5  g21626(new_n6083, new_n6050, new_n23975);
nor_5  g21627(new_n23975, new_n6092, new_n23976);
not_8  g21628(new_n23976, new_n23977);
xnor_4 g21629(new_n23975, new_n6093, new_n23978);
nand_5 g21630(new_n23978, new_n6059, new_n23979);
nand_5 g21631(new_n23979, new_n23977, new_n23980);
not_8  g21632(new_n23980, new_n23981);
nor_5  g21633(new_n23981, new_n23974_1, new_n23982);
nor_5  g21634(new_n23982, new_n23972, new_n23983);
not_8  g21635(new_n23983, new_n23984);
nand_5 g21636(new_n23984, new_n23970, new_n23985);
nand_5 g21637(new_n23985, new_n23969, new_n23986_1);
xnor_4 g21638(new_n23986_1, new_n23968, n10647);
nor_5  g21639(new_n8854, new_n8848, new_n23988);
nor_5  g21640(new_n21101, new_n3722, new_n23989);
not_8  g21641(new_n23989, new_n23990);
not_8  g21642(new_n3737, new_n23991);
nor_5  g21643(new_n3806, new_n23991, new_n23992);
nor_5  g21644(new_n23992, new_n21100, new_n23993);
nand_5 g21645(new_n23993, new_n23990, new_n23994);
nor_5  g21646(new_n23994, new_n14359, new_n23995);
xnor_4 g21647(new_n23995, new_n23988, new_n23996);
xnor_4 g21648(new_n23994, new_n14358, new_n23997);
nor_5  g21649(new_n23997, new_n8857, new_n23998);
not_8  g21650(new_n23998, new_n23999);
not_8  g21651(new_n3807, new_n24000);
nand_5 g21652(new_n24000, new_n3673, new_n24001);
nand_5 g21653(new_n3875, new_n3808, new_n24002_1);
nand_5 g21654(new_n24002_1, new_n24001, new_n24003);
not_8  g21655(new_n24003, new_n24004_1);
xnor_4 g21656(new_n23997, new_n8856_1, new_n24005);
nand_5 g21657(new_n24005, new_n24004_1, new_n24006);
nand_5 g21658(new_n24006, new_n23999, new_n24007);
xnor_4 g21659(new_n24007, new_n23996, n10653);
xnor_4 g21660(new_n9625, new_n9624, n10692);
xor_4  g21661(new_n15692, new_n4491, n10694);
xnor_4 g21662(new_n21556, new_n21530, n10701);
xnor_4 g21663(new_n6463, new_n6445, n10756);
or_5   g21664(new_n19485, n5101, new_n24013);
nand_5 g21665(new_n17005, new_n17001, new_n24014);
nand_5 g21666(new_n24014, new_n24013, new_n24015);
nor_5  g21667(new_n17006_1, n13419, new_n24016);
not_8  g21668(new_n17006_1, new_n24017);
nor_5  g21669(new_n24017, new_n17000, new_n24018);
nor_5  g21670(new_n16950, n4967, new_n24019);
nor_5  g21671(new_n16951_1, new_n16953, new_n24020);
nor_5  g21672(new_n20502, new_n24020, new_n24021);
nor_5  g21673(new_n24021, new_n24019, new_n24022);
nor_5  g21674(new_n24022, new_n24018, new_n24023);
nor_5  g21675(new_n24023, new_n24016, new_n24024);
nand_5 g21676(new_n24024, new_n24015, new_n24025);
xnor_4 g21677(new_n24025, new_n3292, new_n24026);
xnor_4 g21678(new_n24024, new_n24015, new_n24027);
nor_5  g21679(new_n24027, new_n3438, new_n24028);
xnor_4 g21680(new_n24027, new_n3438, new_n24029);
xnor_4 g21681(new_n24022, new_n17007, new_n24030);
nor_5  g21682(new_n24030, new_n3307, new_n24031);
xnor_4 g21683(new_n24030, new_n3307, new_n24032_1);
not_8  g21684(new_n3313, new_n24033);
nand_5 g21685(new_n20503, new_n24033, new_n24034);
nand_5 g21686(new_n20554, new_n20504, new_n24035);
nand_5 g21687(new_n24035, new_n24034, new_n24036);
nor_5  g21688(new_n24036, new_n24032_1, new_n24037);
nor_5  g21689(new_n24037, new_n24031, new_n24038);
nor_5  g21690(new_n24038, new_n24029, new_n24039_1);
nor_5  g21691(new_n24039_1, new_n24028, new_n24040);
xnor_4 g21692(new_n24040, new_n24026, n10775);
xnor_4 g21693(new_n22405, new_n22398, n10780);
xnor_4 g21694(n17095, new_n4301, new_n24043);
nor_5  g21695(n22591, n22274, new_n24044);
nand_5 g21696(n26167, n24129, new_n24045);
xnor_4 g21697(n22591, new_n4303, new_n24046);
nand_5 g21698(new_n24046, new_n24045, new_n24047);
not_8  g21699(new_n24047, new_n24048_1);
nor_5  g21700(new_n24048_1, new_n24044, new_n24049);
xnor_4 g21701(new_n24049, new_n24043, new_n24050);
xnor_4 g21702(new_n24050, n21749, new_n24051);
nand_5 g21703(new_n9483, n21138, new_n24052_1);
nand_5 g21704(new_n24052_1, new_n10133, new_n24053);
not_8  g21705(new_n24053, new_n24054);
xnor_4 g21706(new_n24046, new_n24045, new_n24055);
xnor_4 g21707(new_n24052_1, n7769, new_n24056);
and_5  g21708(new_n24056, new_n24055, new_n24057);
nor_5  g21709(new_n24057, new_n24054, new_n24058);
xnor_4 g21710(new_n24058, new_n24051, new_n24059);
xnor_4 g21711(new_n24059, new_n19632, new_n24060);
not_8  g21712(new_n24056, new_n24061);
xnor_4 g21713(new_n24061, new_n24055, new_n24062);
and_5  g21714(new_n24062, new_n19635, new_n24063);
nor_5  g21715(new_n9484, new_n19639, new_n24064);
not_8  g21716(new_n24064, new_n24065);
xnor_4 g21717(new_n24062, new_n19635, new_n24066);
nor_5  g21718(new_n24066, new_n24065, new_n24067);
nor_5  g21719(new_n24067, new_n24063, new_n24068);
xor_4  g21720(new_n24068, new_n24060, n10817);
nor_5  g21721(new_n23158, new_n23154, new_n24070);
nand_5 g21722(new_n23153, new_n23148, new_n24071);
nand_5 g21723(new_n23158, new_n23154, new_n24072);
nand_5 g21724(new_n23164, new_n24072, new_n24073);
nand_5 g21725(new_n24073, new_n24071, new_n24074);
nor_5  g21726(new_n24074, new_n24070, new_n24075);
nor_5  g21727(new_n24075, new_n12479, new_n24076);
nand_5 g21728(new_n23165, new_n8187, new_n24077);
nand_5 g21729(new_n23169, new_n23166_1, new_n24078);
nand_5 g21730(new_n24078, new_n24077, new_n24079);
xnor_4 g21731(new_n24075, new_n8187, new_n24080);
not_8  g21732(new_n24080, new_n24081);
nor_5  g21733(new_n24081, new_n24079, new_n24082);
nor_5  g21734(new_n24082, new_n24076, n10834);
xnor_4 g21735(new_n23428, new_n23408, n10851);
xnor_4 g21736(new_n22944, new_n22935, n10874);
xnor_4 g21737(new_n23628_1, new_n23619_1, new_n24086);
xnor_4 g21738(new_n24086, new_n23614, n10924);
nor_5  g21739(new_n11903, new_n11837_1, new_n24088);
not_8  g21740(new_n11841_1, new_n24089);
nor_5  g21741(new_n11906, new_n24089, new_n24090);
nor_5  g21742(new_n24090, new_n24088, n10943);
xnor_4 g21743(new_n12688, new_n12648, n10961);
xnor_4 g21744(new_n11275_1, new_n11262, n11005);
xnor_4 g21745(new_n22690, new_n22681, n11023);
nand_5 g21746(new_n19321, new_n7706, new_n24095);
xnor_4 g21747(new_n19290, new_n7706, new_n24096_1);
nor_5  g21748(new_n19292, new_n7713, new_n24097_1);
not_8  g21749(new_n24097_1, new_n24098);
xnor_4 g21750(new_n19292, new_n7710, new_n24099);
nor_5  g21751(new_n19295, new_n7717, new_n24100);
xnor_4 g21752(new_n17919, new_n7716, new_n24101);
not_8  g21753(new_n12879, new_n24102);
nor_5  g21754(new_n24102, new_n7723, new_n24103);
nor_5  g21755(new_n12911, new_n12880, new_n24104);
nor_5  g21756(new_n24104, new_n24103, new_n24105_1);
nor_5  g21757(new_n24105_1, new_n24101, new_n24106);
nor_5  g21758(new_n24106, new_n24100, new_n24107);
nand_5 g21759(new_n24107, new_n24099, new_n24108);
nand_5 g21760(new_n24108, new_n24098, new_n24109);
nand_5 g21761(new_n24109, new_n24096_1, new_n24110);
nand_5 g21762(new_n24110, new_n24095, new_n24111);
nand_5 g21763(new_n24111, new_n7684, new_n24112);
nor_5  g21764(new_n24112, new_n19319, new_n24113);
xnor_4 g21765(new_n24111, new_n7684, new_n24114);
xnor_4 g21766(new_n24114, new_n19320, new_n24115);
not_8  g21767(new_n24115, new_n24116);
nand_5 g21768(new_n24116, new_n23578, new_n24117);
xnor_4 g21769(new_n24115, new_n23578, new_n24118);
not_8  g21770(new_n24096_1, new_n24119_1);
xnor_4 g21771(new_n24109, new_n24119_1, new_n24120);
nand_5 g21772(new_n24120, new_n23586_1, new_n24121);
xnor_4 g21773(new_n24120, new_n23585_1, new_n24122);
not_8  g21774(new_n24099, new_n24123);
xnor_4 g21775(new_n24107, new_n24123, new_n24124);
nand_5 g21776(new_n24124, new_n23590, new_n24125);
xnor_4 g21777(new_n24124, new_n23589, new_n24126);
xnor_4 g21778(new_n24105_1, new_n24101, new_n24127);
nand_5 g21779(new_n24127, new_n23594, new_n24128);
xnor_4 g21780(new_n24127, new_n18735, new_n24129_1);
nand_5 g21781(new_n12912, new_n18737_1, new_n24130);
nand_5 g21782(new_n12959, new_n12913, new_n24131);
nand_5 g21783(new_n24131, new_n24130, new_n24132);
nand_5 g21784(new_n24132, new_n24129_1, new_n24133_1);
nand_5 g21785(new_n24133_1, new_n24128, new_n24134);
nand_5 g21786(new_n24134, new_n24126, new_n24135);
nand_5 g21787(new_n24135, new_n24125, new_n24136);
nand_5 g21788(new_n24136, new_n24122, new_n24137);
nand_5 g21789(new_n24137, new_n24121, new_n24138);
nand_5 g21790(new_n24138, new_n24118, new_n24139);
nand_5 g21791(new_n24139, new_n24117, new_n24140);
nand_5 g21792(new_n24140, new_n24113, new_n24141_1);
xnor_4 g21793(new_n24140, new_n24113, new_n24142);
nand_5 g21794(new_n24142, new_n23610, new_n24143);
nand_5 g21795(new_n24143, new_n24141_1, n11025);
xnor_4 g21796(new_n17544, new_n9196, new_n24145_1);
nand_5 g21797(new_n17547, n13775, new_n24146_1);
xnor_4 g21798(new_n17547, new_n7219, new_n24147);
nand_5 g21799(new_n17550, n1293, new_n24148);
xnor_4 g21800(new_n17550, new_n7223, new_n24149);
nand_5 g21801(new_n17554, n19042, new_n24150_1);
nand_5 g21802(new_n20367, new_n20363, new_n24151);
nand_5 g21803(new_n24151, new_n24150_1, new_n24152);
nand_5 g21804(new_n24152, new_n24149, new_n24153);
nand_5 g21805(new_n24153, new_n24148, new_n24154);
nand_5 g21806(new_n24154, new_n24147, new_n24155_1);
nand_5 g21807(new_n24155_1, new_n24146_1, new_n24156);
xnor_4 g21808(new_n24156, new_n24145_1, new_n24157);
nor_5  g21809(new_n20369, n26752, new_n24158);
nand_5 g21810(new_n24158, new_n6652_1, new_n24159);
nor_5  g21811(new_n24159, n25464, new_n24160_1);
xnor_4 g21812(new_n24160_1, n3795, new_n24161);
xnor_4 g21813(new_n24161, new_n9340, new_n24162);
xnor_4 g21814(new_n24159, n25464, new_n24163);
nand_5 g21815(new_n24163, new_n9348, new_n24164);
not_8  g21816(new_n24163, new_n24165);
xnor_4 g21817(new_n24165, new_n9348, new_n24166);
xnor_4 g21818(new_n24158, n4590, new_n24167_1);
not_8  g21819(new_n24167_1, new_n24168);
nand_5 g21820(new_n24168, new_n9355, new_n24169);
xnor_4 g21821(new_n24167_1, new_n9355, new_n24170_1);
nand_5 g21822(new_n20370, new_n9360, new_n24171);
not_8  g21823(new_n20371, new_n24172_1);
nand_5 g21824(new_n20374, new_n24172_1, new_n24173);
nand_5 g21825(new_n24173, new_n24171, new_n24174);
nand_5 g21826(new_n24174, new_n24170_1, new_n24175);
nand_5 g21827(new_n24175, new_n24169, new_n24176);
nand_5 g21828(new_n24176, new_n24166, new_n24177_1);
nand_5 g21829(new_n24177_1, new_n24164, new_n24178);
xnor_4 g21830(new_n24178, new_n24162, new_n24179);
xnor_4 g21831(new_n24179, new_n24157, new_n24180);
xnor_4 g21832(new_n24154, new_n24147, new_n24181);
xnor_4 g21833(new_n24176, new_n24166, new_n24182);
not_8  g21834(new_n24182, new_n24183);
nand_5 g21835(new_n24183, new_n24181, new_n24184);
xnor_4 g21836(new_n24182, new_n24181, new_n24185);
xnor_4 g21837(new_n24152, new_n24149, new_n24186);
xnor_4 g21838(new_n24174, new_n24170_1, new_n24187);
not_8  g21839(new_n24187, new_n24188);
nand_5 g21840(new_n24188, new_n24186, new_n24189);
xnor_4 g21841(new_n24187, new_n24186, new_n24190);
not_8  g21842(new_n20368, new_n24191);
nand_5 g21843(new_n20375, new_n24191, new_n24192);
nand_5 g21844(new_n20380, new_n20376, new_n24193);
nand_5 g21845(new_n24193, new_n24192, new_n24194);
nand_5 g21846(new_n24194, new_n24190, new_n24195);
nand_5 g21847(new_n24195, new_n24189, new_n24196_1);
nand_5 g21848(new_n24196_1, new_n24185, new_n24197);
nand_5 g21849(new_n24197, new_n24184, new_n24198);
xnor_4 g21850(new_n24198, new_n24180, n11063);
xnor_4 g21851(new_n21710, new_n21700, n11078);
xnor_4 g21852(new_n22409, new_n22396, n11080);
xnor_4 g21853(new_n14735, new_n14721, n11094);
xnor_4 g21854(new_n23836, new_n23835, n11101);
xnor_4 g21855(new_n22489_1, new_n15348, new_n24204);
xnor_4 g21856(new_n24204, new_n22492_1, n11103);
xnor_4 g21857(new_n6936, new_n6906, n11120);
xnor_4 g21858(new_n5275, new_n5271, n11127);
xnor_4 g21859(new_n15967_1, new_n15966, n11132);
xnor_4 g21860(new_n11898_1, new_n11851, n11134);
xnor_4 g21861(new_n3859, new_n3857, n11138);
xnor_4 g21862(new_n11152, new_n11136, n11182);
xnor_4 g21863(new_n14745, new_n14700, n11234);
xnor_4 g21864(new_n23128, new_n19818, new_n24213);
not_8  g21865(new_n19823, new_n24214);
nand_5 g21866(new_n22764_1, new_n24214, new_n24215);
nand_5 g21867(new_n22789, new_n22765, new_n24216);
nand_5 g21868(new_n24216, new_n24215, new_n24217);
xnor_4 g21869(new_n24217, new_n24213, n11245);
xnor_4 g21870(new_n9191_1, new_n9174, n11261);
xnor_4 g21871(new_n24196_1, new_n24185, n11275);
not_8  g21872(new_n14424, new_n24221);
nand_5 g21873(new_n24221, new_n14352, n11290);
xnor_4 g21874(new_n10011, new_n10008, n11313);
xnor_4 g21875(new_n17896, new_n17294, new_n24224);
xnor_4 g21876(new_n24224, new_n17911_1, n11325);
xnor_4 g21877(new_n14793, new_n14792, n11326);
xnor_4 g21878(new_n18156, new_n18120, n11330);
xnor_4 g21879(new_n11892, new_n11863, n11347);
xnor_4 g21880(new_n23909, new_n23901, n11348);
xnor_4 g21881(new_n16084, new_n16076, n11352);
or_5   g21882(new_n8719, n3324, new_n24231);
xnor_4 g21883(n22442, n3324, new_n24232);
or_5   g21884(n17911, new_n7404, new_n24233);
or_5   g21885(n21997, new_n7408_1, new_n24234);
nand_5 g21886(new_n18376, new_n18363, new_n24235);
nand_5 g21887(new_n24235, new_n24234, new_n24236);
xnor_4 g21888(n17911, n468, new_n24237);
nand_5 g21889(new_n24237, new_n24236, new_n24238);
nand_5 g21890(new_n24238, new_n24233, new_n24239);
nand_5 g21891(new_n24239, new_n24232, new_n24240);
nand_5 g21892(new_n24240, new_n24231, new_n24241);
not_8  g21893(new_n24241, new_n24242);
nor_5  g21894(new_n18932, new_n18925, new_n24243);
nor_5  g21895(new_n24243, new_n8140, new_n24244);
nand_5 g21896(new_n18932, new_n18925, new_n24245);
nand_5 g21897(new_n24245, new_n8140, new_n24246);
not_8  g21898(new_n24246, new_n24247);
nor_5  g21899(new_n24247, new_n24244, new_n24248);
xnor_4 g21900(new_n24248, new_n24242, new_n24249);
nand_5 g21901(new_n24242, new_n18934, new_n24250);
not_8  g21902(new_n18934, new_n24251);
nand_5 g21903(new_n24241, new_n24251, new_n24252);
xnor_4 g21904(new_n24239, new_n24232, new_n24253);
nand_5 g21905(new_n24253, new_n18936, new_n24254);
not_8  g21906(new_n24254, new_n24255);
xnor_4 g21907(new_n24253, new_n18936, new_n24256);
xnor_4 g21908(new_n24237, new_n24236, new_n24257);
nor_5  g21909(new_n24257, new_n18940_1, new_n24258_1);
not_8  g21910(new_n24258_1, new_n24259);
xnor_4 g21911(new_n24257, new_n18939, new_n24260_1);
nor_5  g21912(new_n18377_1, new_n18943, new_n24261);
not_8  g21913(new_n24261, new_n24262);
nand_5 g21914(new_n18389, new_n18378, new_n24263);
nand_5 g21915(new_n24263, new_n24262, new_n24264);
nand_5 g21916(new_n24264, new_n24260_1, new_n24265);
nand_5 g21917(new_n24265, new_n24259, new_n24266);
nor_5  g21918(new_n24266, new_n24256, new_n24267);
nor_5  g21919(new_n24267, new_n24255, new_n24268);
nand_5 g21920(new_n24268, new_n24252, new_n24269);
nand_5 g21921(new_n24269, new_n24250, new_n24270);
xnor_4 g21922(new_n24270, new_n24249, n11375);
not_8  g21923(new_n7592, new_n24272);
xnor_4 g21924(new_n13325, new_n24272, n11379);
or_5   g21925(new_n16503, n2570, new_n24274);
nand_5 g21926(new_n17541, new_n17511, new_n24275);
nand_5 g21927(new_n24275, new_n24274, new_n24276);
xnor_4 g21928(new_n24276, new_n12757, new_n24277);
nand_5 g21929(new_n17542, new_n12702_1, new_n24278_1);
nand_5 g21930(new_n17580, new_n17543, new_n24279);
nand_5 g21931(new_n24279, new_n24278_1, new_n24280);
xnor_4 g21932(new_n24280, new_n24277, new_n24281);
xnor_4 g21933(new_n24281, new_n6684_1, new_n24282);
not_8  g21934(new_n17581, new_n24283);
nand_5 g21935(new_n24283, new_n6688, new_n24284);
nand_5 g21936(new_n17620, new_n17582, new_n24285);
nand_5 g21937(new_n24285, new_n24284, new_n24286);
xnor_4 g21938(new_n24286, new_n24282, n11386);
xnor_4 g21939(new_n20543, new_n20529, n11391);
xnor_4 g21940(new_n22749, new_n22748, n11398);
xnor_4 g21941(new_n13650, new_n13649, n11403);
xnor_4 g21942(new_n13040, new_n13033, n11419);
xnor_4 g21943(new_n20351, new_n20333_1, n11439);
xnor_4 g21944(n7569, new_n17368, new_n24293);
nor_5  g21945(n19033, n17037, new_n24294);
xnor_4 g21946(n19033, new_n12174, new_n24295);
not_8  g21947(new_n24295, new_n24296);
nor_5  g21948(n5386, n655, new_n24297_1);
xnor_4 g21949(n5386, new_n17380, new_n24298);
not_8  g21950(new_n24298, new_n24299);
nor_5  g21951(n26191, n18145, new_n24300);
xnor_4 g21952(n26191, new_n17370, new_n24301);
not_8  g21953(new_n24301, new_n24302);
nor_5  g21954(n26512, n10712, new_n24303);
xnor_4 g21955(n26512, new_n16658, new_n24304);
not_8  g21956(new_n24304, new_n24305);
nor_5  g21957(n25126, n19575, new_n24306);
xnor_4 g21958(n25126, new_n12176, new_n24307_1);
not_8  g21959(new_n24307_1, new_n24308);
nand_5 g21960(n19608, n15378, new_n24309);
nor_5  g21961(n19608, n15378, new_n24310);
not_8  g21962(new_n24310, new_n24311);
nor_5  g21963(n17095, n1689, new_n24312);
not_8  g21964(new_n24043, new_n24313);
nor_5  g21965(new_n24049, new_n24313, new_n24314);
nor_5  g21966(new_n24314, new_n24312, new_n24315);
nand_5 g21967(new_n24315, new_n24311, new_n24316);
nand_5 g21968(new_n24316, new_n24309, new_n24317);
nor_5  g21969(new_n24317, new_n24308, new_n24318);
nor_5  g21970(new_n24318, new_n24306, new_n24319_1);
nor_5  g21971(new_n24319_1, new_n24305, new_n24320);
nor_5  g21972(new_n24320, new_n24303, new_n24321);
nor_5  g21973(new_n24321, new_n24302, new_n24322);
nor_5  g21974(new_n24322, new_n24300, new_n24323_1);
nor_5  g21975(new_n24323_1, new_n24299, new_n24324);
nor_5  g21976(new_n24324, new_n24297_1, new_n24325);
nor_5  g21977(new_n24325, new_n24296, new_n24326);
nor_5  g21978(new_n24326, new_n24294, new_n24327_1);
xnor_4 g21979(new_n24327_1, new_n24293, new_n24328);
nor_5  g21980(new_n24328, n10514, new_n24329);
xnor_4 g21981(new_n24328, new_n22097, new_n24330);
not_8  g21982(new_n24330, new_n24331);
xnor_4 g21983(new_n24325, new_n24295, new_n24332);
nand_5 g21984(new_n24332, n18649, new_n24333);
xnor_4 g21985(new_n24332, n18649, new_n24334);
not_8  g21986(new_n24334, new_n24335);
xnor_4 g21987(new_n24323_1, new_n24298, new_n24336);
nand_5 g21988(new_n24336, n6218, new_n24337);
xnor_4 g21989(new_n24336, new_n12116, new_n24338);
xnor_4 g21990(new_n24321, new_n24301, new_n24339);
nand_5 g21991(new_n24339, n20470, new_n24340);
xnor_4 g21992(new_n24339, n20470, new_n24341);
not_8  g21993(new_n24341, new_n24342_1);
xnor_4 g21994(new_n24319_1, new_n24304, new_n24343);
nand_5 g21995(new_n24343, n21222, new_n24344);
xnor_4 g21996(new_n24343, new_n11623, new_n24345_1);
xnor_4 g21997(new_n24317, new_n24307_1, new_n24346);
nand_5 g21998(new_n24346, n9832, new_n24347_1);
xnor_4 g21999(new_n24346, n9832, new_n24348);
not_8  g22000(new_n24348, new_n24349);
xnor_4 g22001(n19608, new_n10171, new_n24350);
xnor_4 g22002(new_n24350, new_n24315, new_n24351);
nor_5  g22003(new_n24351, n1558, new_n24352);
xnor_4 g22004(new_n24351, n1558, new_n24353);
nor_5  g22005(new_n24050, n21749, new_n24354);
nor_5  g22006(new_n24058, new_n24051, new_n24355);
nor_5  g22007(new_n24355, new_n24354, new_n24356);
nor_5  g22008(new_n24356, new_n24353, new_n24357);
nor_5  g22009(new_n24357, new_n24352, new_n24358);
nand_5 g22010(new_n24358, new_n24349, new_n24359);
nand_5 g22011(new_n24359, new_n24347_1, new_n24360);
nand_5 g22012(new_n24360, new_n24345_1, new_n24361);
nand_5 g22013(new_n24361, new_n24344, new_n24362);
nand_5 g22014(new_n24362, new_n24342_1, new_n24363);
nand_5 g22015(new_n24363, new_n24340, new_n24364);
nand_5 g22016(new_n24364, new_n24338, new_n24365);
nand_5 g22017(new_n24365, new_n24337, new_n24366);
nand_5 g22018(new_n24366, new_n24335, new_n24367);
nand_5 g22019(new_n24367, new_n24333, new_n24368);
nor_5  g22020(new_n24368, new_n24331, new_n24369);
nor_5  g22021(new_n24369, new_n24329, new_n24370);
or_5   g22022(n7569, n2570, new_n24371);
not_8  g22023(new_n24327_1, new_n24372);
nand_5 g22024(new_n24372, new_n24293, new_n24373_1);
nand_5 g22025(new_n24373_1, new_n24371, new_n24374_1);
xnor_4 g22026(new_n24374_1, new_n24370, new_n24375);
nand_5 g22027(new_n24160_1, new_n6645, new_n24376);
nor_5  g22028(new_n24376, n6105, new_n24377);
xnor_4 g22029(new_n24377, new_n11840, new_n24378);
xnor_4 g22030(new_n24376, new_n6641, new_n24379);
not_8  g22031(new_n24379, new_n24380);
nand_5 g22032(new_n24380, new_n9273, new_n24381);
xnor_4 g22033(new_n24379, new_n9273, new_n24382);
not_8  g22034(new_n24161, new_n24383);
nand_5 g22035(new_n24383, new_n9340, new_n24384);
nand_5 g22036(new_n24178, new_n24162, new_n24385);
nand_5 g22037(new_n24385, new_n24384, new_n24386);
nand_5 g22038(new_n24386, new_n24382, new_n24387);
nand_5 g22039(new_n24387, new_n24381, new_n24388);
xnor_4 g22040(new_n24388, new_n24378, new_n24389);
xnor_4 g22041(new_n24389, new_n24375, new_n24390);
xnor_4 g22042(new_n24368, new_n24330, new_n24391);
not_8  g22043(new_n24391, new_n24392);
xnor_4 g22044(new_n24386, new_n24382, new_n24393);
not_8  g22045(new_n24393, new_n24394);
nand_5 g22046(new_n24394, new_n24392, new_n24395);
xnor_4 g22047(new_n24394, new_n24391, new_n24396);
not_8  g22048(new_n24179, new_n24397);
xnor_4 g22049(new_n24366, new_n24334, new_n24398);
nand_5 g22050(new_n24398, new_n24397, new_n24399);
xnor_4 g22051(new_n24398, new_n24179, new_n24400);
not_8  g22052(new_n24338, new_n24401);
xnor_4 g22053(new_n24364, new_n24401, new_n24402);
nand_5 g22054(new_n24402, new_n24183, new_n24403);
xnor_4 g22055(new_n24402, new_n24182, new_n24404);
xnor_4 g22056(new_n24362, new_n24341, new_n24405);
nand_5 g22057(new_n24405, new_n24188, new_n24406_1);
xnor_4 g22058(new_n24405, new_n24187, new_n24407);
xnor_4 g22059(new_n24360, new_n24345_1, new_n24408);
not_8  g22060(new_n24408, new_n24409);
nand_5 g22061(new_n24409, new_n20375, new_n24410);
xnor_4 g22062(new_n24408, new_n20375, new_n24411);
xnor_4 g22063(new_n24358, new_n24348, new_n24412);
nand_5 g22064(new_n24412, new_n20377, new_n24413);
xnor_4 g22065(new_n24412, new_n19606, new_n24414);
xnor_4 g22066(new_n24356, new_n24353, new_n24415_1);
not_8  g22067(new_n24415_1, new_n24416);
nor_5  g22068(new_n24416, new_n19626, new_n24417);
not_8  g22069(new_n24417, new_n24418);
nor_5  g22070(new_n24059, new_n19632, new_n24419);
nor_5  g22071(new_n24068, new_n24060, new_n24420);
nor_5  g22072(new_n24420, new_n24419, new_n24421_1);
xnor_4 g22073(new_n24415_1, new_n19626, new_n24422);
nand_5 g22074(new_n24422, new_n24421_1, new_n24423);
nand_5 g22075(new_n24423, new_n24418, new_n24424);
nand_5 g22076(new_n24424, new_n24414, new_n24425);
nand_5 g22077(new_n24425, new_n24413, new_n24426);
nand_5 g22078(new_n24426, new_n24411, new_n24427);
nand_5 g22079(new_n24427, new_n24410, new_n24428);
nand_5 g22080(new_n24428, new_n24407, new_n24429);
nand_5 g22081(new_n24429, new_n24406_1, new_n24430);
nand_5 g22082(new_n24430, new_n24404, new_n24431_1);
nand_5 g22083(new_n24431_1, new_n24403, new_n24432);
nand_5 g22084(new_n24432, new_n24400, new_n24433);
nand_5 g22085(new_n24433, new_n24399, new_n24434);
nand_5 g22086(new_n24434, new_n24396, new_n24435);
nand_5 g22087(new_n24435, new_n24395, new_n24436);
xnor_4 g22088(new_n24436, new_n24390, n11462);
xnor_4 g22089(new_n21716, new_n21688, n11470);
xnor_4 g22090(new_n16430, new_n16414, n11472);
xnor_4 g22091(new_n20173, new_n7766, new_n24440);
xnor_4 g22092(new_n24440, new_n20189, n11496);
xnor_4 g22093(new_n21470, new_n21430, n11506);
xnor_4 g22094(new_n23310, new_n6011, new_n24443);
nand_5 g22095(new_n16797, new_n6017, new_n24444);
xnor_4 g22096(new_n16797, new_n6016, new_n24445);
nand_5 g22097(new_n11306, new_n6022_1, new_n24446);
xnor_4 g22098(new_n11306, new_n6021, new_n24447);
nand_5 g22099(new_n11331, new_n6028, new_n24448);
xnor_4 g22100(new_n5974, new_n5934, new_n24449);
xnor_4 g22101(new_n11331, new_n24449, new_n24450);
nand_5 g22102(new_n11335, new_n6035, new_n24451);
nand_5 g22103(new_n23986_1, new_n23968, new_n24452);
nand_5 g22104(new_n24452, new_n24451, new_n24453);
nand_5 g22105(new_n24453, new_n24450, new_n24454);
nand_5 g22106(new_n24454, new_n24448, new_n24455);
nand_5 g22107(new_n24455, new_n24447, new_n24456);
nand_5 g22108(new_n24456, new_n24446, new_n24457);
nand_5 g22109(new_n24457, new_n24445, new_n24458);
nand_5 g22110(new_n24458, new_n24444, new_n24459);
xnor_4 g22111(new_n24459, new_n24443, n11515);
xnor_4 g22112(new_n22419, new_n22385, n11538);
xnor_4 g22113(new_n19941_1, new_n19940, n11548);
xnor_4 g22114(new_n20223, new_n20216, n11564);
nor_5  g22115(new_n8719, n8856, new_n24464);
not_8  g22116(new_n23191, new_n24465);
nor_5  g22117(new_n23194, new_n24465, new_n24466);
nor_5  g22118(new_n24466, new_n24464, new_n24467);
not_8  g22119(new_n24467, new_n24468);
or_5   g22120(n3324, n2272, new_n24469);
nand_5 g22121(new_n23200_1, new_n23196, new_n24470);
nand_5 g22122(new_n24470, new_n24469, new_n24471);
and_5  g22123(new_n24471, new_n7966, new_n24472_1);
nor_5  g22124(new_n23201, new_n7960, new_n24473);
not_8  g22125(new_n24473, new_n24474);
nand_5 g22126(new_n23207, new_n23202, new_n24475);
nand_5 g22127(new_n24475, new_n24474, new_n24476_1);
xnor_4 g22128(new_n24471, new_n7965, new_n24477);
not_8  g22129(new_n24477, new_n24478);
nor_5  g22130(new_n24478, new_n24476_1, new_n24479);
nor_5  g22131(new_n24479, new_n24472_1, new_n24480);
xnor_4 g22132(new_n24480, new_n24468, new_n24481);
xnor_4 g22133(new_n24478, new_n24476_1, new_n24482);
nor_5  g22134(new_n24482, new_n24467, new_n24483_1);
xnor_4 g22135(new_n24482, new_n24467, new_n24484);
nand_5 g22136(new_n23209, new_n23195, new_n24485_1);
xnor_4 g22137(new_n23208, new_n23195, new_n24486);
nand_5 g22138(new_n23214, new_n24486, new_n24487);
nand_5 g22139(new_n24487, new_n24485_1, new_n24488);
nor_5  g22140(new_n24488, new_n24484, new_n24489);
nor_5  g22141(new_n24489, new_n24483_1, new_n24490);
xnor_4 g22142(new_n24490, new_n24481, n11591);
not_8  g22143(new_n8843, new_n24492);
nand_5 g22144(new_n24492, new_n8836, new_n24493);
not_8  g22145(new_n24493, new_n24494);
nand_5 g22146(new_n8856_1, new_n8844, new_n24495);
nor_5  g22147(new_n8856_1, new_n8844, new_n24496);
nor_5  g22148(new_n8915, new_n24496, new_n24497);
nor_5  g22149(new_n24497, new_n23988, new_n24498);
nand_5 g22150(new_n24498, new_n24495, new_n24499);
nor_5  g22151(new_n24499, new_n24494, n11607);
xnor_4 g22152(new_n19878, new_n19846, n11647);
xor_4  g22153(new_n24264, new_n24260_1, n11674);
xnor_4 g22154(new_n20890, new_n16452, new_n24503);
nor_5  g22155(new_n20902, new_n16452, new_n24504);
nor_5  g22156(new_n22751, new_n22738, new_n24505);
nor_5  g22157(new_n24505, new_n24504, new_n24506);
xnor_4 g22158(new_n24506, new_n24503, n11682);
xnor_4 g22159(new_n23426, new_n23413, n11710);
xnor_4 g22160(new_n14739, new_n14713, n11712);
xnor_4 g22161(new_n23071, new_n23057, n11724);
xnor_4 g22162(new_n19262, new_n19260, n11741);
xor_4  g22163(new_n18990, new_n3138, n11770);
xnor_4 g22164(new_n8902, new_n8901, n11771);
xnor_4 g22165(new_n20063, new_n20029, n11818);
xnor_4 g22166(new_n23980, new_n23973, n11837);
and_5  g22167(new_n17175, new_n3675, new_n24516);
xnor_4 g22168(new_n24516, n2743, new_n24517);
not_8  g22169(new_n24517, new_n24518);
nor_5  g22170(new_n24518, new_n6236, new_n24519);
xnor_4 g22171(new_n24517, new_n6236, new_n24520);
not_8  g22172(new_n24520, new_n24521);
not_8  g22173(new_n17176, new_n24522);
nor_5  g22174(new_n24522, new_n6240, new_n24523);
not_8  g22175(new_n17177, new_n24524);
nor_5  g22176(new_n17220, new_n24524, new_n24525);
nor_5  g22177(new_n24525, new_n24523, new_n24526);
nor_5  g22178(new_n24526, new_n24521, new_n24527);
nor_5  g22179(new_n24527, new_n24519, new_n24528);
and_5  g22180(new_n24516, new_n14355, new_n24529);
xnor_4 g22181(new_n24529, new_n14287, new_n24530);
xnor_4 g22182(new_n24530, new_n24528, new_n24531);
xnor_4 g22183(new_n24531, new_n23132, new_n24532);
xnor_4 g22184(new_n24526, new_n24520, new_n24533);
not_8  g22185(new_n24533, new_n24534);
nand_5 g22186(new_n24534, new_n22677, new_n24535);
xnor_4 g22187(new_n24533, new_n22677, new_n24536);
not_8  g22188(new_n17221, new_n24537);
nand_5 g22189(new_n17231, new_n24537, new_n24538);
nand_5 g22190(new_n17279, new_n17232_1, new_n24539);
nand_5 g22191(new_n24539, new_n24538, new_n24540);
nand_5 g22192(new_n24540, new_n24536, new_n24541);
nand_5 g22193(new_n24541, new_n24535, new_n24542);
xnor_4 g22194(new_n24542, new_n24532, n11842);
xnor_4 g22195(new_n16755, new_n16734, n11843);
xnor_4 g22196(new_n19648_1, new_n19629, n11905);
xnor_4 g22197(new_n12086, new_n12081, n11965);
xnor_4 g22198(new_n19531_1, new_n19527, n12000);
xor_4  g22199(new_n17363, new_n17359_1, n12003);
xnor_4 g22200(new_n17990, new_n17989, n12011);
xnor_4 g22201(new_n18543, new_n18527, n12072);
xor_4  g22202(new_n11387, new_n11386_1, n12131);
and_5  g22203(new_n17334, new_n17300, new_n24552);
nor_5  g22204(new_n24552, new_n17335, n12146);
xnor_4 g22205(new_n17607, new_n17604, n12157);
xnor_4 g22206(new_n10890, new_n10831, n12158);
xnor_4 g22207(new_n23516, new_n23494, n12179);
xnor_4 g22208(new_n6754, new_n6699, n12192);
xnor_4 g22209(new_n23911, new_n23898, n12223);
xnor_4 g22210(new_n10888, new_n10836, n12225);
xnor_4 g22211(new_n23984, new_n23970, n12228);
xnor_4 g22212(new_n14209, new_n10185, n12235);
xnor_4 g22213(new_n9642, new_n9612, n12302);
xnor_4 g22214(new_n17756, new_n17724, n12304);
xnor_4 g22215(n19196, n1742, new_n24564);
or_5   g22216(new_n12714, n4858, new_n24565);
xnor_4 g22217(n23586, n4858, new_n24566);
nor_5  g22218(new_n16517_1, n8244, new_n24567);
xnor_4 g22219(n21226, n8244, new_n24568);
nor_5  g22220(n9493, new_n6497, new_n24569);
not_8  g22221(new_n24569, new_n24570);
nor_5  g22222(n20036, new_n6831, new_n24571);
not_8  g22223(new_n20820, new_n24572);
nor_5  g22224(new_n20826_1, new_n24572, new_n24573);
nor_5  g22225(new_n24573, new_n24571, new_n24574);
xnor_4 g22226(n9493, n4426, new_n24575);
nand_5 g22227(new_n24575, new_n24574, new_n24576_1);
nand_5 g22228(new_n24576_1, new_n24570, new_n24577);
and_5  g22229(new_n24577, new_n24568, new_n24578);
nor_5  g22230(new_n24578, new_n24567, new_n24579_1);
not_8  g22231(new_n24579_1, new_n24580);
nand_5 g22232(new_n24580, new_n24566, new_n24581);
nand_5 g22233(new_n24581, new_n24565, new_n24582);
xnor_4 g22234(new_n24582, new_n24564, new_n24583);
xnor_4 g22235(new_n24583, new_n20774_1, new_n24584);
xnor_4 g22236(new_n24579_1, new_n24566, new_n24585);
not_8  g22237(new_n24585, new_n24586);
nand_5 g22238(new_n24586, new_n19241, new_n24587);
xnor_4 g22239(new_n24585, new_n19241, new_n24588);
not_8  g22240(new_n24568, new_n24589);
xnor_4 g22241(new_n24577, new_n24589, new_n24590);
not_8  g22242(new_n24590, new_n24591);
nand_5 g22243(new_n24591, new_n19245, new_n24592);
xnor_4 g22244(new_n24590, new_n19245, new_n24593);
xnor_4 g22245(new_n24575, new_n24574, new_n24594);
nand_5 g22246(new_n24594, new_n19249, new_n24595);
xnor_4 g22247(new_n24594, new_n19248, new_n24596);
nand_5 g22248(new_n20827, new_n19252, new_n24597);
nand_5 g22249(new_n20838, new_n20828, new_n24598);
nand_5 g22250(new_n24598, new_n24597, new_n24599);
nand_5 g22251(new_n24599, new_n24596, new_n24600);
nand_5 g22252(new_n24600, new_n24595, new_n24601);
nand_5 g22253(new_n24601, new_n24593, new_n24602_1);
nand_5 g22254(new_n24602_1, new_n24592, new_n24603);
nand_5 g22255(new_n24603, new_n24588, new_n24604_1);
nand_5 g22256(new_n24604_1, new_n24587, new_n24605);
xnor_4 g22257(new_n24605, new_n24584, n12324);
xnor_4 g22258(new_n22746, new_n22742, n12325);
xor_4  g22259(new_n11154, new_n11130, n12329);
xnor_4 g22260(new_n9189, new_n9188, n12330);
xnor_4 g22261(new_n6072, new_n6019, n12346);
xnor_4 g22262(new_n8077, new_n8052_1, n12349);
xnor_4 g22263(new_n20539, new_n20537, n12364);
not_8  g22264(new_n5997, new_n24613);
nor_5  g22265(new_n23396, new_n24613, new_n24614);
xnor_4 g22266(new_n23396, new_n5997, new_n24615);
not_8  g22267(new_n24615, new_n24616);
nand_5 g22268(new_n23397, new_n6002, new_n24617);
xnor_4 g22269(new_n23397, new_n6001, new_n24618_1);
nand_5 g22270(new_n23308, new_n6007, new_n24619);
xnor_4 g22271(new_n23308, new_n6006, new_n24620_1);
nand_5 g22272(new_n23310, new_n6012_1, new_n24621);
nand_5 g22273(new_n24459, new_n24443, new_n24622);
nand_5 g22274(new_n24622, new_n24621, new_n24623);
nand_5 g22275(new_n24623, new_n24620_1, new_n24624);
nand_5 g22276(new_n24624, new_n24619, new_n24625);
nand_5 g22277(new_n24625, new_n24618_1, new_n24626_1);
nand_5 g22278(new_n24626_1, new_n24617, new_n24627);
nor_5  g22279(new_n24627, new_n24616, new_n24628);
nor_5  g22280(new_n24628, new_n24614, n12383);
xnor_4 g22281(new_n9093, new_n9092, n12397);
xor_4  g22282(new_n18150, new_n18137, n12408);
nor_5  g22283(new_n20890, new_n16453, new_n24632);
not_8  g22284(new_n24503, new_n24633);
nor_5  g22285(new_n24506, new_n24633, new_n24634);
nor_5  g22286(new_n24634, new_n24632, n12449);
xnor_4 g22287(new_n22506, new_n22470_1, n12461);
nand_5 g22288(new_n22336, new_n12758, new_n24637);
nand_5 g22289(new_n24637, new_n18242, new_n24638_1);
not_8  g22290(new_n24637, new_n24639);
nand_5 g22291(new_n24639, new_n18241_1, new_n24640);
not_8  g22292(new_n22337, new_n24641);
nand_5 g22293(new_n24641, new_n18301_1, new_n24642);
nand_5 g22294(new_n22346, new_n22338, new_n24643);
nand_5 g22295(new_n24643, new_n24642, new_n24644);
nand_5 g22296(new_n24644, new_n24640, new_n24645);
nand_5 g22297(new_n24645, new_n24638_1, n12462);
not_8  g22298(new_n23528, new_n24647);
xnor_4 g22299(new_n24647, new_n23522, n12467);
nand_5 g22300(new_n23161, new_n16856, new_n24649);
nand_5 g22301(new_n16916, new_n16883, new_n24650);
nand_5 g22302(new_n24650, new_n24649, new_n24651);
nor_5  g22303(new_n24651, new_n23159, new_n24652);
not_8  g22304(new_n24652, new_n24653);
not_8  g22305(new_n24015, new_n24654);
nor_5  g22306(new_n17007, new_n16999, new_n24655);
nor_5  g22307(new_n24017, n13419, new_n24656);
nor_5  g22308(new_n24656, new_n24655, new_n24657);
nand_5 g22309(new_n24657, new_n24654, new_n24658);
xnor_4 g22310(new_n24651, new_n23158, new_n24659);
not_8  g22311(new_n24659, new_n24660);
xnor_4 g22312(new_n24657, new_n24015, new_n24661);
not_8  g22313(new_n24661, new_n24662);
nand_5 g22314(new_n24662, new_n24660, new_n24663);
xnor_4 g22315(new_n24661, new_n24660, new_n24664);
nor_5  g22316(new_n17009, new_n16918, new_n24665);
nor_5  g22317(new_n17056, new_n17010, new_n24666);
nor_5  g22318(new_n24666, new_n24665, new_n24667);
nand_5 g22319(new_n24667, new_n24664, new_n24668);
nand_5 g22320(new_n24668, new_n24663, new_n24669);
xnor_4 g22321(new_n24669, new_n24658, new_n24670);
xnor_4 g22322(new_n24670, new_n24653, n12469);
xnor_4 g22323(new_n11671, new_n11642, n12515);
or_5   g22324(new_n16503, n5140, new_n24673);
xnor_4 g22325(n10250, n5140, new_n24674);
or_5   g22326(new_n6481, n6204, new_n24675);
xnor_4 g22327(n7674, n6204, new_n24676);
or_5   g22328(new_n6484, n3349, new_n24677);
xnor_4 g22329(n6397, n3349, new_n24678);
or_5   g22330(new_n6487, n1742, new_n24679);
nand_5 g22331(new_n24582, new_n24564, new_n24680);
nand_5 g22332(new_n24680, new_n24679, new_n24681);
nand_5 g22333(new_n24681, new_n24678, new_n24682);
nand_5 g22334(new_n24682, new_n24677, new_n24683);
nand_5 g22335(new_n24683, new_n24676, new_n24684);
nand_5 g22336(new_n24684, new_n24675, new_n24685);
nand_5 g22337(new_n24685, new_n24674, new_n24686);
nand_5 g22338(new_n24686, new_n24673, new_n24687);
xnor_4 g22339(new_n24687, new_n23243, new_n24688);
nor_5  g22340(new_n24687, new_n23245, new_n24689);
not_8  g22341(new_n24687, new_n24690);
nor_5  g22342(new_n24690, new_n22081, new_n24691);
xnor_4 g22343(new_n24685, new_n24674, new_n24692);
nand_5 g22344(new_n24692, new_n22083, new_n24693);
not_8  g22345(new_n22083, new_n24694);
xnor_4 g22346(new_n24692, new_n24694, new_n24695);
xnor_4 g22347(new_n24683, new_n24676, new_n24696);
nand_5 g22348(new_n24696, new_n20766, new_n24697);
not_8  g22349(new_n20766, new_n24698);
xnor_4 g22350(new_n24696, new_n24698, new_n24699);
xnor_4 g22351(new_n24681, new_n24678, new_n24700);
nand_5 g22352(new_n24700, new_n20770, new_n24701);
xnor_4 g22353(new_n24700, new_n20769, new_n24702);
nand_5 g22354(new_n24583, new_n20775, new_n24703);
nand_5 g22355(new_n24605, new_n24584, new_n24704);
nand_5 g22356(new_n24704, new_n24703, new_n24705);
nand_5 g22357(new_n24705, new_n24702, new_n24706);
nand_5 g22358(new_n24706, new_n24701, new_n24707);
nand_5 g22359(new_n24707, new_n24699, new_n24708);
nand_5 g22360(new_n24708, new_n24697, new_n24709);
nand_5 g22361(new_n24709, new_n24695, new_n24710);
nand_5 g22362(new_n24710, new_n24693, new_n24711);
nor_5  g22363(new_n24711, new_n24691, new_n24712);
nor_5  g22364(new_n24712, new_n24689, new_n24713);
xnor_4 g22365(new_n24713, new_n24688, n12516);
xnor_4 g22366(new_n7866, new_n7852, n12540);
xnor_4 g22367(new_n12437, new_n12436, n12545);
xnor_4 g22368(new_n21714, new_n21692, n12552);
xnor_4 g22369(new_n8701, new_n8676, n12566);
xnor_4 g22370(new_n14162, new_n14142, n12569);
xnor_4 g22371(new_n6758, new_n6687, n12607);
xnor_4 g22372(new_n10694_1, new_n10620, n12620);
xnor_4 g22373(new_n3869_1, new_n3827, n12621);
xnor_4 g22374(new_n19452, new_n19450_1, n12654);
xnor_4 g22375(new_n20829, new_n15984, n12665);
xnor_4 g22376(new_n18189, new_n18177, n12670);
xnor_4 g22377(new_n8064, new_n2547_1, n12707);
xnor_4 g22378(new_n7595, new_n7584, n12725);
xnor_4 g22379(new_n17054, new_n17016, n12727);
xor_4  g22380(new_n10364, new_n10336, n12740);
xnor_4 g22381(new_n22047, new_n22046, n12742);
xnor_4 g22382(new_n22236, new_n2875, n12746);
xnor_4 g22383(new_n9820, new_n9818, n12756);
xnor_4 g22384(new_n7608, new_n7549, n12783);
xnor_4 g22385(new_n24687, new_n22081, new_n24734);
xnor_4 g22386(new_n24734, new_n24711, n12801);
xnor_4 g22387(new_n18876, new_n18873, n12812);
xnor_4 g22388(new_n17277, new_n17237, n12816);
nand_5 g22389(new_n18399, new_n19485, new_n24738);
nand_5 g22390(new_n19509, new_n19486, new_n24739);
nand_5 g22391(new_n24739, new_n24738, new_n24740);
nor_5  g22392(new_n24740, new_n22869, new_n24741);
not_8  g22393(new_n24741, new_n24742);
xnor_4 g22394(new_n24740, new_n22869, new_n24743);
nand_5 g22395(new_n24743, new_n24660, new_n24744);
xnor_4 g22396(new_n24743, new_n24659, new_n24745);
nand_5 g22397(new_n19510, new_n16918, new_n24746);
nand_5 g22398(new_n19539_1, new_n19511, new_n24747);
nand_5 g22399(new_n24747, new_n24746, new_n24748);
nand_5 g22400(new_n24748, new_n24745, new_n24749_1);
nand_5 g22401(new_n24749_1, new_n24744, new_n24750);
nand_5 g22402(new_n24750, new_n24742, new_n24751);
nand_5 g22403(new_n24751, new_n24653, new_n24752);
not_8  g22404(new_n24752, n12843);
xnor_4 g22405(new_n22285, new_n22284, n12864);
not_8  g22406(new_n19931, new_n24755);
nor_5  g22407(new_n23662, new_n5089, new_n24756);
nor_5  g22408(new_n23693, new_n23663_1, new_n24757);
nor_5  g22409(new_n24757, new_n24756, new_n24758_1);
or_5   g22410(n21784, n3740, new_n24759);
nand_5 g22411(new_n23661, new_n23638, new_n24760);
nand_5 g22412(new_n24760, new_n24759, new_n24761);
xnor_4 g22413(new_n24761, new_n5151, new_n24762);
not_8  g22414(new_n24762, new_n24763);
xnor_4 g22415(new_n24763, new_n24758_1, new_n24764);
nor_5  g22416(new_n24764, new_n24755, new_n24765);
not_8  g22417(new_n24765, new_n24766);
nor_5  g22418(new_n23694, new_n23637_1, new_n24767);
not_8  g22419(new_n24767, new_n24768_1);
xnor_4 g22420(new_n23694, new_n18612, new_n24769);
nand_5 g22421(new_n23732, new_n24769, new_n24770);
nand_5 g22422(new_n24770, new_n24768_1, new_n24771);
xnor_4 g22423(new_n24764, new_n19931, new_n24772);
nand_5 g22424(new_n24772, new_n24771, new_n24773);
nand_5 g22425(new_n24773, new_n24766, new_n24774);
nor_5  g22426(new_n24761, new_n15119, new_n24775);
and_5  g22427(new_n24761, new_n15119, new_n24776);
nor_5  g22428(new_n24776, new_n24758_1, new_n24777);
nor_5  g22429(new_n24777, new_n24775, new_n24778);
not_8  g22430(new_n24778, new_n24779);
nor_5  g22431(new_n24779, new_n24774, n12865);
xnor_4 g22432(new_n13743, new_n13720, n12870);
xnor_4 g22433(new_n22245, new_n22224, n12873);
not_8  g22434(new_n19724, new_n24783);
not_8  g22435(new_n23859, new_n24784_1);
nand_5 g22436(new_n24784_1, new_n24783, new_n24785);
xnor_4 g22437(new_n24784_1, new_n19724, new_n24786_1);
nand_5 g22438(new_n23861, new_n19818, new_n24787);
nand_5 g22439(new_n24217, new_n24213, new_n24788);
nand_5 g22440(new_n24788, new_n24787, new_n24789);
nand_5 g22441(new_n24789, new_n24786_1, new_n24790);
nand_5 g22442(new_n24790, new_n24785, n12904);
xnor_4 g22443(new_n11160, new_n11158, n12941);
xnor_4 g22444(new_n11961, new_n11953, n12942);
xnor_4 g22445(new_n6166, new_n6169, new_n24794);
xnor_4 g22446(new_n24794, new_n6172, n12978);
xnor_4 g22447(new_n10377, new_n8384, n12980);
xnor_4 g22448(new_n6921, new_n4935, n12985);
xnor_4 g22449(new_n15506_1, new_n15470_1, n12987);
or_5   g22450(n11220, new_n12514, new_n24799);
nand_5 g22451(new_n17836, new_n17820_1, new_n24800);
nand_5 g22452(new_n24800, new_n24799, new_n24801);
not_8  g22453(new_n24801, new_n24802);
xnor_4 g22454(new_n24802, new_n15778, new_n24803);
nor_5  g22455(new_n17837, new_n15818, new_n24804);
nor_5  g22456(new_n17858, new_n17838, new_n24805);
nor_5  g22457(new_n24805, new_n24804, new_n24806);
xnor_4 g22458(new_n24806, new_n24803, n12992);
or_5   g22459(new_n23452, n6659, new_n24808);
or_5   g22460(new_n22428, n23250, new_n24809);
nand_5 g22461(new_n22464, new_n22429, new_n24810);
nand_5 g22462(new_n24810, new_n24809, new_n24811);
or_5   g22463(new_n23454, new_n19485, new_n24812);
nand_5 g22464(new_n24812, new_n24811, new_n24813);
nand_5 g22465(new_n24813, new_n24808, new_n24814);
nand_5 g22466(new_n24814, new_n23450_1, new_n24815);
xnor_4 g22467(new_n24815, new_n21093_1, new_n24816);
xnor_4 g22468(new_n23452, new_n19485, new_n24817);
xnor_4 g22469(new_n24817, new_n24811, new_n24818);
nand_5 g22470(new_n24818, new_n21109, new_n24819);
nand_5 g22471(new_n22465, new_n15278, new_n24820);
nand_5 g22472(new_n22508, new_n22466, new_n24821);
nand_5 g22473(new_n24821, new_n24820, new_n24822);
xnor_4 g22474(new_n24818, new_n21108, new_n24823);
nand_5 g22475(new_n24823, new_n24822, new_n24824);
nand_5 g22476(new_n24824, new_n24819, new_n24825);
xnor_4 g22477(new_n24825, new_n24816, n13005);
xnor_4 g22478(new_n21213, new_n17698, n13043);
xnor_4 g22479(new_n18963, new_n18961, n13048);
xnor_4 g22480(new_n16381, new_n16380, n13054);
xnor_4 g22481(new_n19142, new_n19128, n13082);
xnor_4 g22482(new_n7600, new_n7570, n13096);
xnor_4 g22483(new_n19144_1, new_n19120, n13116);
xnor_4 g22484(new_n21230, new_n21187, n13122);
xnor_4 g22485(new_n6739, new_n6737, n13141);
xor_4  g22486(new_n21047, new_n21036, n13144);
xnor_4 g22487(new_n21720, new_n21680_1, n13168);
xnor_4 g22488(new_n22413, new_n22391, n13198);
xnor_4 g22489(new_n15500, new_n15479, n13199);
xnor_4 g22490(new_n15626, new_n15611, n13204);
xnor_4 g22491(new_n10880, new_n10850, n13209);
xnor_4 g22492(new_n20816, new_n20806, n13270);
xnor_4 g22493(new_n14036_1, new_n14013, n13273);
xnor_4 g22494(new_n23518, new_n23489, n13285);
xnor_4 g22495(new_n22860, new_n22837, n13338);
xnor_4 g22496(new_n8402, new_n8369, n13407);
xnor_4 g22497(new_n5710, new_n4450, new_n24846);
xnor_4 g22498(new_n24846, new_n17317, n13409);
xnor_4 g22499(new_n5726, new_n5689, n13456);
nand_5 g22500(new_n22825, new_n22096, new_n24849);
not_8  g22501(new_n24849, new_n24850);
nor_5  g22502(new_n22720, new_n23946, new_n24851);
nor_5  g22503(new_n23951, new_n23947, new_n24852);
nor_5  g22504(new_n24852, new_n24851, new_n24853_1);
not_8  g22505(new_n24853_1, new_n24854);
nor_5  g22506(new_n22704, new_n22095, new_n24855);
nor_5  g22507(new_n24855, new_n24854, new_n24856);
nand_5 g22508(new_n24856, new_n24850, new_n24857_1);
xnor_4 g22509(new_n22703, new_n22095, new_n24858);
xnor_4 g22510(new_n24858, new_n24853_1, new_n24859);
not_8  g22511(new_n24859, new_n24860);
nand_5 g22512(new_n24860, new_n21234, new_n24861);
xnor_4 g22513(new_n24859, new_n21234, new_n24862);
nor_5  g22514(new_n23952, new_n12231, new_n24863);
nor_5  g22515(new_n23956, new_n23953, new_n24864);
nor_5  g22516(new_n24864, new_n24863, new_n24865);
nand_5 g22517(new_n24865, new_n24862, new_n24866);
nand_5 g22518(new_n24866, new_n24861, new_n24867);
xnor_4 g22519(new_n22792, new_n22096, new_n24868);
not_8  g22520(new_n24868, new_n24869);
nor_5  g22521(new_n24869, new_n24854, new_n24870);
not_8  g22522(new_n24870, new_n24871);
not_8  g22523(new_n24856, new_n24872);
nand_5 g22524(new_n24869, new_n24872, new_n24873);
nand_5 g22525(new_n24873, new_n24871, new_n24874);
nand_5 g22526(new_n24874, new_n24867, new_n24875);
nand_5 g22527(new_n24875, new_n24857_1, n13457);
xnor_4 g22528(new_n12990, new_n12979, n13477);
xnor_4 g22529(new_n13337, new_n13336, n13484);
xnor_4 g22530(new_n21923, new_n21889, n13486);
xnor_4 g22531(new_n23410, new_n22891_1, new_n24880);
not_8  g22532(new_n24880, new_n24881);
nor_5  g22533(new_n23320, new_n18495, new_n24882);
nor_5  g22534(new_n23352, new_n23321, new_n24883);
nor_5  g22535(new_n24883, new_n24882, new_n24884);
xnor_4 g22536(new_n24884, new_n24881, n13487);
xnor_4 g22537(new_n5481, new_n5461, n13500);
xor_4  g22538(new_n4801, new_n4800, n13501);
xnor_4 g22539(new_n6746, new_n6721, n13506);
xnor_4 g22540(new_n6461, new_n6451, n13548);
xnor_4 g22541(new_n24428, new_n24407, n13551);
xnor_4 g22542(new_n5280, new_n5258, n13602);
xnor_4 g22543(new_n18597, new_n18584_1, n13626);
xnor_4 g22544(new_n8697, new_n8689, n13683);
xnor_4 g22545(new_n21472_1, new_n21426, n13710);
xnor_4 g22546(new_n21051, new_n21029, n13722);
xnor_4 g22547(new_n15115, new_n15052_1, new_n24896);
xnor_4 g22548(new_n24896, new_n15198, n13754);
xor_4  g22549(new_n2889, new_n2853_1, n13764);
xnor_4 g22550(new_n15351, new_n15348, new_n24899);
xnor_4 g22551(new_n24899, new_n15356, n13798);
xnor_4 g22552(new_n18601, new_n18579, n13835);
xnor_4 g22553(new_n16850, new_n16849, n13850);
xnor_4 g22554(new_n19129, new_n8242, n13922);
xnor_4 g22555(new_n20782, new_n20772, n13923);
xnor_4 g22556(new_n12442, new_n12441, n14004);
xnor_4 g22557(new_n12690, new_n12643, n14036);
xnor_4 g22558(new_n22946, new_n22932, n14059);
xor_4  g22559(new_n18387, new_n18384, n14081);
xnor_4 g22560(new_n20185, new_n20182, n14095);
xnor_4 g22561(new_n7095, new_n3488, n14107);
xnor_4 g22562(new_n9470, new_n9433, n14121);
xnor_4 g22563(new_n12943, new_n12942_1, n14126);
xnor_4 g22564(new_n21055, new_n21021, n14136);
nor_5  g22565(new_n24801, new_n15778, new_n24914);
not_8  g22566(new_n15778, new_n24915);
nor_5  g22567(new_n24802, new_n24915, new_n24916);
nor_5  g22568(new_n24806, new_n24916, new_n24917);
nor_5  g22569(new_n24917, new_n24914, new_n24918);
xnor_4 g22570(new_n24802, new_n23751, new_n24919);
xnor_4 g22571(new_n24919, new_n24918, n14147);
xnor_4 g22572(new_n22642, new_n22595, n14174);
xnor_4 g22573(new_n17616, new_n17590, n14190);
xnor_4 g22574(new_n5724, new_n5695, n14211);
xnor_4 g22575(new_n17811, new_n17807, n14222);
xnor_4 g22576(new_n14420, new_n14366, n14267);
xnor_4 g22577(new_n6062, new_n6048, n14271);
xnor_4 g22578(new_n10014, new_n10001, n14277);
xnor_4 g22579(new_n8897, new_n8896, n14294);
xnor_4 g22580(new_n24434, new_n24396, n14310);
xnor_4 g22581(new_n24453, new_n24450, n14326);
xnor_4 g22582(new_n13288, new_n13234, n14342);
xnor_4 g22583(new_n19646, new_n19634, n14353);
nand_5 g22584(new_n22928, new_n12467_1, new_n24933);
not_8  g22585(new_n22928, new_n24934_1);
nand_5 g22586(new_n24934_1, new_n9529, new_n24935);
nand_5 g22587(new_n22948, new_n22929, new_n24936);
nand_5 g22588(new_n24936, new_n24935, new_n24937_1);
nand_5 g22589(new_n24937_1, new_n24933, new_n24938);
nand_5 g22590(new_n24934_1, new_n12466, new_n24939);
nand_5 g22591(new_n24939, new_n24936, new_n24940);
nand_5 g22592(new_n24940, new_n24938, new_n24941);
not_8  g22593(new_n24941, n14364);
xor_4  g22594(new_n23420, new_n23417, n14375);
xnor_4 g22595(new_n23920, new_n23886, n14412);
not_8  g22596(new_n12391, new_n24945);
nor_5  g22597(new_n18826, new_n6570, new_n24946);
not_8  g22598(new_n24946, new_n24947);
nor_5  g22599(new_n18856, new_n24947, new_n24948);
xnor_4 g22600(new_n24948, new_n24945, new_n24949);
not_8  g22601(new_n18857, new_n24950);
nand_5 g22602(new_n24950, new_n12392, new_n24951);
nand_5 g22603(new_n18884, new_n18858_1, new_n24952);
nand_5 g22604(new_n24952, new_n24951, new_n24953);
xnor_4 g22605(new_n24953, new_n24949, n14414);
xnor_4 g22606(new_n16596_1, new_n16594, n14457);
xnor_4 g22607(new_n5284, new_n5246, n14464);
xnor_4 g22608(new_n11669, new_n11647_1, n14471);
nor_5  g22609(new_n21083, new_n8855, new_n24958);
not_8  g22610(new_n24958, new_n24959);
nand_5 g22611(new_n21092, new_n21084, new_n24960);
nand_5 g22612(new_n24960, new_n24959, new_n24961);
xnor_4 g22613(new_n24961, new_n24815, new_n24962);
not_8  g22614(new_n21093_1, new_n24963);
not_8  g22615(new_n24815, new_n24964);
nand_5 g22616(new_n24964, new_n24963, new_n24965);
nand_5 g22617(new_n24815, new_n21093_1, new_n24966);
nand_5 g22618(new_n24825, new_n24966, new_n24967);
nand_5 g22619(new_n24967, new_n24965, new_n24968);
xnor_4 g22620(new_n24968, new_n24962, n14475);
xnor_4 g22621(new_n13276, new_n13275, n14541);
not_8  g22622(new_n23177, new_n24971);
nand_5 g22623(new_n24971, new_n23172, new_n24972);
nand_5 g22624(new_n23186, new_n23178, new_n24973);
nand_5 g22625(new_n24973, new_n24972, n14546);
xnor_4 g22626(new_n11881, new_n11879, n14547);
xnor_4 g22627(new_n13659, new_n13638, n14593);
xnor_4 g22628(new_n10018_1, new_n9989, n14636);
xnor_4 g22629(new_n24603, new_n24588, n14701);
xnor_4 g22630(new_n13044_1, new_n13031, n14734);
xnor_4 g22631(new_n7606, new_n7554, n14746);
xnor_4 g22632(new_n10355, new_n10353, n14763);
xnor_4 g22633(new_n24134, new_n24126, n14772);
xnor_4 g22634(new_n23424, new_n23422, n14801);
xnor_4 g22635(new_n22992, new_n22974, n14819);
xnor_4 g22636(new_n15635, new_n15595, n14827);
xnor_4 g22637(new_n22344, new_n22341_1, n14839);
xnor_4 g22638(new_n18591, new_n18589, n14849);
nand_5 g22639(new_n22202, new_n15580, new_n24988);
nand_5 g22640(new_n22260, new_n22203, new_n24989);
nand_5 g22641(new_n24989, new_n24988, new_n24990);
nand_5 g22642(new_n24990, new_n22197, new_n24991);
not_8  g22643(new_n24991, n14891);
xnor_4 g22644(new_n6883, new_n4971, n14931);
and_5  g22645(new_n24948, new_n24945, new_n24994);
nand_5 g22646(new_n24953, new_n24994, new_n24995);
nor_5  g22647(new_n24948, new_n24945, new_n24996);
not_8  g22648(new_n24953, new_n24997);
nand_5 g22649(new_n24997, new_n24996, new_n24998_1);
nand_5 g22650(new_n24998_1, new_n24995, n14944);
xnor_4 g22651(new_n19640, new_n9481, n14977);
xnor_4 g22652(new_n13667, new_n13616, n14989);
xnor_4 g22653(new_n11555, new_n11546, n15002);
xnor_4 g22654(new_n23978, new_n6059, n15004);
xnor_4 g22655(new_n9646_1, new_n9599, n15011);
xnor_4 g22656(new_n24030, new_n3306_1, new_n25005);
xnor_4 g22657(new_n24036, new_n25005, n15019);
not_8  g22658(new_n16354, new_n25007);
nand_5 g22659(new_n16363, new_n25007, new_n25008);
nand_5 g22660(new_n16387, new_n16364, new_n25009);
nand_5 g22661(new_n25009, new_n25008, n15031);
xnor_4 g22662(new_n19131, new_n19129, n15033);
xnor_4 g22663(new_n12805, new_n7637, n15052);
xnor_4 g22664(new_n20950, new_n20939, n15082);
xnor_4 g22665(new_n8699, new_n8682, n15094);
not_8  g22666(new_n12498, new_n25015);
xnor_4 g22667(new_n12503, new_n25015, n15118);
xnor_4 g22668(new_n24789, new_n24786_1, n15128);
xnor_4 g22669(new_n20067, new_n20021, n15139);
xnor_4 g22670(new_n17901, new_n17896, new_n25019);
xnor_4 g22671(new_n25019, new_n17913, n15145);
xnor_4 g22672(new_n15854, new_n15823, n15165);
xnor_4 g22673(new_n16296, new_n5347, n15176);
xor_4  g22674(new_n21708, new_n21707, n15180);
xnor_4 g22675(new_n17336, new_n17297, n15205);
xnor_4 g22676(new_n5717, new_n4453, n15230);
xnor_4 g22677(new_n18185, new_n18183, n15255);
xnor_4 g22678(new_n10368, new_n10323, n15275);
xnor_4 g22679(new_n14935, new_n14932, n15300);
nor_5  g22680(new_n24529, new_n14286, new_n25029);
nand_5 g22681(new_n25029, new_n24528, new_n25030);
not_8  g22682(new_n24528, new_n25031);
nand_5 g22683(new_n24529, new_n14286, new_n25032_1);
not_8  g22684(new_n25032_1, new_n25033);
nand_5 g22685(new_n25033, new_n25031, new_n25034);
nand_5 g22686(new_n25034, new_n25030, new_n25035);
xnor_4 g22687(new_n25035, new_n23172, new_n25036);
nand_5 g22688(new_n24531, new_n23133, new_n25037);
nand_5 g22689(new_n24542, new_n24532, new_n25038);
nand_5 g22690(new_n25038, new_n25037, new_n25039);
xnor_4 g22691(new_n25039, new_n25036, n15307);
xnor_4 g22692(new_n21474, new_n21422, n15327);
xnor_4 g22693(new_n21460, new_n21450, n15345);
xnor_4 g22694(new_n13657, new_n13644, n15353);
xnor_4 g22695(new_n24627, new_n24615, n15366);
xnor_4 g22696(new_n24779, new_n24774, n15382);
xnor_4 g22697(new_n9826, new_n9806, n15407);
xnor_4 g22698(new_n16216, new_n14493, n15428);
nand_5 g22699(new_n24374_1, new_n24370, new_n25048);
not_8  g22700(new_n24375, new_n25049);
nand_5 g22701(new_n24389, new_n25049, new_n25050);
nand_5 g22702(new_n24436, new_n24390, new_n25051);
nand_5 g22703(new_n25051, new_n25050, new_n25052);
nand_5 g22704(new_n25052, new_n25048, new_n25053);
not_8  g22705(new_n24377, new_n25054);
nand_5 g22706(new_n25054, new_n11840, new_n25055);
not_8  g22707(new_n25055, new_n25056);
nand_5 g22708(new_n24388, new_n25056, new_n25057);
not_8  g22709(new_n25057, new_n25058);
nand_5 g22710(new_n25058, new_n25048, new_n25059);
nand_5 g22711(new_n25059, new_n25051, new_n25060);
nand_5 g22712(new_n25060, new_n25053, new_n25061);
not_8  g22713(new_n25061, n15435);
not_8  g22714(new_n23988, new_n25063);
nor_5  g22715(new_n23995, new_n25063, new_n25064);
nand_5 g22716(new_n24007, new_n25064, new_n25065);
not_8  g22717(new_n23995, new_n25066);
nor_5  g22718(new_n25066, new_n23988, new_n25067);
xnor_4 g22719(new_n23997, new_n8857, new_n25068_1);
nor_5  g22720(new_n25068_1, new_n24003, new_n25069);
nor_5  g22721(new_n25069, new_n23998, new_n25070);
nand_5 g22722(new_n25070, new_n25067, new_n25071);
nand_5 g22723(new_n25071, new_n25065, n15438);
xnor_4 g22724(new_n24430, new_n24404, n15465);
xnor_4 g22725(new_n9091, new_n7023, n15467);
xnor_4 g22726(new_n8412, new_n8340, n15470);
xnor_4 g22727(new_n15639, new_n15589, n15477);
xnor_4 g22728(new_n24707, new_n24699, n15481);
xnor_4 g22729(new_n16082, new_n16079, n15496);
xnor_4 g22730(new_n12957, new_n12918, n15501);
xnor_4 g22731(new_n20187_1, new_n20179_1, n15555);
xnor_4 g22732(new_n22787_1, new_n22769, n15558);
nand_5 g22733(new_n23171, new_n24784_1, new_n25082);
nand_5 g22734(new_n23864, new_n23860, new_n25083_1);
nand_5 g22735(new_n25083_1, new_n25082, n15559);
not_8  g22736(new_n24075, new_n25085);
or_5   g22737(n23895, new_n3384, new_n25086);
nand_5 g22738(new_n21742, new_n21727, new_n25087);
nand_5 g22739(new_n25087, new_n25086, new_n25088);
nor_5  g22740(new_n25088, new_n25085, new_n25089);
nor_5  g22741(new_n21792, new_n21743, new_n25090);
not_8  g22742(new_n25090, new_n25091);
not_8  g22743(new_n21793, new_n25092);
nand_5 g22744(new_n21822, new_n25092, new_n25093);
nand_5 g22745(new_n25093, new_n25091, new_n25094_1);
nand_5 g22746(new_n25088, new_n23165, new_n25095);
nand_5 g22747(new_n25095, new_n25094_1, new_n25096);
not_8  g22748(new_n25096, new_n25097_1);
nand_5 g22749(new_n25097_1, new_n25085, new_n25098);
not_8  g22750(new_n25088, new_n25099);
nand_5 g22751(new_n25099, new_n23165, new_n25100);
nand_5 g22752(new_n25100, new_n25096, new_n25101);
nand_5 g22753(new_n25101, new_n25098, new_n25102);
nor_5  g22754(new_n25102, new_n25089, n15570);
xnor_4 g22755(new_n13294, new_n13219, n15573);
xnor_4 g22756(new_n12454, new_n12452, n15588);
xnor_4 g22757(new_n22988, new_n22980, n15590);
xnor_4 g22758(new_n23599, new_n23588_1, n15598);
xnor_4 g22759(new_n10021_1, new_n9983, n15614);
xnor_4 g22760(new_n24138, new_n24118, n15662);
xnor_4 g22761(new_n3509, new_n3469, n15716);
xnor_4 g22762(new_n15508_1, new_n15467_1, n15749);
xnor_4 g22763(new_n20091, new_n20085, n15762);
xnor_4 g22764(new_n8386, new_n8384, n15793);
xnor_4 g22765(new_n23914, new_n23895_1, n15812);
xnor_4 g22766(new_n13290, new_n13229, n15815);
xnor_4 g22767(new_n8894, new_n8893, n15816);
xnor_4 g22768(new_n12813, new_n12796, n15831);
xnor_4 g22769(new_n10217, new_n10215, n15846);
xnor_4 g22770(new_n8954, new_n8953, n15859);
not_8  g22771(new_n23227, new_n25120_1);
nor_5  g22772(new_n8574, new_n4548, new_n25121);
not_8  g22773(new_n21308, new_n25122);
nor_5  g22774(new_n21323, new_n25122, new_n25123);
nor_5  g22775(new_n25123, new_n25121, new_n25124);
nor_5  g22776(new_n25124, new_n8572, new_n25125);
xnor_4 g22777(new_n25125, new_n25120_1, new_n25126_1);
xnor_4 g22778(new_n25124, new_n8636, new_n25127);
not_8  g22779(new_n25127, new_n25128);
nand_5 g22780(new_n25128, new_n21671, new_n25129);
not_8  g22781(new_n21324, new_n25130);
nand_5 g22782(new_n25130, new_n21307, new_n25131);
nand_5 g22783(new_n21353, new_n21325, new_n25132);
nand_5 g22784(new_n25132, new_n25131, new_n25133_1);
xnor_4 g22785(new_n25127, new_n21671, new_n25134);
nand_5 g22786(new_n25134, new_n25133_1, new_n25135);
nand_5 g22787(new_n25135, new_n25129, new_n25136);
xnor_4 g22788(new_n25136, new_n25126_1, n15869);
xnor_4 g22789(new_n20234, new_n20207, n15885);
not_8  g22790(new_n22591_1, new_n25139);
nor_5  g22791(new_n25139, new_n16624, new_n25140);
nand_5 g22792(new_n22644, new_n25140, new_n25141);
nand_5 g22793(new_n22643, new_n25139, new_n25142);
nand_5 g22794(new_n25142, new_n25141, n15889);
xnor_4 g22795(new_n20219, new_n14791, n15917);
xnor_4 g22796(new_n14785, new_n14784, n15922);
xor_4  g22797(new_n7586, new_n7585_1, n15947);
and_5  g22798(new_n20869_1, new_n7685, new_n25147);
not_8  g22799(new_n22265, new_n25148);
nor_5  g22800(new_n22276, new_n25148, new_n25149);
nor_5  g22801(new_n25149, new_n25147, new_n25150);
xnor_4 g22802(new_n25150, new_n20898, new_n25151);
nand_5 g22803(new_n22277, new_n20899, new_n25152);
nand_5 g22804(new_n22287, new_n22278, new_n25153);
nand_5 g22805(new_n25153, new_n25152, new_n25154);
xnor_4 g22806(new_n25154, new_n25151, n15956);
xnor_4 g22807(new_n14518, new_n14514, n15958);
not_8  g22808(new_n13011, new_n25157);
nor_5  g22809(new_n18222, new_n25157, new_n25158);
not_8  g22810(new_n18222, new_n25159);
nor_5  g22811(new_n25159, new_n18217, new_n25160);
nor_5  g22812(new_n25160, new_n25158, new_n25161);
nand_5 g22813(new_n18218, new_n13011, new_n25162);
not_8  g22814(new_n18219, new_n25163);
nand_5 g22815(new_n25163, new_n25162, new_n25164);
nor_5  g22816(new_n25164, new_n25161, n15986);
xnor_4 g22817(new_n24540, new_n24536, n16013);
not_8  g22818(new_n23374, new_n25167);
nand_5 g22819(new_n25167, new_n22277, new_n25168_1);
not_8  g22820(new_n22277, new_n25169);
nand_5 g22821(new_n23374, new_n25169, new_n25170);
nand_5 g22822(new_n23384, new_n25170, new_n25171);
nand_5 g22823(new_n25171, new_n25168_1, new_n25172);
xnor_4 g22824(new_n25150, new_n23374, new_n25173);
xnor_4 g22825(new_n25173, new_n25172, n16060);
nand_5 g22826(new_n17542, n25972, new_n25175);
xnor_4 g22827(new_n17542, new_n12752, new_n25176);
nand_5 g22828(new_n17544, n21915, new_n25177);
nand_5 g22829(new_n24156, new_n24145_1, new_n25178);
nand_5 g22830(new_n25178, new_n25177, new_n25179);
nand_5 g22831(new_n25179, new_n25176, new_n25180);
nand_5 g22832(new_n25180, new_n25175, new_n25181_1);
nand_5 g22833(new_n25181_1, new_n24276, new_n25182);
not_8  g22834(new_n24276, new_n25183);
xnor_4 g22835(new_n25181_1, new_n25183, new_n25184);
not_8  g22836(new_n25184, new_n25185);
nand_5 g22837(new_n25185, new_n24389, new_n25186);
xnor_4 g22838(new_n25184, new_n24389, new_n25187);
xnor_4 g22839(new_n25179, new_n25176, new_n25188);
nand_5 g22840(new_n25188, new_n24394, new_n25189);
xnor_4 g22841(new_n25188, new_n24393, new_n25190);
nand_5 g22842(new_n24397, new_n24157, new_n25191);
nand_5 g22843(new_n24198, new_n24180, new_n25192);
nand_5 g22844(new_n25192, new_n25191, new_n25193);
nand_5 g22845(new_n25193, new_n25190, new_n25194);
nand_5 g22846(new_n25194, new_n25189, new_n25195);
nand_5 g22847(new_n25195, new_n25187, new_n25196);
nand_5 g22848(new_n25196, new_n25186, new_n25197);
xnor_4 g22849(new_n25197, new_n25182, new_n25198);
xnor_4 g22850(new_n25198, new_n25057, n16062);
xnor_4 g22851(new_n24625, new_n24618_1, n16068);
xnor_4 g22852(new_n24865, new_n24862, n16080);
nand_5 g22853(new_n24281, new_n6685, new_n25202);
nand_5 g22854(new_n24286, new_n24282, new_n25203);
nand_5 g22855(new_n25203, new_n25202, new_n25204);
nand_5 g22856(new_n24276, new_n12757, new_n25205);
not_8  g22857(new_n24277, new_n25206);
nand_5 g22858(new_n24280, new_n25206, new_n25207);
nand_5 g22859(new_n25207, new_n25205, new_n25208);
xnor_4 g22860(new_n25208, new_n25204, n16098);
xnor_4 g22861(new_n18816, new_n18804, n16110);
xnor_4 g22862(new_n16229, new_n16198, n16142);
xnor_4 g22863(new_n17750, new_n17735_1, n16185);
xnor_4 g22864(new_n13334, new_n13314, n16196);
xnor_4 g22865(new_n22302, new_n22301, n16206);
xor_4  g22866(new_n22377, new_n22374, n16215);
xnor_4 g22867(new_n20349_1, new_n20339, n16218);
xnor_4 g22868(new_n12670_1, new_n4079, n16219);
xnor_4 g22869(new_n7340, new_n7337, n16230);
xor_4  g22870(new_n8951, new_n8942, n16243);
xnor_4 g22871(new_n18541, new_n18530, n16275);
xnor_4 g22872(new_n10884, new_n10882, n16279);
nand_5 g22873(new_n21871, new_n19011, new_n25222);
nand_5 g22874(new_n21933, new_n21872, new_n25223);
nand_5 g22875(new_n25223, new_n25222, n16322);
xnor_4 g22876(new_n18549, new_n18510, n16327);
xnor_4 g22877(new_n22783, new_n22774, n16350);
xnor_4 g22878(new_n7024, new_n7023, n16367);
xnor_4 g22879(new_n20456, new_n20455_1, n16379);
xnor_4 g22880(new_n21464, new_n21442, n16398);
xnor_4 g22881(new_n14502, new_n14500, n16406);
xnor_4 g22882(new_n23601, new_n23583, n16407);
xnor_4 g22883(new_n25195, new_n25187, n16419);
xnor_4 g22884(new_n8911_1, new_n8864, n16424);
xnor_4 g22885(new_n14903, new_n14836, new_n25234);
xnor_4 g22886(new_n25234, new_n14948, n16428);
xnor_4 g22887(new_n12830, new_n12762, n16433);
xnor_4 g22888(new_n12826, new_n12770, n16440);
xnor_4 g22889(new_n18818, new_n18800, n16445);
xnor_4 g22890(new_n15193, new_n15128_1, n16460);
xnor_4 g22891(new_n21349_1, new_n21337, n16481);
nor_5  g22892(new_n21982, new_n11837_1, new_n25241);
nand_5 g22893(new_n15815_1, new_n11842_1, new_n25242);
nand_5 g22894(new_n21999, new_n21983, new_n25243);
nand_5 g22895(new_n25243, new_n25242, new_n25244_1);
xnor_4 g22896(new_n15815_1, new_n11837_1, new_n25245);
not_8  g22897(new_n25245, new_n25246);
nor_5  g22898(new_n25246, new_n25244_1, new_n25247);
nor_5  g22899(new_n25247, new_n25241, n16493);
xnor_4 g22900(new_n4987, new_n4956, n16506);
xnor_4 g22901(new_n13733, new_n13731, n16516);
xnor_4 g22902(new_n23722, new_n23721, n16517);
xnor_4 g22903(new_n16748, new_n16747, n16527);
xnor_4 g22904(new_n11548_1, new_n11547, n16554);
xnor_4 g22905(new_n6456_1, new_n6109, n16583);
xnor_4 g22906(new_n23097, new_n10738, new_n25255);
xnor_4 g22907(new_n25255, new_n23102, n16584);
xnor_4 g22908(new_n20548, new_n20519, n16589);
and_5  g22909(new_n20918, new_n20917, new_n25258);
nor_5  g22910(new_n25258, new_n20919, n16596);
xnor_4 g22911(new_n23926, new_n23877, n16617);
xnor_4 g22912(new_n8081, new_n8043, n16630);
xnor_4 g22913(new_n23906, new_n5188, n16640);
xnor_4 g22914(new_n2547_1, new_n2545, n16656);
xnor_4 g22915(new_n7354, new_n7301, n16674);
xnor_4 g22916(new_n15191, new_n15133, n16682);
xnor_4 g22917(new_n23841, new_n23815, n16684);
xnor_4 g22918(new_n11273_1, new_n11269, n16688);
xnor_4 g22919(new_n6742, new_n6733, n16733);
xnor_4 g22920(new_n8398, new_n8395, n16798);
xnor_4 g22921(new_n17854, new_n17852, n16834);
xnor_4 g22922(new_n3157, new_n3111, n16837);
xnor_4 g22923(new_n23382, new_n23378, n16841);
xnor_4 g22924(new_n5352, new_n5351_1, n16885);
xnor_4 g22925(new_n8713, new_n8640, n16905);
nor_5  g22926(new_n23290, new_n23285, new_n25275);
xnor_4 g22927(new_n25275, new_n19390, n16951);
xor_4  g22928(new_n17322, new_n17312, n16954);
xnor_4 g22929(new_n8891, new_n3854, n16989);
xnor_4 g22930(new_n20458, new_n20422, n17006);
xnor_4 g22931(new_n14402, new_n14400, n17068);
xnor_4 g22932(new_n16219_1, new_n16217_1, n17070);
xnor_4 g22933(new_n21929, new_n21878, n17075);
xnor_4 g22934(new_n18152_1, new_n18132, n17084);
xnor_4 g22935(new_n4979, new_n4978, n17104);
xnor_4 g22936(new_n14164, new_n14134, n17106);
xor_4  g22937(new_n10360, new_n10348, n17119);
xnor_4 g22938(new_n14040, new_n14003, n17130);
xnor_4 g22939(new_n24426, new_n24411, n17138);
xnor_4 g22940(new_n23726, new_n23715, n17163);
xor_4  g22941(new_n21554, new_n21553, n17168);
xnor_4 g22942(new_n12262, new_n12251, n17202);
xor_4  g22943(new_n20725, new_n20724, n17219);
xnor_4 g22944(new_n19880, new_n19839, n17232);
xnor_4 g22945(new_n16335, new_n16332, n17236);
not_8  g22946(new_n11165, new_n25295);
xnor_4 g22947(new_n25295, new_n11164, n17243);
xnor_4 g22948(new_n11886, new_n11870, n17263);
nor_5  g22949(new_n20898, new_n20890, new_n25298);
not_8  g22950(new_n20900, new_n25299);
nor_5  g22951(new_n20922, new_n25299, new_n25300);
nor_5  g22952(new_n25300, new_n25298, n17285);
xnor_4 g22953(new_n12446_1, new_n12415, n17320);
xnor_4 g22954(new_n2893, new_n2842, n17337);
xnor_4 g22955(new_n23512, new_n23502, n17344);
xnor_4 g22956(new_n23520, new_n23485, n17359);
xnor_4 g22957(new_n15173, new_n14228, n17387);
xnor_4 g22958(new_n5348, new_n5347, n17391);
xnor_4 g22959(new_n20453, new_n20429_1, n17392);
xnor_4 g22960(new_n23844, new_n23810, n17421);
xnor_4 g22961(new_n12987_1, new_n6925, n17432);
xnor_4 g22962(new_n22633, new_n22611, n17436);
xnor_4 g22963(new_n7585_1, new_n4970, n17440);
xnor_4 g22964(new_n8988, new_n6110, n17450);
not_8  g22965(new_n7808, new_n25314);
not_8  g22966(new_n20195, new_n25315);
nand_5 g22967(new_n25315, new_n25314, new_n25316_1);
nand_5 g22968(new_n7808, new_n20162, new_n25317);
nand_5 g22969(new_n25314, new_n7766, new_n25318);
nand_5 g22970(new_n7884_1, new_n25318, new_n25319);
nand_5 g22971(new_n25319, new_n25317, new_n25320);
nand_5 g22972(new_n25320, new_n25316_1, new_n25321);
nand_5 g22973(new_n20195, new_n7808, new_n25322);
nand_5 g22974(new_n25322, new_n25319, new_n25323);
nand_5 g22975(new_n25323, new_n25321, new_n25324);
not_8  g22976(new_n25324, n17461);
not_8  g22977(new_n24823, new_n25326);
xnor_4 g22978(new_n25326, new_n24822, n17466);
xnor_4 g22979(new_n14418, new_n14370, n17493);
xor_4  g22980(new_n23142, new_n23139, n17500);
xnor_4 g22981(new_n24132, new_n24129_1, n17524);
xnor_4 g22982(new_n6070, new_n6024, n17529);
xnor_4 g22983(new_n16010, new_n6105_1, new_n25332_1);
xnor_4 g22984(new_n25332_1, new_n16014, n17557);
xnor_4 g22985(new_n17758, new_n17721_1, n17583);
xnor_4 g22986(new_n15183, new_n15155, n17592);
xnor_4 g22987(new_n8899, new_n8881, n17638);
xnor_4 g22988(new_n21351, new_n21331, n17687);
xnor_4 g22989(new_n14743, new_n14705, n17721);
xnor_4 g22990(new_n23350, new_n23326, n17735);
not_8  g22991(new_n22715, new_n25340);
nand_5 g22992(new_n22716, new_n10760, new_n25341);
not_8  g22993(new_n25341, new_n25342);
nand_5 g22994(new_n25342, new_n25340, new_n25343);
nor_5  g22995(new_n22716, new_n10760, new_n25344);
nand_5 g22996(new_n25344, new_n22715, new_n25345_1);
nand_5 g22997(new_n25345_1, new_n25343, new_n25346);
nor_5  g22998(new_n25346, new_n22825, new_n25347);
nand_5 g22999(new_n25346, new_n22825, new_n25348);
not_8  g23000(new_n22718, new_n25349);
nor_5  g23001(new_n25349, new_n22703, new_n25350);
nor_5  g23002(new_n22729, new_n22719, new_n25351);
nor_5  g23003(new_n25351, new_n25350, new_n25352);
nand_5 g23004(new_n25352, new_n25348, new_n25353);
nand_5 g23005(new_n25353, new_n25343, new_n25354);
nor_5  g23006(new_n25354, new_n25347, n17738);
xor_4  g23007(new_n16426, new_n16421, n17746);
xnor_4 g23008(new_n24599, new_n24596, n17749);
xnor_4 g23009(new_n20059, new_n20037, n17820);
xnor_4 g23010(new_n15181, new_n15161, n17855);
nor_5  g23011(new_n15119, new_n5148, new_n25360);
nand_5 g23012(new_n5214, new_n25360, new_n25361);
not_8  g23013(new_n25361, new_n25362_1);
nor_5  g23014(new_n5214, new_n23874, new_n25363);
nor_5  g23015(new_n25363, new_n25362_1, new_n25364);
not_8  g23016(new_n25364, new_n25365_1);
not_8  g23017(new_n5215, new_n25366);
nor_5  g23018(new_n25366, new_n5040, new_n25367);
nor_5  g23019(new_n5294, new_n5216, new_n25368);
nor_5  g23020(new_n25368, new_n25367, new_n25369);
nor_5  g23021(new_n25369, new_n25365_1, new_n25370_1);
nor_5  g23022(new_n25370_1, new_n25362_1, n17877);
xnor_4 g23023(new_n16619, new_n16618, n17889);
not_8  g23024(new_n24480, new_n25373);
nor_5  g23025(new_n25373, new_n24468, new_n25374);
nor_5  g23026(new_n24490, new_n25374, new_n25375);
nor_5  g23027(new_n24480, new_n24467, new_n25376);
nor_5  g23028(new_n24489, new_n25376, new_n25377);
nor_5  g23029(new_n25377, new_n25375, n17912);
xnor_4 g23030(new_n23832, new_n23826, n17927);
xnor_4 g23031(new_n23918, new_n23889, n17931);
xnor_4 g23032(new_n8390, new_n8388, n17948);
xor_4  g23033(new_n16847, new_n16844, n17956);
not_8  g23034(new_n13448, new_n25383);
nor_5  g23035(new_n13676, new_n25383, new_n25384);
nor_5  g23036(new_n13596, new_n25383, new_n25385);
nor_5  g23037(new_n13675, new_n25385, new_n25386);
nor_5  g23038(new_n25386, new_n25384, n17963);
or_5   g23039(n25494, new_n19485, new_n25388);
nand_5 g23040(new_n18793, new_n18778, new_n25389);
nand_5 g23041(new_n25389, new_n25388, new_n25390);
not_8  g23042(new_n25390, new_n25391);
nand_5 g23043(new_n25391, new_n13998, new_n25392);
not_8  g23044(new_n25392, new_n25393);
not_8  g23045(new_n14001, new_n25394);
nor_5  g23046(new_n25391, new_n25394, new_n25395);
xnor_4 g23047(new_n25390, new_n14001, new_n25396);
not_8  g23048(new_n18794, new_n25397);
nand_5 g23049(new_n25397, new_n14005, new_n25398);
nand_5 g23050(new_n18820, new_n18795, new_n25399);
nand_5 g23051(new_n25399, new_n25398, new_n25400);
nor_5  g23052(new_n25400, new_n25396, new_n25401);
nor_5  g23053(new_n25401, new_n25395, new_n25402);
nor_5  g23054(new_n25402, new_n25393, new_n25403);
nor_5  g23055(new_n25391, new_n13998, new_n25404);
nor_5  g23056(new_n25404, new_n25401, new_n25405);
nor_5  g23057(new_n25405, new_n25403, n17976);
xnor_4 g23058(new_n7604, new_n7559, n17998);
xnor_4 g23059(new_n15618, new_n2876, n18025);
xnor_4 g23060(new_n22254, new_n22253_1, n18043);
xnor_4 g23061(new_n23742, new_n23739, n18045);
xnor_4 g23062(new_n4085_1, new_n4074, n18059);
xnor_4 g23063(new_n21927, new_n21882, n18061);
xnor_4 g23064(new_n3517, new_n3448, n18071);
xnor_4 g23065(new_n10692_1, new_n10625, n18143);
xnor_4 g23066(new_n23144, new_n23137, n18152);
xnor_4 g23067(new_n8073, new_n8063, n18193);
not_8  g23068(new_n12494, new_n25417);
not_8  g23069(new_n11937, new_n25418);
nor_5  g23070(new_n11969, new_n25418, new_n25419);
nor_5  g23071(new_n25419, new_n12499, new_n25420);
nor_5  g23072(new_n25420, new_n25015, new_n25421);
nor_5  g23073(new_n25421, new_n12496, new_n25422);
nand_5 g23074(new_n25422, new_n25417, new_n25423);
nand_5 g23075(new_n25423, new_n12492, new_n25424);
xnor_4 g23076(new_n12490, new_n12482, new_n25425);
xnor_4 g23077(new_n25425, new_n25424, n18232);
xnor_4 g23078(new_n18154, new_n18126, n18238);
xnor_4 g23079(new_n19866, new_n19862, n18241);
xnor_4 g23080(new_n22629, new_n22619_1, n18254);
xnor_4 g23081(new_n23348, new_n23329, n18288);
xnor_4 g23082(new_n13060, new_n13018, n18301);
xnor_4 g23083(new_n23728, new_n23709, n18304);
xnor_4 g23084(new_n14422, new_n14361, n18310);
xnor_4 g23085(new_n7028, new_n7025, n18311);
xnor_4 g23086(new_n18959, new_n18942, n18323);
xnor_4 g23087(new_n5728, new_n5685, n18332);
xnor_4 g23088(new_n23929, new_n23928, n18343);
xnor_4 g23089(new_n20814, new_n20811, n18350);
xnor_4 g23090(new_n19456, new_n19454_1, n18362);
xnor_4 g23091(new_n5290, new_n5229, n18377);
xnor_4 g23092(new_n4289, new_n4262, n18405);
xnor_4 g23093(new_n17992, new_n17982, n18414);
xnor_4 g23094(new_n15701, new_n15691, n18418);
xnor_4 g23095(new_n8707, new_n8658, n18437);
xnor_4 g23096(new_n21722, new_n21676, n18439);
xnor_4 g23097(new_n11959, new_n11958, n18445);
xnor_4 g23098(new_n7352, new_n7306, n18467);
xnor_4 g23099(new_n19886, new_n19822, n18482);
xnor_4 g23100(new_n20232, new_n20209, n18509);
xnor_4 g23101(new_n14978, new_n9632, n18513);
xnor_4 g23102(new_n16227, new_n16226, n18515);
xnor_4 g23103(new_n17162, new_n17138_1, n18572);
nor_5  g23104(new_n25197, new_n25182, new_n25453);
nor_5  g23105(new_n25453, new_n25057, new_n25454);
nand_5 g23106(new_n25197, new_n25182, new_n25455);
nand_5 g23107(new_n25455, new_n25057, new_n25456);
not_8  g23108(new_n25456, new_n25457);
nor_5  g23109(new_n25457, new_n25454, n18574);
xnor_4 g23110(new_n22781, new_n22776, n18576);
xnor_4 g23111(new_n24266, new_n24256, n18582);
xnor_4 g23112(new_n21462, new_n21446_1, n18583);
xnor_4 g23113(new_n21911, new_n21909, n18610);
xnor_4 g23114(new_n23758, new_n23754, n18635);
xnor_4 g23115(new_n7110, new_n7109, n18653);
xnor_4 g23116(new_n3873, new_n3815, n18679);
xnor_4 g23117(new_n22050_1, new_n22036, n18693);
xnor_4 g23118(new_n3155, new_n3116, n18708);
xnor_4 g23119(new_n24637, new_n18241_1, new_n25468_1);
xnor_4 g23120(new_n25468_1, new_n24644, n18721);
xnor_4 g23121(new_n20065, new_n20025, n18725);
xnor_4 g23122(new_n22415, new_n22389, n18751);
xnor_4 g23123(new_n17752, new_n17732, n18780);
xnor_4 g23124(new_n21061, new_n21009, n18782);
nand_5 g23125(new_n8020, new_n7930, new_n25474);
nand_5 g23126(new_n8091, new_n25474, new_n25475_1);
not_8  g23127(new_n8020, new_n25476);
nand_5 g23128(new_n25476, new_n7929, new_n25477);
nand_5 g23129(new_n8090, new_n25477, new_n25478);
nand_5 g23130(new_n25478, new_n25475_1, new_n25479);
not_8  g23131(new_n25479, n18802);
xor_4  g23132(new_n11664, new_n11663, n18830);
xnor_4 g23133(new_n13768, new_n13762, n18831);
xnor_4 g23134(new_n12811_1, new_n12801_1, n18843);
xnor_4 g23135(new_n3150, new_n3128, n18858);
xnor_4 g23136(new_n10679, new_n10658, n18859);
xnor_4 g23137(new_n18551, new_n18503, n18864);
xnor_4 g23138(new_n4817, new_n4740, n18865);
xnor_4 g23139(new_n23069, new_n23068_1, n18886);
xnor_4 g23140(new_n17748, new_n17747, n18887);
xnor_4 g23141(new_n9472, new_n9427, n18919);
xnor_4 g23142(new_n13278, new_n13265, n18940);
not_8  g23143(new_n24772, new_n25492);
xnor_4 g23144(new_n25492, new_n24771, n18945);
xnor_4 g23145(new_n24457, new_n24445, n18970);
xnor_4 g23146(new_n18218, new_n13016, new_n25495);
xnor_4 g23147(new_n25495, new_n18222, n18977);
xnor_4 g23148(new_n16337, new_n16329, n18982);
xor_4  g23149(new_n22502, new_n22501, n18999);
xnor_4 g23150(new_n6076, new_n6009, n19044);
xor_4  g23151(new_n16017, new_n16007, n19125);
xnor_4 g23152(new_n6074, new_n6014, n19141);
xnor_4 g23153(new_n15044, new_n15003, new_n25502);
xnor_4 g23154(new_n18661, new_n25502, new_n25503);
nand_5 g23155(new_n18665, new_n15131, new_n25504);
xnor_4 g23156(new_n15042, new_n15040, new_n25505);
xnor_4 g23157(new_n18665, new_n25505, new_n25506);
nand_5 g23158(new_n18668, new_n15135, new_n25507);
nand_5 g23159(new_n20097, new_n20079, new_n25508);
nand_5 g23160(new_n25508, new_n25507, new_n25509);
nand_5 g23161(new_n25509, new_n25506, new_n25510);
nand_5 g23162(new_n25510, new_n25504, new_n25511);
xnor_4 g23163(new_n25511, new_n25503, n19164);
xnor_4 g23164(new_n8907, new_n8906, n19174);
xnor_4 g23165(new_n22688, new_n22685, n19176);
xnor_4 g23166(new_n23730, new_n23702, n19202);
xnor_4 g23167(new_n21817, new_n21807, n19220);
and_5  g23168(new_n8410, new_n8346, new_n25517);
nor_5  g23169(new_n25517, new_n8411, n19221);
xnor_4 g23170(new_n12090, new_n12089, n19223);
xnor_4 g23171(new_n18537_1, new_n18535, n19224);
xnor_4 g23172(new_n16787, new_n16775, n19233);
xnor_4 g23173(new_n13749, new_n13713, n19244);
xnor_4 g23174(new_n9474, new_n9422, n19314);
xnor_4 g23175(new_n11558, new_n11557, n19315);
xnor_4 g23176(new_n14414_1, new_n14380, n19323);
xnor_4 g23177(new_n23510, new_n23506, n19333);
nand_5 g23178(new_n19160, new_n18652, new_n25527);
nand_5 g23179(new_n25527, new_n10614_1, new_n25528);
not_8  g23180(new_n25528, new_n25529);
nand_5 g23181(new_n18657, new_n10617_1, new_n25530);
nand_5 g23182(new_n18683, new_n18658, new_n25531);
nand_5 g23183(new_n25531, new_n25530, new_n25532_1);
not_8  g23184(new_n25527, new_n25533);
xnor_4 g23185(new_n25533, new_n10614_1, new_n25534);
not_8  g23186(new_n25534, new_n25535);
nor_5  g23187(new_n25535, new_n25532_1, new_n25536);
nor_5  g23188(new_n25536, new_n25529, n19348);
xnor_4 g23189(new_n18166, new_n18089, n19354);
xnor_4 g23190(new_n11894, new_n11859, n19367);
xnor_4 g23191(new_n20630, new_n20600, n19385);
xnor_4 g23192(new_n18297, new_n18241_1, new_n25541);
xnor_4 g23193(new_n25541, new_n18329, n19389);
xnor_4 g23194(new_n17618, new_n17586, n19401);
not_8  g23195(new_n24029, new_n25544);
xnor_4 g23196(new_n24038, new_n25544, n19414);
xnor_4 g23197(new_n20836, new_n19261, n19424);
xnor_4 g23198(new_n23073, new_n23053, n19450);
nand_5 g23199(new_n25533, new_n15052_1, new_n25548);
xnor_4 g23200(new_n25527, new_n15052_1, new_n25549);
not_8  g23201(new_n15118_1, new_n25550_1);
nand_5 g23202(new_n18657, new_n25550_1, new_n25551);
xnor_4 g23203(new_n18657, new_n15118_1, new_n25552);
nand_5 g23204(new_n18661, new_n15124, new_n25553);
nand_5 g23205(new_n25511, new_n25503, new_n25554);
nand_5 g23206(new_n25554, new_n25553, new_n25555);
nand_5 g23207(new_n25555, new_n25552, new_n25556);
nand_5 g23208(new_n25556, new_n25551, new_n25557);
nand_5 g23209(new_n25557, new_n25549, new_n25558);
nand_5 g23210(new_n25558, new_n25548, n19458);
xnor_4 g23211(new_n16428_1, new_n16418, n19467);
xnor_4 g23212(new_n8709, new_n8652, n19496);
not_8  g23213(new_n16383, new_n25562);
xnor_4 g23214(new_n25562, new_n16373, n19523);
xnor_4 g23215(new_n4809, new_n4765, n19570);
xnor_4 g23216(new_n12951, new_n12937, n19602);
xnor_4 g23217(new_n13327, new_n13321, n19617);
xnor_4 g23218(new_n14741, new_n14709, n19623);
xnor_4 g23219(new_n24080, new_n24079, n19641);
xnor_4 g23220(new_n23846, new_n23806, n19648);
xnor_4 g23221(new_n17160, new_n17142, n19664);
xnor_4 g23222(new_n21551, new_n21537, n19736);
not_8  g23223(new_n24025, new_n25572);
nor_5  g23224(new_n24040, new_n25572, new_n25573);
nor_5  g23225(new_n25572, new_n3293, new_n25574);
nor_5  g23226(new_n24039_1, new_n25574, new_n25575);
nor_5  g23227(new_n25575, new_n25573, n19749);
xnor_4 g23228(new_n16086, new_n16073, n19756);
xnor_4 g23229(new_n12947, new_n12945, n19767);
xnor_4 g23230(new_n3439, new_n3436, new_n25579);
xnor_4 g23231(new_n25579, new_n3519, n19780);
xnor_4 g23232(new_n24667, new_n24664, n19792);
xnor_4 g23233(new_n22243, new_n22227, n19798);
xor_4  g23234(new_n17850, new_n17847, n19873);
nand_5 g23235(new_n19922_1, new_n19899, new_n25584);
nand_5 g23236(new_n19909_1, new_n19899, new_n25585);
nand_5 g23237(new_n19921, new_n25585, new_n25586_1);
nand_5 g23238(new_n25586_1, new_n25584, new_n25587);
not_8  g23239(new_n25587, n19909);
xnor_4 g23240(new_n21549_1, new_n21541, n19916);
xnor_4 g23241(new_n22247, new_n22221, n19923);
xnor_4 g23242(new_n20460, new_n20419, n19930);
xnor_4 g23243(new_n6760, new_n6637, n19968);
xnor_4 g23244(new_n21049, new_n21033, n19988);
nand_5 g23245(new_n23098, new_n22316, new_n25594);
nand_5 g23246(new_n22315, new_n10820, new_n25595);
nand_5 g23247(new_n22320, new_n22317_1, new_n25596);
nand_5 g23248(new_n25596, new_n25595, new_n25597);
nand_5 g23249(new_n25597, new_n25594, new_n25598);
nand_5 g23250(new_n23097, new_n22315, new_n25599);
nand_5 g23251(new_n25599, new_n25596, new_n25600);
nand_5 g23252(new_n25600, new_n25598, new_n25601);
not_8  g23253(new_n25601, n20004);
xnor_4 g23254(new_n22411, new_n22393, n20017);
xnor_4 g23255(new_n19882, new_n19833, n20033);
xnor_4 g23256(new_n14940, new_n14939, n20061);
xnor_4 g23257(new_n19405, new_n19401_1, n20069);
nand_5 g23258(new_n15579, new_n15570_1, new_n25607);
nand_5 g23259(new_n15643, new_n15581, new_n25608);
nand_5 g23260(new_n25608, new_n25607, n20086);
xnor_4 g23261(new_n20915_1, new_n20912, n20096);
xnor_4 g23262(new_n14405, new_n14394, n20103);
xnor_4 g23263(new_n12448, new_n12410, n20126);
xnor_4 g23264(new_n22864, new_n22830, n20149);
xnor_4 g23265(new_n12824, new_n12774, n20187);
xnor_4 g23266(new_n18774, new_n18741, n20279);
nand_5 g23267(new_n24248, new_n24242, new_n25616);
nand_5 g23268(new_n24252, new_n25616, new_n25617);
not_8  g23269(new_n24248, new_n25618);
nand_5 g23270(new_n24268, new_n25618, new_n25619_1);
not_8  g23271(new_n24268, new_n25620);
nand_5 g23272(new_n25620, new_n18934, new_n25621);
nand_5 g23273(new_n25621, new_n25619_1, new_n25622);
nor_5  g23274(new_n25622, new_n25617, n20287);
xnor_4 g23275(new_n22088, new_n22085, n20301);
not_8  g23276(new_n8634, new_n25625);
nand_5 g23277(new_n8715, new_n25625, new_n25626);
nand_5 g23278(new_n25626, new_n23614, new_n25627);
not_8  g23279(new_n25627, n20330);
xnor_4 g23280(new_n12820, new_n12781, n20333);
not_8  g23281(new_n11087, new_n25630);
nor_5  g23282(new_n25630, new_n10941, new_n25631);
not_8  g23283(new_n11092, new_n25632);
not_8  g23284(new_n11170, new_n25633);
nand_5 g23285(new_n25633, new_n25632, new_n25634);
nand_5 g23286(new_n25634, new_n25631, new_n25635);
not_8  g23287(new_n10941, new_n25636);
nor_5  g23288(new_n11087, new_n25636, new_n25637);
nand_5 g23289(new_n11171, new_n25637, new_n25638);
nand_5 g23290(new_n25638, new_n25635, n20355);
xor_4  g23291(new_n8943_1, new_n5469, n20366);
xnor_4 g23292(new_n20667, new_n20663, n20388);
xnor_4 g23293(new_n23916, new_n23892, n20402);
xnor_4 g23294(new_n16606, new_n16578, n20403);
xor_4  g23295(new_n3138, new_n3137, n20424);
xnor_4 g23296(new_n21916, new_n21902, n20436);
xor_4  g23297(new_n8695, new_n8694_1, n20441);
xnor_4 g23298(new_n8089, new_n8025, n20445);
xnor_4 g23299(new_n5292, new_n5224, n20450);
xnor_4 g23300(new_n17764, new_n17762, n20490);
xor_4  g23301(new_n21815, new_n21812, n20495);
nor_5  g23302(new_n16626, new_n16624, new_n25651);
nand_5 g23303(new_n25651, new_n16622, new_n25652);
nand_5 g23304(new_n16626, new_n16624, new_n25653);
not_8  g23305(new_n25653, new_n25654);
nand_5 g23306(new_n25654, new_n16623, new_n25655);
nand_5 g23307(new_n25655, new_n25652, n20515);
nand_5 g23308(new_n24669, new_n24658, new_n25657);
nand_5 g23309(new_n25657, new_n24653, new_n25658);
not_8  g23310(new_n25658, n20533);
xnor_4 g23311(new_n19265, new_n19256, n20582);
xnor_4 g23312(new_n21228, new_n21193_1, n20590);
xnor_4 g23313(new_n3500, new_n3496, n20602);
xnor_4 g23314(new_n17745, new_n17743, n20609);
xnor_4 g23315(new_n6929, new_n6920, n20623);
xnor_4 g23316(new_n22258, new_n22207, n20629);
xnor_4 g23317(new_n14937, new_n14929, n20661);
xnor_4 g23318(new_n8992, new_n8991, n20673);
xnor_4 g23319(new_n22251, new_n22215, n20678);
nor_5  g23320(new_n16060_1, new_n12696, new_n25669);
nor_5  g23321(new_n16092, new_n25669, new_n25670);
not_8  g23322(new_n16056, new_n25671);
nand_5 g23323(new_n16060_1, new_n12696, new_n25672);
nand_5 g23324(new_n25672, new_n25671, new_n25673);
nor_5  g23325(new_n25673, new_n25670, n20680);
xnor_4 g23326(new_n6736_1, new_n4343, n20685);
xnor_4 g23327(new_n25390, new_n13998, new_n25676);
xnor_4 g23328(new_n25676, new_n25402, n20691);
xnor_4 g23329(new_n17158, new_n17147, n20696);
xnor_4 g23330(new_n24424, new_n24414, n20704);
xor_4  g23331(new_n23342_1, new_n23341_1, n20705);
xnor_4 g23332(new_n10690, new_n10630, n20709);
xnor_4 g23333(new_n15971, new_n15946, n20713);
xnor_4 g23334(new_n9183, new_n9182_1, n20722);
not_8  g23335(new_n24961, new_n25684);
nor_5  g23336(new_n25684, new_n21106, new_n25685);
nor_5  g23337(new_n21105, new_n24963, new_n25686);
nor_5  g23338(new_n21106, new_n21093_1, new_n25687);
nor_5  g23339(new_n21118, new_n25687, new_n25688);
nor_5  g23340(new_n25688, new_n25686, new_n25689);
nor_5  g23341(new_n25689, new_n25685, new_n25690);
nor_5  g23342(new_n24961, new_n21105, new_n25691);
nor_5  g23343(new_n25691, new_n25688, new_n25692);
nor_5  g23344(new_n25692, new_n25690, n20723);
xnor_4 g23345(new_n24241, new_n18934, new_n25694_1);
xnor_4 g23346(new_n25694_1, new_n25620, n20748);
xor_4  g23347(new_n5720, new_n5709, n20761);
xnor_4 g23348(new_n21925, new_n21885, n20774);
xnor_4 g23349(new_n25557, new_n25549, n20788);
nor_5  g23350(new_n24802, new_n23751, new_n25699);
nor_5  g23351(new_n25699, new_n24918, new_n25700);
nor_5  g23352(new_n24801, new_n23752, new_n25701);
nor_5  g23353(new_n25701, new_n24917, new_n25702);
nor_5  g23354(new_n25702, new_n25700, n20795);
xnor_4 g23355(new_n21961, new_n21948, new_n25704);
nand_5 g23356(new_n21971, new_n21948, new_n25705);
nand_5 g23357(new_n25705, new_n21966, new_n25706_1);
nand_5 g23358(new_n25706_1, new_n21973, new_n25707);
xnor_4 g23359(new_n25707, new_n25704, n20803);
xnor_4 g23360(new_n25369, new_n25364, n20869);
xnor_4 g23361(new_n24601, new_n24593, n20879);
xnor_4 g23362(new_n6748, new_n6716, n20915);
xnor_4 g23363(n19282, n2160, new_n25712);
or_5   g23364(n12657, new_n17821, new_n25713);
nand_5 g23365(new_n23359, new_n23355_1, new_n25714);
nand_5 g23366(new_n25714, new_n25713, new_n25715);
xnor_4 g23367(new_n25715, new_n25712, new_n25716);
not_8  g23368(new_n25716, new_n25717);
nor_5  g23369(new_n25717, new_n23209, new_n25718);
not_8  g23370(new_n25718, new_n25719_1);
nor_5  g23371(new_n23360, new_n21496, new_n25720);
nor_5  g23372(new_n23364, new_n23361, new_n25721);
nor_5  g23373(new_n25721, new_n25720, new_n25722);
xnor_4 g23374(new_n25716, new_n23208, new_n25723);
nor_5  g23375(new_n25723, new_n25722, new_n25724);
not_8  g23376(new_n25724, new_n25725);
nand_5 g23377(new_n25725, new_n25719_1, new_n25726);
or_5   g23378(n19282, new_n12514, new_n25727);
nand_5 g23379(new_n25715, new_n25712, new_n25728);
nand_5 g23380(new_n25728, new_n25727, new_n25729);
nor_5  g23381(new_n25729, new_n24482, new_n25730);
nand_5 g23382(new_n25730, new_n25726, new_n25731);
not_8  g23383(new_n25731, new_n25732);
nand_5 g23384(new_n25732, new_n24480, new_n25733);
nor_5  g23385(new_n25724, new_n25718, new_n25734);
not_8  g23386(new_n24482, new_n25735);
not_8  g23387(new_n25729, new_n25736);
nor_5  g23388(new_n25736, new_n25735, new_n25737);
nand_5 g23389(new_n25737, new_n25734, new_n25738_1);
not_8  g23390(new_n25738_1, new_n25739);
nand_5 g23391(new_n25739, new_n25373, new_n25740);
nand_5 g23392(new_n25740, new_n25733, n20935);
xnor_4 g23393(new_n23839, new_n23819, n20936);
xnor_4 g23394(new_n18201, new_n18199, n21008);
xnor_4 g23395(new_n21059, new_n21013, n21017);
nor_5  g23396(new_n25035, new_n23171, new_n25745);
nand_5 g23397(new_n25035, new_n23171, new_n25746);
not_8  g23398(new_n25039, new_n25747);
nand_5 g23399(new_n25747, new_n25746, new_n25748);
nand_5 g23400(new_n25748, new_n25034, new_n25749_1);
nor_5  g23401(new_n25749_1, new_n25745, n21034);
xnor_4 g23402(new_n24005, new_n24003, n21046);
xnor_4 g23403(new_n9101, new_n9080, n21062);
xnor_4 g23404(new_n24750, new_n24741, new_n25753);
xnor_4 g23405(new_n25753, new_n24652, n21093);
xnor_4 g23406(new_n10394, new_n8379, n21094);
xnor_4 g23407(new_n15852, new_n15829, n21123);
xnor_4 g23408(new_n20346, new_n19479, n21154);
xnor_4 g23409(new_n16757, new_n16730, n21157);
xnor_4 g23410(new_n22856, new_n22846, n21168);
xnor_4 g23411(new_n7855, new_n7853, n21173);
xnor_4 g23412(new_n4805, new_n4777_1, n21176);
xnor_4 g23413(new_n15496_1, new_n15487, n21182);
nand_5 g23414(new_n23798, new_n22885, new_n25763);
not_8  g23415(new_n23848, new_n25764);
nand_5 g23416(new_n25764, new_n22884, new_n25765);
nand_5 g23417(new_n25765, new_n25763, new_n25766);
not_8  g23418(new_n23802, new_n25767);
nand_5 g23419(new_n23848, new_n22896, new_n25768);
nand_5 g23420(new_n25768, new_n25767, new_n25769);
nor_5  g23421(new_n25769, new_n25766, n21193);
xnor_4 g23422(new_n10112, new_n10110, n21203);
xnor_4 g23423(new_n17742, new_n2570_1, n21225);
xnor_4 g23424(new_n21476, new_n21418, n21238);
xnor_4 g23425(new_n14942, new_n14922, n21254);
xnor_4 g23426(new_n21718, new_n21684, n21298);
xnor_4 g23427(new_n21455, new_n10005, n21302);
xnor_4 g23428(new_n21547, new_n21544, n21349);
xnor_4 g23429(new_n17325, new_n17324, n21365);
xnor_4 g23430(new_n16385, new_n16369, n21367);
xnor_4 g23431(new_n12686, new_n12653, n21396);
xnor_4 g23432(new_n8087, new_n8030, n21399);
not_8  g23433(new_n3528_1, new_n25782);
xnor_4 g23434(new_n25782, new_n3521, n21404);
xnor_4 g23435(new_n8994, new_n8982_1, n21446);
xnor_4 g23436(new_n12505, new_n12494, n21472);
xnor_4 g23437(new_n7878, new_n7824, n21525);
xnor_4 g23438(new_n18603, new_n18576_1, n21549);
xnor_4 g23439(new_n21347, new_n21343, n21615);
nor_5  g23440(new_n24248, new_n14512, new_n25789);
xnor_4 g23441(new_n24248, new_n8331, new_n25790);
not_8  g23442(new_n25790, new_n25791);
nor_5  g23443(new_n24251, new_n8331, new_n25792_1);
nor_5  g23444(new_n18965, new_n18935, new_n25793);
nor_5  g23445(new_n25793, new_n25792_1, new_n25794);
nor_5  g23446(new_n25794, new_n25791, new_n25795);
nor_5  g23447(new_n25795, new_n25789, n21628);
nor_5  g23448(new_n23406, new_n22891_1, new_n25797_1);
xnor_4 g23449(new_n23405, new_n22891_1, new_n25798);
not_8  g23450(new_n25798, new_n25799);
nor_5  g23451(new_n23411, new_n22895, new_n25800);
nor_5  g23452(new_n24884, new_n24880, new_n25801);
nor_5  g23453(new_n25801, new_n25800, new_n25802);
nor_5  g23454(new_n25802, new_n25799, new_n25803);
nor_5  g23455(new_n25803, new_n25797_1, n21637);
xnor_4 g23456(new_n23344, new_n23335, n21645);
xnor_4 g23457(new_n12980_1, new_n6921, n21665);
xnor_4 g23458(new_n16090, new_n16067, n21680);
xnor_4 g23459(new_n23924_1, new_n23880, n21685);
xnor_4 g23460(new_n20061_1, new_n20033_1, n21717);
xnor_4 g23461(new_n18187, new_n18180, n21719);
xnor_4 g23462(new_n20053, new_n20049, n21750);
xnor_4 g23463(new_n23626, new_n23625, n21765);
xnor_4 g23464(new_n25723, new_n25722, n21800);
xnor_4 g23465(new_n4485, new_n4481, new_n25814);
xnor_4 g23466(new_n25814, new_n4492, n21820);
xnor_4 g23467(new_n21053, new_n21025, n21874);
xnor_4 g23468(new_n14407, new_n14391, n21943);
xnor_4 g23469(new_n17329, new_n17305, n21960);
xnor_4 g23470(new_n7593_1, new_n24272, n21976);
xnor_4 g23471(new_n12099, new_n12068, n21986);
xnor_4 g23472(new_n11896, new_n11855, n22016);
xnor_4 g23473(new_n20055, new_n20045, n22027);
xnor_4 g23474(new_n14160, new_n14148_1, n22050);
xnor_4 g23475(new_n4345, new_n4344, n22063);
xnor_4 g23476(new_n22854, new_n22850, n22076);
nor_5  g23477(new_n21958, new_n14900, new_n25826_1);
not_8  g23478(new_n22290_1, new_n25827);
nor_5  g23479(new_n22310, new_n25827, new_n25828);
nor_5  g23480(new_n25828, new_n25826_1, n22090);
xnor_4 g23481(new_n24455, new_n24447, n22107);
xnor_4 g23482(new_n19146, new_n19114, n22113);
not_8  g23483(new_n14900, new_n25832);
nor_5  g23484(new_n25832, new_n14836, new_n25833);
nor_5  g23485(new_n14950, new_n25833, new_n25834);
nor_5  g23486(new_n14900, new_n14837, new_n25835);
nor_5  g23487(new_n14949, new_n25835, new_n25836);
nor_5  g23488(new_n25836, new_n25834, n22124);
not_8  g23489(new_n25150, new_n25838);
nor_5  g23490(new_n25838, new_n20898, new_n25839_1);
not_8  g23491(new_n25151, new_n25840_1);
nor_5  g23492(new_n25154, new_n25840_1, new_n25841);
nor_5  g23493(new_n25841, new_n25839_1, n22126);
nor_5  g23494(new_n25739, new_n25732, new_n25843);
xnor_4 g23495(new_n25843, new_n25373, n22130);
xor_4  g23496(new_n19347, new_n19346, n22144);
xnor_4 g23497(new_n24874, new_n24867, n22150);
xnor_4 g23498(new_n21276_1, new_n21268, n22157);
xnor_4 g23499(new_n25509, new_n25506, n22213);
xnor_4 g23500(new_n11150, new_n11149, n22283);
xor_4  g23501(new_n21993_1, new_n21992, n22311);
xnor_4 g23502(new_n9476, new_n9417, n22317);
xnor_4 g23503(new_n18880_1, new_n18866, n22341);
not_8  g23504(new_n19654, new_n25853);
nor_5  g23505(new_n7631, new_n7617, new_n25854);
not_8  g23506(new_n25854, new_n25855);
nor_5  g23507(new_n25855, new_n7612, new_n25856);
not_8  g23508(new_n25856, new_n25857);
not_8  g23509(new_n7631, new_n25858);
nor_5  g23510(new_n25858, new_n7616_1, new_n25859);
nand_5 g23511(new_n25859, new_n7612, new_n25860);
nand_5 g23512(new_n25860, new_n25857, new_n25861);
xnor_4 g23513(new_n25861, new_n25853, n22353);
xnor_4 g23514(new_n18878, new_n18870, n22444);
xnor_4 g23515(new_n10873, new_n20729, n22467);
xnor_4 g23516(new_n9453, new_n9452, n22484);
xnor_4 g23517(new_n4815, new_n4747_1, n22489);
xnor_4 g23518(new_n8913, new_n8861_1, n22494);
xnor_4 g23519(new_n11156, new_n11125, n22533);
xnor_4 g23520(new_n24422, new_n24421_1, n22584);
not_8  g23521(new_n19353, new_n25870);
nor_5  g23522(new_n25870, new_n19327_1, new_n25871);
nor_5  g23523(new_n25871, new_n19287, n22589);
xnor_4 g23524(new_n25555, new_n25552, n22620);
xnor_4 g23525(new_n8990, new_n8989, n22623);
xnor_4 g23526(new_n18325, new_n18311_1, n22697);
xnor_4 g23527(new_n9466, new_n9445_1, n22714);
xnor_4 g23528(new_n12828, new_n12766, n22761);
xnor_4 g23529(new_n20545, new_n20524, n22779);
xnor_4 g23530(new_n24432, new_n24400, n22787);
xnor_4 g23531(new_n2564, new_n2525, n22819);
xnor_4 g23532(new_n9817, new_n23118, n22858);
xnor_4 g23533(new_n24934_1, new_n12466, new_n25882);
xnor_4 g23534(new_n25882, new_n24937_1, n22870);
xor_4  g23535(new_n10362, new_n10342, n22891);
xor_4  g23536(new_n21220, new_n21205, n22897);
xnor_4 g23537(new_n10892, new_n10826, n22903);
xnor_4 g23538(new_n15510, new_n15464, n22907);
xnor_4 g23539(new_n7598_1, new_n7597, n22910);
xnor_4 g23540(new_n13304, new_n13296, n22914);
xnor_4 g23541(new_n6083, new_n6049, n22939);
xnor_4 g23542(new_n20672, new_n4610, new_n25891);
xnor_4 g23543(new_n25891, new_n20669, n22998);
xnor_4 g23544(new_n9462, new_n9461, n23006);
xnor_4 g23545(new_n13771, new_n13760, n23007);
xnor_4 g23546(new_n19557, new_n19554, n23009);
xnor_4 g23547(new_n18164, new_n18096, n23014);
xnor_4 g23548(new_n25802, new_n25798, n23047);
xnor_4 g23549(new_n18957, new_n18945_1, n23058);
nand_5 g23550(new_n20076, new_n20069_1, new_n25899);
not_8  g23551(new_n25899, n23066);
nor_5  g23552(new_n19951, new_n25636, new_n25901);
nor_5  g23553(new_n25901, new_n19953, new_n25902);
xnor_4 g23554(new_n25902, new_n19947, n23067);
xor_4  g23555(new_n17320_1, new_n17314, n23238);
xnor_4 g23556(new_n18681, new_n18663, n23247);
xnor_4 g23557(new_n16222, new_n16212, n23248);
xnor_4 g23558(new_n18767, new_n18751_1, n23270);
xnor_4 g23559(new_n24488, new_n24484, n23289);
xnor_4 g23560(new_n5730, new_n5681, n23305);
xnor_4 g23561(new_n22627, new_n22623_1, n23341);
xnor_4 g23562(new_n10006, new_n5191, n23342);
nand_5 g23563(new_n22971, new_n8020, new_n25912);
nand_5 g23564(new_n22994, new_n25912, new_n25913);
nand_5 g23565(new_n22970, new_n25476, new_n25914);
nand_5 g23566(new_n22993, new_n25914, new_n25915);
nand_5 g23567(new_n25915, new_n25913, new_n25916);
not_8  g23568(new_n25916, n23355);
xnor_4 g23569(new_n20780, new_n20777, n23371);
xnor_4 g23570(new_n16610, new_n16568, n23401);
xnor_4 g23571(new_n14157, new_n14156, n23414);
xnor_4 g23572(new_n18772, new_n18745_1, n23429);
nand_5 g23573(new_n23232, new_n23223, new_n25922);
nand_5 g23574(new_n23227, new_n23223, new_n25923_1);
nand_5 g23575(new_n25923_1, new_n23231, new_n25924);
nand_5 g23576(new_n25924, new_n25922, new_n25925);
not_8  g23577(new_n25925, n23433);
xnor_4 g23578(new_n19874, new_n19855, n23434);
nand_5 g23579(new_n25150, new_n23374, new_n25928);
nand_5 g23580(new_n25928, new_n25172, new_n25929);
nand_5 g23581(new_n25838, new_n25167, new_n25930);
nand_5 g23582(new_n25930, new_n25171, new_n25931);
nand_5 g23583(new_n25931, new_n25929, new_n25932);
not_8  g23584(new_n25932, n23450);
xnor_4 g23585(new_n18162, new_n18102, n23471);
xnor_4 g23586(new_n22637, new_n22603, n23480);
xnor_4 g23587(new_n19181, new_n19174_1, n23546);
xnor_4 g23588(new_n22241, new_n22232, n23550);
xnor_4 g23589(new_n7872, new_n7841_1, n23585);
xor_4  g23590(new_n21218, new_n21209, n23588);
xor_4  g23591(new_n22499, new_n22498, n23619);
xnor_4 g23592(new_n3148, new_n3136_1, n23624);
xnor_4 g23593(new_n12678, new_n12669, n23628);
xnor_4 g23594(new_n23514, new_n23498, n23637);
xnor_4 g23595(new_n24194, new_n24190, n23663);
xnor_4 g23596(new_n12680, new_n12665_1, n23669);
xnor_4 g23597(new_n14038, new_n14008, n23684);
xnor_4 g23598(new_n20448, new_n20439, n23690);
xnor_4 g23599(new_n23922, new_n23883_1, n23714);
nand_5 g23600(new_n25208, new_n25204, new_n25949);
not_8  g23601(new_n25949, n23719);
xnor_4 g23602(new_n22942, new_n22939_1, n23748);
xnor_4 g23603(new_n11658, new_n7635, n23856);
xnor_4 g23604(new_n7870, new_n7869, n23883);
xnor_4 g23605(new_n15489, new_n11145, new_n25954);
xnor_4 g23606(new_n25954, new_n15492, n23888);
xnor_4 g23607(new_n3507, new_n3474, n23899);
xnor_4 g23608(new_n16013_1, new_n10104, n23903);
xnor_4 g23609(new_n13747, new_n13716, n23924);
xnor_4 g23610(new_n17814, new_n17813, n23935);
xnor_4 g23611(new_n14034, new_n14018, n23942);
xnor_4 g23612(new_n18998, new_n18989, n23954);
xnor_4 g23613(new_n20157, new_n20131, n23958);
xnor_4 g23614(new_n24066, new_n24064, n23986);
xnor_4 g23615(new_n18204, new_n18197, n24002);
xnor_4 g23616(new_n13927, new_n13918, n24039);
xnor_4 g23617(new_n25134, new_n25133_1, n24052);
xnor_4 g23618(new_n21918, new_n21898_1, n24092);
xnor_4 g23619(new_n16753, new_n16752, n24096);
xnor_4 g23620(new_n13052, new_n13023, n24097);
xnor_4 g23621(new_n12684, new_n12657_1, n24105);
xnor_4 g23622(new_n19537, new_n19515_1, n24119);
xnor_4 g23623(new_n16088, new_n16070, n24133);
xnor_4 g23624(new_n21468, new_n21434, n24141);
xnor_4 g23625(new_n22822, new_n22792, new_n25974_1);
xnor_4 g23626(new_n25974_1, new_n22866, n24145);
xnor_4 g23627(new_n23597, new_n23593, n24146);
xnor_4 g23628(new_n13669, new_n13611, n24155);
xnor_4 g23629(new_n25400, new_n25396, n24160);
xnor_4 g23630(new_n9832_1, new_n9795, n24167);
nor_5  g23631(new_n22059, new_n22052, n24172);
xnor_4 g23632(new_n15498, new_n15482, n24177);
xnor_4 g23633(new_n25245, new_n25244_1, n24228);
xnor_4 g23634(new_n18882, new_n18862, n24258);
nor_5  g23635(new_n19654, new_n7617, new_n25984);
nor_5  g23636(new_n25860, new_n19654, new_n25985_1);
nor_5  g23637(new_n25985_1, new_n25856, new_n25986);
nor_5  g23638(new_n25986, new_n25984, n24260);
xnor_4 g23639(new_n20550, new_n20514, n24289);
xnor_4 g23640(new_n4982, new_n4968, n24297);
xnor_4 g23641(new_n12676, new_n4075, n24307);
xnor_4 g23642(new_n2558, new_n2544, n24342);
xnor_4 g23643(new_n17327, new_n17308, n24345);
xnor_4 g23644(new_n10116, new_n10102, n24347);
xnor_4 g23645(new_n5288, new_n5234, n24373);
xor_4  g23646(new_n19468, new_n19467_1, n24406);
xnor_4 g23647(new_n14795, new_n14782, n24415);
xnor_4 g23648(new_n11553, new_n11552, n24421);
xnor_4 g23649(new_n14612, new_n14582, n24431);
xnor_4 g23650(new_n12818, new_n12784, n24472);
nand_5 g23651(new_n24497, new_n23988, new_n26000);
nand_5 g23652(new_n26000, new_n24499, new_n26001);
xnor_4 g23653(new_n26001, new_n24493, n24476);
xnor_4 g23654(new_n10886, new_n10841, n24483);
xnor_4 g23655(new_n14493, new_n14491, n24501);
xnor_4 g23656(new_n19580, new_n19576, n24512);
xnor_4 g23657(new_n4985, new_n4984, n24558);
xnor_4 g23658(new_n2877, new_n2875, n24576);
xnor_4 g23659(new_n2881, new_n2879, n24579);
xnor_4 g23660(new_n21997_1, new_n21985, n24602);
xnor_4 g23661(new_n15365, new_n15329, n24604);
xnor_4 g23662(new_n24623, new_n24620_1, n24626);
xnor_4 g23663(new_n23609, new_n23605, n24629);
xnor_4 g23664(new_n23346, new_n23332, n24636);
xnor_4 g23665(new_n23066_1, new_n23063, n24715);
xnor_4 g23666(new_n21931, new_n21875, n24723);
xnor_4 g23667(new_n18084, new_n18040, new_n26016);
xnor_4 g23668(new_n26016, new_n18168, n24749);
xnor_4 g23669(new_n21921, new_n21892, n24758);
xnor_4 g23670(new_n24705, new_n24702, n24784);
xnor_4 g23671(new_n17506, new_n17505, n24807);
xnor_4 g23672(new_n10388_1, new_n8386, n24826);
xnor_4 g23673(new_n8083, new_n8040, n24840);
xnor_4 g23674(new_n10677, new_n10664, n24841);
xnor_4 g23675(new_n5479, new_n5467, n24853);
xnor_4 g23676(new_n3153, new_n3121, n24857);
xnor_4 g23677(new_n6744, new_n6728, n24887);
xor_4  g23678(new_n9822, new_n9814, n24934);
xnor_4 g23679(new_n7882, new_n7814, n24998);
xnor_4 g23680(new_n12439, new_n12424, n25006);
xnor_4 g23681(new_n22306, new_n22294, n25032);
xnor_4 g23682(new_n17447, new_n17424, n25062);
xnor_4 g23683(new_n21002, new_n18040, new_n26032);
xnor_4 g23684(new_n26032, new_n21065, n25083);
xor_4  g23685(new_n14030, new_n14027, n25097);
xnor_4 g23686(new_n19172, new_n19168, n25133);
xnor_4 g23687(new_n19876, new_n19852, n25155);
xnor_4 g23688(new_n25736, new_n24482, new_n26037);
xnor_4 g23689(new_n26037, new_n25734, n25181);
xnor_4 g23690(new_n22308, new_n22292, n25200);
nor_5  g23691(new_n23082, new_n23079, new_n26040);
xnor_4 g23692(new_n23075, new_n18241_1, new_n26041);
xnor_4 g23693(new_n26041, new_n26040, n25209);
xnor_4 g23694(new_n16302, new_n16300, n25215);
xnor_4 g23695(new_n19660, new_n19656, n25244);
xnor_4 g23696(new_n19269, new_n19247, n25254);
xor_4  g23697(new_n22504, new_n22474, n25256);
nor_5  g23698(new_n25088, new_n23165, new_n26047);
nor_5  g23699(new_n26047, new_n25097_1, new_n26048);
xnor_4 g23700(new_n25088, new_n24075, new_n26049);
xnor_4 g23701(new_n26049, new_n26048, n25293);
xor_4  g23702(new_n22494_1, new_n22486, n25328);
xnor_4 g23703(new_n11875, new_n4490, n25332);
not_8  g23704(new_n23243, new_n26053_1);
nor_5  g23705(new_n24690, new_n26053_1, new_n26054_1);
nor_5  g23706(new_n24713, new_n26054_1, new_n26055);
nor_5  g23707(new_n24687, new_n23243, new_n26056);
nor_5  g23708(new_n24712, new_n26056, new_n26057);
nor_5  g23709(new_n26057, new_n26055, n25337);
xnor_4 g23710(new_n12253, new_n11641, new_n26059);
xnor_4 g23711(new_n26059, new_n12260, n25356);
xnor_4 g23712(new_n9636, new_n9623, n25362);
xnor_4 g23713(new_n15629, new_n15606, n25412);
xnor_4 g23714(new_n16599, new_n16597, n25460);
xnor_4 g23715(new_n7874, new_n7835, n25468);
xnor_4 g23716(new_n15631, new_n15602_1, n25499);
xnor_4 g23717(new_n21458, new_n21457, n25513);
xnor_4 g23718(new_n13050, new_n13025, n25518);
xnor_4 g23719(new_n14416, new_n14375_1, n25532);
xnor_4 g23720(new_n21820_1, new_n21801, n25539);
xnor_4 g23721(new_n18323_1, new_n18314, n25550);
xnor_4 g23722(new_n22631_1, new_n22615, n25611);
xnor_4 g23723(new_n5713, new_n5712, new_n26072);
xnor_4 g23724(new_n26072, new_n5718, n25614);
xnor_4 g23725(new_n13745, new_n13718, n25619);
nand_5 g23726(new_n25684, new_n24815, new_n26075);
nand_5 g23727(new_n24968, new_n26075, new_n26076);
nand_5 g23728(new_n24961, new_n24964, new_n26077);
nand_5 g23729(new_n24967, new_n26077, new_n26078);
nand_5 g23730(new_n26078, new_n26076, new_n26079);
not_8  g23731(new_n26079, n25665);
xnor_4 g23732(new_n9828, new_n9802, n25706);
xnor_4 g23733(new_n24961, new_n21106, new_n26082);
xnor_4 g23734(new_n26082, new_n25689, n25719);
xor_4  g23735(new_n10370, new_n10318, n25756);
nand_5 g23736(new_n13998, new_n13957, new_n26085);
nand_5 g23737(new_n14042, new_n26085, new_n26086);
not_8  g23738(new_n13998, new_n26087);
nand_5 g23739(new_n26087, new_n13956, new_n26088);
nand_5 g23740(new_n14041, new_n26088, new_n26089);
nand_5 g23741(new_n26089, new_n26086, new_n26090);
not_8  g23742(new_n26090, n25758);
xnor_4 g23743(new_n16012, new_n6085, n25773);
xnor_4 g23744(new_n22403, new_n19137, n25784);
xnor_4 g23745(new_n8904, new_n8873, n25792);
xnor_4 g23746(new_n7350, new_n7311, n25816);
xnor_4 g23747(new_n6750, new_n6710, n25826);
xnor_4 g23748(new_n13268, new_n13266, n25839);
xnor_4 g23749(new_n15189, new_n15139_1, n25840);
xnor_4 g23750(new_n8703, new_n8670, n25873);
xnor_4 g23751(new_n25794, new_n25790, n25934);
xnor_4 g23752(new_n22858_1, new_n22842, n25938);
xnor_4 g23753(new_n23184, new_n23181, n25985);
xnor_4 g23754(new_n14971, new_n9625, n25994);
not_8  g23755(new_n19816, new_n26104);
nand_5 g23756(new_n26104, new_n19724, new_n26105);
nand_5 g23757(new_n19888, new_n19817, new_n26106);
nand_5 g23758(new_n26106, new_n26105, n26084);
xnor_4 g23759(new_n24709, new_n24695, n26096);
nand_5 g23760(new_n12458, new_n24945, new_n26109);
nor_5  g23761(new_n26109, new_n12370, n26111);
xnor_4 g23762(new_n12444, new_n12419, n26113);
xor_4  g23763(new_n21941, new_n21937, n26156);
xnor_4 g23764(new_n18545, new_n18522, n26159);
xnor_4 g23765(new_n3871_1, new_n3821, n26179);
xnor_4 g23766(new_n15174, new_n15173, n26220);
xnor_4 g23767(new_n24748, new_n24745, n26229);
xnor_4 g23768(new_n13663, new_n13626_1, n26237);
xnor_4 g23769(new_n17048, new_n17032, n26250);
not_8  g23770(new_n22899, new_n26119);
xnor_4 g23771(new_n22902, new_n26119, n26274);
xnor_4 g23772(new_n17052, new_n17022, n26287);
xnor_4 g23773(new_n23097, new_n22315, new_n26122);
xnor_4 g23774(new_n26122, new_n25597, n26317);
nand_5 g23775(new_n25315, new_n20175, new_n26124);
nand_5 g23776(new_n26124, new_n20191, new_n26125);
nand_5 g23777(new_n20195, new_n20173, new_n26126);
nand_5 g23778(new_n26126, new_n20190, new_n26127);
nand_5 g23779(new_n26127, new_n26125, new_n26128);
not_8  g23780(new_n26128, n26353);
xnor_4 g23781(new_n21995, new_n21988, n26375);
not_8  g23782(new_n25125, new_n26131);
nand_5 g23783(new_n26131, new_n25120_1, new_n26132);
nand_5 g23784(new_n25136, new_n25126_1, new_n26133);
nand_5 g23785(new_n26133, new_n26132, new_n26134);
not_8  g23786(new_n26134, n26396);
xnor_4 g23787(new_n5717, new_n5715, n26429);
xnor_4 g23788(new_n15703, new_n15687, n26431);
xnor_4 g23789(new_n7610_1, new_n7544, n26439);
xnor_4 g23790(new_n22239, new_n22238, n26492);
xnor_4 g23791(new_n10878, new_n10877, n26515);
xnor_4 g23792(new_n2562, new_n2531, n26538);
xnor_4 g23793(new_n16224, new_n16208, n26590);
xnor_4 g23794(new_n21043, new_n23857, n26598);
xnor_4 g23795(new_n25088, new_n23165, new_n26144);
xnor_4 g23796(new_n26144, new_n25094_1, n26605);
xnor_4 g23797(new_n25058, new_n25048, new_n26146);
xnor_4 g23798(new_n26146, new_n25052, n26656);
xnor_4 g23799(new_n12434, new_n12433, n26674);
xnor_4 g23800(new_n10221, new_n10203, n26675);
xnor_4 g23801(new_n22249, new_n22218, n26681);
nor_5  g23802(new_n5997, new_n5786, new_n26151);
nor_5  g23803(new_n6080, new_n26151, new_n26152);
nor_5  g23804(new_n24613, new_n5785, new_n26153);
nor_5  g23805(new_n6079, new_n26153, new_n26154);
nor_5  g23806(new_n26154, new_n26152, n26696);
xnor_4 g23807(new_n15969, new_n15951, n26698);
xnor_4 g23808(new_n16744, new_n6114, n26707);
xnor_4 g23809(new_n25534, new_n25532_1, n26719);
xnor_4 g23810(new_n9824, new_n9810, n26727);
nor_5  g23811(new_n23243, new_n20861, new_n26160);
not_8  g23812(new_n23244, new_n26161);
nor_5  g23813(new_n23248_1, new_n26161, new_n26162);
nor_5  g23814(new_n26162, new_n26160, n26729);
not_8  g23815(new_n23267, new_n26164);
xnor_4 g23816(new_n23271, new_n26164, n26745);
xnor_4 g23817(new_n8404, new_n8363_1, n26775);
xnor_4 g23818(new_n11277, new_n11257, n26780);
xnor_4 g23819(new_n23744, new_n23736, n26794);
xnor_4 g23820(new_n3515, new_n3453, n26795);
xnor_4 g23821(new_n11568, new_n11521, n26801);
xnor_4 g23822(new_n11965_1, new_n11944, n26815);
xnor_4 g23823(new_n25193, new_n25190, n26847);
xnor_4 g23824(new_n20195, new_n7808, new_n26173);
xnor_4 g23825(new_n26173, new_n25320, n26900);
xor_4  g23826(new_n20355_1, new_n20353, n26902);
xor_4  g23827(new_n18814, new_n18809, n26905);
xnor_4 g23828(new_n8705, new_n8664, n26921);
xnor_4 g23829(new_n24136, new_n24122, n26923);
xnor_4 g23830(new_n11661, new_n11660, n26929);
xnor_4 g23831(new_n13674, new_n13601, n26930);
xnor_4 g23832(new_n17050, new_n17027, n26943);
xnor_4 g23833(new_n15633, new_n15598_1, n26970);
xnor_4 g23834(new_n22785, new_n22771, n27004);
xnor_4 g23835(new_n11169, new_n11095, n27011);
xnor_4 g23836(new_n21063, new_n21004, n27019);
xnor_4 g23837(new_n5278, new_n5264, n27031);
xnor_4 g23838(new_n23800, new_n22896, new_n26187);
xnor_4 g23839(new_n26187, new_n23848, n27051);
xor_4  g23840(new_n18675, new_n18671, n27072);
xnor_4 g23841(new_n16614, new_n16558, n27079);
xnor_4 g23842(new_n4491, new_n4489, n27096);
xnor_4 g23843(new_n15358, new_n15346, n27110);
xnor_4 g23844(new_n14731, new_n14728, n27112);
xnor_4 g23845(new_n24142, new_n23609, n27130);
xnor_4 g23846(new_n17443, new_n17432_1, n27145);
nor_5  g23847(new_n17902, new_n17281, new_n26196);
not_8  g23848(new_n23435, new_n26197);
nor_5  g23849(new_n23438, new_n26197, new_n26198);
nor_5  g23850(new_n26198, new_n26196, n27158);
xnor_4 g23851(new_n23016, new_n23013, n27163);
xnor_4 g23852(new_n25346, new_n22825, new_n26201);
xnor_4 g23853(new_n26201, new_n25352, n27194);
endmodule


