// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Thu Jun 27 02:29:38 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095,
    new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269_1, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1318,
    new_n1319, new_n1320, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333_1, new_n1334, new_n1335, new_n1336, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355, new_n1356,
    new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471_1, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1561,
    new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1,
    new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389,
    new_n2390, new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1,
    new_n2432, new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1, new_n2510,
    new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339_1, new_n3340, new_n3341, new_n3342_1, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986_1, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992_1, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005_1,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086_1, new_n4087, new_n4088_1, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094_1, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155_1, new_n4156,
    new_n4157, new_n4158, new_n4159_1, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187_1, new_n4188, new_n4189_1, new_n4190_1, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203_1, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226_1, new_n4227, new_n4228,
    new_n4229, new_n4230_1, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300_1, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312_1, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326_1, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333_1, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370_1, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378_1, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397_1,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436_1, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499_1,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516_1, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553_1,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4609, new_n4610, new_n4611, new_n4612, new_n4613,
    new_n4614, new_n4615, new_n4616, new_n4617, new_n4618, new_n4619,
    new_n4620, new_n4621, new_n4622, new_n4623, new_n4624, new_n4625,
    new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4632,
    new_n4633, new_n4634_1, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686_1, new_n4687, new_n4688, new_n4689_1,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733_1, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757_1, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805_1, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817_1, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826_1, new_n4827,
    new_n4828_1, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212_1, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314_1, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1,
    new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481,
    new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487,
    new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493,
    new_n5494, new_n5495, new_n5496, new_n5497, new_n5498, new_n5499,
    new_n5500, new_n5501, new_n5502, new_n5503, new_n5504, new_n5505,
    new_n5506, new_n5507, new_n5508, new_n5509, new_n5510, new_n5511,
    new_n5512, new_n5513, new_n5514, new_n5515, new_n5516, new_n5517,
    new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523,
    new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529,
    new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535,
    new_n5536, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541,
    new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547,
    new_n5548, new_n5549, new_n5550, new_n5551, new_n5552, new_n5553,
    new_n5554, new_n5555, new_n5556, new_n5557, new_n5558, new_n5559,
    new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565,
    new_n5566, new_n5567, new_n5568, new_n5569, new_n5570, new_n5571,
    new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577,
    new_n5578, new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583,
    new_n5584, new_n5585, new_n5586, new_n5587, new_n5588, new_n5589,
    new_n5590, new_n5591, new_n5592, new_n5593, new_n5594, new_n5595,
    new_n5596, new_n5597, new_n5598, new_n5599, new_n5600, new_n5601,
    new_n5602, new_n5603, new_n5604, new_n5605, new_n5606, new_n5607,
    new_n5608, new_n5609, new_n5610, new_n5611, new_n5612, new_n5613,
    new_n5614, new_n5615, new_n5616, new_n5617, new_n5618, new_n5619,
    new_n5620, new_n5621, new_n5622, new_n5623, new_n5624, new_n5625,
    new_n5626, new_n5627, new_n5628, new_n5629, new_n5630, new_n5631,
    new_n5632, new_n5633, new_n5634, new_n5635, new_n5636, new_n5637,
    new_n5638, new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643,
    new_n5644, new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649,
    new_n5650, new_n5651, new_n5652, new_n5653, new_n5654, new_n5655,
    new_n5656, new_n5657, new_n5658, new_n5659, new_n5660, new_n5661,
    new_n5662, new_n5663, new_n5664, new_n5665, new_n5666, new_n5667,
    new_n5668, new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673,
    new_n5674, new_n5675, new_n5676, new_n5677, new_n5678, new_n5679,
    new_n5680, new_n5681, new_n5682, new_n5683, new_n5684, new_n5685,
    new_n5686, new_n5687, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859, new_n5860_1,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934_1, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6005, new_n6006, new_n6007, new_n6008, new_n6009, new_n6010,
    new_n6011, new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1,
    new_n6017, new_n6018, new_n6019, new_n6020, new_n6021, new_n6022,
    new_n6023, new_n6024, new_n6025, new_n6026, new_n6027, new_n6028,
    new_n6029, new_n6030, new_n6031, new_n6032, new_n6033, new_n6034,
    new_n6035, new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040,
    new_n6041, new_n6042, new_n6043, new_n6044, new_n6045, new_n6046,
    new_n6047, new_n6048, new_n6049, new_n6050, new_n6051, new_n6052,
    new_n6053, new_n6054, new_n6055, new_n6056, new_n6057, new_n6058,
    new_n6059, new_n6060, new_n6061, new_n6062, new_n6063, new_n6064,
    new_n6065, new_n6066, new_n6067, new_n6068, new_n6069, new_n6070,
    new_n6071, new_n6072, new_n6073, new_n6074, new_n6075, new_n6076,
    new_n6077, new_n6078, new_n6079, new_n6080, new_n6081, new_n6082,
    new_n6083, new_n6084, new_n6085, new_n6086, new_n6087, new_n6088,
    new_n6089_1, new_n6090, new_n6091, new_n6092, new_n6093, new_n6094,
    new_n6095, new_n6096, new_n6097, new_n6098, new_n6099, new_n6100,
    new_n6101, new_n6102, new_n6103, new_n6104, new_n6105, new_n6106,
    new_n6107, new_n6108, new_n6109, new_n6110, new_n6111, new_n6112,
    new_n6113, new_n6114, new_n6115, new_n6116, new_n6117, new_n6118,
    new_n6119, new_n6120, new_n6121, new_n6122, new_n6123, new_n6124,
    new_n6125, new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130,
    new_n6131, new_n6132, new_n6133, new_n6134, new_n6135, new_n6136,
    new_n6137, new_n6138, new_n6139, new_n6140, new_n6141, new_n6142,
    new_n6143, new_n6144, new_n6145, new_n6146, new_n6147, new_n6148,
    new_n6149, new_n6150, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160,
    new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166,
    new_n6167, new_n6168, new_n6169, new_n6170, new_n6171, new_n6172,
    new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178,
    new_n6179, new_n6180, new_n6181, new_n6182, new_n6183, new_n6184,
    new_n6185, new_n6186, new_n6187, new_n6188, new_n6189, new_n6190,
    new_n6191, new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204, new_n6205, new_n6206, new_n6207, new_n6208,
    new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214,
    new_n6215, new_n6216, new_n6217, new_n6218, new_n6219, new_n6220,
    new_n6221, new_n6222, new_n6223, new_n6224, new_n6225, new_n6226,
    new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232,
    new_n6233, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238,
    new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254_1, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273_1, new_n6274, new_n6275,
    new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6288, new_n6289, new_n6290, new_n6291, new_n6292, new_n6293,
    new_n6294_1, new_n6295, new_n6296, new_n6297, new_n6298, new_n6299,
    new_n6300, new_n6301, new_n6302, new_n6303, new_n6304, new_n6305,
    new_n6306, new_n6307, new_n6308, new_n6309, new_n6310, new_n6311,
    new_n6312, new_n6313, new_n6314, new_n6315, new_n6316, new_n6317,
    new_n6318, new_n6319, new_n6320, new_n6321, new_n6322, new_n6323,
    new_n6324, new_n6325, new_n6326, new_n6327, new_n6328, new_n6329,
    new_n6330, new_n6331, new_n6332, new_n6333, new_n6334, new_n6335,
    new_n6336, new_n6337, new_n6338, new_n6339, new_n6340, new_n6341,
    new_n6342, new_n6343, new_n6344, new_n6345, new_n6346, new_n6347,
    new_n6348, new_n6349, new_n6350, new_n6351, new_n6352, new_n6353,
    new_n6354, new_n6355, new_n6356, new_n6357, new_n6358_1, new_n6359_1,
    new_n6360, new_n6361, new_n6362, new_n6363, new_n6364, new_n6365,
    new_n6366, new_n6367, new_n6368, new_n6369, new_n6370, new_n6371,
    new_n6372, new_n6373, new_n6374, new_n6375, new_n6376, new_n6377,
    new_n6378, new_n6379, new_n6380, new_n6381, new_n6382, new_n6383,
    new_n6384, new_n6385, new_n6386, new_n6387, new_n6388, new_n6389,
    new_n6390, new_n6391, new_n6392, new_n6393, new_n6394, new_n6395,
    new_n6396, new_n6397, new_n6398, new_n6399, new_n6400, new_n6401,
    new_n6402, new_n6403, new_n6404, new_n6405, new_n6406, new_n6407,
    new_n6408, new_n6409, new_n6410, new_n6411, new_n6412, new_n6413,
    new_n6414, new_n6415, new_n6416, new_n6417, new_n6418, new_n6419,
    new_n6420, new_n6421, new_n6422, new_n6423, new_n6424, new_n6425,
    new_n6426, new_n6427, new_n6428, new_n6429_1, new_n6430, new_n6431_1,
    new_n6432, new_n6433, new_n6434, new_n6435, new_n6436, new_n6437,
    new_n6438, new_n6439, new_n6440, new_n6441_1, new_n6442, new_n6443,
    new_n6444, new_n6445_1, new_n6446, new_n6447, new_n6448, new_n6449,
    new_n6450, new_n6451, new_n6452, new_n6453, new_n6454, new_n6455,
    new_n6456, new_n6457, new_n6458, new_n6459, new_n6460, new_n6461,
    new_n6462, new_n6463, new_n6464, new_n6465, new_n6466, new_n6467,
    new_n6468, new_n6469, new_n6470, new_n6471, new_n6472, new_n6473,
    new_n6474, new_n6475, new_n6476, new_n6477, new_n6478, new_n6479,
    new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502, new_n6503,
    new_n6504, new_n6505, new_n6506, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513, new_n6514, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556, new_n6557,
    new_n6558, new_n6559, new_n6560, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576, new_n6577, new_n6578_1, new_n6579, new_n6580, new_n6581,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604_1, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611_1, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618,
    new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624,
    new_n6625, new_n6626, new_n6627, new_n6628, new_n6629, new_n6630,
    new_n6631, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645_1, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687_1, new_n6688, new_n6689_1, new_n6690,
    new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703_1, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720,
    new_n6721, new_n6722, new_n6723, new_n6724, new_n6725, new_n6726,
    new_n6727, new_n6728, new_n6729, new_n6730, new_n6731, new_n6732,
    new_n6733, new_n6734, new_n6735, new_n6736, new_n6737, new_n6738,
    new_n6739, new_n6740, new_n6741, new_n6742_1, new_n6743, new_n6744,
    new_n6745, new_n6746, new_n6747, new_n6748, new_n6749, new_n6750,
    new_n6751, new_n6752, new_n6753, new_n6754, new_n6755, new_n6756,
    new_n6757, new_n6758, new_n6759, new_n6760, new_n6761, new_n6762,
    new_n6763, new_n6764, new_n6765, new_n6766, new_n6767, new_n6768,
    new_n6769, new_n6770_1, new_n6771, new_n6772, new_n6773, new_n6774,
    new_n6775, new_n6776_1, new_n6777, new_n6778, new_n6779, new_n6780,
    new_n6781, new_n6782, new_n6783, new_n6784, new_n6785, new_n6786,
    new_n6787, new_n6788, new_n6789, new_n6790, new_n6791, new_n6792,
    new_n6793, new_n6794, new_n6795, new_n6796, new_n6797_1, new_n6798,
    new_n6800, new_n6801, new_n6802, new_n6803, new_n6804, new_n6805,
    new_n6806_1, new_n6807, new_n6808, new_n6809_1, new_n6810, new_n6811,
    new_n6812, new_n6813, new_n6814, new_n6815, new_n6816, new_n6817,
    new_n6818, new_n6819, new_n6820, new_n6821, new_n6822_1, new_n6823,
    new_n6824, new_n6825, new_n6826_1, new_n6827, new_n6828, new_n6829,
    new_n6830, new_n6831, new_n6832, new_n6833, new_n6834, new_n6835,
    new_n6836, new_n6837, new_n6838, new_n6839, new_n6840, new_n6841,
    new_n6842, new_n6843, new_n6844, new_n6845, new_n6846, new_n6847,
    new_n6849, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860_1, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877_1, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986_1, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159_1, new_n7160_1, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193_1, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233,
    new_n7234, new_n7235, new_n7236_1, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265_1, new_n7266, new_n7267, new_n7268, new_n7269,
    new_n7270_1, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277, new_n7278, new_n7279, new_n7280, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294_1, new_n7295, new_n7296, new_n7297, new_n7298, new_n7299,
    new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305,
    new_n7306, new_n7307, new_n7308, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320_1, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523_1,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8006, new_n8010, new_n8012, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028_1, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100_1, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202_1, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261,
    new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267,
    new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273,
    new_n8274, new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279,
    new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285,
    new_n8286, new_n8287, new_n8288, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303_1,
    new_n8304, new_n8305, new_n8306, new_n8307, new_n8308, new_n8309,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321,
    new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336_1, new_n8337, new_n8338, new_n8339,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381,
    new_n8382, new_n8383, new_n8384_1, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398_1, new_n8399,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405,
    new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417,
    new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423,
    new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432, new_n8433_1, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595_1, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8639, new_n8640,
    new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646,
    new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652,
    new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658,
    new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664,
    new_n8665_1, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717_1, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759_1, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819_1, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8825, new_n8827, new_n8829,
    new_n8830, new_n8831, new_n8832, new_n8833, new_n8834, new_n8835,
    new_n8836, new_n8837, new_n8838, new_n8839, new_n8841, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927,
    new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933,
    new_n8934, new_n8935, new_n8936, new_n8937, new_n8938, new_n8939,
    new_n8940, new_n8941, new_n8942, new_n8943, new_n8944, new_n8945,
    new_n8946, new_n8947, new_n8948, new_n8949, new_n8950, new_n8951,
    new_n8952, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080_1,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111_1, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137_1, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189_1, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195_1, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241_1, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338,
    new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9344,
    new_n9345, new_n9346, new_n9347, new_n9348, new_n9349, new_n9350,
    new_n9351, new_n9352, new_n9353, new_n9354, new_n9355, new_n9356,
    new_n9357, new_n9358, new_n9359, new_n9360, new_n9361, new_n9362,
    new_n9363, new_n9364, new_n9365, new_n9366, new_n9367, new_n9368,
    new_n9369, new_n9370, new_n9371, new_n9372, new_n9373, new_n9374,
    new_n9375, new_n9376, new_n9377, new_n9378, new_n9379, new_n9380,
    new_n9381, new_n9382, new_n9383, new_n9384, new_n9385, new_n9386,
    new_n9387_1, new_n9388, new_n9389, new_n9390, new_n9391, new_n9392,
    new_n9393, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398,
    new_n9399, new_n9400_1, new_n9401, new_n9402, new_n9403, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422,
    new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457_1, new_n9458,
    new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9568, new_n9569, new_n9570, new_n9571_1, new_n9572,
    new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578_1,
    new_n9579, new_n9580, new_n9581, new_n9582, new_n9583_1, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633, new_n9634, new_n9635, new_n9636, new_n9637_1, new_n9638,
    new_n9639, new_n9640_1, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668,
    new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674,
    new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680,
    new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686,
    new_n9687, new_n9688, new_n9689, new_n9690, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706_1, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725_1,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756_1, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820_1, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920_1, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956_1, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022_1, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174_1, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217_1, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223_1, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277,
    new_n10278_1, new_n10279, new_n10280, new_n10281, new_n10282,
    new_n10283, new_n10284, new_n10285, new_n10286, new_n10287, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300,
    new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306,
    new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312,
    new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318,
    new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326, new_n10327_1, new_n10328, new_n10329,
    new_n10330, new_n10331, new_n10332, new_n10333, new_n10334, new_n10335,
    new_n10336, new_n10337, new_n10338, new_n10339, new_n10340, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345, new_n10346, new_n10347,
    new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383,
    new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389,
    new_n10390, new_n10391_1, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400,
    new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406,
    new_n10407, new_n10408, new_n10409, new_n10410, new_n10411, new_n10412,
    new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418,
    new_n10419, new_n10420, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432, new_n10433, new_n10434, new_n10435, new_n10436,
    new_n10437, new_n10438, new_n10439_1, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451_1, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475,
    new_n10476_1, new_n10477, new_n10478, new_n10479, new_n10480,
    new_n10481, new_n10482, new_n10483, new_n10484, new_n10485, new_n10486,
    new_n10487, new_n10488, new_n10489, new_n10490, new_n10491, new_n10492,
    new_n10493, new_n10494, new_n10495, new_n10496, new_n10497, new_n10498,
    new_n10499, new_n10500, new_n10501, new_n10502, new_n10503, new_n10504,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509,
    new_n10510_1, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520,
    new_n10521, new_n10522, new_n10523, new_n10524, new_n10525, new_n10526,
    new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545_1, new_n10546, new_n10547_1, new_n10548, new_n10549,
    new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555,
    new_n10556, new_n10557, new_n10558, new_n10559, new_n10560, new_n10561,
    new_n10562, new_n10563, new_n10564, new_n10565, new_n10566, new_n10567,
    new_n10568, new_n10569, new_n10570, new_n10571, new_n10572, new_n10573,
    new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579,
    new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585,
    new_n10586, new_n10587, new_n10588, new_n10589_1, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644_1, new_n10645, new_n10646, new_n10647, new_n10648,
    new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654,
    new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10677, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685_1,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695_1, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789_1, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848_1, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898_1, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913_1,
    new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10928_1, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949_1, new_n10950, new_n10951, new_n10952, new_n10953,
    new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959,
    new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965_1, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10990_1, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023_1, new_n11024, new_n11025, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045,
    new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051,
    new_n11052, new_n11053, new_n11054, new_n11055, new_n11056, new_n11057,
    new_n11058, new_n11059, new_n11060, new_n11061, new_n11062, new_n11063,
    new_n11064, new_n11065, new_n11066, new_n11067, new_n11068, new_n11069,
    new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11095, new_n11096, new_n11097, new_n11098, new_n11099,
    new_n11100, new_n11101, new_n11102, new_n11103, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120, new_n11121, new_n11122, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129,
    new_n11130, new_n11131, new_n11132, new_n11133, new_n11134, new_n11135,
    new_n11136, new_n11137, new_n11138, new_n11139, new_n11140, new_n11141,
    new_n11142, new_n11143, new_n11144, new_n11145, new_n11146, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153_1, new_n11154, new_n11155, new_n11156, new_n11157,
    new_n11158, new_n11159, new_n11160, new_n11161, new_n11162, new_n11163,
    new_n11164, new_n11165, new_n11166, new_n11167, new_n11168, new_n11169,
    new_n11170, new_n11171, new_n11172, new_n11173, new_n11174, new_n11175,
    new_n11176, new_n11177, new_n11178, new_n11179, new_n11180, new_n11181,
    new_n11182, new_n11183, new_n11184, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201, new_n11202, new_n11203, new_n11204, new_n11205,
    new_n11206, new_n11207, new_n11208, new_n11209, new_n11210, new_n11211,
    new_n11212, new_n11213, new_n11214, new_n11215, new_n11216_1,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221,
    new_n11222_1, new_n11223, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238,
    new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244,
    new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257_1, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311_1, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326_1, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407_1,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423_1, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478_1, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536_1, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11592, new_n11594, new_n11596, new_n11597,
    new_n11598, new_n11599, new_n11600, new_n11601, new_n11602, new_n11603,
    new_n11604, new_n11605, new_n11606, new_n11607, new_n11608, new_n11609,
    new_n11610, new_n11611, new_n11612, new_n11613, new_n11614, new_n11615,
    new_n11616, new_n11617, new_n11618, new_n11619, new_n11620, new_n11621,
    new_n11622, new_n11623, new_n11624, new_n11625, new_n11626, new_n11627,
    new_n11628, new_n11629, new_n11630, new_n11631, new_n11632, new_n11633,
    new_n11634, new_n11635, new_n11636, new_n11637, new_n11638, new_n11639,
    new_n11640, new_n11641, new_n11642, new_n11643, new_n11644, new_n11645,
    new_n11646, new_n11647, new_n11648, new_n11649, new_n11650, new_n11651,
    new_n11652, new_n11653, new_n11654, new_n11655, new_n11656, new_n11657,
    new_n11658, new_n11659, new_n11660, new_n11661, new_n11662_1,
    new_n11663, new_n11664, new_n11665, new_n11666, new_n11667, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673, new_n11674,
    new_n11675, new_n11676, new_n11677, new_n11678, new_n11679, new_n11680,
    new_n11681, new_n11682, new_n11683, new_n11684, new_n11685, new_n11686,
    new_n11687, new_n11688, new_n11689, new_n11690, new_n11691, new_n11692,
    new_n11693, new_n11694, new_n11695, new_n11696, new_n11697, new_n11698,
    new_n11699, new_n11700, new_n11701, new_n11702, new_n11703, new_n11704,
    new_n11705, new_n11706, new_n11707_1, new_n11708, new_n11709,
    new_n11710, new_n11711, new_n11712, new_n11713, new_n11715, new_n11716,
    new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722,
    new_n11723, new_n11724, new_n11725, new_n11726, new_n11727,
    new_n11728_1, new_n11729, new_n11730, new_n11731, new_n11732,
    new_n11733, new_n11734, new_n11735, new_n11736, new_n11737, new_n11738,
    new_n11739, new_n11740, new_n11741, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749, new_n11750,
    new_n11751, new_n11752, new_n11753, new_n11754, new_n11755_1,
    new_n11756, new_n11757_1, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780_1, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11790, new_n11791_1, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11817, new_n11818,
    new_n11819, new_n11820, new_n11821_1, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876_1,
    new_n11877_1, new_n11878, new_n11879, new_n11880, new_n11881,
    new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887,
    new_n11888, new_n11889, new_n11890, new_n11891, new_n11892_1,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917_1, new_n11918, new_n11919_1, new_n11920, new_n11921,
    new_n11922_1, new_n11923, new_n11924, new_n11925, new_n11926,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956,
    new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962,
    new_n11963, new_n11964, new_n11965, new_n11966, new_n11967_1,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999_1, new_n12000_1, new_n12001, new_n12002,
    new_n12003, new_n12004, new_n12005_1, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014_1, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020_1, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025_1, new_n12026, new_n12027, new_n12028,
    new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044_1, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069_1, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076_1, new_n12077, new_n12078,
    new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108,
    new_n12109, new_n12110, new_n12111_1, new_n12112, new_n12113,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121, new_n12122, new_n12123, new_n12124, new_n12125,
    new_n12126, new_n12127, new_n12128, new_n12129, new_n12130, new_n12131,
    new_n12132, new_n12133, new_n12134, new_n12135, new_n12136, new_n12137,
    new_n12138, new_n12139, new_n12140, new_n12141, new_n12142, new_n12143,
    new_n12144, new_n12145_1, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221_1, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247_1, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299_1, new_n12300, new_n12301,
    new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315, new_n12316, new_n12317, new_n12318, new_n12319,
    new_n12320, new_n12321, new_n12322, new_n12323, new_n12324, new_n12325,
    new_n12326, new_n12327, new_n12328, new_n12329, new_n12330, new_n12331,
    new_n12332, new_n12333, new_n12334, new_n12335, new_n12336, new_n12337,
    new_n12338, new_n12339, new_n12340, new_n12341, new_n12342, new_n12343,
    new_n12344, new_n12345, new_n12346, new_n12347, new_n12348, new_n12349,
    new_n12350, new_n12351, new_n12352, new_n12353, new_n12354, new_n12355,
    new_n12356, new_n12357, new_n12358, new_n12359, new_n12360, new_n12361,
    new_n12362, new_n12363, new_n12364, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380, new_n12381, new_n12382, new_n12383, new_n12384, new_n12385,
    new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391_1, new_n12392, new_n12393, new_n12394, new_n12395,
    new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413,
    new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444_1, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489_1,
    new_n12490, new_n12491, new_n12492, new_n12493, new_n12494, new_n12495,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506, new_n12507,
    new_n12508, new_n12509, new_n12510, new_n12511_1, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540, new_n12541, new_n12542,
    new_n12543, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554,
    new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560,
    new_n12561, new_n12562, new_n12563, new_n12564, new_n12565, new_n12566,
    new_n12567, new_n12568, new_n12569, new_n12570, new_n12571, new_n12572,
    new_n12573, new_n12574, new_n12575, new_n12576, new_n12577, new_n12578,
    new_n12579, new_n12580, new_n12581, new_n12582, new_n12583, new_n12584,
    new_n12585, new_n12586, new_n12587, new_n12588, new_n12589, new_n12590,
    new_n12591_1, new_n12592, new_n12593, new_n12594, new_n12595,
    new_n12596, new_n12597, new_n12598, new_n12599, new_n12600, new_n12601,
    new_n12602, new_n12603, new_n12604, new_n12605, new_n12606, new_n12607,
    new_n12608, new_n12609, new_n12610, new_n12611, new_n12618, new_n12623,
    new_n12625, new_n12626, new_n12627, new_n12628, new_n12629, new_n12630,
    new_n12631, new_n12632, new_n12633, new_n12634, new_n12635, new_n12636,
    new_n12637, new_n12638, new_n12639, new_n12640, new_n12641, new_n12642,
    new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648_1, new_n12649, new_n12650, new_n12651, new_n12652,
    new_n12653, new_n12654, new_n12655, new_n12656, new_n12657, new_n12658,
    new_n12659, new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665, new_n12666, new_n12667, new_n12668, new_n12669, new_n12670,
    new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676,
    new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682,
    new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688,
    new_n12689, new_n12690, new_n12691, new_n12692, new_n12693, new_n12694,
    new_n12695, new_n12696, new_n12697, new_n12698, new_n12699, new_n12700,
    new_n12701, new_n12702, new_n12703, new_n12704_1, new_n12705_1,
    new_n12706_1, new_n12707, new_n12708, new_n12709_1, new_n12710,
    new_n12711, new_n12712, new_n12713, new_n12714, new_n12715, new_n12716,
    new_n12717, new_n12718, new_n12719, new_n12720_1, new_n12721,
    new_n12722, new_n12723, new_n12724, new_n12725, new_n12726, new_n12727,
    new_n12728, new_n12729, new_n12730, new_n12731, new_n12732, new_n12733,
    new_n12734, new_n12735, new_n12736, new_n12737, new_n12738, new_n12739,
    new_n12740, new_n12741, new_n12742, new_n12743, new_n12744, new_n12745,
    new_n12746, new_n12747, new_n12748, new_n12749, new_n12750, new_n12751,
    new_n12752, new_n12753_1, new_n12754, new_n12755, new_n12756,
    new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762,
    new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768,
    new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774,
    new_n12775, new_n12776, new_n12777_1, new_n12778, new_n12779,
    new_n12780, new_n12781, new_n12782, new_n12783, new_n12784, new_n12785,
    new_n12786, new_n12787, new_n12788, new_n12789, new_n12790, new_n12791,
    new_n12792, new_n12793, new_n12794, new_n12795, new_n12796, new_n12797,
    new_n12798, new_n12799, new_n12800, new_n12801, new_n12802, new_n12803,
    new_n12804, new_n12805, new_n12806, new_n12807_1, new_n12808,
    new_n12809, new_n12810, new_n12811, new_n12812, new_n12813, new_n12814,
    new_n12815, new_n12816, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925_1,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947_1, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12995, new_n12996, new_n12997, new_n12998,
    new_n12999, new_n13000, new_n13001, new_n13002, new_n13003, new_n13004,
    new_n13005, new_n13006, new_n13007, new_n13008, new_n13009, new_n13010,
    new_n13011, new_n13012, new_n13013, new_n13014, new_n13015, new_n13016,
    new_n13017, new_n13018, new_n13019, new_n13020, new_n13021, new_n13022,
    new_n13023, new_n13024, new_n13025, new_n13026, new_n13027, new_n13028,
    new_n13029, new_n13030, new_n13031, new_n13032, new_n13033, new_n13034,
    new_n13035, new_n13036, new_n13037, new_n13038, new_n13039, new_n13040,
    new_n13041, new_n13042, new_n13043, new_n13044, new_n13045, new_n13046,
    new_n13047, new_n13048, new_n13049, new_n13050, new_n13051, new_n13052,
    new_n13053, new_n13054, new_n13055, new_n13056, new_n13057, new_n13058,
    new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064,
    new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13072, new_n13073, new_n13074, new_n13075, new_n13076,
    new_n13077, new_n13078, new_n13079, new_n13080, new_n13081, new_n13082,
    new_n13083, new_n13084, new_n13085, new_n13086, new_n13087, new_n13088,
    new_n13089, new_n13090, new_n13091, new_n13092, new_n13093, new_n13094,
    new_n13095, new_n13096, new_n13097, new_n13098, new_n13099, new_n13100,
    new_n13101, new_n13102, new_n13103, new_n13104, new_n13105, new_n13106,
    new_n13107, new_n13108, new_n13109, new_n13110, new_n13111, new_n13112,
    new_n13113, new_n13114, new_n13115, new_n13116, new_n13117, new_n13118,
    new_n13119, new_n13120, new_n13121, new_n13122, new_n13123, new_n13124,
    new_n13125, new_n13126, new_n13127, new_n13128, new_n13129, new_n13130,
    new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137, new_n13138, new_n13139, new_n13140, new_n13141, new_n13142,
    new_n13143, new_n13144, new_n13145, new_n13146, new_n13147, new_n13148,
    new_n13149, new_n13150, new_n13151, new_n13152, new_n13153, new_n13154,
    new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160,
    new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166,
    new_n13167, new_n13168, new_n13169, new_n13170, new_n13171, new_n13172,
    new_n13173, new_n13174, new_n13175, new_n13176, new_n13177, new_n13178,
    new_n13179, new_n13180, new_n13181, new_n13184, new_n13188, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198,
    new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210,
    new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13216,
    new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222,
    new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228,
    new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234,
    new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240,
    new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252,
    new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258,
    new_n13259, new_n13260, new_n13261, new_n13262, new_n13263, new_n13264,
    new_n13265, new_n13266, new_n13267, new_n13268, new_n13269, new_n13270,
    new_n13271, new_n13272, new_n13273, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294,
    new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312,
    new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318,
    new_n13319, new_n13320, new_n13321, new_n13322, new_n13323, new_n13324,
    new_n13325, new_n13326, new_n13327, new_n13328, new_n13329, new_n13330,
    new_n13331, new_n13332, new_n13333, new_n13334, new_n13335, new_n13336,
    new_n13337, new_n13338, new_n13339, new_n13340, new_n13341, new_n13342,
    new_n13343, new_n13344, new_n13345, new_n13346, new_n13347, new_n13348,
    new_n13349, new_n13350, new_n13351, new_n13352, new_n13353, new_n13354,
    new_n13355, new_n13356, new_n13357, new_n13358, new_n13359, new_n13360,
    new_n13361, new_n13362, new_n13363, new_n13364, new_n13365, new_n13366,
    new_n13367, new_n13368, new_n13369, new_n13370, new_n13371, new_n13372,
    new_n13373, new_n13374, new_n13375, new_n13376, new_n13377, new_n13378,
    new_n13379, new_n13380, new_n13381, new_n13382, new_n13383, new_n13384,
    new_n13385, new_n13386, new_n13387, new_n13388, new_n13389, new_n13390,
    new_n13391, new_n13392, new_n13393, new_n13394, new_n13395, new_n13396,
    new_n13397, new_n13398, new_n13399, new_n13400, new_n13401, new_n13402,
    new_n13403, new_n13404, new_n13405, new_n13406, new_n13407, new_n13408,
    new_n13409, new_n13410, new_n13411, new_n13412, new_n13413, new_n13414,
    new_n13415, new_n13416, new_n13417, new_n13418, new_n13419, new_n13420,
    new_n13421, new_n13422, new_n13423, new_n13424, new_n13425, new_n13426,
    new_n13427, new_n13428, new_n13429, new_n13430, new_n13431, new_n13432,
    new_n13433, new_n13434, new_n13435, new_n13436, new_n13437, new_n13438,
    new_n13439, new_n13440, new_n13441, new_n13442, new_n13443, new_n13444,
    new_n13445, new_n13446, new_n13447, new_n13448, new_n13449, new_n13450,
    new_n13451, new_n13452, new_n13453, new_n13454, new_n13455, new_n13456,
    new_n13457, new_n13458, new_n13459, new_n13460, new_n13461, new_n13462,
    new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468,
    new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474,
    new_n13475, new_n13476, new_n13477, new_n13478, new_n13479, new_n13480,
    new_n13481, new_n13482, new_n13483, new_n13484, new_n13485, new_n13486,
    new_n13487, new_n13488, new_n13489, new_n13490, new_n13491, new_n13492,
    new_n13493, new_n13494, new_n13495, new_n13496, new_n13497, new_n13498,
    new_n13499, new_n13500, new_n13501, new_n13502, new_n13503, new_n13504,
    new_n13505, new_n13506, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534,
    new_n13535, new_n13536, new_n13537, new_n13538, new_n13539, new_n13540,
    new_n13541, new_n13542, new_n13543, new_n13544, new_n13545, new_n13546,
    new_n13547, new_n13548, new_n13549, new_n13550, new_n13551, new_n13552,
    new_n13553, new_n13554, new_n13555, new_n13556, new_n13557, new_n13558,
    new_n13559, new_n13560, new_n13561, new_n13562, new_n13563, new_n13564,
    new_n13565, new_n13566, new_n13567, new_n13568, new_n13569, new_n13570,
    new_n13571, new_n13572, new_n13573, new_n13574, new_n13575, new_n13576,
    new_n13577, new_n13578, new_n13579, new_n13580, new_n13581, new_n13582,
    new_n13583, new_n13586, new_n13589, new_n13594, new_n13596, new_n13599,
    new_n13601, new_n13602, new_n13603, new_n13604, new_n13605, new_n13606,
    new_n13607, new_n13608, new_n13609, new_n13610, new_n13611, new_n13612,
    new_n13613, new_n13614, new_n13615, new_n13616, new_n13617, new_n13618,
    new_n13619, new_n13620, new_n13621, new_n13622, new_n13623, new_n13624,
    new_n13625, new_n13626, new_n13627, new_n13628, new_n13629, new_n13630,
    new_n13631, new_n13632, new_n13633, new_n13634, new_n13635, new_n13636,
    new_n13637, new_n13638, new_n13639, new_n13640, new_n13641, new_n13642,
    new_n13643, new_n13644, new_n13645, new_n13646, new_n13647, new_n13648,
    new_n13649, new_n13650, new_n13651, new_n13652, new_n13653, new_n13654,
    new_n13655, new_n13656, new_n13657, new_n13658, new_n13659, new_n13660,
    new_n13661, new_n13662, new_n13663, new_n13664, new_n13665, new_n13666,
    new_n13667, new_n13668, new_n13669, new_n13670, new_n13671, new_n13672,
    new_n13673, new_n13674, new_n13675, new_n13676, new_n13677, new_n13678,
    new_n13679, new_n13680, new_n13681, new_n13682, new_n13683, new_n13684,
    new_n13685, new_n13686, new_n13687, new_n13688, new_n13689, new_n13690,
    new_n13691, new_n13692, new_n13693, new_n13694, new_n13695, new_n13696,
    new_n13697, new_n13698, new_n13699, new_n13700, new_n13701, new_n13702,
    new_n13703, new_n13704, new_n13705, new_n13706, new_n13707, new_n13708,
    new_n13709, new_n13710, new_n13711, new_n13712, new_n13713, new_n13714,
    new_n13715, new_n13716, new_n13717, new_n13718, new_n13719, new_n13720,
    new_n13721, new_n13722, new_n13723, new_n13724, new_n13725, new_n13726,
    new_n13727, new_n13728, new_n13729, new_n13730, new_n13731, new_n13732,
    new_n13733, new_n13734, new_n13735, new_n13736, new_n13737, new_n13738,
    new_n13739, new_n13740, new_n13741, new_n13742, new_n13743, new_n13744,
    new_n13745, new_n13746, new_n13747, new_n13748, new_n13749, new_n13750,
    new_n13751, new_n13752, new_n13753, new_n13754, new_n13755, new_n13756,
    new_n13757, new_n13758, new_n13759, new_n13760, new_n13761, new_n13762,
    new_n13763, new_n13764, new_n13765, new_n13766, new_n13767, new_n13768,
    new_n13769, new_n13770, new_n13771, new_n13772, new_n13773, new_n13774,
    new_n13775, new_n13776, new_n13777, new_n13778, new_n13779, new_n13780,
    new_n13781, new_n13782, new_n13783, new_n13784, new_n13785, new_n13786,
    new_n13788, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806,
    new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812,
    new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818,
    new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824,
    new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830,
    new_n13831, new_n13832, new_n13833, new_n13834, new_n13835, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872,
    new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878,
    new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884,
    new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890,
    new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13911, new_n13912, new_n13913, new_n13914,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922, new_n13923, new_n13924, new_n13925, new_n13926,
    new_n13927, new_n13928, new_n13929, new_n13930, new_n13931, new_n13932,
    new_n13933, new_n13934, new_n13935, new_n13936, new_n13937, new_n13938,
    new_n13939, new_n13940, new_n13941, new_n13942, new_n13943, new_n13944,
    new_n13945, new_n13946, new_n13947, new_n13948, new_n13949, new_n13950,
    new_n13951, new_n13952, new_n13953, new_n13954, new_n13955, new_n13956,
    new_n13957, new_n13958, new_n13959, new_n13960, new_n13961, new_n13962,
    new_n13963, new_n13964, new_n13965, new_n13966, new_n13967, new_n13968,
    new_n13969, new_n13970, new_n13971, new_n13972, new_n13974, new_n13976,
    new_n13979, new_n13981, new_n13983, new_n13985, new_n13987, new_n13991,
    new_n13992, new_n13993, new_n13994, new_n13995, new_n13996, new_n13997,
    new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003,
    new_n14004, new_n14005, new_n14006, new_n14007, new_n14008, new_n14009,
    new_n14010, new_n14011, new_n14012, new_n14013, new_n14014, new_n14015,
    new_n14016, new_n14017, new_n14018, new_n14019, new_n14020, new_n14021,
    new_n14022, new_n14023, new_n14024, new_n14025, new_n14026, new_n14027,
    new_n14028, new_n14029, new_n14030, new_n14031, new_n14032, new_n14033,
    new_n14034, new_n14035, new_n14036, new_n14037, new_n14038, new_n14039,
    new_n14040, new_n14041, new_n14042, new_n14043, new_n14044, new_n14045,
    new_n14046, new_n14047, new_n14048, new_n14049, new_n14050, new_n14051,
    new_n14052, new_n14053, new_n14054, new_n14055, new_n14056, new_n14057,
    new_n14058, new_n14059, new_n14060, new_n14061, new_n14062, new_n14063,
    new_n14064, new_n14065, new_n14066, new_n14067, new_n14068, new_n14069,
    new_n14070, new_n14071, new_n14072, new_n14073, new_n14074, new_n14075,
    new_n14076, new_n14077, new_n14078, new_n14079, new_n14080, new_n14081,
    new_n14082, new_n14083, new_n14084, new_n14085, new_n14086, new_n14087,
    new_n14088, new_n14089, new_n14090, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095, new_n14096, new_n14097, new_n14098, new_n14099,
    new_n14100, new_n14101, new_n14102, new_n14103, new_n14104, new_n14105,
    new_n14106, new_n14107, new_n14108, new_n14109, new_n14110, new_n14111,
    new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117,
    new_n14118, new_n14119, new_n14120, new_n14121, new_n14122, new_n14123,
    new_n14124, new_n14125, new_n14126, new_n14127, new_n14128, new_n14129,
    new_n14130, new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136, new_n14137, new_n14138, new_n14139, new_n14140, new_n14141,
    new_n14142, new_n14143, new_n14144, new_n14145, new_n14146, new_n14147,
    new_n14148, new_n14149, new_n14150, new_n14151, new_n14152, new_n14153,
    new_n14154, new_n14155, new_n14156, new_n14157, new_n14158, new_n14159,
    new_n14160, new_n14161, new_n14162, new_n14163, new_n14164, new_n14165,
    new_n14166, new_n14167, new_n14168, new_n14169, new_n14170, new_n14171,
    new_n14172, new_n14173, new_n14174, new_n14175, new_n14176, new_n14177,
    new_n14178, new_n14179, new_n14180, new_n14181, new_n14182, new_n14183,
    new_n14184, new_n14185, new_n14186, new_n14187, new_n14188, new_n14189,
    new_n14190, new_n14191, new_n14192, new_n14193, new_n14194, new_n14195,
    new_n14196, new_n14198, new_n14200, new_n14202, new_n14206, new_n14207,
    new_n14210, new_n14213, new_n14216, new_n14217, new_n14218, new_n14219,
    new_n14220, new_n14221, new_n14222, new_n14223, new_n14224, new_n14225,
    new_n14226, new_n14227, new_n14228, new_n14229, new_n14230, new_n14231,
    new_n14232, new_n14233, new_n14234, new_n14235, new_n14236, new_n14237,
    new_n14238, new_n14239, new_n14240, new_n14241, new_n14242, new_n14243,
    new_n14244, new_n14245, new_n14246, new_n14247, new_n14248, new_n14249,
    new_n14250, new_n14251, new_n14252, new_n14253, new_n14254, new_n14255,
    new_n14256, new_n14257, new_n14258, new_n14259, new_n14260, new_n14261,
    new_n14262, new_n14263, new_n14264, new_n14265, new_n14266, new_n14267,
    new_n14268, new_n14269, new_n14270, new_n14271, new_n14272, new_n14273,
    new_n14274, new_n14275, new_n14276, new_n14277, new_n14278, new_n14279,
    new_n14280, new_n14281, new_n14282, new_n14283, new_n14284, new_n14285,
    new_n14286, new_n14287, new_n14288, new_n14289, new_n14290, new_n14291,
    new_n14292, new_n14293, new_n14294, new_n14295, new_n14296, new_n14297,
    new_n14298, new_n14299, new_n14300, new_n14301, new_n14302, new_n14303,
    new_n14304, new_n14305, new_n14306, new_n14307, new_n14308, new_n14309,
    new_n14310, new_n14311, new_n14312, new_n14313, new_n14314, new_n14315,
    new_n14316, new_n14317, new_n14318, new_n14319, new_n14320, new_n14321,
    new_n14322, new_n14323, new_n14324, new_n14325, new_n14326, new_n14327,
    new_n14328, new_n14329, new_n14330, new_n14331, new_n14332, new_n14333,
    new_n14334, new_n14335, new_n14336, new_n14337, new_n14338, new_n14339,
    new_n14340, new_n14341, new_n14342, new_n14343, new_n14344, new_n14345,
    new_n14346, new_n14347, new_n14348, new_n14349, new_n14350, new_n14351,
    new_n14352, new_n14353, new_n14354, new_n14355, new_n14356, new_n14357,
    new_n14358, new_n14359, new_n14360, new_n14361, new_n14362, new_n14363,
    new_n14364, new_n14365, new_n14366, new_n14367, new_n14368, new_n14369,
    new_n14370, new_n14371, new_n14372, new_n14373, new_n14374, new_n14375,
    new_n14376, new_n14377, new_n14378, new_n14379, new_n14380, new_n14381,
    new_n14382, new_n14383, new_n14384, new_n14385, new_n14386, new_n14387,
    new_n14388, new_n14389, new_n14390, new_n14391, new_n14392, new_n14393,
    new_n14394, new_n14395, new_n14396, new_n14397, new_n14398, new_n14399,
    new_n14400, new_n14401, new_n14402, new_n14403, new_n14404, new_n14405,
    new_n14406, new_n14407, new_n14409, new_n14411, new_n14419, new_n14421;
nand_1 g00000(n6687, n6038, new_n377);
nand_1 g00001(n8336, n7354, new_n378);
nand_1 g00002(n11222, n8028, new_n379);
not_4  g00003(new_n379, new_n380);
nand_1 g00004(n12069, n1564, new_n381_1);
not_4  g00005(new_n381_1, new_n382);
nand_1 g00006(new_n382, new_n380, new_n383);
nand_1 g00007(new_n381_1, new_n379, new_n384);
nand_1 g00008(new_n384, new_n383, new_n385);
not_4  g00009(new_n385, new_n386);
xnor_1 g00010(new_n386, new_n378, new_n387);
xnor_1 g00011(new_n387, new_n377, n112);
nand_1 g00012(n12720, n4312, new_n389);
nand_1 g00013(n12025, n6038, new_n390);
nand_1 g00014(n12705, n2509, new_n391);
not_4  g00015(new_n391, new_n392);
xnor_1 g00016(new_n392, new_n390, new_n393);
xnor_1 g00017(new_n393, new_n389, new_n394);
nand_1 g00018(n12705, n6038, new_n395);
nand_1 g00019(n12720, n1097, new_n396);
nand_1 g00020(new_n396, new_n395, new_n397_1);
nand_1 g00021(n4312, n2509, new_n398);
not_4  g00022(new_n396, new_n399);
xnor_1 g00023(new_n399, new_n395, new_n400);
nand_1 g00024(new_n400, new_n398, new_n401);
nand_1 g00025(new_n401, new_n397_1, new_n402);
xnor_1 g00026(new_n402, new_n394, new_n403);
not_4  g00027(new_n403, new_n404);
nand_1 g00028(n2508, n1097, new_n405_1);
nand_1 g00029(n5964, n2585, new_n406);
nand_1 g00030(new_n406, new_n405_1, new_n407);
not_4  g00031(new_n405_1, new_n408);
not_4  g00032(new_n406, new_n409);
nand_1 g00033(new_n409, new_n408, new_n410);
nand_1 g00034(new_n410, new_n407, new_n411);
not_4  g00035(new_n411, new_n412);
xnor_1 g00036(new_n412, new_n404, new_n413);
nand_1 g00037(n5964, n2508, new_n414);
not_4  g00038(new_n400, new_n415);
xnor_1 g00039(new_n415, new_n398, new_n416);
nand_1 g00040(new_n416, new_n414, new_n417);
not_4  g00041(new_n414, new_n418);
xnor_1 g00042(new_n416, new_n418, new_n419);
nand_1 g00043(n6038, n4312, new_n420);
nand_1 g00044(n12720, n5964, new_n421);
nand_1 g00045(new_n421, new_n420, new_n422);
not_4  g00046(new_n420, new_n423);
not_4  g00047(new_n421, new_n424);
nand_1 g00048(new_n424, new_n423, new_n425);
nand_1 g00049(n2509, n1097, new_n426);
nand_1 g00050(new_n426, new_n425, new_n427);
nand_1 g00051(new_n427, new_n422, new_n428);
nand_1 g00052(new_n428, new_n419, new_n429);
nand_1 g00053(new_n429, new_n417, new_n430);
xnor_1 g00054(new_n430, new_n413, new_n431);
nand_1 g00055(n5305, n2585, new_n432);
xnor_1 g00056(new_n428, new_n419, new_n433);
not_4  g00057(new_n433, new_n434);
nand_1 g00058(new_n434, new_n432, new_n435);
xnor_1 g00059(new_n433, new_n432, new_n436);
not_4  g00060(new_n436, new_n437);
nand_1 g00061(n5305, n2508, new_n438);
not_4  g00062(new_n438, new_n439);
nand_1 g00063(n6038, n1097, new_n440);
not_4  g00064(new_n440, new_n441);
nand_1 g00065(n12720, n5305, new_n442);
not_4  g00066(new_n442, new_n443);
nand_1 g00067(new_n443, new_n441, new_n444);
nand_1 g00068(new_n442, new_n440, new_n445);
nand_1 g00069(n5964, n2509, new_n446);
not_4  g00070(new_n446, new_n447_1);
nand_1 g00071(new_n447_1, new_n445, new_n448);
nand_1 g00072(new_n448, new_n444, new_n449);
nand_1 g00073(new_n449, new_n439, new_n450);
xnor_1 g00074(new_n449, new_n438, new_n451);
not_4  g00075(new_n451, new_n452);
nand_1 g00076(new_n425, new_n422, new_n453);
xnor_1 g00077(new_n453, new_n426, new_n454);
nor_1  g00078(new_n454, new_n452, new_n455);
not_4  g00079(new_n455, new_n456);
nand_1 g00080(new_n456, new_n450, new_n457);
nor_1  g00081(new_n457, new_n437, new_n458);
not_4  g00082(new_n458, new_n459);
nand_1 g00083(new_n459, new_n435, new_n460);
not_4  g00084(new_n460, new_n461);
nand_1 g00085(new_n461, new_n431, new_n462);
not_4  g00086(new_n389, new_n463);
nand_1 g00087(new_n393, new_n463, new_n464);
not_4  g00088(new_n394, new_n465);
nor_1  g00089(new_n402, new_n465, new_n466);
not_4  g00090(new_n466, new_n467);
nand_1 g00091(new_n467, new_n464, new_n468);
nand_1 g00092(n5964, n4005, new_n469);
nand_1 g00093(n2585, n1097, new_n470);
nand_1 g00094(n12706, n5305, new_n471);
nand_1 g00095(new_n471, new_n470, new_n472);
not_4  g00096(new_n470, new_n473);
not_4  g00097(new_n471, new_n474);
nand_1 g00098(new_n474, new_n473, new_n475);
nand_1 g00099(new_n475, new_n472, new_n476);
xnor_1 g00100(new_n476, new_n469, new_n477);
xnor_1 g00101(new_n477, new_n468, new_n478);
not_4  g00102(new_n390, new_n479);
nand_1 g00103(new_n392, new_n479, new_n480);
not_4  g00104(new_n480, new_n481);
nand_1 g00105(n4312, n2508, new_n482);
not_4  g00106(new_n482, new_n483);
nand_1 g00107(new_n483, new_n481, new_n484);
nand_1 g00108(new_n482, new_n480, new_n485);
nand_1 g00109(new_n485, new_n484, new_n486);
nand_1 g00110(n12025, n2509, new_n487);
nand_1 g00111(n12720, n12705, new_n488);
nand_1 g00112(n11257, n6038, new_n489);
not_4  g00113(new_n489, new_n490);
xnor_1 g00114(new_n490, new_n488, new_n491);
xnor_1 g00115(new_n491, new_n487, new_n492);
xnor_1 g00116(new_n492, new_n486, new_n493);
not_4  g00117(new_n493, new_n494);
xnor_1 g00118(new_n494, new_n478, new_n495);
nand_1 g00119(new_n412, new_n403, new_n496);
not_4  g00120(new_n410, new_n497);
not_4  g00121(new_n413, new_n498);
nor_1  g00122(new_n430, new_n498, new_n499);
xnor_1 g00123(new_n499, new_n497, new_n500);
nand_1 g00124(new_n500, new_n496, new_n501);
not_4  g00125(new_n501, new_n502);
xnor_1 g00126(new_n502, new_n495, new_n503_1);
xnor_1 g00127(new_n503_1, new_n462, new_n504);
nand_1 g00128(n5305, n4005, new_n505);
not_4  g00129(new_n505, new_n506);
xnor_1 g00130(new_n460, new_n431, new_n507);
nand_1 g00131(new_n507, new_n506, new_n508);
not_4  g00132(new_n507, new_n509);
nand_1 g00133(new_n509, new_n505, new_n510);
xnor_1 g00134(new_n454, new_n451, new_n511);
nand_1 g00135(new_n445, new_n444, new_n512);
not_4  g00136(new_n512, new_n513);
nand_1 g00137(n6038, n5964, new_n514);
not_4  g00138(new_n514, new_n515);
nand_1 g00139(n5305, n2509, new_n516);
not_4  g00140(new_n516, new_n517);
nand_1 g00141(new_n517, new_n515, new_n518);
nor_1  g00142(new_n518, new_n513, new_n519);
nand_1 g00143(new_n519, new_n511, new_n520);
xnor_1 g00144(new_n457, new_n436, new_n521_1);
nor_1  g00145(new_n521_1, new_n520, new_n522);
nand_1 g00146(new_n522, new_n510, new_n523);
nand_1 g00147(new_n523, new_n508, new_n524);
xnor_1 g00148(new_n524, new_n504, new_n525);
nand_1 g00149(n8759, n5105, new_n526);
nand_1 g00150(n12299, n7354, new_n527);
nand_1 g00151(n8759, n1209, new_n528);
nand_1 g00152(new_n528, new_n527, new_n529);
nor_1  g00153(new_n528, new_n527, new_n530);
not_4  g00154(new_n530, new_n531);
nand_1 g00155(n7500, n6776, new_n532);
nand_1 g00156(new_n532, new_n531, new_n533_1);
nand_1 g00157(new_n533_1, new_n529, new_n534);
nor_1  g00158(new_n534, new_n526, new_n535);
not_4  g00159(new_n535, new_n536);
nand_1 g00160(new_n534, new_n526, new_n537);
nand_1 g00161(new_n537, new_n536, new_n538);
nand_1 g00162(n12299, n7500, new_n539);
nand_1 g00163(n7436, n7354, new_n540);
nand_1 g00164(n6776, n1209, new_n541);
not_4  g00165(new_n541, new_n542);
xnor_1 g00166(new_n542, new_n540, new_n543);
xnor_1 g00167(new_n543, new_n539, new_n544);
not_4  g00168(new_n544, new_n545);
xnor_1 g00169(new_n545, new_n538, new_n546);
not_4  g00170(new_n532, new_n547);
not_4  g00171(new_n529, new_n548);
nand_1 g00172(n8759, n7354, new_n549);
nand_1 g00173(new_n549, new_n547, new_n550);
nand_1 g00174(new_n550, new_n548, new_n551);
nand_1 g00175(new_n551, new_n531, new_n552);
nand_1 g00176(new_n552, new_n547, new_n553);
nor_1  g00177(new_n553, new_n546, new_n554);
nand_1 g00178(n8759, n4141, new_n555);
nand_1 g00179(n6776, n5105, new_n556);
nand_1 g00180(new_n541, new_n540, new_n557);
nand_1 g00181(new_n543, new_n539, new_n558);
nand_1 g00182(new_n558, new_n557, new_n559);
not_4  g00183(new_n559, new_n560);
xnor_1 g00184(new_n560, new_n556, new_n561);
nand_1 g00185(n7500, n7436, new_n562);
nand_1 g00186(n12299, n1209, new_n563);
nand_1 g00187(n8276, n7354, new_n564);
not_4  g00188(new_n564, new_n565);
xnor_1 g00189(new_n565, new_n563, new_n566);
not_4  g00190(new_n566, new_n567);
xnor_1 g00191(new_n567, new_n562, new_n568);
xnor_1 g00192(new_n568, new_n561, new_n569);
xnor_1 g00193(new_n569, new_n555, new_n570);
not_4  g00194(new_n538, new_n571);
nand_1 g00195(new_n544, new_n571, new_n572);
nand_1 g00196(new_n572, new_n536, new_n573);
xnor_1 g00197(new_n573, new_n570, new_n574);
not_4  g00198(new_n574, new_n575);
nand_1 g00199(new_n575, new_n554, new_n576);
nand_1 g00200(n8759, n4928, new_n577);
nand_1 g00201(n7436, n1209, new_n578);
not_4  g00202(new_n578, new_n579);
nand_1 g00203(n8276, n7500, new_n580);
nand_1 g00204(n9241, n7354, new_n581);
not_4  g00205(new_n581, new_n582);
xnor_1 g00206(new_n582, new_n580, new_n583);
xnor_1 g00207(new_n583, new_n579, new_n584);
nand_1 g00208(new_n564, new_n563, new_n585);
nand_1 g00209(new_n566, new_n562, new_n586);
nand_1 g00210(new_n586, new_n585, new_n587);
nor_1  g00211(new_n587, new_n584, new_n588);
not_4  g00212(new_n588, new_n589);
nand_1 g00213(new_n587, new_n584, new_n590);
nand_1 g00214(new_n590, new_n589, new_n591);
nand_1 g00215(n6776, n4141, new_n592);
nand_1 g00216(n12299, n5105, new_n593);
not_4  g00217(new_n593, new_n594);
xnor_1 g00218(new_n594, new_n592, new_n595);
xnor_1 g00219(new_n595, new_n591, new_n596);
nor_1  g00220(new_n559, new_n556, new_n597);
not_4  g00221(new_n561, new_n598);
nor_1  g00222(new_n568, new_n598, new_n599);
nor_1  g00223(new_n599, new_n597, new_n600);
xnor_1 g00224(new_n600, new_n596, new_n601);
not_4  g00225(new_n555, new_n602);
nand_1 g00226(new_n569, new_n602, new_n603);
nand_1 g00227(new_n573, new_n570, new_n604);
nand_1 g00228(new_n604, new_n603, new_n605);
nand_1 g00229(new_n605, new_n601, new_n606);
not_4  g00230(new_n606, new_n607);
nor_1  g00231(new_n605, new_n601, new_n608);
nor_1  g00232(new_n608, new_n607, new_n609);
xnor_1 g00233(new_n609, new_n577, new_n610);
xnor_1 g00234(new_n610, new_n576, new_n611);
not_4  g00235(new_n611, new_n612);
xnor_1 g00236(new_n574, new_n554, new_n613);
not_4  g00237(new_n613, new_n614);
xnor_1 g00238(new_n553, new_n546, new_n615_1);
not_4  g00239(new_n549, new_n616);
nand_1 g00240(n5331, n1564, new_n617);
nand_1 g00241(n8028, n7965, new_n618);
not_4  g00242(new_n618, new_n619);
xnor_1 g00243(new_n619, new_n617, new_n620);
nand_1 g00244(new_n620, new_n616, new_n621);
not_4  g00245(new_n621, new_n622);
nand_1 g00246(n7354, n6776, new_n623);
nand_1 g00247(n8759, n7500, new_n624);
not_4  g00248(new_n624, new_n625);
xnor_1 g00249(new_n625, new_n623, new_n626);
nor_1  g00250(new_n626, new_n622, new_n627);
not_4  g00251(new_n627, new_n628);
not_4  g00252(new_n617, new_n629);
nand_1 g00253(new_n619, new_n629, new_n630);
nand_1 g00254(n5331, n1512, new_n631);
nand_1 g00255(n8476, n1564, new_n632);
not_4  g00256(new_n632, new_n633);
xnor_1 g00257(new_n633, new_n631, new_n634);
xnor_1 g00258(new_n634, new_n630, new_n635);
nand_1 g00259(n8028, n7388, new_n636);
nand_1 g00260(n10848, n7965, new_n637);
not_4  g00261(new_n637, new_n638);
xnor_1 g00262(new_n638, new_n636, new_n639);
xnor_1 g00263(new_n639, new_n635, new_n640);
xnor_1 g00264(new_n626, new_n621, new_n641);
nand_1 g00265(new_n641, new_n640, new_n642);
nand_1 g00266(new_n642, new_n628, new_n643);
nor_1  g00267(new_n550, new_n548, new_n644);
nor_1  g00268(new_n644, new_n552, new_n645);
not_4  g00269(new_n645, new_n646);
nand_1 g00270(new_n646, new_n643, new_n647);
nand_1 g00271(n10848, n7388, new_n648);
not_4  g00272(new_n648, new_n649);
nand_1 g00273(new_n649, new_n618, new_n650);
nand_1 g00274(n11892, n8028, new_n651);
nand_1 g00275(n7965, n1980, new_n652);
nand_1 g00276(new_n652, new_n651, new_n653);
nand_1 g00277(n11892, n1980, new_n654);
not_4  g00278(new_n654, new_n655);
nand_1 g00279(new_n655, new_n619, new_n656);
nand_1 g00280(new_n656, new_n653, new_n657);
nand_1 g00281(new_n657, new_n650, new_n658_1);
not_4  g00282(new_n653, new_n659);
nor_1  g00283(new_n659, new_n650, new_n660);
not_4  g00284(new_n660, new_n661);
nand_1 g00285(new_n661, new_n658_1, new_n662);
nand_1 g00286(n8476, n1512, new_n663);
not_4  g00287(new_n663, new_n664);
nand_1 g00288(new_n664, new_n617, new_n665);
nand_1 g00289(n2530, n1564, new_n666);
nand_1 g00290(n5331, n533, new_n667);
nand_1 g00291(new_n667, new_n666, new_n668);
not_4  g00292(new_n668, new_n669);
nand_1 g00293(new_n669, new_n665, new_n670);
not_4  g00294(new_n666, new_n671_1);
not_4  g00295(new_n667, new_n672);
nand_1 g00296(new_n672, new_n671_1, new_n673);
nand_1 g00297(new_n673, new_n670, new_n674);
nor_1  g00298(new_n669, new_n665, new_n675);
nor_1  g00299(new_n675, new_n674, new_n676);
xnor_1 g00300(new_n676, new_n662, new_n677);
not_4  g00301(new_n630, new_n678);
nand_1 g00302(new_n634, new_n678, new_n679);
nand_1 g00303(new_n639, new_n635, new_n680);
nand_1 g00304(new_n680, new_n679, new_n681);
xnor_1 g00305(new_n681, new_n677, new_n682);
xnor_1 g00306(new_n645, new_n643, new_n683);
nand_1 g00307(new_n683, new_n682, new_n684);
nand_1 g00308(new_n684, new_n647, new_n685);
nand_1 g00309(new_n685, new_n615_1, new_n686);
nand_1 g00310(n5331, n2802, new_n687);
nand_1 g00311(new_n673, new_n663, new_n688);
nand_1 g00312(new_n688, new_n668, new_n689);
nor_1  g00313(new_n689, new_n687, new_n690);
not_4  g00314(new_n690, new_n691);
nand_1 g00315(new_n689, new_n687, new_n692);
nand_1 g00316(new_n692, new_n691, new_n693);
nand_1 g00317(n2530, n1512, new_n694);
nand_1 g00318(n12648, n1564, new_n695);
nand_1 g00319(n8476, n533, new_n696);
not_4  g00320(new_n696, new_n697);
xnor_1 g00321(new_n697, new_n695, new_n698);
not_4  g00322(new_n698, new_n699);
xnor_1 g00323(new_n699, new_n694, new_n700);
nor_1  g00324(new_n700, new_n693, new_n701);
not_4  g00325(new_n701, new_n702);
nand_1 g00326(new_n700, new_n693, new_n703);
nand_1 g00327(new_n703, new_n702, new_n704);
nand_1 g00328(new_n674, new_n664, new_n705);
not_4  g00329(new_n705, new_n706);
xnor_1 g00330(new_n706, new_n704, new_n707);
nand_1 g00331(n7965, n7294, new_n708);
nand_1 g00332(new_n656, new_n648, new_n709);
nand_1 g00333(new_n709, new_n653, new_n710);
not_4  g00334(new_n710, new_n711);
xnor_1 g00335(new_n711, new_n708, new_n712);
nand_1 g00336(n11892, n10848, new_n713);
not_4  g00337(new_n713, new_n714);
nand_1 g00338(n7388, n1980, new_n715);
nand_1 g00339(n8028, n2393, new_n716);
nand_1 g00340(new_n716, new_n715, new_n717);
not_4  g00341(new_n715, new_n718);
not_4  g00342(new_n716, new_n719);
nand_1 g00343(new_n719, new_n718, new_n720);
nand_1 g00344(new_n720, new_n717, new_n721);
xnor_1 g00345(new_n721, new_n714, new_n722);
xnor_1 g00346(new_n722, new_n712, new_n723);
nor_1  g00347(new_n658_1, new_n648, new_n724);
xnor_1 g00348(new_n724, new_n723, new_n725);
nand_1 g00349(new_n725, new_n707, new_n726);
nor_1  g00350(new_n725, new_n707, new_n727);
not_4  g00351(new_n727, new_n728);
nand_1 g00352(new_n728, new_n726, new_n729);
not_4  g00353(new_n676, new_n730);
nor_1  g00354(new_n730, new_n662, new_n731);
not_4  g00355(new_n731, new_n732);
nand_1 g00356(new_n681, new_n677, new_n733);
nand_1 g00357(new_n733, new_n732, new_n734);
not_4  g00358(new_n734, new_n735);
xnor_1 g00359(new_n735, new_n729, new_n736);
not_4  g00360(new_n686, new_n737);
nor_1  g00361(new_n685, new_n615_1, new_n738);
nor_1  g00362(new_n738, new_n737, new_n739);
nand_1 g00363(new_n739, new_n736, new_n740);
nand_1 g00364(new_n740, new_n686, new_n741);
nand_1 g00365(new_n741, new_n614, new_n742);
not_4  g00366(new_n723, new_n743);
nand_1 g00367(new_n724, new_n743, new_n744);
nor_1  g00368(new_n710, new_n708, new_n745);
not_4  g00369(new_n745, new_n746);
nand_1 g00370(new_n722, new_n712, new_n747);
nand_1 g00371(new_n747, new_n746, new_n748);
nand_1 g00372(n12704, n7965, new_n749);
nand_1 g00373(n7388, n7294, new_n750);
nand_1 g00374(new_n720, new_n713, new_n751);
nand_1 g00375(new_n751, new_n717, new_n752);
nor_1  g00376(new_n752, new_n750, new_n753_1);
not_4  g00377(new_n753_1, new_n754);
nand_1 g00378(new_n752, new_n750, new_n755);
nand_1 g00379(new_n755, new_n754, new_n756);
nand_1 g00380(n10848, n2393, new_n757);
not_4  g00381(new_n757, new_n758);
nand_1 g00382(n8028, n5860, new_n759);
nand_1 g00383(new_n759, new_n654, new_n760);
nor_1  g00384(new_n759, new_n654, new_n761);
not_4  g00385(new_n761, new_n762);
nand_1 g00386(new_n762, new_n760, new_n763);
xnor_1 g00387(new_n763, new_n758, new_n764);
xnor_1 g00388(new_n764, new_n756, new_n765);
not_4  g00389(new_n765, new_n766);
nand_1 g00390(new_n766, new_n749, new_n767);
nor_1  g00391(new_n766, new_n749, new_n768);
not_4  g00392(new_n768, new_n769);
nand_1 g00393(new_n769, new_n767, new_n770);
xnor_1 g00394(new_n770, new_n748, new_n771);
xnor_1 g00395(new_n771, new_n744, new_n772);
nor_1  g00396(new_n705, new_n704, new_n773);
nand_1 g00397(n6806, n5331, new_n774);
nand_1 g00398(n8476, n2802, new_n775);
nand_1 g00399(new_n696, new_n695, new_n776);
nand_1 g00400(new_n698, new_n694, new_n777);
nand_1 g00401(new_n777, new_n776, new_n778);
not_4  g00402(new_n778, new_n779);
xnor_1 g00403(new_n779, new_n775, new_n780);
nand_1 g00404(n12648, n1512, new_n781);
nand_1 g00405(n2530, n533, new_n782);
nand_1 g00406(n10545, n1564, new_n783_1);
xnor_1 g00407(new_n783_1, new_n782, new_n784);
xnor_1 g00408(new_n784, new_n781, new_n785);
xnor_1 g00409(new_n785, new_n780, new_n786);
xnor_1 g00410(new_n786, new_n774, new_n787);
not_4  g00411(new_n787, new_n788);
nand_1 g00412(new_n702, new_n691, new_n789);
xnor_1 g00413(new_n789, new_n788, new_n790);
xnor_1 g00414(new_n790, new_n773, new_n791);
not_4  g00415(new_n791, new_n792);
nor_1  g00416(new_n734, new_n729, new_n793);
nor_1  g00417(new_n793, new_n727, new_n794);
nand_1 g00418(new_n794, new_n792, new_n795);
nor_1  g00419(new_n794, new_n792, new_n796);
not_4  g00420(new_n796, new_n797);
nand_1 g00421(new_n797, new_n795, new_n798);
nand_1 g00422(new_n798, new_n772, new_n799);
nor_1  g00423(new_n798, new_n772, new_n800);
not_4  g00424(new_n800, new_n801);
nand_1 g00425(new_n801, new_n799, new_n802);
not_4  g00426(new_n802, new_n803);
xnor_1 g00427(new_n741, new_n613, new_n804);
nand_1 g00428(new_n804, new_n803, new_n805);
nand_1 g00429(new_n805, new_n742, new_n806_1);
nand_1 g00430(new_n806_1, new_n612, new_n807);
not_4  g00431(new_n742, new_n808);
xnor_1 g00432(new_n741, new_n614, new_n809);
nor_1  g00433(new_n809, new_n802, new_n810);
nor_1  g00434(new_n810, new_n808, new_n811);
nand_1 g00435(new_n811, new_n611, new_n812);
nand_1 g00436(new_n812, new_n807, new_n813);
not_4  g00437(new_n813, new_n814);
nand_1 g00438(new_n801, new_n797, new_n815);
nand_1 g00439(new_n790, new_n773, new_n816);
nand_1 g00440(n5331, n5069, new_n817);
not_4  g00441(new_n817, new_n818);
nand_1 g00442(n12648, n533, new_n819);
nand_1 g00443(n10545, n1512, new_n820);
nand_1 g00444(n7690, n1564, new_n821);
not_4  g00445(new_n821, new_n822);
xnor_1 g00446(new_n822, new_n820, new_n823);
xnor_1 g00447(new_n823, new_n819, new_n824);
nand_1 g00448(new_n783_1, new_n782, new_n825);
not_4  g00449(new_n825, new_n826);
not_4  g00450(new_n781, new_n827);
nor_1  g00451(new_n784, new_n827, new_n828);
nor_1  g00452(new_n828, new_n826, new_n829);
nand_1 g00453(new_n829, new_n824, new_n830);
not_4  g00454(new_n830, new_n831);
nor_1  g00455(new_n829, new_n824, new_n832);
nor_1  g00456(new_n832, new_n831, new_n833);
nand_1 g00457(n8476, n6806, new_n834);
nand_1 g00458(n2802, n2530, new_n835);
nand_1 g00459(new_n835, new_n834, new_n836);
not_4  g00460(new_n834, new_n837_1);
not_4  g00461(new_n835, new_n838);
nand_1 g00462(new_n838, new_n837_1, new_n839);
nand_1 g00463(new_n839, new_n836, new_n840);
xnor_1 g00464(new_n840, new_n833, new_n841);
nor_1  g00465(new_n778, new_n775, new_n842);
not_4  g00466(new_n780, new_n843);
nor_1  g00467(new_n785, new_n843, new_n844_1);
nor_1  g00468(new_n844_1, new_n842, new_n845);
xnor_1 g00469(new_n845, new_n841, new_n846);
not_4  g00470(new_n774, new_n847);
nand_1 g00471(new_n786, new_n847, new_n848);
nand_1 g00472(new_n789, new_n787, new_n849);
nand_1 g00473(new_n849, new_n848, new_n850);
xnor_1 g00474(new_n850, new_n846, new_n851);
not_4  g00475(new_n851, new_n852);
nand_1 g00476(new_n852, new_n818, new_n853);
nand_1 g00477(new_n851, new_n817, new_n854);
nand_1 g00478(new_n854, new_n853, new_n855);
xnor_1 g00479(new_n855, new_n816, new_n856);
nor_1  g00480(new_n856, new_n815, new_n857);
not_4  g00481(new_n815, new_n858);
not_4  g00482(new_n856, new_n859);
nor_1  g00483(new_n859, new_n858, new_n860);
nor_1  g00484(new_n860, new_n857, new_n861);
not_4  g00485(new_n744, new_n862);
nand_1 g00486(new_n771, new_n862, new_n863);
nand_1 g00487(n7965, n5814, new_n864);
not_4  g00488(new_n864, new_n865);
nand_1 g00489(n2393, n1980, new_n866);
not_4  g00490(new_n866, new_n867);
nand_1 g00491(n8028, n3986, new_n868);
nand_1 g00492(n10848, n5860, new_n869);
not_4  g00493(new_n869, new_n870);
xnor_1 g00494(new_n870, new_n868, new_n871);
xnor_1 g00495(new_n871, new_n867, new_n872);
nand_1 g00496(new_n762, new_n757, new_n873);
nand_1 g00497(new_n873, new_n760, new_n874);
nor_1  g00498(new_n874, new_n872, new_n875);
not_4  g00499(new_n875, new_n876);
nand_1 g00500(new_n874, new_n872, new_n877);
nand_1 g00501(new_n877, new_n876, new_n878);
nand_1 g00502(n12704, n7388, new_n879);
nand_1 g00503(n11892, n7294, new_n880);
not_4  g00504(new_n880, new_n881);
xnor_1 g00505(new_n881, new_n879, new_n882);
xnor_1 g00506(new_n882, new_n878, new_n883);
not_4  g00507(new_n756, new_n884);
nand_1 g00508(new_n764, new_n884, new_n885);
nand_1 g00509(new_n885, new_n754, new_n886);
xnor_1 g00510(new_n886, new_n883, new_n887);
nor_1  g00511(new_n768, new_n748, new_n888);
not_4  g00512(new_n888, new_n889);
nand_1 g00513(new_n889, new_n767, new_n890);
nor_1  g00514(new_n890, new_n887, new_n891);
not_4  g00515(new_n891, new_n892);
nand_1 g00516(new_n890, new_n887, new_n893);
nand_1 g00517(new_n893, new_n892, new_n894);
not_4  g00518(new_n894, new_n895);
nand_1 g00519(new_n895, new_n865, new_n896);
nand_1 g00520(new_n894, new_n864, new_n897);
nand_1 g00521(new_n897, new_n896, new_n898);
xnor_1 g00522(new_n898, new_n863, new_n899);
xnor_1 g00523(new_n899, new_n861, new_n900);
xnor_1 g00524(new_n900, new_n814, new_n901);
not_4  g00525(new_n901, new_n902);
nand_1 g00526(new_n510, new_n508, new_n903);
xnor_1 g00527(new_n903, new_n522, new_n904);
nand_1 g00528(new_n904, new_n902, new_n905);
xnor_1 g00529(new_n521_1, new_n520, new_n906);
xnor_1 g00530(new_n804, new_n802, new_n907);
nor_1  g00531(new_n907, new_n906, new_n908);
not_4  g00532(new_n908, new_n909);
not_4  g00533(new_n907, new_n910);
xnor_1 g00534(new_n910, new_n906, new_n911_1);
xnor_1 g00535(new_n519, new_n511, new_n912);
not_4  g00536(new_n736, new_n913);
xnor_1 g00537(new_n739, new_n913, new_n914);
nor_1  g00538(new_n914, new_n912, new_n915);
xnor_1 g00539(new_n683, new_n682, new_n916);
not_4  g00540(new_n916, new_n917);
nand_1 g00541(n6038, n5305, new_n918);
nand_1 g00542(new_n918, new_n447_1, new_n919);
nand_1 g00543(new_n919, new_n512, new_n920);
not_4  g00544(new_n918, new_n921);
nor_1  g00545(new_n921, new_n448, new_n922);
not_4  g00546(new_n922, new_n923);
nand_1 g00547(new_n923, new_n920, new_n924);
nand_1 g00548(new_n924, new_n917, new_n925);
xnor_1 g00549(new_n924, new_n916, new_n926);
xnor_1 g00550(new_n620, new_n549, new_n927);
nand_1 g00551(new_n927, new_n921, new_n928);
nand_1 g00552(new_n516, new_n514, new_n929);
nand_1 g00553(new_n929, new_n518, new_n930);
nand_1 g00554(new_n930, new_n928, new_n931);
xnor_1 g00555(new_n641, new_n640, new_n932);
xnor_1 g00556(new_n930, new_n928, new_n933);
nor_1  g00557(new_n933, new_n932, new_n934);
not_4  g00558(new_n934, new_n935);
nand_1 g00559(new_n935, new_n931, new_n936);
nand_1 g00560(new_n936, new_n926, new_n937);
nand_1 g00561(new_n937, new_n925, new_n938);
xnor_1 g00562(new_n914, new_n912, new_n939);
nor_1  g00563(new_n939, new_n938, new_n940);
nor_1  g00564(new_n940, new_n915, new_n941);
not_4  g00565(new_n941, new_n942);
nand_1 g00566(new_n942, new_n911_1, new_n943);
nand_1 g00567(new_n943, new_n909, new_n944);
not_4  g00568(new_n905, new_n945);
nor_1  g00569(new_n904, new_n902, new_n946);
nor_1  g00570(new_n946, new_n945, new_n947);
nand_1 g00571(new_n947, new_n944, new_n948);
nand_1 g00572(new_n948, new_n905, new_n949);
not_4  g00573(new_n949, new_n950);
nand_1 g00574(new_n950, new_n525, new_n951);
nor_1  g00575(new_n950, new_n525, new_n952);
not_4  g00576(new_n952, new_n953);
nand_1 g00577(new_n953, new_n951, new_n954);
nand_1 g00578(new_n583, new_n579, new_n955);
nand_1 g00579(new_n589, new_n955, new_n956);
nand_1 g00580(n6776, n4928, new_n957);
nand_1 g00581(n12299, n4141, new_n958);
nand_1 g00582(n8759, n8236, new_n959);
not_4  g00583(new_n959, new_n960);
xnor_1 g00584(new_n960, new_n958, new_n961);
xnor_1 g00585(new_n961, new_n957, new_n962);
not_4  g00586(new_n962, new_n963);
xnor_1 g00587(new_n963, new_n956, new_n964);
not_4  g00588(new_n580, new_n965);
nand_1 g00589(new_n582, new_n965, new_n966);
not_4  g00590(new_n966, new_n967);
nand_1 g00591(n7436, n5105, new_n968);
not_4  g00592(new_n968, new_n969);
nand_1 g00593(new_n969, new_n967, new_n970);
nand_1 g00594(new_n968, new_n966, new_n971);
nand_1 g00595(new_n971, new_n970, new_n972);
nand_1 g00596(n9241, n7500, new_n973);
nand_1 g00597(n8276, n1209, new_n974);
nand_1 g00598(n10510, n7354, new_n975);
nand_1 g00599(new_n975, new_n974, new_n976);
not_4  g00600(new_n974, new_n977);
not_4  g00601(new_n975, new_n978);
nand_1 g00602(new_n978, new_n977, new_n979);
nand_1 g00603(new_n979, new_n976, new_n980);
xnor_1 g00604(new_n980, new_n973, new_n981);
not_4  g00605(new_n981, new_n982);
xnor_1 g00606(new_n982, new_n972, new_n983);
xnor_1 g00607(new_n983, new_n964, new_n984);
not_4  g00608(new_n591, new_n985);
nand_1 g00609(new_n595, new_n985, new_n986);
nor_1  g00610(new_n593, new_n592, new_n987);
not_4  g00611(new_n600, new_n988);
nand_1 g00612(new_n988, new_n596, new_n989);
not_4  g00613(new_n989, new_n990);
xnor_1 g00614(new_n990, new_n987, new_n991);
nand_1 g00615(new_n991, new_n986, new_n992_1);
xnor_1 g00616(new_n992_1, new_n984, new_n993);
xnor_1 g00617(new_n993, new_n606, new_n994);
not_4  g00618(new_n577, new_n995);
nand_1 g00619(new_n609, new_n995, new_n996_1);
not_4  g00620(new_n576, new_n997);
nand_1 g00621(new_n610, new_n997, new_n998);
nand_1 g00622(new_n998, new_n996_1, new_n999);
xnor_1 g00623(new_n999, new_n994, new_n1000);
nand_1 g00624(new_n850, new_n846, new_n1001);
not_4  g00625(new_n819, new_n1002);
nand_1 g00626(new_n823, new_n1002, new_n1003);
nand_1 g00627(new_n830, new_n1003, new_n1004);
nand_1 g00628(n8476, n5069, new_n1005);
not_4  g00629(new_n1005, new_n1006);
nand_1 g00630(n6806, n2530, new_n1007);
nand_1 g00631(n12044, n5331, new_n1008);
not_4  g00632(new_n1008, new_n1009);
xnor_1 g00633(new_n1009, new_n1007, new_n1010);
xnor_1 g00634(new_n1010, new_n1006, new_n1011);
xnor_1 g00635(new_n1011, new_n1004, new_n1012);
not_4  g00636(new_n820, new_n1013);
nand_1 g00637(new_n822, new_n1013, new_n1014);
nand_1 g00638(n12648, n2802, new_n1015);
nand_1 g00639(new_n1015, new_n1014, new_n1016);
not_4  g00640(new_n1014, new_n1017);
not_4  g00641(new_n1015, new_n1018);
nand_1 g00642(new_n1018, new_n1017, new_n1019);
nand_1 g00643(new_n1019, new_n1016, new_n1020_1);
not_4  g00644(new_n1020_1, new_n1021);
nand_1 g00645(n7690, n1512, new_n1022);
nand_1 g00646(n10545, n533, new_n1023);
nand_1 g00647(n3616, n1564, new_n1024);
not_4  g00648(new_n1024, new_n1025);
xnor_1 g00649(new_n1025, new_n1023, new_n1026);
xnor_1 g00650(new_n1026, new_n1022, new_n1027);
not_4  g00651(new_n1027, new_n1028);
xnor_1 g00652(new_n1028, new_n1021, new_n1029);
xnor_1 g00653(new_n1029, new_n1012, new_n1030);
not_4  g00654(new_n1030, new_n1031);
not_4  g00655(new_n840, new_n1032);
nand_1 g00656(new_n1032, new_n833, new_n1033);
not_4  g00657(new_n1033, new_n1034);
not_4  g00658(new_n845, new_n1035);
nand_1 g00659(new_n1035, new_n841, new_n1036);
not_4  g00660(new_n1036, new_n1037);
xnor_1 g00661(new_n1037, new_n839, new_n1038);
nor_1  g00662(new_n1038, new_n1034, new_n1039);
xnor_1 g00663(new_n1039, new_n1031, new_n1040);
xnor_1 g00664(new_n1040, new_n1001, new_n1041);
not_4  g00665(new_n1041, new_n1042);
not_4  g00666(new_n816, new_n1043);
nand_1 g00667(new_n854, new_n1043, new_n1044);
nand_1 g00668(new_n1044, new_n853, new_n1045);
xnor_1 g00669(new_n1045, new_n1042, new_n1046);
nand_1 g00670(new_n871, new_n867, new_n1047);
nand_1 g00671(new_n876, new_n1047, new_n1048);
nand_1 g00672(n7388, n5814, new_n1049);
nand_1 g00673(n12704, n11892, new_n1050);
nand_1 g00674(n7965, n4903, new_n1051);
not_4  g00675(new_n1051, new_n1052);
xnor_1 g00676(new_n1052, new_n1050, new_n1053);
xnor_1 g00677(new_n1053, new_n1049, new_n1054);
xnor_1 g00678(new_n1054, new_n1048, new_n1055);
not_4  g00679(new_n868, new_n1056);
nand_1 g00680(new_n870, new_n1056, new_n1057);
nand_1 g00681(n7294, n2393, new_n1058);
not_4  g00682(new_n1058, new_n1059);
xnor_1 g00683(new_n1059, new_n1057, new_n1060);
nand_1 g00684(n10848, n3986, new_n1061);
nand_1 g00685(n5860, n1980, new_n1062);
nand_1 g00686(n8028, n5857, new_n1063);
not_4  g00687(new_n1063, new_n1064);
xnor_1 g00688(new_n1064, new_n1062, new_n1065);
xnor_1 g00689(new_n1065, new_n1061, new_n1066);
not_4  g00690(new_n1066, new_n1067_1);
xnor_1 g00691(new_n1067_1, new_n1060, new_n1068);
xnor_1 g00692(new_n1068, new_n1055, new_n1069);
not_4  g00693(new_n1069, new_n1070);
not_4  g00694(new_n878, new_n1071);
nand_1 g00695(new_n882, new_n1071, new_n1072);
nor_1  g00696(new_n880, new_n879, new_n1073);
nand_1 g00697(new_n886, new_n883, new_n1074);
not_4  g00698(new_n1074, new_n1075);
xnor_1 g00699(new_n1075, new_n1073, new_n1076);
nand_1 g00700(new_n1076, new_n1072, new_n1077);
xnor_1 g00701(new_n1077, new_n1070, new_n1078);
xnor_1 g00702(new_n1078, new_n892, new_n1079);
nand_1 g00703(new_n896, new_n863, new_n1080);
nand_1 g00704(new_n1080, new_n897, new_n1081);
xnor_1 g00705(new_n1081, new_n1079, new_n1082);
nand_1 g00706(new_n1082, new_n1046, new_n1083);
nor_1  g00707(new_n1082, new_n1046, new_n1084);
not_4  g00708(new_n1084, new_n1085);
nand_1 g00709(new_n1085, new_n1083, new_n1086);
nor_1  g00710(new_n899, new_n860, new_n1087);
nor_1  g00711(new_n1087, new_n857, new_n1088);
xnor_1 g00712(new_n1088, new_n1086, new_n1089);
not_4  g00713(new_n1089, new_n1090);
xnor_1 g00714(new_n1090, new_n1000, new_n1091);
not_4  g00715(new_n900, new_n1092);
nand_1 g00716(new_n1092, new_n814, new_n1093);
nand_1 g00717(new_n1093, new_n807, new_n1094_1);
xnor_1 g00718(new_n1094_1, new_n1091, new_n1095);
xnor_1 g00719(new_n1095, new_n954, n226);
nand_1 g00720(n5305, n4634, new_n1097_1);
nand_1 g00721(n10223, n5305, new_n1098);
nand_1 g00722(n7265, n1097, new_n1099);
nand_1 g00723(new_n1099, new_n1098, new_n1100);
nand_1 g00724(n7265, n5305, new_n1101);
not_4  g00725(new_n1101, new_n1102);
nand_1 g00726(n10223, n1097, new_n1103);
not_4  g00727(new_n1103, new_n1104);
nand_1 g00728(new_n1104, new_n1102, new_n1105);
nand_1 g00729(n5964, n2879, new_n1106);
nand_1 g00730(new_n1106, new_n1105, new_n1107);
nand_1 g00731(new_n1107, new_n1100, new_n1108);
nor_1  g00732(new_n1108, new_n1097_1, new_n1109);
not_4  g00733(new_n1109, new_n1110);
nand_1 g00734(new_n1108, new_n1097_1, new_n1111);
nand_1 g00735(new_n1111, new_n1110, new_n1112);
nand_1 g00736(n2879, n1097, new_n1113);
not_4  g00737(new_n1113, new_n1114);
nand_1 g00738(n10223, n5964, new_n1115);
nand_1 g00739(n7265, n4312, new_n1116);
nand_1 g00740(new_n1116, new_n1115, new_n1117);
nor_1  g00741(new_n1116, new_n1115, new_n1118);
not_4  g00742(new_n1118, new_n1119);
nand_1 g00743(new_n1119, new_n1117, new_n1120);
xnor_1 g00744(new_n1120, new_n1114, new_n1121);
xnor_1 g00745(new_n1121, new_n1112, new_n1122);
not_4  g00746(new_n1106, new_n1123);
nand_1 g00747(new_n1123, new_n1101, new_n1124);
nand_1 g00748(new_n1105, new_n1100, new_n1125);
nand_1 g00749(new_n1125, new_n1124, new_n1126);
not_4  g00750(new_n1126, new_n1127);
nand_1 g00751(new_n1127, new_n1123, new_n1128);
xnor_1 g00752(new_n1128, new_n1122, new_n1129);
not_4  g00753(new_n1124, new_n1130);
nand_1 g00754(new_n1130, new_n1100, new_n1131);
nand_1 g00755(new_n1131, new_n1126, new_n1132);
nand_1 g00756(n8759, n7946, new_n1133);
not_4  g00757(new_n1133, new_n1134);
nand_1 g00758(n5331, n2558, new_n1135);
not_4  g00759(new_n1135, new_n1136_1);
nand_1 g00760(n9763, n7965, new_n1137);
not_4  g00761(new_n1137, new_n1138_1);
nand_1 g00762(new_n1138_1, new_n1136_1, new_n1139);
nand_1 g00763(new_n1137, new_n1135, new_n1140);
nand_1 g00764(new_n1140, new_n1139, new_n1141);
not_4  g00765(new_n1141, new_n1142);
nand_1 g00766(new_n1142, new_n1134, new_n1143);
not_4  g00767(new_n1143, new_n1144);
nand_1 g00768(n7946, n6776, new_n1145);
nand_1 g00769(n8759, n2024, new_n1146);
xnor_1 g00770(new_n1146, new_n1145, new_n1147);
not_4  g00771(new_n1147, new_n1148);
nand_1 g00772(new_n1148, new_n1144, new_n1149);
nand_1 g00773(n9111, n7965, new_n1150);
nand_1 g00774(n9763, n7388, new_n1151);
not_4  g00775(new_n1151, new_n1152);
xnor_1 g00776(new_n1152, new_n1150, new_n1153);
xnor_1 g00777(new_n1153, new_n1139, new_n1154);
nand_1 g00778(n5331, n2498, new_n1155);
nand_1 g00779(n8476, n2558, new_n1156);
nand_1 g00780(new_n1156, new_n1155, new_n1157);
not_4  g00781(new_n1155, new_n1158);
not_4  g00782(new_n1156, new_n1159);
nand_1 g00783(new_n1159, new_n1158, new_n1160);
nand_1 g00784(new_n1160, new_n1157, new_n1161);
xnor_1 g00785(new_n1161, new_n1154, new_n1162);
xnor_1 g00786(new_n1148, new_n1143, new_n1163);
nand_1 g00787(new_n1163, new_n1162, new_n1164);
nand_1 g00788(new_n1164, new_n1149, new_n1165);
not_4  g00789(new_n1165, new_n1166);
nand_1 g00790(n6776, n2024, new_n1167);
not_4  g00791(new_n1167, new_n1168);
nand_1 g00792(new_n1168, new_n1133, new_n1169);
nand_1 g00793(n12299, n7946, new_n1170);
nand_1 g00794(n9189, n8759, new_n1171);
nand_1 g00795(new_n1171, new_n1170, new_n1172);
not_4  g00796(new_n1170, new_n1173);
not_4  g00797(new_n1171, new_n1174);
nand_1 g00798(new_n1174, new_n1173, new_n1175);
nand_1 g00799(new_n1175, new_n1172, new_n1176);
nand_1 g00800(new_n1176, new_n1169, new_n1177);
not_4  g00801(new_n1177, new_n1178);
not_4  g00802(new_n1172, new_n1179);
nor_1  g00803(new_n1179, new_n1169, new_n1180);
nor_1  g00804(new_n1180, new_n1178, new_n1181);
xnor_1 g00805(new_n1181, new_n1166, new_n1182);
not_4  g00806(new_n1139, new_n1183);
nor_1  g00807(new_n1153, new_n1183, new_n1184);
not_4  g00808(new_n1184, new_n1185);
nand_1 g00809(new_n1161, new_n1154, new_n1186);
nand_1 g00810(new_n1186, new_n1185, new_n1187);
nand_1 g00811(n9111, n7388, new_n1188);
not_4  g00812(new_n1188, new_n1189);
nand_1 g00813(new_n1189, new_n1137, new_n1190);
nand_1 g00814(n11892, n3342, new_n1191);
not_4  g00815(new_n1191, new_n1192);
nand_1 g00816(new_n1192, new_n1138_1, new_n1193);
nand_1 g00817(n11892, n9763, new_n1194);
nand_1 g00818(n7965, n3342, new_n1195);
nand_1 g00819(new_n1195, new_n1194, new_n1196);
nand_1 g00820(new_n1196, new_n1193, new_n1197);
nand_1 g00821(new_n1197, new_n1190, new_n1198_1);
not_4  g00822(new_n1198_1, new_n1199_1);
not_4  g00823(new_n1196, new_n1200);
nor_1  g00824(new_n1200, new_n1190, new_n1201);
nor_1  g00825(new_n1201, new_n1199_1, new_n1202);
xnor_1 g00826(new_n1202, new_n1187, new_n1203);
nand_1 g00827(n8476, n2498, new_n1204);
not_4  g00828(new_n1204, new_n1205);
nand_1 g00829(new_n1205, new_n1135, new_n1206);
not_4  g00830(new_n1206, new_n1207);
nand_1 g00831(n2558, n2530, new_n1208);
nand_1 g00832(n5579, n5331, new_n1209_1);
nand_1 g00833(new_n1209_1, new_n1208, new_n1210);
not_4  g00834(new_n1210, new_n1211);
nand_1 g00835(new_n1211, new_n1207, new_n1212);
nand_1 g00836(n5579, n2530, new_n1213);
not_4  g00837(new_n1213, new_n1214);
nand_1 g00838(new_n1214, new_n1136_1, new_n1215);
nand_1 g00839(new_n1215, new_n1210, new_n1216);
not_4  g00840(new_n1216, new_n1217);
nand_1 g00841(new_n1217, new_n1206, new_n1218);
nand_1 g00842(new_n1218, new_n1212, new_n1219);
xnor_1 g00843(new_n1219, new_n1203, new_n1220);
xnor_1 g00844(new_n1220, new_n1182, new_n1221);
not_4  g00845(new_n1221, new_n1222);
nor_1  g00846(new_n1222, new_n1132, new_n1223);
not_4  g00847(new_n1223, new_n1224);
xnor_1 g00848(new_n1142, new_n1133, new_n1225);
nand_1 g00849(new_n1225, new_n1102, new_n1226);
nand_1 g00850(n7265, n5964, new_n1227);
nand_1 g00851(n5305, n2879, new_n1228);
xnor_1 g00852(new_n1228, new_n1227, new_n1229);
nand_1 g00853(new_n1229, new_n1226, new_n1230);
xnor_1 g00854(new_n1163, new_n1162, new_n1231);
not_4  g00855(new_n1231, new_n1232);
xnor_1 g00856(new_n1229, new_n1226, new_n1233);
nor_1  g00857(new_n1233, new_n1232, new_n1234);
not_4  g00858(new_n1234, new_n1235);
nand_1 g00859(new_n1235, new_n1230, new_n1236);
not_4  g00860(new_n1236, new_n1237);
xnor_1 g00861(new_n1221, new_n1132, new_n1238);
nand_1 g00862(new_n1238, new_n1237, new_n1239);
nand_1 g00863(new_n1239, new_n1224, new_n1240);
xnor_1 g00864(new_n1240, new_n1129, new_n1241);
not_4  g00865(new_n1241, new_n1242);
nand_1 g00866(n8759, n2522, new_n1243);
nand_1 g00867(new_n1175, new_n1167, new_n1244);
nand_1 g00868(new_n1244, new_n1172, new_n1245);
xnor_1 g00869(new_n1245, new_n1243, new_n1246);
nand_1 g00870(n12299, n2024, new_n1247);
not_4  g00871(new_n1247, new_n1248);
nand_1 g00872(n7946, n7436, new_n1249);
nand_1 g00873(n9189, n6776, new_n1250);
nand_1 g00874(new_n1250, new_n1249, new_n1251);
not_4  g00875(new_n1249, new_n1252);
not_4  g00876(new_n1250, new_n1253);
nand_1 g00877(new_n1253, new_n1252, new_n1254);
nand_1 g00878(new_n1254, new_n1251, new_n1255);
xnor_1 g00879(new_n1255, new_n1248, new_n1256);
not_4  g00880(new_n1256, new_n1257);
nor_1  g00881(new_n1257, new_n1246, new_n1258);
not_4  g00882(new_n1258, new_n1259);
nand_1 g00883(new_n1257, new_n1246, new_n1260);
nand_1 g00884(new_n1260, new_n1259, new_n1261);
nand_1 g00885(new_n1178, new_n1168, new_n1262);
nand_1 g00886(new_n1262, new_n1261, new_n1263);
not_4  g00887(new_n1261, new_n1264);
not_4  g00888(new_n1262, new_n1265);
nand_1 g00889(new_n1265, new_n1264, new_n1266);
nand_1 g00890(new_n1266, new_n1263, new_n1267);
not_4  g00891(new_n1181, new_n1268);
nand_1 g00892(new_n1268, new_n1166, new_n1269_1);
nand_1 g00893(new_n1220, new_n1182, new_n1270);
nand_1 g00894(new_n1270, new_n1269_1, new_n1271);
not_4  g00895(new_n1271, new_n1272);
xnor_1 g00896(new_n1272, new_n1267, new_n1273);
nand_1 g00897(n5331, n521, new_n1274);
nand_1 g00898(new_n1215, new_n1204, new_n1275);
nand_1 g00899(new_n1275, new_n1210, new_n1276);
not_4  g00900(new_n1276, new_n1277);
xnor_1 g00901(new_n1277, new_n1274, new_n1278);
nand_1 g00902(n2530, n2498, new_n1279);
nand_1 g00903(n12648, n2558, new_n1280);
nand_1 g00904(n8476, n5579, new_n1281);
nand_1 g00905(new_n1281, new_n1280, new_n1282);
not_4  g00906(new_n1280, new_n1283);
not_4  g00907(new_n1281, new_n1284);
nand_1 g00908(new_n1284, new_n1283, new_n1285);
nand_1 g00909(new_n1285, new_n1282, new_n1286);
xnor_1 g00910(new_n1286, new_n1279, new_n1287);
not_4  g00911(new_n1287, new_n1288);
xnor_1 g00912(new_n1288, new_n1278, new_n1289);
nor_1  g00913(new_n1217, new_n1160, new_n1290);
xnor_1 g00914(new_n1290, new_n1289, new_n1291);
nand_1 g00915(n7965, n806, new_n1292);
nand_1 g00916(new_n1196, new_n1189, new_n1293);
nand_1 g00917(new_n1293, new_n1193, new_n1294);
xnor_1 g00918(new_n1294, new_n1292, new_n1295);
not_4  g00919(new_n1295, new_n1296);
nand_1 g00920(n11892, n9111, new_n1297);
nand_1 g00921(n9763, n2393, new_n1298);
nand_1 g00922(n7388, n3342, new_n1299);
nand_1 g00923(new_n1299, new_n1298, new_n1300);
not_4  g00924(new_n1298, new_n1301);
not_4  g00925(new_n1299, new_n1302);
nand_1 g00926(new_n1302, new_n1301, new_n1303);
nand_1 g00927(new_n1303, new_n1300, new_n1304);
xnor_1 g00928(new_n1304, new_n1297, new_n1305);
xnor_1 g00929(new_n1305, new_n1296, new_n1306);
not_4  g00930(new_n1306, new_n1307);
nand_1 g00931(new_n1199_1, new_n1189, new_n1308);
xnor_1 g00932(new_n1308, new_n1307, new_n1309);
nand_1 g00933(new_n1309, new_n1291, new_n1310);
nor_1  g00934(new_n1309, new_n1291, new_n1311);
not_4  g00935(new_n1311, new_n1312);
nand_1 g00936(new_n1312, new_n1310, new_n1313);
not_4  g00937(new_n1202, new_n1314);
nand_1 g00938(new_n1314, new_n1187, new_n1315);
not_4  g00939(new_n1219, new_n1316);
nand_1 g00940(new_n1316, new_n1203, new_n1317);
nand_1 g00941(new_n1317, new_n1315, new_n1318);
not_4  g00942(new_n1318, new_n1319);
nand_1 g00943(new_n1319, new_n1313, new_n1320);
nor_1  g00944(new_n1319, new_n1313, new_n1321);
not_4  g00945(new_n1321, new_n1322);
nand_1 g00946(new_n1322, new_n1320, new_n1323);
xnor_1 g00947(new_n1323, new_n1273, new_n1324);
xnor_1 g00948(new_n1324, new_n1242, n381);
nand_1 g00949(n7862, n6038, new_n1326);
nand_1 g00950(n7354, n6877, new_n1327);
nand_1 g00951(n4805, n1564, new_n1328);
not_4  g00952(new_n1328, new_n1329);
nand_1 g00953(n8028, n7236, new_n1330);
not_4  g00954(new_n1330, new_n1331);
nand_1 g00955(new_n1331, new_n1329, new_n1332);
nand_1 g00956(new_n1330, new_n1328, new_n1333_1);
nand_1 g00957(new_n1333_1, new_n1332, new_n1334);
not_4  g00958(new_n1334, new_n1335);
xnor_1 g00959(new_n1335, new_n1327, new_n1336);
xnor_1 g00960(new_n1336, new_n1326, n397);
nand_1 g00961(n6687, n4370, new_n1338);
nand_1 g00962(n11407, n4189, new_n1339);
nand_1 g00963(n11877, n6687, new_n1340);
nand_1 g00964(new_n1340, new_n1339, new_n1341);
not_4  g00965(new_n1339, new_n1342);
not_4  g00966(new_n1340, new_n1343);
nand_1 g00967(new_n1343, new_n1342, new_n1344);
nand_1 g00968(n5212, n2564, new_n1345);
nand_1 g00969(new_n1345, new_n1344, new_n1346);
nand_1 g00970(new_n1346, new_n1341, new_n1347);
xnor_1 g00971(new_n1347, new_n1338, new_n1348);
nand_1 g00972(n5212, n4189, new_n1349);
nand_1 g00973(n11407, n6770, new_n1350);
nand_1 g00974(n11877, n2564, new_n1351);
xnor_1 g00975(new_n1351, new_n1350, new_n1352);
xnor_1 g00976(new_n1352, new_n1349, new_n1353_1);
xnor_1 g00977(new_n1353_1, new_n1348, new_n1354);
not_4  g00978(new_n1345, new_n1355);
not_4  g00979(new_n1341, new_n1356);
nand_1 g00980(n11407, n6687, new_n1357_1);
nand_1 g00981(new_n1357_1, new_n1355, new_n1358);
nand_1 g00982(new_n1358, new_n1356, new_n1359);
nand_1 g00983(new_n1359, new_n1344, new_n1360);
nand_1 g00984(new_n1360, new_n1355, new_n1361);
nor_1  g00985(new_n1361, new_n1354, new_n1362);
not_4  g00986(new_n1362, new_n1363);
nand_1 g00987(new_n1361, new_n1354, new_n1364);
nand_1 g00988(new_n1364, new_n1363, new_n1365);
nand_1 g00989(n12709, n8336, new_n1366);
not_4  g00990(new_n1366, new_n1367);
nand_1 g00991(n11222, n10990, new_n1368);
not_4  g00992(new_n1368, new_n1369);
nand_1 g00993(n12489, n12069, new_n1370);
not_4  g00994(new_n1370, new_n1371);
nand_1 g00995(new_n1371, new_n1369, new_n1372);
nand_1 g00996(new_n1370, new_n1368, new_n1373);
nand_1 g00997(new_n1373, new_n1372, new_n1374);
not_4  g00998(new_n1374, new_n1375);
nand_1 g00999(new_n1375, new_n1367, new_n1376);
nand_1 g01000(n11728, n8336, new_n1377);
nand_1 g01001(n12709, n10928, new_n1378);
xnor_1 g01002(new_n1378, new_n1377, new_n1379);
nand_1 g01003(new_n1379, new_n1376, new_n1380);
nand_1 g01004(n11222, n5760, new_n1381);
nand_1 g01005(n11153, n10990, new_n1382);
not_4  g01006(new_n1382, new_n1383);
xnor_1 g01007(new_n1383, new_n1381, new_n1384);
xnor_1 g01008(new_n1384, new_n1372, new_n1385);
not_4  g01009(new_n1385, new_n1386);
nand_1 g01010(n12069, n7159, new_n1387);
nand_1 g01011(n12489, n12391, new_n1388);
xnor_1 g01012(new_n1388, new_n1387, new_n1389);
not_4  g01013(new_n1389, new_n1390);
xnor_1 g01014(new_n1390, new_n1386, new_n1391);
not_4  g01015(new_n1391, new_n1392);
xnor_1 g01016(new_n1379, new_n1376, new_n1393);
not_4  g01017(new_n1393, new_n1394);
nand_1 g01018(new_n1394, new_n1392, new_n1395);
nand_1 g01019(new_n1395, new_n1380, new_n1396);
nand_1 g01020(n11728, n10928, new_n1397);
not_4  g01021(new_n1397, new_n1398);
nand_1 g01022(new_n1398, new_n1366, new_n1399);
nand_1 g01023(n6986, n6429, new_n1400);
not_4  g01024(new_n1400, new_n1401);
nand_1 g01025(new_n1401, new_n1367, new_n1402);
nand_1 g01026(n12709, n6986, new_n1403);
nand_1 g01027(n8336, n6429, new_n1404);
nand_1 g01028(new_n1404, new_n1403, new_n1405);
nand_1 g01029(new_n1405, new_n1402, new_n1406);
nand_1 g01030(new_n1406, new_n1399, new_n1407);
not_4  g01031(new_n1407, new_n1408);
not_4  g01032(new_n1405, new_n1409);
nor_1  g01033(new_n1409, new_n1399, new_n1410);
nor_1  g01034(new_n1410, new_n1408, new_n1411);
xnor_1 g01035(new_n1411, new_n1396, new_n1412);
nand_1 g01036(n12391, n7159, new_n1413);
not_4  g01037(new_n1413, new_n1414);
nand_1 g01038(new_n1414, new_n1370, new_n1415);
nand_1 g01039(n12489, n7891, new_n1416);
nand_1 g01040(n12777, n12069, new_n1417);
nand_1 g01041(new_n1417, new_n1416, new_n1418);
not_4  g01042(new_n1418, new_n1419);
nand_1 g01043(new_n1419, new_n1415, new_n1420);
not_4  g01044(new_n1416, new_n1421);
not_4  g01045(new_n1417, new_n1422);
nand_1 g01046(new_n1422, new_n1421, new_n1423);
nand_1 g01047(new_n1423, new_n1420, new_n1424);
nor_1  g01048(new_n1419, new_n1415, new_n1425);
nor_1  g01049(new_n1425, new_n1424, new_n1426);
nand_1 g01050(n11153, n5760, new_n1427);
not_4  g01051(new_n1427, new_n1428);
nand_1 g01052(new_n1428, new_n1368, new_n1429);
nand_1 g01053(n10990, n5314, new_n1430);
nand_1 g01054(n11222, n1478, new_n1431);
nand_1 g01055(new_n1431, new_n1430, new_n1432);
not_4  g01056(new_n1430, new_n1433);
not_4  g01057(new_n1431, new_n1434);
nand_1 g01058(new_n1434, new_n1433, new_n1435);
nand_1 g01059(new_n1435, new_n1432, new_n1436);
nand_1 g01060(new_n1436, new_n1429, new_n1437);
not_4  g01061(new_n1437, new_n1438);
not_4  g01062(new_n1432, new_n1439);
nor_1  g01063(new_n1439, new_n1429, new_n1440);
nor_1  g01064(new_n1440, new_n1438, new_n1441);
xnor_1 g01065(new_n1441, new_n1426, new_n1442);
not_4  g01066(new_n1372, new_n1443);
nand_1 g01067(new_n1384, new_n1443, new_n1444);
nand_1 g01068(new_n1390, new_n1385, new_n1445);
nand_1 g01069(new_n1445, new_n1444, new_n1446);
xnor_1 g01070(new_n1446, new_n1442, new_n1447);
xnor_1 g01071(new_n1447, new_n1412, new_n1448);
not_4  g01072(new_n1448, new_n1449);
nor_1  g01073(new_n1358, new_n1356, new_n1450);
nor_1  g01074(new_n1450, new_n1360, new_n1451);
nor_1  g01075(new_n1451, new_n1449, new_n1452);
xnor_1 g01076(new_n1451, new_n1449, new_n1453);
not_4  g01077(new_n1357_1, new_n1454);
xnor_1 g01078(new_n1375, new_n1366, new_n1455);
nand_1 g01079(new_n1455, new_n1454, new_n1456);
nand_1 g01080(n11407, n2564, new_n1457);
nand_1 g01081(n6687, n5212, new_n1458);
xnor_1 g01082(new_n1458, new_n1457, new_n1459);
nand_1 g01083(new_n1459, new_n1456, new_n1460);
xnor_1 g01084(new_n1394, new_n1391, new_n1461);
not_4  g01085(new_n1461, new_n1462);
xnor_1 g01086(new_n1459, new_n1456, new_n1463);
nor_1  g01087(new_n1463, new_n1462, new_n1464);
not_4  g01088(new_n1464, new_n1465);
nand_1 g01089(new_n1465, new_n1460, new_n1466);
not_4  g01090(new_n1466, new_n1467);
nor_1  g01091(new_n1467, new_n1453, new_n1468);
nor_1  g01092(new_n1468, new_n1452, new_n1469);
xnor_1 g01093(new_n1469, new_n1365, new_n1470);
not_4  g01094(new_n1470, new_n1471_1);
nand_1 g01095(n8819, n8336, new_n1472);
nand_1 g01096(n11728, n6986, new_n1473);
not_4  g01097(new_n1473, new_n1474);
nand_1 g01098(n10928, n6429, new_n1475);
nand_1 g01099(n12709, n2226, new_n1476);
nand_1 g01100(new_n1476, new_n1475, new_n1477);
not_4  g01101(new_n1475, new_n1478_1);
not_4  g01102(new_n1476, new_n1479);
nand_1 g01103(new_n1479, new_n1478_1, new_n1480);
nand_1 g01104(new_n1480, new_n1477, new_n1481);
xnor_1 g01105(new_n1481, new_n1474, new_n1482);
xnor_1 g01106(new_n1482, new_n1472, new_n1483);
nand_1 g01107(new_n1405, new_n1398, new_n1484);
nand_1 g01108(new_n1484, new_n1402, new_n1485);
not_4  g01109(new_n1485, new_n1486);
xnor_1 g01110(new_n1486, new_n1483, new_n1487);
nand_1 g01111(new_n1408, new_n1398, new_n1488);
xnor_1 g01112(new_n1488, new_n1487, new_n1489);
nand_1 g01113(n12069, n6254, new_n1490);
nand_1 g01114(new_n1423, new_n1413, new_n1491);
nand_1 g01115(new_n1491, new_n1418, new_n1492);
nor_1  g01116(new_n1492, new_n1490, new_n1493);
not_4  g01117(new_n1493, new_n1494);
nand_1 g01118(new_n1492, new_n1490, new_n1495);
nand_1 g01119(new_n1495, new_n1494, new_n1496);
nand_1 g01120(n12489, n7160, new_n1497);
nand_1 g01121(n12777, n12391, new_n1498);
nand_1 g01122(n7891, n7159, new_n1499);
not_4  g01123(new_n1499, new_n1500);
xnor_1 g01124(new_n1500, new_n1498, new_n1501);
not_4  g01125(new_n1501, new_n1502);
xnor_1 g01126(new_n1502, new_n1497, new_n1503);
nor_1  g01127(new_n1503, new_n1496, new_n1504);
not_4  g01128(new_n1504, new_n1505);
nand_1 g01129(new_n1503, new_n1496, new_n1506);
nand_1 g01130(new_n1506, new_n1505, new_n1507);
nand_1 g01131(new_n1424, new_n1414, new_n1508);
nand_1 g01132(new_n1508, new_n1507, new_n1509);
nor_1  g01133(new_n1508, new_n1507, new_n1510_1);
not_4  g01134(new_n1510_1, new_n1511);
nand_1 g01135(new_n1511, new_n1509, new_n1512_1);
not_4  g01136(new_n1512_1, new_n1513);
nand_1 g01137(n11791, n11222, new_n1514);
nand_1 g01138(new_n1435, new_n1427, new_n1515);
nand_1 g01139(new_n1515, new_n1432, new_n1516);
nor_1  g01140(new_n1516, new_n1514, new_n1517);
not_4  g01141(new_n1517, new_n1518);
nand_1 g01142(new_n1516, new_n1514, new_n1519);
nand_1 g01143(new_n1519, new_n1518, new_n1520);
nand_1 g01144(n5760, n5314, new_n1521);
not_4  g01145(new_n1521, new_n1522);
nand_1 g01146(n10990, n996, new_n1523_1);
nand_1 g01147(n11153, n1478, new_n1524);
nand_1 g01148(new_n1524, new_n1523_1, new_n1525);
not_4  g01149(new_n1525, new_n1526);
nor_1  g01150(new_n1524, new_n1523_1, new_n1527);
nor_1  g01151(new_n1527, new_n1526, new_n1528);
xnor_1 g01152(new_n1528, new_n1522, new_n1529);
nor_1  g01153(new_n1529, new_n1520, new_n1530);
not_4  g01154(new_n1530, new_n1531);
nand_1 g01155(new_n1529, new_n1520, new_n1532);
nand_1 g01156(new_n1532, new_n1531, new_n1533);
not_4  g01157(new_n1533, new_n1534);
nand_1 g01158(new_n1438, new_n1428, new_n1535);
not_4  g01159(new_n1535, new_n1536);
nand_1 g01160(new_n1536, new_n1534, new_n1537);
nand_1 g01161(new_n1535, new_n1533, new_n1538);
nand_1 g01162(new_n1538, new_n1537, new_n1539);
not_4  g01163(new_n1539, new_n1540);
nand_1 g01164(new_n1540, new_n1513, new_n1541);
nand_1 g01165(new_n1539, new_n1512_1, new_n1542);
nand_1 g01166(new_n1542, new_n1541, new_n1543);
nand_1 g01167(new_n1441, new_n1426, new_n1544);
not_4  g01168(new_n1442, new_n1545);
nand_1 g01169(new_n1446, new_n1545, new_n1546);
nand_1 g01170(new_n1546, new_n1544, new_n1547);
nor_1  g01171(new_n1547, new_n1543, new_n1548);
not_4  g01172(new_n1548, new_n1549);
nand_1 g01173(new_n1547, new_n1543, new_n1550);
nand_1 g01174(new_n1550, new_n1549, new_n1551);
xnor_1 g01175(new_n1551, new_n1489, new_n1552);
not_4  g01176(new_n1552, new_n1553);
not_4  g01177(new_n1411, new_n1554);
nand_1 g01178(new_n1554, new_n1396, new_n1555);
not_4  g01179(new_n1447, new_n1556);
nand_1 g01180(new_n1556, new_n1412, new_n1557);
nand_1 g01181(new_n1557, new_n1555, new_n1558);
xnor_1 g01182(new_n1558, new_n1553, new_n1559);
xnor_1 g01183(new_n1559, new_n1471_1, n658);
nand_1 g01184(n7862, n2585, new_n1561);
nand_1 g01185(n2508, n1333, new_n1562);
nand_1 g01186(n11757, n6038, new_n1563);
nand_1 g01187(n12720, n1333, new_n1564_1);
nand_1 g01188(new_n1564_1, new_n1563, new_n1565);
not_4  g01189(new_n1563, new_n1566);
not_4  g01190(new_n1564_1, new_n1567);
nand_1 g01191(new_n1567, new_n1566, new_n1568);
nand_1 g01192(n3172, n2509, new_n1569);
nand_1 g01193(new_n1569, new_n1568, new_n1570);
nand_1 g01194(new_n1570, new_n1565, new_n1571);
not_4  g01195(new_n1571, new_n1572);
xnor_1 g01196(new_n1572, new_n1562, new_n1573);
not_4  g01197(new_n1573, new_n1574);
nand_1 g01198(n11757, n2509, new_n1575);
nand_1 g01199(n6038, n5240, new_n1576_1);
nand_1 g01200(n12720, n3172, new_n1577);
not_4  g01201(new_n1577, new_n1578);
xnor_1 g01202(new_n1578, new_n1576_1, new_n1579);
not_4  g01203(new_n1579, new_n1580);
xnor_1 g01204(new_n1580, new_n1575, new_n1581);
xnor_1 g01205(new_n1581, new_n1574, new_n1582);
nand_1 g01206(new_n1582, new_n1561, new_n1583);
xnor_1 g01207(new_n1582, new_n1561, new_n1584);
nand_1 g01208(n7862, n2508, new_n1585);
not_4  g01209(new_n1585, new_n1586);
nand_1 g01210(n2509, n1333, new_n1587);
not_4  g01211(new_n1587, new_n1588);
nand_1 g01212(n6038, n3172, new_n1589);
nand_1 g01213(n12720, n7862, new_n1590);
nand_1 g01214(new_n1590, new_n1589, new_n1591);
nand_1 g01215(new_n1591, new_n1588, new_n1592);
nor_1  g01216(new_n1590, new_n1589, new_n1593);
not_4  g01217(new_n1593, new_n1594);
nand_1 g01218(new_n1594, new_n1592, new_n1595);
nand_1 g01219(new_n1595, new_n1586, new_n1596);
xnor_1 g01220(new_n1595, new_n1585, new_n1597);
not_4  g01221(new_n1597, new_n1598);
nand_1 g01222(new_n1568, new_n1565, new_n1599);
xnor_1 g01223(new_n1599, new_n1569, new_n1600);
nor_1  g01224(new_n1600, new_n1598, new_n1601);
not_4  g01225(new_n1601, new_n1602);
nand_1 g01226(new_n1602, new_n1596, new_n1603);
nor_1  g01227(new_n1603, new_n1584, new_n1604);
not_4  g01228(new_n1604, new_n1605);
nand_1 g01229(new_n1605, new_n1583, new_n1606);
not_4  g01230(new_n1606, new_n1607);
nand_1 g01231(n12720, n11757, new_n1608);
nand_1 g01232(n5240, n2509, new_n1609);
not_4  g01233(new_n1609, new_n1610);
nand_1 g01234(n11821, n6038, new_n1611);
not_4  g01235(new_n1611, new_n1612);
nand_1 g01236(new_n1612, new_n1610, new_n1613);
nand_1 g01237(new_n1611, new_n1609, new_n1614);
nand_1 g01238(new_n1614, new_n1613, new_n1615);
not_4  g01239(new_n1615, new_n1616);
xnor_1 g01240(new_n1616, new_n1608, new_n1617);
not_4  g01241(new_n1617, new_n1618);
nand_1 g01242(new_n1577, new_n1576_1, new_n1619);
nand_1 g01243(new_n1579, new_n1575, new_n1620);
nand_1 g01244(new_n1620, new_n1619, new_n1621);
nor_1  g01245(new_n1621, new_n1618, new_n1622);
not_4  g01246(new_n1622, new_n1623);
nand_1 g01247(new_n1621, new_n1618, new_n1624);
nand_1 g01248(new_n1624, new_n1623, new_n1625);
not_4  g01249(new_n1625, new_n1626);
nor_1  g01250(new_n1571, new_n1562, new_n1627);
nor_1  g01251(new_n1581, new_n1574, new_n1628);
nor_1  g01252(new_n1628, new_n1627, new_n1629);
nand_1 g01253(n2585, n1333, new_n1630);
not_4  g01254(new_n1630, new_n1631);
nand_1 g01255(n3172, n2508, new_n1632);
not_4  g01256(new_n1632, new_n1633);
nand_1 g01257(new_n1633, new_n1631, new_n1634);
nand_1 g01258(new_n1632, new_n1630, new_n1635);
nand_1 g01259(new_n1635, new_n1634, new_n1636);
nand_1 g01260(new_n1636, new_n1629, new_n1637);
nor_1  g01261(new_n1636, new_n1629, new_n1638);
not_4  g01262(new_n1638, new_n1639);
nand_1 g01263(new_n1639, new_n1637, new_n1640);
xnor_1 g01264(new_n1640, new_n1626, new_n1641);
nand_1 g01265(new_n1641, new_n1607, new_n1642);
nand_1 g01266(new_n1637, new_n1626, new_n1643);
xnor_1 g01267(new_n1643, new_n1634, new_n1644);
nand_1 g01268(new_n1644, new_n1639, new_n1645);
nand_1 g01269(n11757, n2508, new_n1646);
xnor_1 g01270(new_n1646, new_n1613, new_n1647);
nand_1 g01271(n11821, n2509, new_n1648);
not_4  g01272(new_n1648, new_n1649);
nand_1 g01273(n12720, n5240, new_n1650);
nand_1 g01274(n9080, n6038, new_n1651);
not_4  g01275(new_n1651, new_n1652);
xnor_1 g01276(new_n1652, new_n1650, new_n1653);
xnor_1 g01277(new_n1653, new_n1649, new_n1654);
xnor_1 g01278(new_n1654, new_n1647, new_n1655);
not_4  g01279(new_n1655, new_n1656);
not_4  g01280(new_n1608, new_n1657);
nand_1 g01281(new_n1616, new_n1657, new_n1658_1);
nand_1 g01282(new_n1623, new_n1658_1, new_n1659);
nand_1 g01283(n4005, n1333, new_n1660);
nand_1 g01284(n3172, n2585, new_n1661);
nand_1 g01285(n12706, n7862, new_n1662);
nand_1 g01286(new_n1662, new_n1661, new_n1663);
not_4  g01287(new_n1661, new_n1664);
not_4  g01288(new_n1662, new_n1665);
nand_1 g01289(new_n1665, new_n1664, new_n1666);
nand_1 g01290(new_n1666, new_n1663, new_n1667);
xnor_1 g01291(new_n1667, new_n1660, new_n1668);
xnor_1 g01292(new_n1668, new_n1659, new_n1669);
xnor_1 g01293(new_n1669, new_n1656, new_n1670);
xnor_1 g01294(new_n1670, new_n1645, new_n1671);
xnor_1 g01295(new_n1671, new_n1642, new_n1672);
nand_1 g01296(n7862, n4005, new_n1673);
not_4  g01297(new_n1673, new_n1674);
xnor_1 g01298(new_n1641, new_n1606, new_n1675);
nand_1 g01299(new_n1675, new_n1674, new_n1676);
xnor_1 g01300(new_n1600, new_n1597, new_n1677);
nand_1 g01301(new_n1594, new_n1591, new_n1678);
not_4  g01302(new_n1678, new_n1679);
nand_1 g01303(n6038, n1333, new_n1680);
not_4  g01304(new_n1680, new_n1681);
nand_1 g01305(n7862, n2509, new_n1682);
not_4  g01306(new_n1682, new_n1683);
nand_1 g01307(new_n1683, new_n1681, new_n1684);
nor_1  g01308(new_n1684, new_n1679, new_n1685);
nand_1 g01309(new_n1685, new_n1677, new_n1686);
not_4  g01310(new_n1686, new_n1687);
nand_1 g01311(new_n1603, new_n1584, new_n1688);
nand_1 g01312(new_n1688, new_n1605, new_n1689);
nand_1 g01313(new_n1689, new_n1687, new_n1690);
not_4  g01314(new_n1690, new_n1691);
xnor_1 g01315(new_n1675, new_n1673, new_n1692);
nand_1 g01316(new_n1692, new_n1691, new_n1693);
nand_1 g01317(new_n1693, new_n1676, new_n1694);
xnor_1 g01318(new_n1694, new_n1672, new_n1695);
nand_1 g01319(n6877, n5105, new_n1696);
nand_1 g01320(n6877, n1209, new_n1697);
not_4  g01321(new_n1697, new_n1698);
nand_1 g01322(n7354, n2464, new_n1699);
not_4  g01323(new_n1699, new_n1700);
nand_1 g01324(new_n1700, new_n1698, new_n1701);
nand_1 g01325(new_n1699, new_n1697, new_n1702);
nand_1 g01326(n9400, n7500, new_n1703);
not_4  g01327(new_n1703, new_n1704);
nand_1 g01328(new_n1704, new_n1702, new_n1705);
nand_1 g01329(new_n1705, new_n1701, new_n1706);
xnor_1 g01330(new_n1706, new_n1696, new_n1707);
nand_1 g01331(n7500, n2464, new_n1708);
not_4  g01332(new_n1708, new_n1709);
nand_1 g01333(n9400, n1209, new_n1710);
nand_1 g01334(n11311, n7354, new_n1711);
nand_1 g01335(new_n1711, new_n1710, new_n1712);
not_4  g01336(new_n1710, new_n1713);
not_4  g01337(new_n1711, new_n1714);
nand_1 g01338(new_n1714, new_n1713, new_n1715);
nand_1 g01339(new_n1715, new_n1712, new_n1716);
xnor_1 g01340(new_n1716, new_n1709, new_n1717);
xnor_1 g01341(new_n1717, new_n1707, new_n1718);
not_4  g01342(new_n1718, new_n1719);
nand_1 g01343(new_n1702, new_n1701, new_n1720);
not_4  g01344(new_n1720, new_n1721);
nand_1 g01345(n9400, n7354, new_n1722);
not_4  g01346(new_n1722, new_n1723);
nand_1 g01347(n7500, n6877, new_n1724);
not_4  g01348(new_n1724, new_n1725);
nand_1 g01349(new_n1725, new_n1723, new_n1726);
nor_1  g01350(new_n1726, new_n1721, new_n1727);
nand_1 g01351(new_n1727, new_n1719, new_n1728);
not_4  g01352(new_n1728, new_n1729);
nand_1 g01353(n11311, n7500, new_n1730);
nand_1 g01354(n2464, n1209, new_n1731);
nand_1 g01355(n7354, n4187, new_n1732);
not_4  g01356(new_n1732, new_n1733);
xnor_1 g01357(new_n1733, new_n1731, new_n1734);
xnor_1 g01358(new_n1734, new_n1730, new_n1735);
nand_1 g01359(n9400, n5105, new_n1736);
nand_1 g01360(new_n1715, new_n1708, new_n1737);
nand_1 g01361(new_n1737, new_n1712, new_n1738);
not_4  g01362(new_n1738, new_n1739);
xnor_1 g01363(new_n1739, new_n1736, new_n1740);
xnor_1 g01364(new_n1740, new_n1735, new_n1741);
nand_1 g01365(n6877, n4141, new_n1742);
not_4  g01366(new_n1696, new_n1743);
nand_1 g01367(new_n1706, new_n1743, new_n1744);
nand_1 g01368(new_n1717, new_n1707, new_n1745);
nand_1 g01369(new_n1745, new_n1744, new_n1746);
xnor_1 g01370(new_n1746, new_n1742, new_n1747);
xnor_1 g01371(new_n1747, new_n1741, new_n1748);
nand_1 g01372(new_n1748, new_n1729, new_n1749);
nand_1 g01373(n6877, n4928, new_n1750);
not_4  g01374(new_n1742, new_n1751);
nor_1  g01375(new_n1746, new_n1751, new_n1752);
not_4  g01376(new_n1752, new_n1753);
nand_1 g01377(new_n1747, new_n1741, new_n1754);
nand_1 g01378(new_n1754, new_n1753, new_n1755);
nand_1 g01379(n11311, n1209, new_n1756);
nand_1 g01380(n7500, n4187, new_n1757);
nand_1 g01381(n7354, n4203, new_n1758);
nand_1 g01382(new_n1758, new_n1757, new_n1759);
not_4  g01383(new_n1757, new_n1760);
not_4  g01384(new_n1758, new_n1761);
nand_1 g01385(new_n1761, new_n1760, new_n1762);
nand_1 g01386(new_n1762, new_n1759, new_n1763);
not_4  g01387(new_n1763, new_n1764);
xnor_1 g01388(new_n1764, new_n1756, new_n1765);
not_4  g01389(new_n1765, new_n1766);
nand_1 g01390(new_n1732, new_n1731, new_n1767);
nand_1 g01391(new_n1734, new_n1730, new_n1768);
nand_1 g01392(new_n1768, new_n1767, new_n1769);
nor_1  g01393(new_n1769, new_n1766, new_n1770);
not_4  g01394(new_n1770, new_n1771);
nand_1 g01395(new_n1769, new_n1766, new_n1772);
nand_1 g01396(new_n1772, new_n1771, new_n1773);
not_4  g01397(new_n1773, new_n1774);
nor_1  g01398(new_n1738, new_n1736, new_n1775);
not_4  g01399(new_n1775, new_n1776);
nand_1 g01400(new_n1740, new_n1735, new_n1777);
nand_1 g01401(new_n1777, new_n1776, new_n1778);
nand_1 g01402(n9400, n4141, new_n1779);
not_4  g01403(new_n1779, new_n1780);
nand_1 g01404(n5105, n2464, new_n1781);
not_4  g01405(new_n1781, new_n1782);
nand_1 g01406(new_n1782, new_n1780, new_n1783);
nand_1 g01407(new_n1781, new_n1779, new_n1784);
nand_1 g01408(new_n1784, new_n1783, new_n1785);
not_4  g01409(new_n1785, new_n1786);
nor_1  g01410(new_n1786, new_n1778, new_n1787);
not_4  g01411(new_n1787, new_n1788);
nand_1 g01412(new_n1786, new_n1778, new_n1789);
nand_1 g01413(new_n1789, new_n1788, new_n1790);
xnor_1 g01414(new_n1790, new_n1774, new_n1791);
xnor_1 g01415(new_n1791, new_n1755, new_n1792);
xnor_1 g01416(new_n1792, new_n1750, new_n1793);
xnor_1 g01417(new_n1793, new_n1749, new_n1794);
not_4  g01418(new_n1794, new_n1795);
nand_1 g01419(n7294, n7236, new_n1796);
nand_1 g01420(n10848, n3992, new_n1797);
not_4  g01421(new_n1797, new_n1798_1);
nand_1 g01422(n8384, n8028, new_n1799);
nand_1 g01423(n7236, n1980, new_n1800);
nand_1 g01424(new_n1800, new_n1799, new_n1801);
nand_1 g01425(new_n1801, new_n1798_1, new_n1802);
not_4  g01426(new_n1799, new_n1803);
not_4  g01427(new_n1800, new_n1804);
nand_1 g01428(new_n1804, new_n1803, new_n1805);
nand_1 g01429(new_n1805, new_n1802, new_n1806);
xnor_1 g01430(new_n1806, new_n1796, new_n1807);
nand_1 g01431(n8028, n6358, new_n1808);
not_4  g01432(new_n1808, new_n1809);
nand_1 g01433(n10848, n8384, new_n1810);
nand_1 g01434(n3992, n1980, new_n1811);
xnor_1 g01435(new_n1811, new_n1810, new_n1812);
xnor_1 g01436(new_n1812, new_n1809, new_n1813);
xnor_1 g01437(new_n1813, new_n1807, new_n1814);
not_4  g01438(new_n1814, new_n1815);
nand_1 g01439(new_n1805, new_n1801, new_n1816);
not_4  g01440(new_n1816, new_n1817);
nand_1 g01441(n10848, n7236, new_n1818);
not_4  g01442(new_n1818, new_n1819);
nand_1 g01443(n8028, n3992, new_n1820);
not_4  g01444(new_n1820, new_n1821);
nand_1 g01445(new_n1821, new_n1819, new_n1822);
nor_1  g01446(new_n1822, new_n1817, new_n1823);
nand_1 g01447(new_n1823, new_n1815, new_n1824);
nand_1 g01448(n10848, n6358, new_n1825);
nand_1 g01449(n8384, n1980, new_n1826);
nand_1 g01450(n8028, n5198, new_n1827);
not_4  g01451(new_n1827, new_n1828);
xnor_1 g01452(new_n1828, new_n1826, new_n1829);
xnor_1 g01453(new_n1829, new_n1825, new_n1830);
not_4  g01454(new_n1830, new_n1831);
nand_1 g01455(n7294, n3992, new_n1832);
nand_1 g01456(new_n1811, new_n1810, new_n1833);
not_4  g01457(new_n1833, new_n1834);
nor_1  g01458(new_n1812, new_n1809, new_n1835_1);
nor_1  g01459(new_n1835_1, new_n1834, new_n1836);
xnor_1 g01460(new_n1836, new_n1832, new_n1837);
xnor_1 g01461(new_n1837, new_n1831, new_n1838);
not_4  g01462(new_n1838, new_n1839);
nand_1 g01463(n12704, n7236, new_n1840);
not_4  g01464(new_n1840, new_n1841);
not_4  g01465(new_n1796, new_n1842);
nand_1 g01466(new_n1806, new_n1842, new_n1843);
nand_1 g01467(new_n1813, new_n1807, new_n1844);
nand_1 g01468(new_n1844, new_n1843, new_n1845);
xnor_1 g01469(new_n1845, new_n1841, new_n1846);
xnor_1 g01470(new_n1846, new_n1839, new_n1847_1);
nor_1  g01471(new_n1847_1, new_n1824, new_n1848);
nand_1 g01472(n7236, n5814, new_n1849);
not_4  g01473(new_n1832, new_n1850);
nand_1 g01474(new_n1836, new_n1850, new_n1851);
nand_1 g01475(new_n1837, new_n1830, new_n1852);
nand_1 g01476(new_n1852, new_n1851, new_n1853);
nand_1 g01477(n8384, n7294, new_n1854);
nand_1 g01478(n12704, n3992, new_n1855);
xnor_1 g01479(new_n1855, new_n1854, new_n1856);
xnor_1 g01480(new_n1856, new_n1853, new_n1857);
nand_1 g01481(n6358, n1980, new_n1858);
not_4  g01482(new_n1858, new_n1859);
nand_1 g01483(new_n1827, new_n1826, new_n1860);
nand_1 g01484(new_n1829, new_n1825, new_n1861);
nand_1 g01485(new_n1861, new_n1860, new_n1862);
xnor_1 g01486(new_n1862, new_n1859, new_n1863);
nand_1 g01487(n10848, n5198, new_n1864);
nand_1 g01488(n8028, n1471, new_n1865);
nand_1 g01489(new_n1865, new_n1864, new_n1866);
not_4  g01490(new_n1864, new_n1867);
not_4  g01491(new_n1865, new_n1868);
nand_1 g01492(new_n1868, new_n1867, new_n1869);
nand_1 g01493(new_n1869, new_n1866, new_n1870);
not_4  g01494(new_n1870, new_n1871);
xnor_1 g01495(new_n1871, new_n1863, new_n1872);
xnor_1 g01496(new_n1872, new_n1857, new_n1873);
nor_1  g01497(new_n1845, new_n1841, new_n1874);
nor_1  g01498(new_n1846, new_n1838, new_n1875);
nor_1  g01499(new_n1875, new_n1874, new_n1876);
nand_1 g01500(new_n1876, new_n1873, new_n1877);
not_4  g01501(new_n1877, new_n1878);
nor_1  g01502(new_n1876, new_n1873, new_n1879);
nor_1  g01503(new_n1879, new_n1878, new_n1880);
xnor_1 g01504(new_n1880, new_n1849, new_n1881);
nand_1 g01505(new_n1881, new_n1848, new_n1882);
not_4  g01506(new_n1848, new_n1883);
not_4  g01507(new_n1849, new_n1884);
xnor_1 g01508(new_n1880, new_n1884, new_n1885);
nand_1 g01509(new_n1885, new_n1883, new_n1886);
nand_1 g01510(new_n1886, new_n1882, new_n1887);
not_4  g01511(new_n1887, new_n1888);
nand_1 g01512(n4805, n2802, new_n1889);
nand_1 g01513(n5283, n1564, new_n1890);
not_4  g01514(new_n1890, new_n1891);
nand_1 g01515(n4805, n533, new_n1892);
not_4  g01516(new_n1892, new_n1893);
nand_1 g01517(new_n1893, new_n1891, new_n1894);
nand_1 g01518(new_n1892, new_n1890, new_n1895);
nand_1 g01519(n11478, n1512, new_n1896);
not_4  g01520(new_n1896, new_n1897);
nand_1 g01521(new_n1897, new_n1895, new_n1898);
nand_1 g01522(new_n1898, new_n1894, new_n1899);
xnor_1 g01523(new_n1899, new_n1889, new_n1900);
nand_1 g01524(n1564, n137, new_n1901);
nand_1 g01525(n5283, n1512, new_n1902);
nand_1 g01526(n11478, n533, new_n1903);
not_4  g01527(new_n1903, new_n1904);
xnor_1 g01528(new_n1904, new_n1902, new_n1905);
not_4  g01529(new_n1905, new_n1906_1);
xnor_1 g01530(new_n1906_1, new_n1901, new_n1907);
xnor_1 g01531(new_n1907, new_n1900, new_n1908);
nand_1 g01532(new_n1895, new_n1894, new_n1909);
not_4  g01533(new_n1909, new_n1910);
nand_1 g01534(n4805, n1512, new_n1911);
not_4  g01535(new_n1911, new_n1912);
nand_1 g01536(n11478, n1564, new_n1913);
not_4  g01537(new_n1913, new_n1914);
nand_1 g01538(new_n1914, new_n1912, new_n1915);
nor_1  g01539(new_n1915, new_n1910, new_n1916);
nand_1 g01540(new_n1916, new_n1908, new_n1917);
not_4  g01541(new_n1917, new_n1918);
nand_1 g01542(n6806, n4805, new_n1919);
not_4  g01543(new_n1919, new_n1920);
nand_1 g01544(n11478, n2802, new_n1921);
nand_1 g01545(new_n1903, new_n1902, new_n1922);
nand_1 g01546(new_n1905, new_n1901, new_n1923);
nand_1 g01547(new_n1923, new_n1922, new_n1924);
not_4  g01548(new_n1924, new_n1925);
xnor_1 g01549(new_n1925, new_n1921, new_n1926);
not_4  g01550(new_n1926, new_n1927);
nand_1 g01551(n1512, n137, new_n1928);
not_4  g01552(new_n1928, new_n1929);
nand_1 g01553(n5283, n533, new_n1930);
nand_1 g01554(n6294, n1564, new_n1931);
xnor_1 g01555(new_n1931, new_n1930, new_n1932);
xnor_1 g01556(new_n1932, new_n1929, new_n1933);
xnor_1 g01557(new_n1933, new_n1927, new_n1934);
xnor_1 g01558(new_n1934, new_n1920, new_n1935);
not_4  g01559(new_n1889, new_n1936);
nand_1 g01560(new_n1899, new_n1936, new_n1937);
not_4  g01561(new_n1900, new_n1938);
nor_1  g01562(new_n1907, new_n1938, new_n1939);
not_4  g01563(new_n1939, new_n1940);
nand_1 g01564(new_n1940, new_n1937, new_n1941);
nor_1  g01565(new_n1941, new_n1935, new_n1942);
not_4  g01566(new_n1942, new_n1943);
nand_1 g01567(new_n1941, new_n1935, new_n1944);
nand_1 g01568(new_n1944, new_n1943, new_n1945);
nand_1 g01569(new_n1945, new_n1918, new_n1946);
nand_1 g01570(n5069, n4805, new_n1947);
nand_1 g01571(n533, n137, new_n1948);
nand_1 g01572(n6294, n1512, new_n1949);
nand_1 g01573(n6797, n1564, new_n1950);
not_4  g01574(new_n1950, new_n1951);
xnor_1 g01575(new_n1951, new_n1949, new_n1952);
xnor_1 g01576(new_n1952, new_n1948, new_n1953);
nand_1 g01577(new_n1931, new_n1930, new_n1954);
not_4  g01578(new_n1954, new_n1955);
nor_1  g01579(new_n1932, new_n1929, new_n1956);
nor_1  g01580(new_n1956, new_n1955, new_n1957);
xnor_1 g01581(new_n1957, new_n1953, new_n1958);
nand_1 g01582(n11478, n6806, new_n1959);
nand_1 g01583(n5283, n2802, new_n1960);
not_4  g01584(new_n1960, new_n1961);
xnor_1 g01585(new_n1961, new_n1959, new_n1962);
xnor_1 g01586(new_n1962, new_n1958, new_n1963);
nor_1  g01587(new_n1924, new_n1921, new_n1964);
not_4  g01588(new_n1964, new_n1965);
nand_1 g01589(new_n1933, new_n1926, new_n1966);
nand_1 g01590(new_n1966, new_n1965, new_n1967);
xnor_1 g01591(new_n1967, new_n1963, new_n1968);
nor_1  g01592(new_n1934, new_n1920, new_n1969);
nor_1  g01593(new_n1942, new_n1969, new_n1970);
xnor_1 g01594(new_n1970, new_n1968, new_n1971);
xnor_1 g01595(new_n1971, new_n1947, new_n1972);
xnor_1 g01596(new_n1972, new_n1946, new_n1973);
xnor_1 g01597(new_n1973, new_n1888, new_n1974);
not_4  g01598(new_n1974, new_n1975);
not_4  g01599(new_n1847_1, new_n1976);
xnor_1 g01600(new_n1976, new_n1824, new_n1977);
not_4  g01601(new_n1977, new_n1978);
xnor_1 g01602(new_n1916, new_n1908, new_n1979);
not_4  g01603(new_n1979, new_n1980_1);
xnor_1 g01604(new_n1823, new_n1814, new_n1981);
nor_1  g01605(new_n1981, new_n1980_1, new_n1982);
not_4  g01606(new_n1982, new_n1983);
nand_1 g01607(new_n1913, new_n1911, new_n1984);
nand_1 g01608(new_n1984, new_n1915, new_n1985);
nand_1 g01609(new_n1985, new_n1332, new_n1986);
xnor_1 g01610(new_n1985, new_n1332, new_n1987);
not_4  g01611(new_n1987, new_n1988);
nand_1 g01612(new_n1820, new_n1818, new_n1989);
nand_1 g01613(new_n1989, new_n1822, new_n1990);
nand_1 g01614(new_n1990, new_n1988, new_n1991);
nand_1 g01615(new_n1991, new_n1986, new_n1992);
nand_1 g01616(new_n1897, new_n1328, new_n1993);
nand_1 g01617(new_n1993, new_n1909, new_n1994);
nor_1  g01618(new_n1898, new_n1329, new_n1995);
not_4  g01619(new_n1995, new_n1996);
nand_1 g01620(new_n1996, new_n1994, new_n1997);
nand_1 g01621(new_n1997, new_n1992, new_n1998);
xnor_1 g01622(new_n1997, new_n1992, new_n1999);
not_4  g01623(new_n1999, new_n2000);
nand_1 g01624(new_n1798_1, new_n1330, new_n2001);
nand_1 g01625(new_n2001, new_n1816, new_n2002);
nor_1  g01626(new_n1802, new_n1331, new_n2003);
not_4  g01627(new_n2003, new_n2004);
nand_1 g01628(new_n2004, new_n2002, new_n2005);
nand_1 g01629(new_n2005, new_n2000, new_n2006);
nand_1 g01630(new_n2006, new_n1998, new_n2007);
xnor_1 g01631(new_n1981, new_n1979, new_n2008);
nand_1 g01632(new_n2008, new_n2007, new_n2009);
nand_1 g01633(new_n2009, new_n1983, new_n2010);
nand_1 g01634(new_n2010, new_n1978, new_n2011);
xnor_1 g01635(new_n1945, new_n1918, new_n2012);
xnor_1 g01636(new_n2010, new_n1977, new_n2013);
nand_1 g01637(new_n2013, new_n2012, new_n2014);
nand_1 g01638(new_n2014, new_n2011, new_n2015);
nand_1 g01639(new_n2015, new_n1975, new_n2016);
not_4  g01640(new_n2016, new_n2017);
nor_1  g01641(new_n2015, new_n1975, new_n2018);
nor_1  g01642(new_n2018, new_n2017, new_n2019);
nand_1 g01643(new_n2019, new_n1795, new_n2020);
not_4  g01644(new_n2020, new_n2021);
nor_1  g01645(new_n2019, new_n1795, new_n2022);
nor_1  g01646(new_n2022, new_n2021, new_n2023);
not_4  g01647(new_n1748, new_n2024_1);
xnor_1 g01648(new_n2024_1, new_n1729, new_n2025);
not_4  g01649(new_n2025, new_n2026);
not_4  g01650(new_n2013, new_n2027);
xnor_1 g01651(new_n2027, new_n2012, new_n2028);
nor_1  g01652(new_n2028, new_n2026, new_n2029);
not_4  g01653(new_n2029, new_n2030);
xnor_1 g01654(new_n2028, new_n2025, new_n2031);
xnor_1 g01655(new_n1727, new_n1718, new_n2032);
xnor_1 g01656(new_n2008, new_n2007, new_n2033);
nand_1 g01657(new_n2033, new_n2032, new_n2034);
xnor_1 g01658(new_n2033, new_n2032, new_n2035);
not_4  g01659(new_n2035, new_n2036);
xnor_1 g01660(new_n2005, new_n1999, new_n2037);
nand_1 g01661(new_n1704, new_n1327, new_n2038);
nor_1  g01662(new_n2038, new_n1702, new_n2039);
not_4  g01663(new_n2039, new_n2040);
nand_1 g01664(new_n2038, new_n1721, new_n2041);
nand_1 g01665(new_n2041, new_n2040, new_n2042);
not_4  g01666(new_n2042, new_n2043);
nor_1  g01667(new_n2043, new_n2037, new_n2044);
not_4  g01668(new_n2044, new_n2045);
nand_1 g01669(new_n2043, new_n2037, new_n2046);
nand_1 g01670(new_n2046, new_n2045, new_n2047);
not_4  g01671(new_n2047, new_n2048);
xnor_1 g01672(new_n1990, new_n1987, new_n2049);
not_4  g01673(new_n2049, new_n2050);
nand_1 g01674(new_n1724, new_n1722, new_n2051);
nand_1 g01675(new_n2051, new_n1726, new_n2052);
not_4  g01676(new_n2052, new_n2053);
nand_1 g01677(new_n2053, new_n2050, new_n2054);
not_4  g01678(new_n1327, new_n2055);
nand_1 g01679(new_n1335, new_n2055, new_n2056);
not_4  g01680(new_n2056, new_n2057);
xnor_1 g01681(new_n2052, new_n2050, new_n2058);
nand_1 g01682(new_n2058, new_n2057, new_n2059);
nand_1 g01683(new_n2059, new_n2054, new_n2060);
nand_1 g01684(new_n2060, new_n2048, new_n2061);
nand_1 g01685(new_n2061, new_n2045, new_n2062);
nand_1 g01686(new_n2062, new_n2036, new_n2063);
nand_1 g01687(new_n2063, new_n2034, new_n2064);
nand_1 g01688(new_n2064, new_n2031, new_n2065);
nand_1 g01689(new_n2065, new_n2030, new_n2066);
not_4  g01690(new_n2066, new_n2067);
nand_1 g01691(new_n2067, new_n2023, new_n2068);
nand_1 g01692(new_n2068, new_n2020, new_n2069);
not_4  g01693(new_n2069, new_n2070);
not_4  g01694(new_n1755, new_n2071);
nand_1 g01695(new_n1791, new_n2071, new_n2072);
not_4  g01696(new_n1756, new_n2073);
nand_1 g01697(new_n1764, new_n2073, new_n2074);
nand_1 g01698(new_n1771, new_n2074, new_n2075);
nand_1 g01699(n9400, n4928, new_n2076);
nand_1 g01700(n4141, n2464, new_n2077);
not_4  g01701(new_n2077, new_n2078);
nand_1 g01702(n8236, n6877, new_n2079);
not_4  g01703(new_n2079, new_n2080);
nand_1 g01704(new_n2080, new_n2078, new_n2081);
nand_1 g01705(new_n2079, new_n2077, new_n2082);
nand_1 g01706(new_n2082, new_n2081, new_n2083);
xnor_1 g01707(new_n2083, new_n2076, new_n2084);
xnor_1 g01708(new_n2084, new_n2075, new_n2085);
not_4  g01709(new_n1762, new_n2086);
nand_1 g01710(n11311, n5105, new_n2087_1);
not_4  g01711(new_n2087_1, new_n2088);
nand_1 g01712(new_n2088, new_n2086, new_n2089);
nand_1 g01713(new_n2087_1, new_n1762, new_n2090);
nand_1 g01714(new_n2090, new_n2089, new_n2091);
not_4  g01715(new_n2091, new_n2092);
nand_1 g01716(n7500, n4203, new_n2093);
nand_1 g01717(n4187, n1209, new_n2094);
nand_1 g01718(n12753, n7354, new_n2095);
not_4  g01719(new_n2095, new_n2096_1);
xnor_1 g01720(new_n2096_1, new_n2094, new_n2097);
xnor_1 g01721(new_n2097, new_n2093, new_n2098);
not_4  g01722(new_n2098, new_n2099);
xnor_1 g01723(new_n2099, new_n2092, new_n2100);
xnor_1 g01724(new_n2100, new_n2085, new_n2101);
nand_1 g01725(new_n1788, new_n1774, new_n2102);
xnor_1 g01726(new_n2102, new_n1783, new_n2103);
nand_1 g01727(new_n2103, new_n1789, new_n2104);
xnor_1 g01728(new_n2104, new_n2101, new_n2105);
xnor_1 g01729(new_n2105, new_n2072, new_n2106);
not_4  g01730(new_n1750, new_n2107);
nand_1 g01731(new_n1792, new_n2107, new_n2108);
not_4  g01732(new_n1749, new_n2109);
nand_1 g01733(new_n1793, new_n2109, new_n2110);
nand_1 g01734(new_n2110, new_n2108, new_n2111);
xnor_1 g01735(new_n2111, new_n2106, new_n2112);
nand_1 g01736(new_n1862, new_n1858, new_n2113);
nand_1 g01737(new_n1870, new_n1863, new_n2114);
nand_1 g01738(new_n2114, new_n2113, new_n2115);
nand_1 g01739(n5814, n3992, new_n2116);
nand_1 g01740(n12704, n8384, new_n2117);
nand_1 g01741(n7236, n4903, new_n2118);
not_4  g01742(new_n2118, new_n2119);
xnor_1 g01743(new_n2119, new_n2117, new_n2120);
xnor_1 g01744(new_n2120, new_n2116, new_n2121);
xnor_1 g01745(new_n2121, new_n2115, new_n2122);
not_4  g01746(new_n1869, new_n2123);
nand_1 g01747(n7294, n6358, new_n2124);
not_4  g01748(new_n2124, new_n2125);
nand_1 g01749(new_n2125, new_n2123, new_n2126);
nand_1 g01750(new_n2124, new_n1869, new_n2127);
nand_1 g01751(new_n2127, new_n2126, new_n2128);
not_4  g01752(new_n2128, new_n2129);
nand_1 g01753(n10848, n1471, new_n2130);
nand_1 g01754(n5198, n1980, new_n2131_1);
nand_1 g01755(n8028, n7646, new_n2132);
not_4  g01756(new_n2132, new_n2133);
xnor_1 g01757(new_n2133, new_n2131_1, new_n2134);
xnor_1 g01758(new_n2134, new_n2130, new_n2135);
not_4  g01759(new_n2135, new_n2136);
xnor_1 g01760(new_n2136, new_n2129, new_n2137);
xnor_1 g01761(new_n2137, new_n2122, new_n2138);
not_4  g01762(new_n1856, new_n2139);
nand_1 g01763(new_n2139, new_n1853, new_n2140);
nor_1  g01764(new_n1855, new_n1854, new_n2141);
xnor_1 g01765(new_n2139, new_n1853, new_n2142);
nor_1  g01766(new_n1872, new_n2142, new_n2143);
xnor_1 g01767(new_n2143, new_n2141, new_n2144);
nand_1 g01768(new_n2144, new_n2140, new_n2145);
xnor_1 g01769(new_n2145, new_n2138, new_n2146);
nand_1 g01770(new_n2146, new_n1878, new_n2147);
not_4  g01771(new_n2138, new_n2148);
xnor_1 g01772(new_n2145, new_n2148, new_n2149);
nand_1 g01773(new_n2149, new_n1877, new_n2150);
nand_1 g01774(new_n2150, new_n2147, new_n2151);
nand_1 g01775(new_n1880, new_n1884, new_n2152);
nand_1 g01776(new_n1882, new_n2152, new_n2153);
not_4  g01777(new_n2153, new_n2154);
xnor_1 g01778(new_n2154, new_n2151, new_n2155);
not_4  g01779(new_n1947, new_n2156);
nand_1 g01780(new_n1971, new_n2156, new_n2157);
not_4  g01781(new_n1972, new_n2158);
nor_1  g01782(new_n2158, new_n1946, new_n2159);
not_4  g01783(new_n2159, new_n2160);
nand_1 g01784(new_n2160, new_n2157, new_n2161);
not_4  g01785(new_n1968, new_n2162);
nand_1 g01786(new_n1970, new_n2162, new_n2163);
not_4  g01787(new_n1948, new_n2164);
nand_1 g01788(new_n1952, new_n2164, new_n2165);
nand_1 g01789(new_n1957, new_n1953, new_n2166);
nand_1 g01790(new_n2166, new_n2165, new_n2167);
not_4  g01791(new_n2167, new_n2168);
nand_1 g01792(n11478, n5069, new_n2169);
nand_1 g01793(n6806, n5283, new_n2170);
nand_1 g01794(n12044, n4805, new_n2171);
nand_1 g01795(new_n2171, new_n2170, new_n2172);
not_4  g01796(new_n2170, new_n2173);
not_4  g01797(new_n2171, new_n2174);
nand_1 g01798(new_n2174, new_n2173, new_n2175);
nand_1 g01799(new_n2175, new_n2172, new_n2176);
xnor_1 g01800(new_n2176, new_n2169, new_n2177);
xnor_1 g01801(new_n2177, new_n2168, new_n2178);
not_4  g01802(new_n1949, new_n2179);
nand_1 g01803(new_n1951, new_n2179, new_n2180);
nand_1 g01804(n2802, n137, new_n2181);
nand_1 g01805(new_n2181, new_n2180, new_n2182);
not_4  g01806(new_n2180, new_n2183);
not_4  g01807(new_n2181, new_n2184);
nand_1 g01808(new_n2184, new_n2183, new_n2185);
nand_1 g01809(new_n2185, new_n2182, new_n2186);
nand_1 g01810(n6797, n1512, new_n2187);
nand_1 g01811(n6294, n533, new_n2188);
nand_1 g01812(n3146, n1564, new_n2189);
not_4  g01813(new_n2189, new_n2190);
xnor_1 g01814(new_n2190, new_n2188, new_n2191);
not_4  g01815(new_n2191, new_n2192);
xnor_1 g01816(new_n2192, new_n2187, new_n2193);
nand_1 g01817(new_n2193, new_n2186, new_n2194);
not_4  g01818(new_n2186, new_n2195);
not_4  g01819(new_n2193, new_n2196);
nand_1 g01820(new_n2196, new_n2195, new_n2197);
nand_1 g01821(new_n2197, new_n2194, new_n2198);
xnor_1 g01822(new_n2198, new_n2178, new_n2199);
not_4  g01823(new_n1958, new_n2200);
nand_1 g01824(new_n1962, new_n2200, new_n2201);
nor_1  g01825(new_n1960, new_n1959, new_n2202);
nand_1 g01826(new_n1967, new_n1963, new_n2203);
not_4  g01827(new_n2203, new_n2204);
xnor_1 g01828(new_n2204, new_n2202, new_n2205);
nand_1 g01829(new_n2205, new_n2201, new_n2206);
xnor_1 g01830(new_n2206, new_n2199, new_n2207);
xnor_1 g01831(new_n2207, new_n2163, new_n2208);
xnor_1 g01832(new_n2208, new_n2161, new_n2209);
nand_1 g01833(new_n2209, new_n2155, new_n2210);
xnor_1 g01834(new_n2153, new_n2151, new_n2211);
not_4  g01835(new_n2209, new_n2212);
nand_1 g01836(new_n2212, new_n2211, new_n2213);
nand_1 g01837(new_n2213, new_n2210, new_n2214);
nor_1  g01838(new_n1973, new_n1888, new_n2215);
nor_1  g01839(new_n2017, new_n2215, new_n2216);
nor_1  g01840(new_n2216, new_n2214, new_n2217);
nor_1  g01841(new_n2212, new_n2211, new_n2218);
nor_1  g01842(new_n2209, new_n2155, new_n2219);
nor_1  g01843(new_n2219, new_n2218, new_n2220);
not_4  g01844(new_n2216, new_n2221);
nor_1  g01845(new_n2221, new_n2220, new_n2222);
nor_1  g01846(new_n2222, new_n2217, new_n2223);
nand_1 g01847(new_n2223, new_n2112, new_n2224);
not_4  g01848(new_n2112, new_n2225);
nand_1 g01849(new_n2221, new_n2220, new_n2226_1);
nand_1 g01850(new_n2216, new_n2214, new_n2227);
nand_1 g01851(new_n2227, new_n2226_1, new_n2228);
nand_1 g01852(new_n2228, new_n2225, new_n2229);
nand_1 g01853(new_n2229, new_n2224, new_n2230);
nor_1  g01854(new_n2230, new_n2070, new_n2231);
nor_1  g01855(new_n2228, new_n2225, new_n2232);
nor_1  g01856(new_n2223, new_n2112, new_n2233);
nor_1  g01857(new_n2233, new_n2232, new_n2234);
nor_1  g01858(new_n2234, new_n2069, new_n2235);
nor_1  g01859(new_n2235, new_n2231, new_n2236);
nor_1  g01860(new_n2236, new_n1695, new_n2237);
not_4  g01861(new_n1695, new_n2238);
nand_1 g01862(new_n2234, new_n2069, new_n2239);
nand_1 g01863(new_n2230, new_n2070, new_n2240);
nand_1 g01864(new_n2240, new_n2239, new_n2241);
nand_1 g01865(new_n2241, new_n2238, new_n2242);
nand_1 g01866(new_n2236, new_n1695, new_n2243);
nand_1 g01867(new_n2243, new_n2242, new_n2244);
xnor_1 g01868(new_n1692, new_n1690, new_n2245);
nor_1  g01869(new_n2067, new_n2023, new_n2246);
not_4  g01870(new_n2246, new_n2247);
nand_1 g01871(new_n2247, new_n2068, new_n2248);
nand_1 g01872(new_n2248, new_n2245, new_n2249);
xnor_1 g01873(new_n1689, new_n1687, new_n2250);
xnor_1 g01874(new_n2064, new_n2031, new_n2251);
nand_1 g01875(new_n2251, new_n2250, new_n2252);
xnor_1 g01876(new_n2251, new_n2250, new_n2253_1);
xnor_1 g01877(new_n1685, new_n1677, new_n2254);
not_4  g01878(new_n2254, new_n2255);
xnor_1 g01879(new_n2062, new_n2035, new_n2256);
nor_1  g01880(new_n2256, new_n2255, new_n2257);
not_4  g01881(new_n2060, new_n2258);
nand_1 g01882(new_n2258, new_n2047, new_n2259);
nand_1 g01883(new_n2259, new_n2061, new_n2260);
nand_1 g01884(new_n1588, new_n1326, new_n2261);
nand_1 g01885(new_n2261, new_n1678, new_n2262);
not_4  g01886(new_n1326, new_n2263);
nor_1  g01887(new_n1592, new_n2263, new_n2264);
not_4  g01888(new_n2264, new_n2265);
nand_1 g01889(new_n2265, new_n2262, new_n2266);
nand_1 g01890(new_n2266, new_n2260, new_n2267);
xnor_1 g01891(new_n2266, new_n2260, new_n2268);
nand_1 g01892(new_n1336, new_n2263, new_n2269);
nand_1 g01893(new_n1682, new_n1680, new_n2270);
nand_1 g01894(new_n2270, new_n1684, new_n2271);
nand_1 g01895(new_n2271, new_n2269, new_n2272);
xnor_1 g01896(new_n2058, new_n2056, new_n2273);
xnor_1 g01897(new_n2271, new_n2269, new_n2274);
nor_1  g01898(new_n2274, new_n2273, new_n2275);
not_4  g01899(new_n2275, new_n2276);
nand_1 g01900(new_n2276, new_n2272, new_n2277);
not_4  g01901(new_n2277, new_n2278_1);
nor_1  g01902(new_n2278_1, new_n2268, new_n2279);
not_4  g01903(new_n2279, new_n2280);
nand_1 g01904(new_n2280, new_n2267, new_n2281);
not_4  g01905(new_n2281, new_n2282);
xnor_1 g01906(new_n2256, new_n2255, new_n2283);
nor_1  g01907(new_n2283, new_n2282, new_n2284);
nor_1  g01908(new_n2284, new_n2257, new_n2285);
nor_1  g01909(new_n2285, new_n2253_1, new_n2286);
not_4  g01910(new_n2286, new_n2287);
nand_1 g01911(new_n2287, new_n2252, new_n2288);
not_4  g01912(new_n2288, new_n2289);
not_4  g01913(new_n2249, new_n2290);
nor_1  g01914(new_n2248, new_n2245, new_n2291);
nor_1  g01915(new_n2291, new_n2290, new_n2292);
nand_1 g01916(new_n2292, new_n2289, new_n2293);
nand_1 g01917(new_n2293, new_n2249, new_n2294);
not_4  g01918(new_n2294, new_n2295);
nor_1  g01919(new_n2295, new_n2244, new_n2296);
nor_1  g01920(new_n2296, new_n2237, new_n2297);
nand_1 g01921(new_n2239, new_n2224, new_n2298);
nand_1 g01922(new_n2226_1, new_n2210, new_n2299);
not_4  g01923(new_n1642, new_n2300);
nand_1 g01924(new_n1671, new_n2300, new_n2301_1);
nand_1 g01925(new_n1694, new_n1672, new_n2302);
nand_1 g01926(new_n2302, new_n2301_1, new_n2303);
not_4  g01927(new_n2147, new_n2304);
nor_1  g01928(new_n2154, new_n2151, new_n2305);
nor_1  g01929(new_n2305, new_n2304, new_n2306);
xnor_1 g01930(new_n2306, new_n2303, new_n2307);
nand_1 g01931(new_n2143, new_n2141, new_n2308);
nand_1 g01932(new_n2145, new_n2148, new_n2309);
nand_1 g01933(new_n2309, new_n2308, new_n2310);
nand_1 g01934(new_n2197, new_n2185, new_n2311);
nand_1 g01935(n7862, n615, new_n2312);
nand_1 g01936(n4903, n3992, new_n2313);
nand_1 g01937(n6806, n137, new_n2314);
xnor_1 g01938(new_n2314, new_n2313, new_n2315);
xnor_1 g01939(new_n2315, new_n2312, new_n2316_1);
xnor_1 g01940(new_n2316_1, new_n2311, new_n2317);
nand_1 g01941(n6797, n533, new_n2318);
nand_1 g01942(n8384, n5814, new_n2319);
xnor_1 g01943(new_n2319, new_n2318, new_n2320);
nand_1 g01944(n12044, n11478, new_n2321);
nand_1 g01945(n7294, n5198, new_n2322);
xnor_1 g01946(new_n2322, new_n2321, new_n2323);
xnor_1 g01947(new_n2323, new_n2320, new_n2324);
not_4  g01948(new_n2169, new_n2325);
nand_1 g01949(new_n2172, new_n2325, new_n2326);
nand_1 g01950(new_n2326, new_n2175, new_n2327);
xnor_1 g01951(new_n2327, new_n2324, new_n2328);
nand_1 g01952(n10174, n7354, new_n2329);
nand_1 g01953(n4928, n2464, new_n2330);
nand_1 g01954(n11311, n4141, new_n2331);
xnor_1 g01955(new_n2331, new_n2330, new_n2332);
nand_1 g01956(n4005, n3172, new_n2333);
nand_1 g01957(n7236, n1906, new_n2334);
xnor_1 g01958(new_n2334, new_n2333, new_n2335);
xnor_1 g01959(new_n2335, new_n2332, new_n2336);
xnor_1 g01960(new_n2336, new_n2329, new_n2337);
xnor_1 g01961(new_n2337, new_n2328, new_n2338);
xnor_1 g01962(new_n2338, new_n2317, new_n2339);
xnor_1 g01963(new_n2339, new_n2310, new_n2340);
not_4  g01964(new_n2121, new_n2341);
nand_1 g01965(new_n2341, new_n2115, new_n2342);
not_4  g01966(new_n2137, new_n2343);
nand_1 g01967(new_n2343, new_n2122, new_n2344);
nand_1 g01968(new_n2344, new_n2342, new_n2345);
nand_1 g01969(n9080, n2509, new_n2346);
nand_1 g01970(new_n1651, new_n1650, new_n2347_1);
nand_1 g01971(new_n1653, new_n1648, new_n2348);
nand_1 g01972(new_n2348, new_n2347_1, new_n2349);
nand_1 g01973(n5240, n2508, new_n2350);
nand_1 g01974(n11757, n2585, new_n2351);
nand_1 g01975(n12706, n1333, new_n2352);
xnor_1 g01976(new_n2352, new_n2351, new_n2353);
xnor_1 g01977(new_n2353, new_n2350, new_n2354);
xnor_1 g01978(new_n2354, new_n2349, new_n2355);
xnor_1 g01979(new_n2355, new_n2346, new_n2356);
xnor_1 g01980(new_n2356, new_n2345, new_n2357);
xnor_1 g01981(new_n2357, new_n2340, new_n2358);
not_4  g01982(new_n1783, new_n2359);
not_4  g01983(new_n2102, new_n2360);
nand_1 g01984(new_n2360, new_n2359, new_n2361);
not_4  g01985(new_n2101, new_n2362);
nand_1 g01986(new_n2104, new_n2362, new_n2363);
nand_1 g01987(new_n2363, new_n2361, new_n2364);
nor_1  g01988(new_n1643, new_n1634, new_n2365);
not_4  g01989(new_n1645, new_n2366);
nor_1  g01990(new_n1670, new_n2366, new_n2367);
nor_1  g01991(new_n2367, new_n2365, new_n2368);
xnor_1 g01992(new_n2368, new_n2364, new_n2369);
not_4  g01993(new_n2075, new_n2370);
nand_1 g01994(new_n2084, new_n2370, new_n2371);
not_4  g01995(new_n2100, new_n2372);
nand_1 g01996(new_n2372, new_n2085, new_n2373);
nand_1 g01997(new_n2373, new_n2371, new_n2374);
nand_1 g01998(n12704, n6358, new_n2375);
nand_1 g01999(n3146, n1512, new_n2376);
xnor_1 g02000(new_n2376, new_n2375, new_n2377);
nand_1 g02001(n5105, n4187, new_n2378);
nand_1 g02002(n6294, n2802, new_n2379);
xnor_1 g02003(new_n2379, new_n2378, new_n2380);
nand_1 g02004(n9400, n8236, new_n2381);
nand_1 g02005(n1980, n1471, new_n2382);
not_4  g02006(new_n2382, new_n2383_1);
xnor_1 g02007(new_n2383_1, new_n2381, new_n2384);
xnor_1 g02008(new_n2384, new_n2380, new_n2385);
xnor_1 g02009(new_n2385, new_n2377, new_n2386);
nand_1 g02010(n12720, n11821, new_n2387);
nand_1 g02011(n4938, n1564, new_n2388);
nand_1 g02012(n5694, n4805, new_n2389);
xnor_1 g02013(new_n2389, new_n2388, new_n2390);
xnor_1 g02014(new_n2390, new_n2387, new_n2391);
xnor_1 g02015(new_n2391, new_n2386, new_n2392);
nand_1 g02016(new_n2118, new_n2117, new_n2393_1);
nand_1 g02017(new_n2120, new_n2116, new_n2394);
nand_1 g02018(new_n2394, new_n2393_1, new_n2395);
nor_1  g02019(new_n1646, new_n1613, new_n2396);
nor_1  g02020(new_n1654, new_n1647, new_n2397);
nor_1  g02021(new_n2397, new_n2396, new_n2398);
xnor_1 g02022(new_n2398, new_n2395, new_n2399);
xnor_1 g02023(new_n2399, new_n2392, new_n2400);
xnor_1 g02024(new_n2400, new_n2374, new_n2401);
nand_1 g02025(new_n2204, new_n2202, new_n2402);
not_4  g02026(new_n2199, new_n2403);
nand_1 g02027(new_n2206, new_n2403, new_n2404);
nand_1 g02028(new_n2404, new_n2402, new_n2405);
nand_1 g02029(new_n2177, new_n2168, new_n2406);
not_4  g02030(new_n2178, new_n2407);
nand_1 g02031(new_n2198, new_n2407, new_n2408);
nand_1 g02032(new_n2408, new_n2406, new_n2409);
nand_1 g02033(new_n2135, new_n2129, new_n2410);
nand_1 g02034(new_n2410, new_n2126, new_n2411);
nand_1 g02035(n4203, n1209, new_n2412);
nand_1 g02036(n6826, n6038, new_n2413);
nand_1 g02037(n5283, n5069, new_n2414);
xnor_1 g02038(new_n2414, new_n2413, new_n2415);
xnor_1 g02039(new_n2415, new_n2412, new_n2416);
xnor_1 g02040(new_n2416, new_n2411, new_n2417);
nand_1 g02041(new_n2189, new_n2188, new_n2418);
nand_1 g02042(new_n2191, new_n2187, new_n2419);
nand_1 g02043(new_n2419, new_n2418, new_n2420);
nand_1 g02044(new_n2132, new_n2131_1, new_n2421);
nand_1 g02045(new_n2134, new_n2130, new_n2422);
nand_1 g02046(new_n2422, new_n2421, new_n2423);
not_4  g02047(new_n2076, new_n2424);
nand_1 g02048(new_n2082, new_n2424, new_n2425_1);
nand_1 g02049(new_n2425_1, new_n2081, new_n2426);
xnor_1 g02050(new_n2426, new_n2423, new_n2427);
xnor_1 g02051(new_n2427, new_n2420, new_n2428);
xnor_1 g02052(new_n2428, new_n2417, new_n2429);
xnor_1 g02053(new_n2429, new_n2409, new_n2430);
xnor_1 g02054(new_n2430, new_n2405, new_n2431_1);
xnor_1 g02055(new_n2431_1, new_n2401, new_n2432);
xnor_1 g02056(new_n2432, new_n2369, new_n2433_1);
xnor_1 g02057(new_n2433_1, new_n2358, new_n2434_1);
xnor_1 g02058(new_n2434_1, new_n2307, new_n2435);
xnor_1 g02059(new_n2435, new_n2299, new_n2436);
nand_1 g02060(new_n2098, new_n2092, new_n2437);
nand_1 g02061(new_n2437, new_n2089, new_n2438);
nand_1 g02062(n6877, n783, new_n2439);
nand_1 g02063(n8028, n4722, new_n2440);
xnor_1 g02064(new_n2440, new_n2439, new_n2441);
xnor_1 g02065(new_n2441, new_n2438, new_n2442);
not_4  g02066(new_n2072, new_n2443);
nand_1 g02067(new_n2105, new_n2443, new_n2444);
nand_1 g02068(new_n2111, new_n2106, new_n2445);
nand_1 g02069(new_n2445, new_n2444, new_n2446);
nand_1 g02070(n10848, n7646, new_n2447);
xnor_1 g02071(new_n2447, new_n2446, new_n2448);
xnor_1 g02072(new_n2448, new_n2442, new_n2449);
not_4  g02073(new_n2163, new_n2450);
nand_1 g02074(new_n2207, new_n2450, new_n2451);
nand_1 g02075(new_n2208, new_n2161, new_n2452);
nand_1 g02076(new_n2452, new_n2451, new_n2453);
not_4  g02077(new_n1659, new_n2454);
nand_1 g02078(new_n1668, new_n2454, new_n2455);
nand_1 g02079(new_n1669, new_n1655, new_n2456);
nand_1 g02080(new_n2456, new_n2455, new_n2457);
nand_1 g02081(new_n2095, new_n2094, new_n2458);
nand_1 g02082(new_n2097, new_n2093, new_n2459);
nand_1 g02083(new_n2459, new_n2458, new_n2460);
nand_1 g02084(n12753, n7500, new_n2461);
not_4  g02085(new_n1660, new_n2462);
nand_1 g02086(new_n1663, new_n2462, new_n2463);
nand_1 g02087(new_n2463, new_n1666, new_n2464_1);
xnor_1 g02088(new_n2464_1, new_n2461, new_n2465);
xnor_1 g02089(new_n2465, new_n2460, new_n2466);
xnor_1 g02090(new_n2466, new_n2457, new_n2467);
xnor_1 g02091(new_n2467, new_n2453, new_n2468);
xnor_1 g02092(new_n2468, new_n2449, new_n2469);
xnor_1 g02093(new_n2469, new_n2436, new_n2470);
xnor_1 g02094(new_n2470, new_n2298, new_n2471);
nand_1 g02095(new_n2471, new_n2297, new_n2472);
nor_1  g02096(new_n2241, new_n2238, new_n2473);
nor_1  g02097(new_n2473, new_n2237, new_n2474);
nand_1 g02098(new_n2294, new_n2474, new_n2475);
nand_1 g02099(new_n2475, new_n2242, new_n2476);
not_4  g02100(new_n2471, new_n2477);
nand_1 g02101(new_n2477, new_n2476, new_n2478);
nand_1 g02102(new_n2478, new_n2472, n671);
nand_1 g02103(n11917, n4312, new_n2480);
nand_1 g02104(n12705, n4921, new_n2481);
nand_1 g02105(n12025, n9956, new_n2482);
nand_1 g02106(new_n2482, new_n2481, new_n2483);
not_4  g02107(new_n2481, new_n2484);
not_4  g02108(new_n2482, new_n2485);
nand_1 g02109(new_n2485, new_n2484, new_n2486);
nand_1 g02110(new_n2486, new_n2483, new_n2487);
xnor_1 g02111(new_n2487, new_n2480, new_n2488);
nand_1 g02112(n12705, n9956, new_n2489);
nand_1 g02113(n11917, n1097, new_n2490);
nand_1 g02114(new_n2490, new_n2489, new_n2491);
not_4  g02115(new_n2489, new_n2492);
not_4  g02116(new_n2490, new_n2493);
nand_1 g02117(new_n2493, new_n2492, new_n2494);
nand_1 g02118(n4921, n4312, new_n2495);
nand_1 g02119(new_n2495, new_n2494, new_n2496);
nand_1 g02120(new_n2496, new_n2491, new_n2497);
xnor_1 g02121(new_n2497, new_n2488, new_n2498_1);
not_4  g02122(new_n2498_1, new_n2499);
nand_1 g02123(n5964, n2577, new_n2500);
not_4  g02124(new_n2500, new_n2501);
nand_1 g02125(n3842, n1097, new_n2502);
not_4  g02126(new_n2502, new_n2503);
nand_1 g02127(new_n2503, new_n2501, new_n2504);
nand_1 g02128(new_n2502, new_n2500, new_n2505);
nand_1 g02129(new_n2505, new_n2504, new_n2506);
xnor_1 g02130(new_n2506, new_n2499, new_n2507_1);
not_4  g02131(new_n2507_1, new_n2508_1);
nand_1 g02132(n5964, n3842, new_n2509_1);
nand_1 g02133(n9956, n4312, new_n2510);
nand_1 g02134(n11917, n5964, new_n2511);
nand_1 g02135(new_n2511, new_n2510, new_n2512_1);
nor_1  g02136(new_n2511, new_n2510, new_n2513);
not_4  g02137(new_n2513, new_n2514);
nand_1 g02138(n4921, n1097, new_n2515_1);
nand_1 g02139(new_n2515_1, new_n2514, new_n2516);
nand_1 g02140(new_n2516, new_n2512_1, new_n2517);
nor_1  g02141(new_n2517, new_n2509_1, new_n2518);
xnor_1 g02142(new_n2517, new_n2509_1, new_n2519);
nand_1 g02143(new_n2494, new_n2491, new_n2520);
xnor_1 g02144(new_n2520, new_n2495, new_n2521);
nor_1  g02145(new_n2521, new_n2519, new_n2522_1);
nor_1  g02146(new_n2522_1, new_n2518, new_n2523);
nor_1  g02147(new_n2523, new_n2508_1, new_n2524);
not_4  g02148(new_n2524, new_n2525);
nand_1 g02149(new_n2523, new_n2508_1, new_n2526);
nand_1 g02150(new_n2526, new_n2525, new_n2527);
not_4  g02151(new_n2527, new_n2528);
nand_1 g02152(n5305, n2577, new_n2529);
xnor_1 g02153(new_n2521, new_n2519, new_n2530_1);
nand_1 g02154(new_n2530_1, new_n2529, new_n2531);
xnor_1 g02155(new_n2530_1, new_n2529, new_n2532);
nand_1 g02156(n5305, n3842, new_n2533);
not_4  g02157(new_n2533, new_n2534);
nand_1 g02158(n9956, n1097, new_n2535);
not_4  g02159(new_n2535, new_n2536);
nand_1 g02160(n11917, n5305, new_n2537);
not_4  g02161(new_n2537, new_n2538);
nand_1 g02162(new_n2538, new_n2536, new_n2539);
nand_1 g02163(new_n2537, new_n2535, new_n2540);
nand_1 g02164(n5964, n4921, new_n2541);
not_4  g02165(new_n2541, new_n2542);
nand_1 g02166(new_n2542, new_n2540, new_n2543);
nand_1 g02167(new_n2543, new_n2539, new_n2544);
nand_1 g02168(new_n2544, new_n2534, new_n2545);
xnor_1 g02169(new_n2544, new_n2533, new_n2546);
not_4  g02170(new_n2546, new_n2547);
nand_1 g02171(new_n2514, new_n2512_1, new_n2548);
xnor_1 g02172(new_n2548, new_n2515_1, new_n2549);
nor_1  g02173(new_n2549, new_n2547, new_n2550);
not_4  g02174(new_n2550, new_n2551_1);
nand_1 g02175(new_n2551_1, new_n2545, new_n2552);
nor_1  g02176(new_n2552, new_n2532, new_n2553);
not_4  g02177(new_n2553, new_n2554);
nand_1 g02178(new_n2554, new_n2531, new_n2555);
not_4  g02179(new_n2555, new_n2556);
nand_1 g02180(new_n2556, new_n2528, new_n2557);
not_4  g02181(new_n2557, new_n2558_1);
nand_1 g02182(new_n2487, new_n2480, new_n2559);
not_4  g02183(new_n2488, new_n2560);
nand_1 g02184(new_n2497, new_n2560, new_n2561);
nand_1 g02185(new_n2561, new_n2559, new_n2562);
nand_1 g02186(n9637, n5964, new_n2563);
nand_1 g02187(n2577, n1097, new_n2564_1);
nand_1 g02188(n5305, n1835, new_n2565);
not_4  g02189(new_n2565, new_n2566);
xnor_1 g02190(new_n2566, new_n2564_1, new_n2567);
xnor_1 g02191(new_n2567, new_n2563, new_n2568);
xnor_1 g02192(new_n2568, new_n2562, new_n2569);
nand_1 g02193(n4312, n3842, new_n2570);
xnor_1 g02194(new_n2570, new_n2486, new_n2571);
nand_1 g02195(n12025, n4921, new_n2572);
not_4  g02196(new_n2572, new_n2573);
nand_1 g02197(n12705, n11917, new_n2574);
nand_1 g02198(n11257, n9956, new_n2575);
not_4  g02199(new_n2575, new_n2576);
xnor_1 g02200(new_n2576, new_n2574, new_n2577_1);
xnor_1 g02201(new_n2577_1, new_n2573, new_n2578);
xnor_1 g02202(new_n2578, new_n2571, new_n2579);
xnor_1 g02203(new_n2579, new_n2569, new_n2580);
not_4  g02204(new_n2506, new_n2581_1);
nand_1 g02205(new_n2581_1, new_n2499, new_n2582);
xnor_1 g02206(new_n2524, new_n2504, new_n2583);
not_4  g02207(new_n2583, new_n2584);
nand_1 g02208(new_n2584, new_n2582, new_n2585_1);
xnor_1 g02209(new_n2585_1, new_n2580, new_n2586);
not_4  g02210(new_n2586, new_n2587);
nand_1 g02211(new_n2587, new_n2558_1, new_n2588);
nand_1 g02212(new_n2586, new_n2557, new_n2589);
nand_1 g02213(new_n2589, new_n2588, new_n2590);
nand_1 g02214(n9637, n5305, new_n2591);
not_4  g02215(new_n2591, new_n2592);
xnor_1 g02216(new_n2555, new_n2528, new_n2593);
nand_1 g02217(new_n2593, new_n2592, new_n2594);
xnor_1 g02218(new_n2549, new_n2546, new_n2595);
nand_1 g02219(new_n2540, new_n2539, new_n2596);
not_4  g02220(new_n2596, new_n2597);
nand_1 g02221(n9956, n5964, new_n2598);
not_4  g02222(new_n2598, new_n2599);
nand_1 g02223(n5305, n4921, new_n2600);
not_4  g02224(new_n2600, new_n2601);
nand_1 g02225(new_n2601, new_n2599, new_n2602);
nor_1  g02226(new_n2602, new_n2597, new_n2603);
nand_1 g02227(new_n2603, new_n2595, new_n2604);
not_4  g02228(new_n2604, new_n2605);
nand_1 g02229(new_n2552, new_n2532, new_n2606);
nand_1 g02230(new_n2606, new_n2554, new_n2607);
nand_1 g02231(new_n2607, new_n2605, new_n2608);
not_4  g02232(new_n2608, new_n2609);
xnor_1 g02233(new_n2593, new_n2591, new_n2610);
nand_1 g02234(new_n2610, new_n2609, new_n2611);
nand_1 g02235(new_n2611, new_n2594, new_n2612);
xnor_1 g02236(new_n2612, new_n2590, new_n2613);
nand_1 g02237(n8759, n8065, new_n2614);
not_4  g02238(new_n2614, new_n2615);
nand_1 g02239(n7436, n6126, new_n2616);
not_4  g02240(new_n2616, new_n2617);
nand_1 g02241(n9241, n3719, new_n2618);
nand_1 g02242(n8276, n3602, new_n2619);
not_4  g02243(new_n2619, new_n2620);
xnor_1 g02244(new_n2620, new_n2618, new_n2621);
xnor_1 g02245(new_n2621, new_n2617, new_n2622);
nand_1 g02246(n8276, n3719, new_n2623);
nand_1 g02247(n12299, n6126, new_n2624_1);
nand_1 g02248(new_n2624_1, new_n2623, new_n2625);
not_4  g02249(new_n2623, new_n2626);
not_4  g02250(new_n2624_1, new_n2627);
nand_1 g02251(new_n2627, new_n2626, new_n2628);
nand_1 g02252(n7436, n3602, new_n2629);
nand_1 g02253(new_n2629, new_n2628, new_n2630);
nand_1 g02254(new_n2630, new_n2625, new_n2631);
nor_1  g02255(new_n2631, new_n2622, new_n2632);
not_4  g02256(new_n2632, new_n2633);
nand_1 g02257(new_n2631, new_n2622, new_n2634);
nand_1 g02258(new_n2634, new_n2633, new_n2635);
nand_1 g02259(n10439, n6776, new_n2636);
nand_1 g02260(n12299, n8595, new_n2637);
not_4  g02261(new_n2637, new_n2638);
xnor_1 g02262(new_n2638, new_n2636, new_n2639);
xnor_1 g02263(new_n2639, new_n2635, new_n2640);
nand_1 g02264(n8595, n6776, new_n2641);
nand_1 g02265(n7436, n3719, new_n2642);
nand_1 g02266(n6776, n6126, new_n2643);
nand_1 g02267(new_n2643, new_n2642, new_n2644);
not_4  g02268(new_n2642, new_n2645);
not_4  g02269(new_n2643, new_n2646);
nand_1 g02270(new_n2646, new_n2645, new_n2647);
nand_1 g02271(n12299, n3602, new_n2648);
nand_1 g02272(new_n2648, new_n2647, new_n2649);
nand_1 g02273(new_n2649, new_n2644, new_n2650);
nor_1  g02274(new_n2650, new_n2641, new_n2651);
not_4  g02275(new_n2650, new_n2652);
xnor_1 g02276(new_n2652, new_n2641, new_n2653);
not_4  g02277(new_n2653, new_n2654);
nand_1 g02278(new_n2628, new_n2625, new_n2655);
xnor_1 g02279(new_n2655, new_n2629, new_n2656);
nor_1  g02280(new_n2656, new_n2654, new_n2657);
nor_1  g02281(new_n2657, new_n2651, new_n2658);
not_4  g02282(new_n2658, new_n2659);
xnor_1 g02283(new_n2659, new_n2640, new_n2660);
nand_1 g02284(n10439, n8759, new_n2661);
not_4  g02285(new_n2661, new_n2662);
xnor_1 g02286(new_n2656, new_n2653, new_n2663);
nor_1  g02287(new_n2663, new_n2662, new_n2664);
xnor_1 g02288(new_n2663, new_n2662, new_n2665);
nand_1 g02289(n8759, n8595, new_n2666);
not_4  g02290(new_n2666, new_n2667);
nand_1 g02291(n12299, n3719, new_n2668);
not_4  g02292(new_n2668, new_n2669);
nand_1 g02293(n8759, n6126, new_n2670);
not_4  g02294(new_n2670, new_n2671);
nand_1 g02295(new_n2671, new_n2669, new_n2672);
nand_1 g02296(new_n2670, new_n2668, new_n2673);
nand_1 g02297(n6776, n3602, new_n2674);
not_4  g02298(new_n2674, new_n2675);
nand_1 g02299(new_n2675, new_n2673, new_n2676);
nand_1 g02300(new_n2676, new_n2672, new_n2677);
nand_1 g02301(new_n2677, new_n2667, new_n2678);
xnor_1 g02302(new_n2677, new_n2666, new_n2679_1);
not_4  g02303(new_n2679_1, new_n2680);
nand_1 g02304(new_n2647, new_n2644, new_n2681);
xnor_1 g02305(new_n2681, new_n2648, new_n2682);
nor_1  g02306(new_n2682, new_n2680, new_n2683);
not_4  g02307(new_n2683, new_n2684);
nand_1 g02308(new_n2684, new_n2678, new_n2685);
nor_1  g02309(new_n2685, new_n2665, new_n2686);
nor_1  g02310(new_n2686, new_n2664, new_n2687);
xnor_1 g02311(new_n2687, new_n2660, new_n2688);
nand_1 g02312(new_n2688, new_n2615, new_n2689);
xnor_1 g02313(new_n2682, new_n2679_1, new_n2690);
nand_1 g02314(new_n2673, new_n2672, new_n2691);
not_4  g02315(new_n2691, new_n2692);
nand_1 g02316(n6776, n3719, new_n2693);
not_4  g02317(new_n2693, new_n2694);
nand_1 g02318(n8759, n3602, new_n2695);
not_4  g02319(new_n2695, new_n2696);
nand_1 g02320(new_n2696, new_n2694, new_n2697);
nor_1  g02321(new_n2697, new_n2692, new_n2698);
nand_1 g02322(new_n2698, new_n2690, new_n2699);
not_4  g02323(new_n2699, new_n2700);
xnor_1 g02324(new_n2685, new_n2665, new_n2701);
nand_1 g02325(new_n2701, new_n2700, new_n2702);
not_4  g02326(new_n2702, new_n2703);
xnor_1 g02327(new_n2688, new_n2614, new_n2704);
nand_1 g02328(new_n2704, new_n2703, new_n2705);
nand_1 g02329(new_n2705, new_n2689, new_n2706);
not_4  g02330(new_n2660, new_n2707);
nand_1 g02331(new_n2687, new_n2707, new_n2708_1);
nand_1 g02332(new_n2621, new_n2617, new_n2709);
nand_1 g02333(new_n2633, new_n2709, new_n2710);
nand_1 g02334(n8065, n6776, new_n2711);
not_4  g02335(new_n2711, new_n2712);
nand_1 g02336(n12299, n10439, new_n2713);
nand_1 g02337(n10391, n8759, new_n2714);
not_4  g02338(new_n2714, new_n2715);
xnor_1 g02339(new_n2715, new_n2713, new_n2716);
xnor_1 g02340(new_n2716, new_n2712, new_n2717);
xnor_1 g02341(new_n2717, new_n2710, new_n2718);
not_4  g02342(new_n2618, new_n2719);
nand_1 g02343(new_n2620, new_n2719, new_n2720);
not_4  g02344(new_n2720, new_n2721);
nand_1 g02345(n8595, n7436, new_n2722);
not_4  g02346(new_n2722, new_n2723);
nand_1 g02347(new_n2723, new_n2721, new_n2724);
nand_1 g02348(new_n2722, new_n2720, new_n2725);
nand_1 g02349(new_n2725, new_n2724, new_n2726);
nand_1 g02350(n9241, n3602, new_n2727);
nand_1 g02351(n8276, n6126, new_n2728);
nand_1 g02352(n10510, n3719, new_n2729);
nand_1 g02353(new_n2729, new_n2728, new_n2730);
not_4  g02354(new_n2728, new_n2731);
not_4  g02355(new_n2729, new_n2732);
nand_1 g02356(new_n2732, new_n2731, new_n2733);
nand_1 g02357(new_n2733, new_n2730, new_n2734);
xnor_1 g02358(new_n2734, new_n2727, new_n2735);
not_4  g02359(new_n2735, new_n2736);
xnor_1 g02360(new_n2736, new_n2726, new_n2737);
xnor_1 g02361(new_n2737, new_n2718, new_n2738);
not_4  g02362(new_n2635, new_n2739);
nand_1 g02363(new_n2639, new_n2739, new_n2740);
nor_1  g02364(new_n2637, new_n2636, new_n2741);
nand_1 g02365(new_n2659, new_n2640, new_n2742);
not_4  g02366(new_n2742, new_n2743);
xnor_1 g02367(new_n2743, new_n2741, new_n2744);
nand_1 g02368(new_n2744, new_n2740, new_n2745);
xnor_1 g02369(new_n2745, new_n2738, new_n2746);
xnor_1 g02370(new_n2746, new_n2708_1, new_n2747);
xnor_1 g02371(new_n2747, new_n2706, new_n2748);
nand_1 g02372(n12648, n4826, new_n2749_1);
nand_1 g02373(n10545, n7733, new_n2750);
nand_1 g02374(n12925, n7690, new_n2751);
not_4  g02375(new_n2751, new_n2752);
xnor_1 g02376(new_n2752, new_n2750, new_n2753);
xnor_1 g02377(new_n2753, new_n2749_1, new_n2754);
nand_1 g02378(n12925, n10545, new_n2755);
nand_1 g02379(n4826, n2530, new_n2756);
nand_1 g02380(new_n2756, new_n2755, new_n2757);
nand_1 g02381(n12648, n7733, new_n2758);
not_4  g02382(new_n2756, new_n2759);
xnor_1 g02383(new_n2759, new_n2755, new_n2760);
nand_1 g02384(new_n2760, new_n2758, new_n2761);
nand_1 g02385(new_n2761, new_n2757, new_n2762);
xnor_1 g02386(new_n2762, new_n2754, new_n2763);
not_4  g02387(new_n2763, new_n2764);
nand_1 g02388(n8476, n4970, new_n2765);
nand_1 g02389(n7610, n2530, new_n2766);
not_4  g02390(new_n2766, new_n2767);
xnor_1 g02391(new_n2767, new_n2765, new_n2768);
xnor_1 g02392(new_n2768, new_n2764, new_n2769);
nand_1 g02393(n8476, n7610, new_n2770);
nand_1 g02394(n12925, n12648, new_n2771);
nand_1 g02395(n8476, n4826, new_n2772);
nand_1 g02396(new_n2772, new_n2771, new_n2773);
nand_1 g02397(n7733, n2530, new_n2774);
not_4  g02398(new_n2772, new_n2775);
xnor_1 g02399(new_n2775, new_n2771, new_n2776);
nand_1 g02400(new_n2776, new_n2774, new_n2777);
nand_1 g02401(new_n2777, new_n2773, new_n2778);
nor_1  g02402(new_n2778, new_n2770, new_n2779);
not_4  g02403(new_n2779, new_n2780);
not_4  g02404(new_n2778, new_n2781);
xnor_1 g02405(new_n2781, new_n2770, new_n2782);
xnor_1 g02406(new_n2760, new_n2758, new_n2783);
nand_1 g02407(new_n2783, new_n2782, new_n2784);
nand_1 g02408(new_n2784, new_n2780, new_n2785);
nand_1 g02409(new_n2785, new_n2769, new_n2786);
not_4  g02410(new_n2786, new_n2787);
nor_1  g02411(new_n2785, new_n2769, new_n2788);
nor_1  g02412(new_n2788, new_n2787, new_n2789);
nand_1 g02413(n5331, n4970, new_n2790);
nand_1 g02414(n7610, n5331, new_n2791);
nand_1 g02415(n12925, n2530, new_n2792);
nand_1 g02416(n5331, n4826, new_n2793);
nand_1 g02417(new_n2793, new_n2792, new_n2794);
not_4  g02418(new_n2792, new_n2795);
not_4  g02419(new_n2793, new_n2796);
nand_1 g02420(new_n2796, new_n2795, new_n2797);
nand_1 g02421(n8476, n7733, new_n2798);
nand_1 g02422(new_n2798, new_n2797, new_n2799);
nand_1 g02423(new_n2799, new_n2794, new_n2800);
nor_1  g02424(new_n2800, new_n2791, new_n2801);
xnor_1 g02425(new_n2800, new_n2791, new_n2802_1);
not_4  g02426(new_n2776, new_n2803);
xnor_1 g02427(new_n2803, new_n2774, new_n2804);
nor_1  g02428(new_n2804, new_n2802_1, new_n2805);
nor_1  g02429(new_n2805, new_n2801, new_n2806);
nand_1 g02430(new_n2806, new_n2790, new_n2807);
xnor_1 g02431(new_n2783, new_n2782, new_n2808);
not_4  g02432(new_n2806, new_n2809);
xnor_1 g02433(new_n2809, new_n2790, new_n2810);
nand_1 g02434(new_n2810, new_n2808, new_n2811);
nand_1 g02435(new_n2811, new_n2807, new_n2812);
not_4  g02436(new_n2812, new_n2813);
nand_1 g02437(new_n2813, new_n2789, new_n2814);
nand_1 g02438(new_n2768, new_n2763, new_n2815);
nor_1  g02439(new_n2766, new_n2765, new_n2816);
xnor_1 g02440(new_n2787, new_n2816, new_n2817);
nand_1 g02441(new_n2817, new_n2815, new_n2818_1);
nor_1  g02442(new_n2751, new_n2750, new_n2819);
nand_1 g02443(n12648, n7610, new_n2820);
xnor_1 g02444(new_n2820, new_n2819, new_n2821);
nand_1 g02445(n7733, n7690, new_n2822);
nand_1 g02446(n10545, n4826, new_n2823);
nand_1 g02447(n12925, n3616, new_n2824);
not_4  g02448(new_n2824, new_n2825);
xnor_1 g02449(new_n2825, new_n2823, new_n2826);
xnor_1 g02450(new_n2826, new_n2822, new_n2827);
xnor_1 g02451(new_n2827, new_n2821, new_n2828);
not_4  g02452(new_n2749_1, new_n2829);
nand_1 g02453(new_n2753, new_n2829, new_n2830);
not_4  g02454(new_n2762, new_n2831);
nand_1 g02455(new_n2831, new_n2754, new_n2832);
nand_1 g02456(new_n2832, new_n2830, new_n2833);
nand_1 g02457(n8476, n503, new_n2834);
nand_1 g02458(n4970, n2530, new_n2835);
nand_1 g02459(n10965, n5331, new_n2836);
not_4  g02460(new_n2836, new_n2837);
xnor_1 g02461(new_n2837, new_n2835, new_n2838);
xnor_1 g02462(new_n2838, new_n2834, new_n2839);
not_4  g02463(new_n2839, new_n2840);
xnor_1 g02464(new_n2840, new_n2833, new_n2841);
xnor_1 g02465(new_n2841, new_n2828, new_n2842);
not_4  g02466(new_n2842, new_n2843);
xnor_1 g02467(new_n2843, new_n2818_1, new_n2844);
xnor_1 g02468(new_n2844, new_n2814, new_n2845);
nand_1 g02469(n5331, n503, new_n2846);
not_4  g02470(new_n2846, new_n2847);
xnor_1 g02471(new_n2812, new_n2789, new_n2848);
nand_1 g02472(new_n2848, new_n2847, new_n2849);
xnor_1 g02473(new_n2804, new_n2802_1, new_n2850);
not_4  g02474(new_n2798, new_n2851);
not_4  g02475(new_n2794, new_n2852);
nand_1 g02476(n12925, n5331, new_n2853);
nand_1 g02477(new_n2853, new_n2851, new_n2854);
nand_1 g02478(new_n2854, new_n2852, new_n2855);
nand_1 g02479(new_n2855, new_n2797, new_n2856);
nand_1 g02480(new_n2856, new_n2851, new_n2857);
nor_1  g02481(new_n2857, new_n2850, new_n2858);
xnor_1 g02482(new_n2810, new_n2808, new_n2859);
nand_1 g02483(new_n2859, new_n2858, new_n2860);
not_4  g02484(new_n2860, new_n2861);
xnor_1 g02485(new_n2848, new_n2846, new_n2862);
nand_1 g02486(new_n2862, new_n2861, new_n2863);
nand_1 g02487(new_n2863, new_n2849, new_n2864);
xnor_1 g02488(new_n2864, new_n2845, new_n2865);
nand_1 g02489(n4086, n2393, new_n2866);
not_4  g02490(new_n2866, new_n2867);
nand_1 g02491(n5860, n405, new_n2868);
nand_1 g02492(n8433, n3986, new_n2869);
not_4  g02493(new_n2869, new_n2870);
xnor_1 g02494(new_n2870, new_n2868, new_n2871);
xnor_1 g02495(new_n2871, new_n2867, new_n2872);
nand_1 g02496(n8433, n5860, new_n2873);
nand_1 g02497(n11892, n4086, new_n2874);
nand_1 g02498(new_n2874, new_n2873, new_n2875);
nand_1 g02499(n2393, n405, new_n2876);
not_4  g02500(new_n2874, new_n2877);
xnor_1 g02501(new_n2877, new_n2873, new_n2878);
nand_1 g02502(new_n2878, new_n2876, new_n2879_1);
nand_1 g02503(new_n2879_1, new_n2875, new_n2880);
nor_1  g02504(new_n2880, new_n2872, new_n2881);
not_4  g02505(new_n2881, new_n2882);
nand_1 g02506(new_n2880, new_n2872, new_n2883);
nand_1 g02507(new_n2883, new_n2882, new_n2884);
nand_1 g02508(n7388, n6611, new_n2885);
nand_1 g02509(n11892, n217, new_n2886);
not_4  g02510(new_n2886, new_n2887);
xnor_1 g02511(new_n2887, new_n2885, new_n2888);
xnor_1 g02512(new_n2888, new_n2884, new_n2889);
nand_1 g02513(n7388, n217, new_n2890);
nand_1 g02514(n8433, n2393, new_n2891);
nand_1 g02515(n7388, n4086, new_n2892);
nand_1 g02516(new_n2892, new_n2891, new_n2893);
nand_1 g02517(n11892, n405, new_n2894);
not_4  g02518(new_n2892, new_n2895);
xnor_1 g02519(new_n2895, new_n2891, new_n2896);
nand_1 g02520(new_n2896, new_n2894, new_n2897);
nand_1 g02521(new_n2897, new_n2893, new_n2898);
nor_1  g02522(new_n2898, new_n2890, new_n2899);
not_4  g02523(new_n2898, new_n2900);
xnor_1 g02524(new_n2900, new_n2890, new_n2901);
not_4  g02525(new_n2901, new_n2902_1);
not_4  g02526(new_n2878, new_n2903);
xnor_1 g02527(new_n2903, new_n2876, new_n2904);
nor_1  g02528(new_n2904, new_n2902_1, new_n2905);
nor_1  g02529(new_n2905, new_n2899, new_n2906);
xnor_1 g02530(new_n2906, new_n2889, new_n2907);
nand_1 g02531(n7965, n6611, new_n2908);
not_4  g02532(new_n2908, new_n2909);
xnor_1 g02533(new_n2904, new_n2901, new_n2910);
nand_1 g02534(new_n2910, new_n2909, new_n2911);
xnor_1 g02535(new_n2910, new_n2908, new_n2912);
nand_1 g02536(n7965, n217, new_n2913);
not_4  g02537(new_n2913, new_n2914);
nand_1 g02538(n11892, n8433, new_n2915);
not_4  g02539(new_n2915, new_n2916);
nand_1 g02540(n7965, n4086, new_n2917);
not_4  g02541(new_n2917, new_n2918);
nand_1 g02542(new_n2918, new_n2916, new_n2919);
nand_1 g02543(new_n2917, new_n2915, new_n2920);
nand_1 g02544(n7388, n405, new_n2921);
not_4  g02545(new_n2921, new_n2922);
nand_1 g02546(new_n2922, new_n2920, new_n2923);
nand_1 g02547(new_n2923, new_n2919, new_n2924);
nand_1 g02548(new_n2924, new_n2914, new_n2925);
xnor_1 g02549(new_n2924, new_n2914, new_n2926);
not_4  g02550(new_n2896, new_n2927);
xnor_1 g02551(new_n2927, new_n2894, new_n2928);
nor_1  g02552(new_n2928, new_n2926, new_n2929);
not_4  g02553(new_n2929, new_n2930);
nand_1 g02554(new_n2930, new_n2925, new_n2931);
nand_1 g02555(new_n2931, new_n2912, new_n2932);
nand_1 g02556(new_n2932, new_n2911, new_n2933);
nand_1 g02557(new_n2933, new_n2907, new_n2934);
not_4  g02558(new_n2884, new_n2935);
nand_1 g02559(new_n2888, new_n2935, new_n2936);
nor_1  g02560(new_n2886, new_n2885, new_n2937);
not_4  g02561(new_n2906, new_n2938);
nand_1 g02562(new_n2938, new_n2889, new_n2939);
not_4  g02563(new_n2939, new_n2940);
xnor_1 g02564(new_n2940, new_n2937, new_n2941);
nand_1 g02565(new_n2941, new_n2936, new_n2942);
not_4  g02566(new_n2868, new_n2943);
nand_1 g02567(new_n2870, new_n2943, new_n2944);
not_4  g02568(new_n2944, new_n2945);
nand_1 g02569(n2393, n217, new_n2946);
not_4  g02570(new_n2946, new_n2947);
nand_1 g02571(new_n2947, new_n2945, new_n2948);
nand_1 g02572(new_n2946, new_n2944, new_n2949);
nand_1 g02573(new_n2949, new_n2948, new_n2950);
not_4  g02574(new_n2950, new_n2951);
nand_1 g02575(n3986, n405, new_n2952);
nand_1 g02576(n5860, n4086, new_n2953);
nand_1 g02577(n8433, n5857, new_n2954);
not_4  g02578(new_n2954, new_n2955);
xnor_1 g02579(new_n2955, new_n2953, new_n2956);
xnor_1 g02580(new_n2956, new_n2952, new_n2957);
not_4  g02581(new_n2957, new_n2958);
xnor_1 g02582(new_n2958, new_n2951, new_n2959);
nand_1 g02583(new_n2871, new_n2867, new_n2960);
nand_1 g02584(new_n2882, new_n2960, new_n2961);
nand_1 g02585(n11296, n7965, new_n2962);
nand_1 g02586(n11892, n6611, new_n2963);
nand_1 g02587(n7388, n6359, new_n2964);
not_4  g02588(new_n2964, new_n2965);
xnor_1 g02589(new_n2965, new_n2963, new_n2966);
not_4  g02590(new_n2966, new_n2967);
xnor_1 g02591(new_n2967, new_n2962, new_n2968);
xnor_1 g02592(new_n2968, new_n2961, new_n2969);
xnor_1 g02593(new_n2969, new_n2959, new_n2970);
xnor_1 g02594(new_n2970, new_n2942, new_n2971);
xnor_1 g02595(new_n2971, new_n2934, new_n2972);
nand_1 g02596(n7965, n6359, new_n2973);
not_4  g02597(new_n2973, new_n2974);
not_4  g02598(new_n2907, new_n2975);
xnor_1 g02599(new_n2933, new_n2975, new_n2976);
nand_1 g02600(new_n2976, new_n2974, new_n2977);
nand_1 g02601(new_n2928, new_n2926, new_n2978);
nand_1 g02602(new_n2978, new_n2930, new_n2979);
not_4  g02603(new_n2979, new_n2980);
nand_1 g02604(new_n2920, new_n2919, new_n2981);
not_4  g02605(new_n2981, new_n2982);
nand_1 g02606(n8433, n7388, new_n2983);
not_4  g02607(new_n2983, new_n2984);
nand_1 g02608(n7965, n405, new_n2985);
not_4  g02609(new_n2985, new_n2986);
nand_1 g02610(new_n2986, new_n2984, new_n2987);
nor_1  g02611(new_n2987, new_n2982, new_n2988);
nand_1 g02612(new_n2988, new_n2980, new_n2989);
not_4  g02613(new_n2989, new_n2990);
not_4  g02614(new_n2931, new_n2991);
xnor_1 g02615(new_n2991, new_n2912, new_n2992);
nand_1 g02616(new_n2992, new_n2990, new_n2993);
not_4  g02617(new_n2993, new_n2994);
xnor_1 g02618(new_n2976, new_n2973, new_n2995);
nand_1 g02619(new_n2995, new_n2994, new_n2996);
nand_1 g02620(new_n2996, new_n2977, new_n2997);
nand_1 g02621(new_n2997, new_n2972, new_n2998);
not_4  g02622(new_n2998, new_n2999);
nor_1  g02623(new_n2997, new_n2972, new_n3000);
nor_1  g02624(new_n3000, new_n2999, new_n3001);
xnor_1 g02625(new_n3001, new_n2865, new_n3002);
xnor_1 g02626(new_n2862, new_n2860, new_n3003);
not_4  g02627(new_n3003, new_n3004);
nor_1  g02628(new_n2995, new_n2994, new_n3005);
not_4  g02629(new_n3005, new_n3006);
nand_1 g02630(new_n3006, new_n2996, new_n3007);
nand_1 g02631(new_n3007, new_n3004, new_n3008);
xnor_1 g02632(new_n2992, new_n2989, new_n3009);
not_4  g02633(new_n3009, new_n3010);
not_4  g02634(new_n2858, new_n3011);
nand_1 g02635(new_n2857, new_n2850, new_n3012);
nand_1 g02636(new_n3012, new_n3011, new_n3013);
not_4  g02637(new_n3013, new_n3014);
xnor_1 g02638(new_n2988, new_n2979, new_n3015);
nor_1  g02639(new_n3015, new_n3014, new_n3016);
not_4  g02640(new_n3016, new_n3017);
not_4  g02641(new_n2853, new_n3018);
nand_1 g02642(n8433, n7965, new_n3019);
not_4  g02643(new_n3019, new_n3020);
nand_1 g02644(new_n3020, new_n3018, new_n3021);
nand_1 g02645(new_n2985, new_n2983, new_n3022_1);
nand_1 g02646(new_n3022_1, new_n2987, new_n3023);
nand_1 g02647(new_n3023, new_n3021, new_n3024);
xnor_1 g02648(new_n3023, new_n3021, new_n3025);
not_4  g02649(new_n3025, new_n3026);
nand_1 g02650(n12925, n8476, new_n3027);
nand_1 g02651(n7733, n5331, new_n3028);
xnor_1 g02652(new_n3028, new_n3027, new_n3029);
nand_1 g02653(new_n3029, new_n3026, new_n3030);
nand_1 g02654(new_n3030, new_n3024, new_n3031);
nor_1  g02655(new_n2854, new_n2852, new_n3032);
nor_1  g02656(new_n3032, new_n2856, new_n3033);
not_4  g02657(new_n3033, new_n3034);
nand_1 g02658(new_n3034, new_n3031, new_n3035);
xnor_1 g02659(new_n3033, new_n3031, new_n3036);
nand_1 g02660(new_n3019, new_n2922, new_n3037);
nand_1 g02661(new_n3037, new_n2981, new_n3038);
not_4  g02662(new_n3037, new_n3039);
nand_1 g02663(new_n3039, new_n2920, new_n3040);
nand_1 g02664(new_n3040, new_n3038, new_n3041);
nand_1 g02665(new_n3041, new_n3036, new_n3042);
nand_1 g02666(new_n3042, new_n3035, new_n3043);
xnor_1 g02667(new_n3015, new_n3013, new_n3044);
nand_1 g02668(new_n3044, new_n3043, new_n3045);
nand_1 g02669(new_n3045, new_n3017, new_n3046);
nand_1 g02670(new_n3046, new_n3010, new_n3047);
not_4  g02671(new_n2859, new_n3048);
xnor_1 g02672(new_n3048, new_n2858, new_n3049);
not_4  g02673(new_n3049, new_n3050);
xnor_1 g02674(new_n3046, new_n3009, new_n3051);
nand_1 g02675(new_n3051, new_n3050, new_n3052);
nand_1 g02676(new_n3052, new_n3047, new_n3053);
not_4  g02677(new_n3053, new_n3054);
not_4  g02678(new_n3007, new_n3055);
nand_1 g02679(new_n3055, new_n3003, new_n3056);
nand_1 g02680(new_n3056, new_n3008, new_n3057);
nor_1  g02681(new_n3057, new_n3054, new_n3058);
not_4  g02682(new_n3058, new_n3059);
nand_1 g02683(new_n3059, new_n3008, new_n3060);
xnor_1 g02684(new_n3060, new_n3002, new_n3061);
xnor_1 g02685(new_n3061, new_n2748, new_n3062);
not_4  g02686(new_n3062, new_n3063);
xnor_1 g02687(new_n2704, new_n2702, new_n3064);
nand_1 g02688(new_n3057, new_n3054, new_n3065);
nand_1 g02689(new_n3065, new_n3059, new_n3066);
nor_1  g02690(new_n3066, new_n3064, new_n3067);
not_4  g02691(new_n3067, new_n3068);
nand_1 g02692(new_n3066, new_n3064, new_n3069);
nand_1 g02693(new_n3069, new_n3068, new_n3070);
xnor_1 g02694(new_n2701, new_n2699, new_n3071_1);
not_4  g02695(new_n3071_1, new_n3072);
xnor_1 g02696(new_n3051, new_n3049, new_n3073);
nor_1  g02697(new_n3073, new_n3072, new_n3074);
not_4  g02698(new_n3074, new_n3075);
nand_1 g02699(new_n3073, new_n3072, new_n3076);
nand_1 g02700(new_n3076, new_n3075, new_n3077);
not_4  g02701(new_n3077, new_n3078);
xnor_1 g02702(new_n2698, new_n2690, new_n3079);
not_4  g02703(new_n3079, new_n3080);
xnor_1 g02704(new_n3044, new_n3043, new_n3081);
nand_1 g02705(new_n3081, new_n3080, new_n3082);
xnor_1 g02706(new_n3081, new_n3079, new_n3083);
xnor_1 g02707(new_n3041, new_n3036, new_n3084);
not_4  g02708(new_n3084, new_n3085);
nand_1 g02709(n8759, n3719, new_n3086);
nand_1 g02710(new_n3086, new_n2675, new_n3087);
nand_1 g02711(new_n3087, new_n2691, new_n3088);
not_4  g02712(new_n3087, new_n3089);
nand_1 g02713(new_n3089, new_n2673, new_n3090);
nand_1 g02714(new_n3090, new_n3088, new_n3091);
nor_1  g02715(new_n3091, new_n3085, new_n3092);
not_4  g02716(new_n3092, new_n3093);
xnor_1 g02717(new_n3091, new_n3084, new_n3094);
xnor_1 g02718(new_n3029, new_n3025, new_n3095);
not_4  g02719(new_n3095, new_n3096);
nand_1 g02720(new_n2695, new_n2693, new_n3097);
nand_1 g02721(new_n3097, new_n2697, new_n3098);
not_4  g02722(new_n3098, new_n3099);
nand_1 g02723(new_n3099, new_n3096, new_n3100);
not_4  g02724(new_n3086, new_n3101);
nand_1 g02725(new_n3019, new_n2853, new_n3102);
nand_1 g02726(new_n3102, new_n3021, new_n3103);
not_4  g02727(new_n3103, new_n3104);
nand_1 g02728(new_n3104, new_n3101, new_n3105);
not_4  g02729(new_n3105, new_n3106);
xnor_1 g02730(new_n3098, new_n3096, new_n3107);
nand_1 g02731(new_n3107, new_n3106, new_n3108);
nand_1 g02732(new_n3108, new_n3100, new_n3109);
nand_1 g02733(new_n3109, new_n3094, new_n3110);
nand_1 g02734(new_n3110, new_n3093, new_n3111);
nand_1 g02735(new_n3111, new_n3083, new_n3112);
nand_1 g02736(new_n3112, new_n3082, new_n3113);
nand_1 g02737(new_n3113, new_n3078, new_n3114);
nand_1 g02738(new_n3114, new_n3075, new_n3115);
nor_1  g02739(new_n3115, new_n3070, new_n3116);
not_4  g02740(new_n3116, new_n3117);
nand_1 g02741(new_n3117, new_n3068, new_n3118);
not_4  g02742(new_n3118, new_n3119);
xnor_1 g02743(new_n3119, new_n3063, new_n3120);
nand_1 g02744(new_n3120, new_n2613, new_n3121);
xnor_1 g02745(new_n3120, new_n2613, new_n3122);
not_4  g02746(new_n3122, new_n3123);
xnor_1 g02747(new_n2610, new_n2608, new_n3124_1);
nand_1 g02748(new_n3115, new_n3070, new_n3125);
nand_1 g02749(new_n3125, new_n3117, new_n3126);
nand_1 g02750(new_n3126, new_n3124_1, new_n3127);
not_4  g02751(new_n2607, new_n3128);
nand_1 g02752(new_n3128, new_n2604, new_n3129);
nand_1 g02753(new_n3129, new_n2608, new_n3130);
not_4  g02754(new_n3130, new_n3131);
xnor_1 g02755(new_n3113, new_n3077, new_n3132);
nor_1  g02756(new_n3132, new_n3131, new_n3133);
not_4  g02757(new_n3133, new_n3134);
nand_1 g02758(new_n3132, new_n3131, new_n3135);
nand_1 g02759(new_n3135, new_n3134, new_n3136);
xnor_1 g02760(new_n2603, new_n2595, new_n3137);
xnor_1 g02761(new_n3111, new_n3083, new_n3138);
nand_1 g02762(new_n3138, new_n3137, new_n3139);
xnor_1 g02763(new_n3109, new_n3094, new_n3140);
nand_1 g02764(n9956, n5305, new_n3141);
nand_1 g02765(new_n3141, new_n2542, new_n3142);
nand_1 g02766(new_n3142, new_n2596, new_n3143);
not_4  g02767(new_n3142, new_n3144);
nand_1 g02768(new_n3144, new_n2540, new_n3145);
nand_1 g02769(new_n3145, new_n3143, new_n3146_1);
nand_1 g02770(new_n3146_1, new_n3140, new_n3147);
xnor_1 g02771(new_n3146_1, new_n3140, new_n3148);
not_4  g02772(new_n3141, new_n3149);
xnor_1 g02773(new_n3104, new_n3086, new_n3150);
nand_1 g02774(new_n3150, new_n3149, new_n3151);
nand_1 g02775(new_n2600, new_n2598, new_n3152);
nand_1 g02776(new_n3152, new_n2602, new_n3153);
nand_1 g02777(new_n3153, new_n3151, new_n3154);
xnor_1 g02778(new_n3107, new_n3105, new_n3155);
xnor_1 g02779(new_n3153, new_n3151, new_n3156);
nor_1  g02780(new_n3156, new_n3155, new_n3157);
not_4  g02781(new_n3157, new_n3158);
nand_1 g02782(new_n3158, new_n3154, new_n3159);
not_4  g02783(new_n3159, new_n3160);
nor_1  g02784(new_n3160, new_n3148, new_n3161);
not_4  g02785(new_n3161, new_n3162);
nand_1 g02786(new_n3162, new_n3147, new_n3163);
not_4  g02787(new_n3163, new_n3164);
xnor_1 g02788(new_n3138, new_n3137, new_n3165);
nor_1  g02789(new_n3165, new_n3164, new_n3166);
not_4  g02790(new_n3166, new_n3167);
nand_1 g02791(new_n3167, new_n3139, new_n3168);
not_4  g02792(new_n3168, new_n3169);
nor_1  g02793(new_n3169, new_n3136, new_n3170);
nor_1  g02794(new_n3170, new_n3133, new_n3171);
xnor_1 g02795(new_n3126, new_n3124_1, new_n3172_1);
not_4  g02796(new_n3172_1, new_n3173);
nand_1 g02797(new_n3173, new_n3171, new_n3174);
nand_1 g02798(new_n3174, new_n3127, new_n3175);
nand_1 g02799(new_n3175, new_n3123, new_n3176);
nand_1 g02800(new_n3176, new_n3121, new_n3177);
not_4  g02801(new_n3177, new_n3178);
not_4  g02802(new_n2748, new_n3179);
nand_1 g02803(new_n3061, new_n3179, new_n3180);
nand_1 g02804(new_n3119, new_n3062, new_n3181);
nand_1 g02805(new_n3181, new_n3180, new_n3182);
not_4  g02806(new_n2820, new_n3183);
nand_1 g02807(new_n3183, new_n2819, new_n3184);
nand_1 g02808(new_n2827, new_n2821, new_n3185);
nand_1 g02809(new_n3185, new_n3184, new_n3186);
nand_1 g02810(new_n2824, new_n2823, new_n3187);
nand_1 g02811(new_n2826, new_n2822, new_n3188);
nand_1 g02812(new_n3188, new_n3187, new_n3189);
nand_1 g02813(n12648, n4970, new_n3190);
nand_1 g02814(n11296, n7388, new_n3191);
nand_1 g02815(n9241, n6126, new_n3192);
not_4  g02816(new_n3192, new_n3193);
xnor_1 g02817(new_n3193, new_n3191, new_n3194);
xnor_1 g02818(new_n3194, new_n3190, new_n3195);
xnor_1 g02819(new_n3195, new_n3189, new_n3196);
xnor_1 g02820(new_n3196, new_n3186, new_n3197);
nand_1 g02821(new_n2954, new_n2953, new_n3198);
nand_1 g02822(new_n2956, new_n2952, new_n3199);
nand_1 g02823(new_n3199, new_n3198, new_n3200);
nand_1 g02824(new_n2964, new_n2963, new_n3201);
nand_1 g02825(new_n2966, new_n2962, new_n3202);
nand_1 g02826(new_n3202, new_n3201, new_n3203);
xnor_1 g02827(new_n3203, new_n3200, new_n3204);
nand_1 g02828(n11892, n6359, new_n3205);
nand_1 g02829(n7546, n5331, new_n3206);
xnor_1 g02830(new_n3206, new_n3205, new_n3207);
xnor_1 g02831(new_n3207, new_n3204, new_n3208);
nor_1  g02832(new_n2722, new_n2720, new_n3209);
nor_1  g02833(new_n2735, new_n2726, new_n3210);
nor_1  g02834(new_n3210, new_n3209, new_n3211);
nand_1 g02835(n8595, n8276, new_n3212);
nand_1 g02836(n6611, n2393, new_n3213);
xnor_1 g02837(new_n3213, new_n3212, new_n3214_1);
nand_1 g02838(n12925, n4499, new_n3215);
nand_1 g02839(n11536, n5305, new_n3216);
xnor_1 g02840(new_n3216, new_n3215, new_n3217);
xnor_1 g02841(new_n3217, new_n3214_1, new_n3218);
xnor_1 g02842(new_n3218, new_n3211, new_n3219);
xnor_1 g02843(new_n3219, new_n3208, new_n3220);
nand_1 g02844(new_n2957, new_n2951, new_n3221);
nand_1 g02845(new_n3221, new_n2948, new_n3222);
nand_1 g02846(new_n2836, new_n2835, new_n3223);
nand_1 g02847(new_n2838, new_n2834, new_n3224);
nand_1 g02848(new_n3224, new_n3223, new_n3225);
nand_1 g02849(n4086, n3986, new_n3226);
nand_1 g02850(n7733, n3616, new_n3227);
not_4  g02851(new_n3227, new_n3228);
xnor_1 g02852(new_n3228, new_n3226, new_n3229);
xnor_1 g02853(new_n3229, new_n3225, new_n3230_1);
xnor_1 g02854(new_n3230_1, new_n3222, new_n3231);
xnor_1 g02855(new_n3231, new_n3220, new_n3232);
xnor_1 g02856(new_n3232, new_n3197, new_n3233);
not_4  g02857(new_n2971, new_n3234);
nor_1  g02858(new_n3234, new_n2934, new_n3235);
nor_1  g02859(new_n2999, new_n3235, new_n3236);
nand_1 g02860(n5860, n217, new_n3237);
xnor_1 g02861(new_n3237, new_n3236, new_n3238);
not_4  g02862(new_n2708_1, new_n3239);
nand_1 g02863(new_n2746, new_n3239, new_n3240);
nand_1 g02864(new_n2747, new_n2706, new_n3241);
nand_1 g02865(new_n3241, new_n3240, new_n3242);
nand_1 g02866(new_n2839, new_n2833, new_n3243);
not_4  g02867(new_n2828, new_n3244);
nand_1 g02868(new_n2841, new_n3244, new_n3245);
nand_1 g02869(new_n3245, new_n3243, new_n3246);
nand_1 g02870(n12299, n8065, new_n3247);
nand_1 g02871(n10510, n3602, new_n3248);
xnor_1 g02872(new_n3248, new_n3247, new_n3249);
nand_1 g02873(n10644, n3719, new_n3250);
nand_1 g02874(n7965, n1357, new_n3251);
xnor_1 g02875(new_n3251, new_n3250, new_n3252);
nand_1 g02876(n10439, n7436, new_n3253);
nand_1 g02877(n8759, n4190, new_n3254);
xnor_1 g02878(new_n3254, new_n3253, new_n3255);
xnor_1 g02879(new_n3255, new_n3252, new_n3256);
xnor_1 g02880(new_n3256, new_n3249, new_n3257);
not_4  g02881(new_n3257, new_n3258);
nand_1 g02882(new_n2565, new_n2564_1, new_n3259);
nand_1 g02883(new_n2567, new_n2563, new_n3260);
nand_1 g02884(new_n3260, new_n3259, new_n3261);
nand_1 g02885(n9637, n1097, new_n3262);
xnor_1 g02886(new_n3262, new_n3261, new_n3263);
xnor_1 g02887(new_n3263, new_n3258, new_n3264);
xnor_1 g02888(new_n3264, new_n3246, new_n3265);
not_4  g02889(new_n2710, new_n3266);
nand_1 g02890(new_n2717, new_n3266, new_n3267);
not_4  g02891(new_n2737, new_n3268);
nand_1 g02892(new_n3268, new_n2718, new_n3269);
nand_1 g02893(new_n3269, new_n3267, new_n3270);
not_4  g02894(new_n2568, new_n3271);
nand_1 g02895(new_n3271, new_n2562, new_n3272_1);
nand_1 g02896(new_n2579, new_n2569, new_n3273);
nand_1 g02897(new_n3273, new_n3272_1, new_n3274);
xnor_1 g02898(new_n3274, new_n3270, new_n3275);
xnor_1 g02899(new_n3275, new_n3265, new_n3276);
nand_1 g02900(new_n2743, new_n2741, new_n3277);
not_4  g02901(new_n2738, new_n3278);
nand_1 g02902(new_n2745, new_n3278, new_n3279);
nand_1 g02903(new_n3279, new_n3277, new_n3280);
nand_1 g02904(new_n2714, new_n2713, new_n3281);
nand_1 g02905(new_n2716, new_n2711, new_n3282);
nand_1 g02906(new_n3282, new_n3281, new_n3283);
nand_1 g02907(n4312, n2577, new_n3284);
not_4  g02908(new_n3284, new_n3285);
xnor_1 g02909(new_n3285, new_n3283, new_n3286);
not_4  g02910(new_n2727, new_n3287_1);
nand_1 g02911(new_n2730, new_n3287_1, new_n3288);
nand_1 g02912(new_n3288, new_n2733, new_n3289);
nand_1 g02913(n11257, n4921, new_n3290);
nand_1 g02914(n12705, n3842, new_n3291);
xnor_1 g02915(new_n3291, new_n3290, new_n3292);
xnor_1 g02916(new_n3292, new_n3289, new_n3293);
xnor_1 g02917(new_n3293, new_n3286, new_n3294);
nand_1 g02918(n8433, n45, new_n3295);
nand_1 g02919(n12025, n11917, new_n3296);
xnor_1 g02920(new_n3296, new_n3295, new_n3297);
nand_1 g02921(new_n2575, new_n2574, new_n3298);
nand_1 g02922(new_n2577_1, new_n2572, new_n3299);
nand_1 g02923(new_n3299, new_n3298, new_n3300);
nand_1 g02924(n5964, n1835, new_n3301);
nand_1 g02925(n5857, n405, new_n3302);
xnor_1 g02926(new_n3302, new_n3301, new_n3303);
xnor_1 g02927(new_n3303, new_n3300, new_n3304);
xnor_1 g02928(new_n3304, new_n3297, new_n3305);
nand_1 g02929(new_n2570, new_n2486, new_n3306);
not_4  g02930(new_n2571, new_n3307);
nand_1 g02931(new_n2578, new_n3307, new_n3308);
nand_1 g02932(new_n3308, new_n3306, new_n3309);
nand_1 g02933(n10391, n6776, new_n3310);
xnor_1 g02934(new_n3310, new_n3309, new_n3311);
xnor_1 g02935(new_n3311, new_n3305, new_n3312);
xnor_1 g02936(new_n3312, new_n3294, new_n3313);
xnor_1 g02937(new_n3313, new_n3280, new_n3314);
xnor_1 g02938(new_n3314, new_n3276, new_n3315);
not_4  g02939(new_n3315, new_n3316);
xnor_1 g02940(new_n3316, new_n3242, new_n3317);
xnor_1 g02941(new_n3317, new_n3238, new_n3318);
xnor_1 g02942(new_n3318, new_n3233, new_n3319);
not_4  g02943(new_n2865, new_n3320);
nor_1  g02944(new_n3001, new_n3320, new_n3321);
not_4  g02945(new_n3321, new_n3322);
nand_1 g02946(new_n3060, new_n3002, new_n3323);
nand_1 g02947(new_n3323, new_n3322, new_n3324);
nand_1 g02948(new_n2940, new_n2937, new_n3325);
not_4  g02949(new_n2970, new_n3326);
nand_1 g02950(new_n3326, new_n2942, new_n3327);
nand_1 g02951(new_n3327, new_n3325, new_n3328);
nor_1  g02952(new_n2525, new_n2504, new_n3329);
not_4  g02953(new_n3329, new_n3330);
nand_1 g02954(new_n2585_1, new_n2580, new_n3331);
nand_1 g02955(new_n3331, new_n3330, new_n3332);
xnor_1 g02956(new_n3332, new_n3328, new_n3333);
xnor_1 g02957(new_n3333, new_n3324, new_n3334);
xnor_1 g02958(new_n3334, new_n3319, new_n3335);
xnor_1 g02959(new_n3335, new_n3182, new_n3336);
not_4  g02960(new_n2814, new_n3337);
nand_1 g02961(new_n2844, new_n3337, new_n3338);
nand_1 g02962(new_n2864, new_n2845, new_n3339_1);
nand_1 g02963(new_n3339_1, new_n3338, new_n3340);
not_4  g02964(new_n2590, new_n3341);
nand_1 g02965(new_n2612, new_n3341, new_n3342_1);
nand_1 g02966(new_n3342_1, new_n2588, new_n3343);
xnor_1 g02967(new_n3343, new_n3340, new_n3344);
nand_1 g02968(new_n2787, new_n2816, new_n3345);
nand_1 g02969(new_n2842, new_n2818_1, new_n3346);
nand_1 g02970(new_n3346, new_n3345, new_n3347);
not_4  g02971(new_n2961, new_n3348);
nand_1 g02972(new_n2968, new_n3348, new_n3349);
not_4  g02973(new_n2959, new_n3350);
nand_1 g02974(new_n2969, new_n3350, new_n3351);
nand_1 g02975(new_n3351, new_n3349, new_n3352);
nand_1 g02976(n10547, n9956, new_n3353);
nand_1 g02977(n10965, n8476, new_n3354);
nand_1 g02978(n7690, n4826, new_n3355);
xnor_1 g02979(new_n3355, new_n3354, new_n3356);
nand_1 g02980(n10545, n7610, new_n3357);
nand_1 g02981(n2530, n503, new_n3358);
xnor_1 g02982(new_n3358, new_n3357, new_n3359);
xnor_1 g02983(new_n3359, new_n3356, new_n3360);
xnor_1 g02984(new_n3360, new_n3353, new_n3361);
xnor_1 g02985(new_n3361, new_n3352, new_n3362);
xnor_1 g02986(new_n3362, new_n3347, new_n3363);
xnor_1 g02987(new_n3363, new_n3344, new_n3364);
xnor_1 g02988(new_n3364, new_n3336, new_n3365);
nand_1 g02989(new_n3365, new_n3178, new_n3366);
not_4  g02990(new_n3364, new_n3367);
xnor_1 g02991(new_n3367, new_n3336, new_n3368);
nand_1 g02992(new_n3368, new_n3177, new_n3369);
nand_1 g02993(new_n3369, new_n3366, n837);
nand_1 g02994(n11917, n11757, new_n3371);
nand_1 g02995(n9956, n5240, new_n3372);
not_4  g02996(new_n3372, new_n3373);
nand_1 g02997(n11757, n4921, new_n3374);
nand_1 g02998(n11917, n3172, new_n3375);
not_4  g02999(new_n3375, new_n3376);
xnor_1 g03000(new_n3376, new_n3372, new_n3377);
nand_1 g03001(new_n3377, new_n3374, new_n3378);
nand_1 g03002(new_n3378, new_n3373, new_n3379);
nand_1 g03003(new_n3379, new_n3371, new_n3380);
not_4  g03004(new_n3371, new_n3381);
nand_1 g03005(n4921, n3172, new_n3382);
nand_1 g03006(new_n3382, new_n3379, new_n3383);
nand_1 g03007(new_n3383, new_n3381, new_n3384);
nand_1 g03008(new_n3384, new_n3380, new_n3385);
not_4  g03009(new_n3385, new_n3386);
nand_1 g03010(n5240, n4921, new_n3387);
nand_1 g03011(n11821, n9956, new_n3388);
nand_1 g03012(new_n3388, new_n3387, new_n3389);
not_4  g03013(new_n3387, new_n3390);
not_4  g03014(new_n3388, new_n3391);
nand_1 g03015(new_n3391, new_n3390, new_n3392);
nand_1 g03016(new_n3392, new_n3389, new_n3393);
xnor_1 g03017(new_n3393, new_n3386, new_n3394);
not_4  g03018(new_n3394, new_n3395);
nand_1 g03019(n2577, n1333, new_n3396);
nand_1 g03020(n3842, n3172, new_n3397);
not_4  g03021(new_n3397, new_n3398);
xnor_1 g03022(new_n3398, new_n3396, new_n3399);
xnor_1 g03023(new_n3399, new_n3395, new_n3400);
nand_1 g03024(n3842, n1333, new_n3401);
nand_1 g03025(n11757, n9956, new_n3402);
nand_1 g03026(n11917, n1333, new_n3403);
nand_1 g03027(new_n3403, new_n3402, new_n3404);
nor_1  g03028(new_n3403, new_n3402, new_n3405);
not_4  g03029(new_n3405, new_n3406);
nand_1 g03030(new_n3406, new_n3382, new_n3407);
nand_1 g03031(new_n3407, new_n3404, new_n3408);
nor_1  g03032(new_n3408, new_n3401, new_n3409);
not_4  g03033(new_n3409, new_n3410);
not_4  g03034(new_n3374, new_n3411);
not_4  g03035(new_n3377, new_n3412);
nand_1 g03036(new_n3412, new_n3411, new_n3413);
nand_1 g03037(new_n3413, new_n3378, new_n3414);
nand_1 g03038(new_n3408, new_n3401, new_n3415);
nand_1 g03039(new_n3415, new_n3410, new_n3416);
not_4  g03040(new_n3416, new_n3417);
nand_1 g03041(new_n3417, new_n3414, new_n3418);
nand_1 g03042(new_n3418, new_n3410, new_n3419);
xnor_1 g03043(new_n3419, new_n3400, new_n3420);
not_4  g03044(new_n3420, new_n3421);
nand_1 g03045(n7862, n2577, new_n3422);
not_4  g03046(new_n3422, new_n3423);
xnor_1 g03047(new_n3416, new_n3414, new_n3424);
nand_1 g03048(new_n3424, new_n3423, new_n3425);
nand_1 g03049(n7862, n3842, new_n3426);
not_4  g03050(new_n3426, new_n3427);
nand_1 g03051(n9956, n3172, new_n3428);
not_4  g03052(new_n3428, new_n3429);
nand_1 g03053(n11917, n7862, new_n3430);
not_4  g03054(new_n3430, new_n3431);
nand_1 g03055(new_n3431, new_n3429, new_n3432);
nand_1 g03056(new_n3430, new_n3428, new_n3433);
nand_1 g03057(n4921, n1333, new_n3434);
not_4  g03058(new_n3434, new_n3435);
nand_1 g03059(new_n3435, new_n3433, new_n3436);
nand_1 g03060(new_n3436, new_n3432, new_n3437);
nand_1 g03061(new_n3437, new_n3427, new_n3438);
xnor_1 g03062(new_n3437, new_n3426, new_n3439);
not_4  g03063(new_n3439, new_n3440);
nand_1 g03064(new_n3406, new_n3404, new_n3441);
xnor_1 g03065(new_n3441, new_n3382, new_n3442);
nor_1  g03066(new_n3442, new_n3440, new_n3443);
not_4  g03067(new_n3443, new_n3444);
nand_1 g03068(new_n3444, new_n3438, new_n3445);
xnor_1 g03069(new_n3424, new_n3422, new_n3446);
nand_1 g03070(new_n3446, new_n3445, new_n3447);
nand_1 g03071(new_n3447, new_n3425, new_n3448);
nand_1 g03072(new_n3448, new_n3421, new_n3449);
not_4  g03073(new_n3393, new_n3450);
nand_1 g03074(new_n3450, new_n3386, new_n3451);
nand_1 g03075(new_n3451, new_n3384, new_n3452);
nand_1 g03076(n9637, n1333, new_n3453);
nand_1 g03077(n3172, n2577, new_n3454);
nand_1 g03078(n7862, n1835, new_n3455);
nand_1 g03079(new_n3455, new_n3454, new_n3456_1);
not_4  g03080(new_n3454, new_n3457);
not_4  g03081(new_n3455, new_n3458);
nand_1 g03082(new_n3458, new_n3457, new_n3459);
nand_1 g03083(new_n3459, new_n3456_1, new_n3460);
xnor_1 g03084(new_n3460, new_n3453, new_n3461);
xnor_1 g03085(new_n3461, new_n3452, new_n3462);
not_4  g03086(new_n3392, new_n3463);
nand_1 g03087(n11757, n3842, new_n3464);
not_4  g03088(new_n3464, new_n3465);
nand_1 g03089(new_n3465, new_n3463, new_n3466);
nand_1 g03090(new_n3464, new_n3392, new_n3467);
nand_1 g03091(new_n3467, new_n3466, new_n3468);
not_4  g03092(new_n3468, new_n3469);
nand_1 g03093(n11821, n4921, new_n3470);
nand_1 g03094(n9956, n9080, new_n3471);
nand_1 g03095(n11917, n5240, new_n3472);
not_4  g03096(new_n3472, new_n3473);
xnor_1 g03097(new_n3473, new_n3471, new_n3474);
xnor_1 g03098(new_n3474, new_n3470, new_n3475);
not_4  g03099(new_n3475, new_n3476);
xnor_1 g03100(new_n3476, new_n3469, new_n3477);
xnor_1 g03101(new_n3477, new_n3462, new_n3478);
nand_1 g03102(new_n3399, new_n3394, new_n3479);
nor_1  g03103(new_n3397, new_n3396, new_n3480);
nand_1 g03104(new_n3419, new_n3400, new_n3481);
not_4  g03105(new_n3481, new_n3482);
xnor_1 g03106(new_n3482, new_n3480, new_n3483);
nand_1 g03107(new_n3483, new_n3479, new_n3484);
xnor_1 g03108(new_n3484, new_n3478, new_n3485);
xnor_1 g03109(new_n3485, new_n3449, new_n3486);
nand_1 g03110(n9637, n7862, new_n3487);
not_4  g03111(new_n3487, new_n3488);
xnor_1 g03112(new_n3448, new_n3420, new_n3489);
nand_1 g03113(new_n3489, new_n3488, new_n3490);
xnor_1 g03114(new_n3442, new_n3439, new_n3491);
nand_1 g03115(new_n3433, new_n3432, new_n3492);
not_4  g03116(new_n3492, new_n3493);
nand_1 g03117(n9956, n1333, new_n3494);
not_4  g03118(new_n3494, new_n3495);
nand_1 g03119(n7862, n4921, new_n3496);
not_4  g03120(new_n3496, new_n3497);
nand_1 g03121(new_n3497, new_n3495, new_n3498);
nor_1  g03122(new_n3498, new_n3493, new_n3499);
nand_1 g03123(new_n3499, new_n3491, new_n3500);
not_4  g03124(new_n3500, new_n3501);
xnor_1 g03125(new_n3446, new_n3445, new_n3502);
not_4  g03126(new_n3502, new_n3503);
nand_1 g03127(new_n3503, new_n3501, new_n3504);
not_4  g03128(new_n3504, new_n3505);
xnor_1 g03129(new_n3489, new_n3487, new_n3506);
nand_1 g03130(new_n3506, new_n3505, new_n3507);
nand_1 g03131(new_n3507, new_n3490, new_n3508);
xnor_1 g03132(new_n3508, new_n3486, new_n3509);
xnor_1 g03133(new_n3506, new_n3504, new_n3510);
not_4  g03134(new_n3510, new_n3511);
nand_1 g03135(n8595, n6877, new_n3512);
nand_1 g03136(n6877, n6126, new_n3513);
nand_1 g03137(n3719, n2464, new_n3514);
nand_1 g03138(new_n3514, new_n3513, new_n3515);
nand_1 g03139(n6877, n3719, new_n3516);
not_4  g03140(new_n3516, new_n3517);
nand_1 g03141(n6126, n2464, new_n3518);
not_4  g03142(new_n3518, new_n3519);
nand_1 g03143(new_n3519, new_n3517, new_n3520);
nand_1 g03144(n9400, n3602, new_n3521);
nand_1 g03145(new_n3521, new_n3520, new_n3522);
nand_1 g03146(new_n3522, new_n3515, new_n3523);
nor_1  g03147(new_n3523, new_n3512, new_n3524);
not_4  g03148(new_n3524, new_n3525);
nand_1 g03149(new_n3523, new_n3512, new_n3526);
nand_1 g03150(new_n3526, new_n3525, new_n3527);
nand_1 g03151(n3602, n2464, new_n3528);
not_4  g03152(new_n3528, new_n3529);
nand_1 g03153(n9400, n6126, new_n3530);
nand_1 g03154(n11311, n3719, new_n3531);
nand_1 g03155(new_n3531, new_n3530, new_n3532);
not_4  g03156(new_n3530, new_n3533);
not_4  g03157(new_n3531, new_n3534);
nand_1 g03158(new_n3534, new_n3533, new_n3535);
nand_1 g03159(new_n3535, new_n3532, new_n3536);
xnor_1 g03160(new_n3536, new_n3529, new_n3537);
xnor_1 g03161(new_n3537, new_n3527, new_n3538);
not_4  g03162(new_n3521, new_n3539);
nand_1 g03163(new_n3539, new_n3516, new_n3540);
nand_1 g03164(new_n3520, new_n3515, new_n3541);
nand_1 g03165(new_n3541, new_n3540, new_n3542);
not_4  g03166(new_n3542, new_n3543);
nand_1 g03167(new_n3543, new_n3539, new_n3544);
not_4  g03168(new_n3544, new_n3545);
nand_1 g03169(new_n3545, new_n3538, new_n3546);
not_4  g03170(new_n3546, new_n3547);
nand_1 g03171(n10439, n6877, new_n3548);
nand_1 g03172(n9400, n8595, new_n3549);
nand_1 g03173(new_n3535, new_n3528, new_n3550);
nand_1 g03174(new_n3550, new_n3532, new_n3551);
not_4  g03175(new_n3551, new_n3552);
xnor_1 g03176(new_n3552, new_n3549, new_n3553);
nand_1 g03177(n11311, n3602, new_n3554);
nand_1 g03178(n4187, n3719, new_n3555);
xnor_1 g03179(new_n3555, new_n3519, new_n3556);
not_4  g03180(new_n3556, new_n3557);
xnor_1 g03181(new_n3557, new_n3554, new_n3558);
xnor_1 g03182(new_n3558, new_n3553, new_n3559);
xnor_1 g03183(new_n3559, new_n3548, new_n3560);
not_4  g03184(new_n3527, new_n3561);
nand_1 g03185(new_n3537, new_n3561, new_n3562);
nand_1 g03186(new_n3562, new_n3525, new_n3563);
xnor_1 g03187(new_n3563, new_n3560, new_n3564);
not_4  g03188(new_n3564, new_n3565);
nand_1 g03189(new_n3565, new_n3547, new_n3566);
not_4  g03190(new_n3566, new_n3567);
nand_1 g03191(n8065, n6877, new_n3568);
not_4  g03192(new_n3568, new_n3569);
nand_1 g03193(n11311, n6126, new_n3570);
not_4  g03194(new_n3570, new_n3571);
nand_1 g03195(n4203, n3719, new_n3572);
nand_1 g03196(n4187, n3602, new_n3573);
not_4  g03197(new_n3573, new_n3574);
xnor_1 g03198(new_n3574, new_n3572, new_n3575);
xnor_1 g03199(new_n3575, new_n3571, new_n3576);
nand_1 g03200(new_n3555, new_n3518, new_n3577);
nand_1 g03201(new_n3556, new_n3554, new_n3578);
nand_1 g03202(new_n3578, new_n3577, new_n3579);
nor_1  g03203(new_n3579, new_n3576, new_n3580);
not_4  g03204(new_n3580, new_n3581);
nand_1 g03205(new_n3579, new_n3576, new_n3582);
nand_1 g03206(new_n3582, new_n3581, new_n3583);
nand_1 g03207(n10439, n9400, new_n3584);
nand_1 g03208(n8595, n2464, new_n3585);
not_4  g03209(new_n3585, new_n3586);
xnor_1 g03210(new_n3586, new_n3584, new_n3587);
xnor_1 g03211(new_n3587, new_n3583, new_n3588);
nor_1  g03212(new_n3551, new_n3549, new_n3589);
not_4  g03213(new_n3553, new_n3590);
nor_1  g03214(new_n3558, new_n3590, new_n3591);
nor_1  g03215(new_n3591, new_n3589, new_n3592);
not_4  g03216(new_n3592, new_n3593);
xnor_1 g03217(new_n3593, new_n3588, new_n3594);
not_4  g03218(new_n3548, new_n3595);
nand_1 g03219(new_n3559, new_n3595, new_n3596);
nand_1 g03220(new_n3563, new_n3560, new_n3597);
nand_1 g03221(new_n3597, new_n3596, new_n3598);
xnor_1 g03222(new_n3598, new_n3594, new_n3599);
xnor_1 g03223(new_n3599, new_n3569, new_n3600);
xnor_1 g03224(new_n3600, new_n3567, new_n3601);
not_4  g03225(new_n3601, new_n3602_1);
xnor_1 g03226(new_n3565, new_n3546, new_n3603);
not_4  g03227(new_n3603, new_n3604);
not_4  g03228(new_n3538, new_n3605);
xnor_1 g03229(new_n3545, new_n3605, new_n3606);
not_4  g03230(new_n3540, new_n3607);
nand_1 g03231(new_n3607, new_n3515, new_n3608);
nand_1 g03232(new_n3608, new_n3542, new_n3609);
not_4  g03233(new_n3609, new_n3610);
nand_1 g03234(n8433, n7236, new_n3611);
not_4  g03235(new_n3611, new_n3612);
nand_1 g03236(n12925, n4805, new_n3613);
not_4  g03237(new_n3613, new_n3614);
nand_1 g03238(new_n3614, new_n3612, new_n3615);
nand_1 g03239(n7733, n4805, new_n3616_1);
nand_1 g03240(n12925, n11478, new_n3617);
nand_1 g03241(new_n3617, new_n3616_1, new_n3618);
not_4  g03242(new_n3616_1, new_n3619);
not_4  g03243(new_n3617, new_n3620);
nand_1 g03244(new_n3620, new_n3619, new_n3621);
nand_1 g03245(new_n3621, new_n3618, new_n3622);
nand_1 g03246(new_n3622, new_n3615, new_n3623);
not_4  g03247(new_n3615, new_n3624);
xnor_1 g03248(new_n3622, new_n3624, new_n3625);
nand_1 g03249(n7236, n405, new_n3626);
nand_1 g03250(n8433, n3992, new_n3627_1);
xnor_1 g03251(new_n3627_1, new_n3626, new_n3628);
nand_1 g03252(new_n3628, new_n3625, new_n3629);
nand_1 g03253(new_n3629, new_n3623, new_n3630);
nand_1 g03254(n3992, n405, new_n3631);
nor_1  g03255(new_n3631, new_n3612, new_n3632);
nand_1 g03256(n8433, n8384, new_n3633);
nand_1 g03257(n7236, n4086, new_n3634);
nand_1 g03258(new_n3634, new_n3633, new_n3635);
nor_1  g03259(new_n3635, new_n3632, new_n3636);
not_4  g03260(new_n3633, new_n3637);
not_4  g03261(new_n3634, new_n3638);
nand_1 g03262(new_n3638, new_n3637, new_n3639);
not_4  g03263(new_n3639, new_n3640);
nor_1  g03264(new_n3640, new_n3636, new_n3641);
nand_1 g03265(new_n3635, new_n3632, new_n3642);
nand_1 g03266(new_n3642, new_n3641, new_n3643);
not_4  g03267(new_n3643, new_n3644);
xnor_1 g03268(new_n3644, new_n3630, new_n3645);
nand_1 g03269(n11478, n7733, new_n3646);
not_4  g03270(new_n3646, new_n3647);
nand_1 g03271(new_n3647, new_n3613, new_n3648);
not_4  g03272(new_n3648, new_n3649);
nand_1 g03273(n12925, n5283, new_n3650);
nand_1 g03274(n4826, n4805, new_n3651);
nand_1 g03275(new_n3651, new_n3650, new_n3652);
not_4  g03276(new_n3652, new_n3653);
nand_1 g03277(new_n3653, new_n3649, new_n3654_1);
nor_1  g03278(new_n3651, new_n3650, new_n3655);
not_4  g03279(new_n3655, new_n3656);
nand_1 g03280(new_n3656, new_n3652, new_n3657);
not_4  g03281(new_n3657, new_n3658);
nand_1 g03282(new_n3658, new_n3648, new_n3659);
nand_1 g03283(new_n3659, new_n3654_1, new_n3660);
not_4  g03284(new_n3660, new_n3661_1);
xnor_1 g03285(new_n3661_1, new_n3645, new_n3662);
nand_1 g03286(new_n3662, new_n3610, new_n3663);
xnor_1 g03287(new_n3662, new_n3609, new_n3664);
not_4  g03288(new_n3625, new_n3665);
xnor_1 g03289(new_n3628, new_n3665, new_n3666);
not_4  g03290(new_n3666, new_n3667);
nand_1 g03291(n9400, n3719, new_n3668);
nand_1 g03292(n6877, n3602, new_n3669);
xnor_1 g03293(new_n3669, new_n3668, new_n3670);
not_4  g03294(new_n3670, new_n3671);
nand_1 g03295(new_n3671, new_n3667, new_n3672);
nand_1 g03296(new_n3613, new_n3611, new_n3673);
nand_1 g03297(new_n3673, new_n3615, new_n3674);
not_4  g03298(new_n3674, new_n3675);
nand_1 g03299(new_n3675, new_n3517, new_n3676);
not_4  g03300(new_n3676, new_n3677_1);
xnor_1 g03301(new_n3671, new_n3666, new_n3678);
nand_1 g03302(new_n3678, new_n3677_1, new_n3679);
nand_1 g03303(new_n3679, new_n3672, new_n3680);
nand_1 g03304(new_n3680, new_n3664, new_n3681);
nand_1 g03305(new_n3681, new_n3663, new_n3682);
nor_1  g03306(new_n3682, new_n3606, new_n3683);
nand_1 g03307(n7610, n4805, new_n3684);
nand_1 g03308(new_n3652, new_n3647, new_n3685);
nand_1 g03309(new_n3685, new_n3656, new_n3686);
xnor_1 g03310(new_n3686, new_n3684, new_n3687);
not_4  g03311(new_n3687, new_n3688);
nand_1 g03312(n7733, n5283, new_n3689);
nand_1 g03313(n12925, n137, new_n3690);
nand_1 g03314(n11478, n4826, new_n3691);
not_4  g03315(new_n3691, new_n3692);
xnor_1 g03316(new_n3692, new_n3690, new_n3693);
xnor_1 g03317(new_n3693, new_n3689, new_n3694);
xnor_1 g03318(new_n3694, new_n3688, new_n3695);
nor_1  g03319(new_n3658, new_n3621, new_n3696);
xnor_1 g03320(new_n3696, new_n3695, new_n3697);
nand_1 g03321(n7236, n217, new_n3698);
nand_1 g03322(new_n3639, new_n3631, new_n3699);
nand_1 g03323(new_n3699, new_n3635, new_n3700);
not_4  g03324(new_n3700, new_n3701);
xnor_1 g03325(new_n3701, new_n3698, new_n3702);
nand_1 g03326(n8384, n405, new_n3703);
nand_1 g03327(n8433, n6358, new_n3704);
nand_1 g03328(n4086, n3992, new_n3705);
not_4  g03329(new_n3705, new_n3706);
xnor_1 g03330(new_n3706, new_n3704, new_n3707);
xnor_1 g03331(new_n3707, new_n3703, new_n3708);
xnor_1 g03332(new_n3708, new_n3702, new_n3709);
nor_1  g03333(new_n3641, new_n3631, new_n3710);
xnor_1 g03334(new_n3710, new_n3709, new_n3711);
xnor_1 g03335(new_n3711, new_n3697, new_n3712);
nand_1 g03336(new_n3643, new_n3630, new_n3713);
nand_1 g03337(new_n3661_1, new_n3645, new_n3714);
nand_1 g03338(new_n3714, new_n3713, new_n3715);
xnor_1 g03339(new_n3715, new_n3712, new_n3716);
not_4  g03340(new_n3683, new_n3717);
nand_1 g03341(new_n3682, new_n3606, new_n3718);
nand_1 g03342(new_n3718, new_n3717, new_n3719_1);
nor_1  g03343(new_n3719_1, new_n3716, new_n3720);
nor_1  g03344(new_n3720, new_n3683, new_n3721);
not_4  g03345(new_n3721, new_n3722);
nand_1 g03346(new_n3722, new_n3604, new_n3723);
nand_1 g03347(new_n3721, new_n3603, new_n3724);
not_4  g03348(new_n3709, new_n3725);
nand_1 g03349(new_n3710, new_n3725, new_n3726);
nand_1 g03350(n7236, n6611, new_n3727);
nand_1 g03351(n3992, n217, new_n3728);
nand_1 g03352(new_n3705, new_n3704, new_n3729);
nand_1 g03353(new_n3707, new_n3703, new_n3730);
nand_1 g03354(new_n3730, new_n3729, new_n3731);
not_4  g03355(new_n3731, new_n3732);
xnor_1 g03356(new_n3732, new_n3728, new_n3733);
nand_1 g03357(n6358, n405, new_n3734);
nand_1 g03358(n8384, n4086, new_n3735);
nand_1 g03359(n8433, n5198, new_n3736);
not_4  g03360(new_n3736, new_n3737);
xnor_1 g03361(new_n3737, new_n3735, new_n3738);
not_4  g03362(new_n3738, new_n3739);
xnor_1 g03363(new_n3739, new_n3734, new_n3740);
xnor_1 g03364(new_n3740, new_n3733, new_n3741);
xnor_1 g03365(new_n3741, new_n3727, new_n3742);
nor_1  g03366(new_n3700, new_n3698, new_n3743);
not_4  g03367(new_n3743, new_n3744);
nand_1 g03368(new_n3708, new_n3702, new_n3745);
nand_1 g03369(new_n3745, new_n3744, new_n3746);
xnor_1 g03370(new_n3746, new_n3742, new_n3747);
not_4  g03371(new_n3747, new_n3748);
xnor_1 g03372(new_n3748, new_n3726, new_n3749);
nand_1 g03373(new_n3696, new_n3695, new_n3750);
nand_1 g03374(n4970, n4805, new_n3751);
nand_1 g03375(n11478, n7610, new_n3752);
nand_1 g03376(new_n3691, new_n3690, new_n3753);
nand_1 g03377(new_n3693, new_n3689, new_n3754_1);
nand_1 g03378(new_n3754_1, new_n3753, new_n3755);
not_4  g03379(new_n3755, new_n3756);
xnor_1 g03380(new_n3756, new_n3752, new_n3757);
nand_1 g03381(n7733, n137, new_n3758);
nand_1 g03382(n5283, n4826, new_n3759);
nand_1 g03383(n12925, n6294, new_n3760);
not_4  g03384(new_n3760, new_n3761);
xnor_1 g03385(new_n3761, new_n3759, new_n3762);
not_4  g03386(new_n3762, new_n3763);
xnor_1 g03387(new_n3763, new_n3758, new_n3764);
xnor_1 g03388(new_n3764, new_n3757, new_n3765);
xnor_1 g03389(new_n3765, new_n3751, new_n3766);
not_4  g03390(new_n3684, new_n3767);
nand_1 g03391(new_n3686, new_n3767, new_n3768);
nand_1 g03392(new_n3694, new_n3687, new_n3769);
nand_1 g03393(new_n3769, new_n3768, new_n3770);
not_4  g03394(new_n3770, new_n3771);
xnor_1 g03395(new_n3771, new_n3766, new_n3772);
xnor_1 g03396(new_n3772, new_n3750, new_n3773);
not_4  g03397(new_n3711, new_n3774);
nand_1 g03398(new_n3774, new_n3697, new_n3775);
nand_1 g03399(new_n3715, new_n3712, new_n3776);
nand_1 g03400(new_n3776, new_n3775, new_n3777);
xnor_1 g03401(new_n3777, new_n3773, new_n3778);
xnor_1 g03402(new_n3778, new_n3749, new_n3779);
nand_1 g03403(new_n3779, new_n3724, new_n3780);
nand_1 g03404(new_n3780, new_n3723, new_n3781);
nand_1 g03405(new_n3781, new_n3602_1, new_n3782);
nor_1  g03406(new_n3781, new_n3602_1, new_n3783);
not_4  g03407(new_n3783, new_n3784);
nand_1 g03408(new_n3784, new_n3782, new_n3785);
not_4  g03409(new_n3726, new_n3786);
nand_1 g03410(new_n3748, new_n3786, new_n3787);
not_4  g03411(new_n3787, new_n3788);
nand_1 g03412(n7236, n6359, new_n3789);
not_4  g03413(new_n3789, new_n3790);
nand_1 g03414(n6358, n4086, new_n3791);
nand_1 g03415(new_n3736, new_n3735, new_n3792);
nand_1 g03416(new_n3738, new_n3734, new_n3793);
nand_1 g03417(new_n3793, new_n3792, new_n3794);
not_4  g03418(new_n3794, new_n3795);
xnor_1 g03419(new_n3795, new_n3791, new_n3796);
nand_1 g03420(n5198, n405, new_n3797);
nand_1 g03421(n8433, n1471, new_n3798);
not_4  g03422(new_n3798, new_n3799);
xnor_1 g03423(new_n3799, new_n3797, new_n3800);
xnor_1 g03424(new_n3800, new_n3796, new_n3801);
nand_1 g03425(n8384, n217, new_n3802);
nand_1 g03426(n6611, n3992, new_n3803);
not_4  g03427(new_n3803, new_n3804);
xnor_1 g03428(new_n3804, new_n3802, new_n3805);
xnor_1 g03429(new_n3805, new_n3801, new_n3806);
nor_1  g03430(new_n3731, new_n3728, new_n3807);
not_4  g03431(new_n3733, new_n3808);
nor_1  g03432(new_n3740, new_n3808, new_n3809);
nor_1  g03433(new_n3809, new_n3807, new_n3810);
xnor_1 g03434(new_n3810, new_n3806, new_n3811);
not_4  g03435(new_n3727, new_n3812);
nand_1 g03436(new_n3741, new_n3812, new_n3813);
nand_1 g03437(new_n3746, new_n3742, new_n3814);
nand_1 g03438(new_n3814, new_n3813, new_n3815);
nand_1 g03439(new_n3815, new_n3811, new_n3816);
not_4  g03440(new_n3816, new_n3817);
nor_1  g03441(new_n3815, new_n3811, new_n3818);
nor_1  g03442(new_n3818, new_n3817, new_n3819);
nand_1 g03443(new_n3819, new_n3790, new_n3820);
nor_1  g03444(new_n3819, new_n3790, new_n3821);
not_4  g03445(new_n3821, new_n3822);
nand_1 g03446(new_n3822, new_n3820, new_n3823);
nand_1 g03447(new_n3823, new_n3788, new_n3824);
not_4  g03448(new_n3823, new_n3825);
nand_1 g03449(new_n3825, new_n3787, new_n3826);
nand_1 g03450(new_n3826, new_n3824, new_n3827);
not_4  g03451(new_n3750, new_n3828);
nand_1 g03452(new_n3772, new_n3828, new_n3829);
nand_1 g03453(n4805, n503, new_n3830);
nand_1 g03454(n4826, n137, new_n3831);
not_4  g03455(new_n3831, new_n3832);
nand_1 g03456(n7733, n6294, new_n3833);
nand_1 g03457(n12925, n6797, new_n3834);
not_4  g03458(new_n3834, new_n3835);
xnor_1 g03459(new_n3835, new_n3833, new_n3836);
xnor_1 g03460(new_n3836, new_n3832, new_n3837);
nand_1 g03461(new_n3760, new_n3759, new_n3838);
nand_1 g03462(new_n3762, new_n3758, new_n3839);
nand_1 g03463(new_n3839, new_n3838, new_n3840);
nor_1  g03464(new_n3840, new_n3837, new_n3841);
not_4  g03465(new_n3841, new_n3842_1);
nand_1 g03466(new_n3840, new_n3837, new_n3843);
nand_1 g03467(new_n3843, new_n3842_1, new_n3844);
not_4  g03468(new_n3844, new_n3845);
nand_1 g03469(n11478, n4970, new_n3846);
nand_1 g03470(n7610, n5283, new_n3847);
nand_1 g03471(new_n3847, new_n3846, new_n3848);
not_4  g03472(new_n3846, new_n3849_1);
not_4  g03473(new_n3847, new_n3850);
nand_1 g03474(new_n3850, new_n3849_1, new_n3851);
nand_1 g03475(new_n3851, new_n3848, new_n3852);
not_4  g03476(new_n3852, new_n3853);
nand_1 g03477(new_n3853, new_n3845, new_n3854);
nand_1 g03478(new_n3852, new_n3844, new_n3855);
nand_1 g03479(new_n3855, new_n3854, new_n3856);
nor_1  g03480(new_n3755, new_n3752, new_n3857);
not_4  g03481(new_n3757, new_n3858);
nor_1  g03482(new_n3764, new_n3858, new_n3859);
nor_1  g03483(new_n3859, new_n3857, new_n3860);
nor_1  g03484(new_n3860, new_n3856, new_n3861);
not_4  g03485(new_n3861, new_n3862);
nand_1 g03486(new_n3860, new_n3856, new_n3863);
nand_1 g03487(new_n3863, new_n3862, new_n3864);
not_4  g03488(new_n3751, new_n3865_1);
nand_1 g03489(new_n3765, new_n3865_1, new_n3866);
nand_1 g03490(new_n3770, new_n3766, new_n3867);
nand_1 g03491(new_n3867, new_n3866, new_n3868);
xnor_1 g03492(new_n3868, new_n3864, new_n3869);
xnor_1 g03493(new_n3869, new_n3830, new_n3870);
not_4  g03494(new_n3870, new_n3871);
xnor_1 g03495(new_n3871, new_n3829, new_n3872);
xnor_1 g03496(new_n3872, new_n3827, new_n3873);
not_4  g03497(new_n3773, new_n3874);
nand_1 g03498(new_n3777, new_n3874, new_n3875);
not_4  g03499(new_n3749, new_n3876);
nand_1 g03500(new_n3778, new_n3876, new_n3877);
nand_1 g03501(new_n3877, new_n3875, new_n3878);
xnor_1 g03502(new_n3878, new_n3873, new_n3879);
not_4  g03503(new_n3879, new_n3880);
nor_1  g03504(new_n3880, new_n3785, new_n3881);
not_4  g03505(new_n3881, new_n3882);
nand_1 g03506(new_n3880, new_n3785, new_n3883);
nand_1 g03507(new_n3883, new_n3882, new_n3884);
nand_1 g03508(new_n3884, new_n3511, new_n3885);
nor_1  g03509(new_n3884, new_n3511, new_n3886);
not_4  g03510(new_n3886, new_n3887);
xnor_1 g03511(new_n3503, new_n3500, new_n3888);
not_4  g03512(new_n3888, new_n3889);
nand_1 g03513(new_n3724, new_n3723, new_n3890);
xnor_1 g03514(new_n3890, new_n3779, new_n3891);
nor_1  g03515(new_n3891, new_n3889, new_n3892);
xnor_1 g03516(new_n3499, new_n3491, new_n3893);
not_4  g03517(new_n3716, new_n3894);
xnor_1 g03518(new_n3719_1, new_n3894, new_n3895);
nor_1  g03519(new_n3895, new_n3893, new_n3896);
xnor_1 g03520(new_n3680, new_n3664, new_n3897);
nand_1 g03521(n9956, n7862, new_n3898);
nand_1 g03522(new_n3898, new_n3435, new_n3899);
nand_1 g03523(new_n3899, new_n3492, new_n3900);
not_4  g03524(new_n3899, new_n3901);
nand_1 g03525(new_n3901, new_n3433, new_n3902);
nand_1 g03526(new_n3902, new_n3900, new_n3903);
nand_1 g03527(new_n3903, new_n3897, new_n3904);
xnor_1 g03528(new_n3903, new_n3897, new_n3905);
not_4  g03529(new_n3898, new_n3906);
xnor_1 g03530(new_n3675, new_n3516, new_n3907);
nand_1 g03531(new_n3907, new_n3906, new_n3908);
nand_1 g03532(new_n3496, new_n3494, new_n3909);
nand_1 g03533(new_n3909, new_n3498, new_n3910);
nand_1 g03534(new_n3910, new_n3908, new_n3911);
xnor_1 g03535(new_n3678, new_n3676, new_n3912);
xnor_1 g03536(new_n3910, new_n3908, new_n3913);
nor_1  g03537(new_n3913, new_n3912, new_n3914);
not_4  g03538(new_n3914, new_n3915);
nand_1 g03539(new_n3915, new_n3911, new_n3916);
not_4  g03540(new_n3916, new_n3917);
nor_1  g03541(new_n3917, new_n3905, new_n3918);
not_4  g03542(new_n3918, new_n3919);
nand_1 g03543(new_n3919, new_n3904, new_n3920);
xnor_1 g03544(new_n3895, new_n3893, new_n3921);
nor_1  g03545(new_n3921, new_n3920, new_n3922);
nor_1  g03546(new_n3922, new_n3896, new_n3923);
not_4  g03547(new_n3892, new_n3924);
nand_1 g03548(new_n3891, new_n3889, new_n3925);
nand_1 g03549(new_n3925, new_n3924, new_n3926);
nor_1  g03550(new_n3926, new_n3923, new_n3927);
nor_1  g03551(new_n3927, new_n3892, new_n3928);
nand_1 g03552(new_n3928, new_n3887, new_n3929);
nand_1 g03553(new_n3929, new_n3885, new_n3930);
nand_1 g03554(new_n3930, new_n3509, new_n3931);
not_4  g03555(new_n3509, new_n3932_1);
not_4  g03556(new_n3930, new_n3933);
nand_1 g03557(new_n3933, new_n3932_1, new_n3934);
nand_1 g03558(new_n3934, new_n3931, new_n3935);
not_4  g03559(new_n3594, new_n3936);
nand_1 g03560(new_n3598, new_n3936, new_n3937);
nand_1 g03561(n9400, n8065, new_n3938);
not_4  g03562(new_n3938, new_n3939);
nand_1 g03563(n10439, n2464, new_n3940);
nand_1 g03564(n10391, n6877, new_n3941);
not_4  g03565(new_n3941, new_n3942);
xnor_1 g03566(new_n3942, new_n3940, new_n3943);
not_4  g03567(new_n3943, new_n3944);
nand_1 g03568(new_n3944, new_n3939, new_n3945);
nand_1 g03569(new_n3943, new_n3938, new_n3946);
nand_1 g03570(new_n3946, new_n3945, new_n3947);
not_4  g03571(new_n3947, new_n3948);
nand_1 g03572(new_n3575, new_n3571, new_n3949);
nand_1 g03573(new_n3581, new_n3949, new_n3950);
xnor_1 g03574(new_n3950, new_n3948, new_n3951);
not_4  g03575(new_n3572, new_n3952);
nand_1 g03576(new_n3574, new_n3952, new_n3953);
not_4  g03577(new_n3953, new_n3954);
nand_1 g03578(n11311, n8595, new_n3955);
not_4  g03579(new_n3955, new_n3956);
nand_1 g03580(new_n3956, new_n3954, new_n3957);
nand_1 g03581(new_n3955, new_n3953, new_n3958);
nand_1 g03582(new_n3958, new_n3957, new_n3959);
nand_1 g03583(n4203, n3602, new_n3960);
nand_1 g03584(n6126, n4187, new_n3961);
nand_1 g03585(n12753, n3719, new_n3962);
not_4  g03586(new_n3962, new_n3963);
xnor_1 g03587(new_n3963, new_n3961, new_n3964);
xnor_1 g03588(new_n3964, new_n3960, new_n3965);
xnor_1 g03589(new_n3965, new_n3959, new_n3966);
xnor_1 g03590(new_n3966, new_n3951, new_n3967);
not_4  g03591(new_n3583, new_n3968);
nand_1 g03592(new_n3587, new_n3968, new_n3969);
nor_1  g03593(new_n3585, new_n3584, new_n3970);
nand_1 g03594(new_n3593, new_n3588, new_n3971);
not_4  g03595(new_n3971, new_n3972);
xnor_1 g03596(new_n3972, new_n3970, new_n3973);
nand_1 g03597(new_n3973, new_n3969, new_n3974);
xnor_1 g03598(new_n3974, new_n3967, new_n3975);
xnor_1 g03599(new_n3975, new_n3937, new_n3976);
nor_1  g03600(new_n3599, new_n3569, new_n3977);
nor_1  g03601(new_n3600, new_n3567, new_n3978);
nor_1  g03602(new_n3978, new_n3977, new_n3979);
xnor_1 g03603(new_n3979, new_n3976, new_n3980);
not_4  g03604(new_n3980, new_n3981);
not_4  g03605(new_n3864, new_n3982);
nand_1 g03606(new_n3868, new_n3982, new_n3983);
nand_1 g03607(n10965, n4805, new_n3984);
nand_1 g03608(n5283, n4970, new_n3985);
nand_1 g03609(n11478, n503, new_n3986_1);
not_4  g03610(new_n3986_1, new_n3987);
xnor_1 g03611(new_n3987, new_n3985, new_n3988);
xnor_1 g03612(new_n3988, new_n3984, new_n3989);
not_4  g03613(new_n3989, new_n3990);
nand_1 g03614(new_n3836, new_n3832, new_n3991);
nand_1 g03615(new_n3842_1, new_n3991, new_n3992_1);
xnor_1 g03616(new_n3992_1, new_n3990, new_n3993);
not_4  g03617(new_n3833, new_n3994);
nand_1 g03618(new_n3835, new_n3994, new_n3995);
nand_1 g03619(n7610, n137, new_n3996);
nand_1 g03620(new_n3996, new_n3995, new_n3997);
not_4  g03621(new_n3995, new_n3998);
not_4  g03622(new_n3996, new_n3999);
nand_1 g03623(new_n3999, new_n3998, new_n4000);
nand_1 g03624(new_n4000, new_n3997, new_n4001);
nand_1 g03625(n7733, n6797, new_n4002);
nand_1 g03626(n6294, n4826, new_n4003);
nand_1 g03627(n12925, n3146, new_n4004);
nand_1 g03628(new_n4004, new_n4003, new_n4005_1);
not_4  g03629(new_n4003, new_n4006);
not_4  g03630(new_n4004, new_n4007);
nand_1 g03631(new_n4007, new_n4006, new_n4008);
nand_1 g03632(new_n4008, new_n4005_1, new_n4009);
xnor_1 g03633(new_n4009, new_n4002, new_n4010);
not_4  g03634(new_n4010, new_n4011);
xnor_1 g03635(new_n4011, new_n4001, new_n4012);
xnor_1 g03636(new_n4012, new_n3993, new_n4013);
not_4  g03637(new_n4013, new_n4014);
not_4  g03638(new_n3854, new_n4015);
xnor_1 g03639(new_n3861, new_n3851, new_n4016);
nor_1  g03640(new_n4016, new_n4015, new_n4017);
xnor_1 g03641(new_n4017, new_n4014, new_n4018);
xnor_1 g03642(new_n4018, new_n3983, new_n4019);
not_4  g03643(new_n3830, new_n4020);
nor_1  g03644(new_n3869, new_n4020, new_n4021);
not_4  g03645(new_n4021, new_n4022);
nand_1 g03646(new_n3870, new_n3829, new_n4023);
nand_1 g03647(new_n4023, new_n4022, new_n4024);
not_4  g03648(new_n4024, new_n4025);
xnor_1 g03649(new_n4025, new_n4019, new_n4026);
nand_1 g03650(n11296, n7236, new_n4027);
nand_1 g03651(n8384, n6611, new_n4028);
nand_1 g03652(n6359, n3992, new_n4029);
not_4  g03653(new_n4029, new_n4030);
xnor_1 g03654(new_n4030, new_n4028, new_n4031);
xnor_1 g03655(new_n4031, new_n4027, new_n4032);
not_4  g03656(new_n3791, new_n4033);
nand_1 g03657(new_n3795, new_n4033, new_n4034);
nand_1 g03658(new_n3800, new_n3796, new_n4035);
nand_1 g03659(new_n4035, new_n4034, new_n4036);
xnor_1 g03660(new_n4036, new_n4032, new_n4037);
nor_1  g03661(new_n3798, new_n3797, new_n4038);
nand_1 g03662(n6358, n217, new_n4039);
xnor_1 g03663(new_n4039, new_n4038, new_n4040);
nand_1 g03664(n1471, n405, new_n4041);
nand_1 g03665(n5198, n4086, new_n4042);
nand_1 g03666(n8433, n7646, new_n4043);
nand_1 g03667(new_n4043, new_n4042, new_n4044);
not_4  g03668(new_n4042, new_n4045);
not_4  g03669(new_n4043, new_n4046);
nand_1 g03670(new_n4046, new_n4045, new_n4047);
nand_1 g03671(new_n4047, new_n4044, new_n4048);
xnor_1 g03672(new_n4048, new_n4041, new_n4049);
xnor_1 g03673(new_n4049, new_n4040, new_n4050);
xnor_1 g03674(new_n4050, new_n4037, new_n4051);
not_4  g03675(new_n4051, new_n4052);
not_4  g03676(new_n3801, new_n4053);
nand_1 g03677(new_n3805, new_n4053, new_n4054);
nor_1  g03678(new_n3803, new_n3802, new_n4055);
not_4  g03679(new_n3810, new_n4056);
nand_1 g03680(new_n4056, new_n3806, new_n4057);
not_4  g03681(new_n4057, new_n4058);
xnor_1 g03682(new_n4058, new_n4055, new_n4059);
nand_1 g03683(new_n4059, new_n4054, new_n4060);
xnor_1 g03684(new_n4060, new_n4052, new_n4061);
xnor_1 g03685(new_n4061, new_n3816, new_n4062);
nand_1 g03686(new_n3826, new_n3822, new_n4063);
xnor_1 g03687(new_n4063, new_n4062, new_n4064);
xnor_1 g03688(new_n4064, new_n4026, new_n4065);
not_4  g03689(new_n3827, new_n4066);
nand_1 g03690(new_n3872, new_n4066, new_n4067);
nand_1 g03691(new_n3878, new_n3873, new_n4068);
nand_1 g03692(new_n4068, new_n4067, new_n4069);
xnor_1 g03693(new_n4069, new_n4065, new_n4070);
nand_1 g03694(new_n4070, new_n3981, new_n4071);
nor_1  g03695(new_n4070, new_n3981, new_n4072);
not_4  g03696(new_n4072, new_n4073);
nand_1 g03697(new_n4073, new_n4071, new_n4074);
not_4  g03698(new_n4074, new_n4075);
nand_1 g03699(new_n3882, new_n3784, new_n4076);
not_4  g03700(new_n4076, new_n4077);
nand_1 g03701(new_n4077, new_n4075, new_n4078);
nand_1 g03702(new_n4076, new_n4074, new_n4079);
nand_1 g03703(new_n4079, new_n4078, new_n4080);
xnor_1 g03704(new_n4080, new_n3935, n844);
nand_1 g03705(n7456, n6687, new_n4082);
nand_1 g03706(n12591, n6687, new_n4083);
nand_1 g03707(n4189, n1798, new_n4084);
nand_1 g03708(new_n4084, new_n4083, new_n4085);
nand_1 g03709(n6687, n1798, new_n4086_1);
not_4  g03710(new_n4086_1, new_n4087);
nand_1 g03711(n12591, n4189, new_n4088_1);
not_4  g03712(new_n4088_1, new_n4089);
nand_1 g03713(new_n4089, new_n4087, new_n4090);
nand_1 g03714(n3932, n2564, new_n4091);
nand_1 g03715(new_n4091, new_n4090, new_n4092);
nand_1 g03716(new_n4092, new_n4085, new_n4093);
xnor_1 g03717(new_n4093, new_n4082, new_n4094_1);
nand_1 g03718(n4189, n3932, new_n4095);
nand_1 g03719(n12591, n2564, new_n4096);
nand_1 g03720(n6770, n1798, new_n4097);
nand_1 g03721(new_n4097, new_n4096, new_n4098);
nor_1  g03722(new_n4097, new_n4096, new_n4099);
not_4  g03723(new_n4099, new_n4100);
nand_1 g03724(new_n4100, new_n4098, new_n4101);
xnor_1 g03725(new_n4101, new_n4095, new_n4102);
nor_1  g03726(new_n4102, new_n4094_1, new_n4103);
not_4  g03727(new_n4103, new_n4104);
nand_1 g03728(new_n4102, new_n4094_1, new_n4105);
nand_1 g03729(new_n4105, new_n4104, new_n4106);
not_4  g03730(new_n4106, new_n4107);
not_4  g03731(new_n4091, new_n4108);
nand_1 g03732(new_n4108, new_n4086_1, new_n4109);
nand_1 g03733(new_n4090, new_n4085, new_n4110);
nand_1 g03734(new_n4110, new_n4109, new_n4111);
not_4  g03735(new_n4111, new_n4112);
nand_1 g03736(new_n4112, new_n4108, new_n4113);
not_4  g03737(new_n4113, new_n4114);
nand_1 g03738(new_n4114, new_n4107, new_n4115);
nand_1 g03739(new_n4113, new_n4106, new_n4116);
nand_1 g03740(new_n4116, new_n4115, new_n4117);
not_4  g03741(new_n4109, new_n4118);
nand_1 g03742(new_n4118, new_n4085, new_n4119);
nand_1 g03743(new_n4119, new_n4111, new_n4120);
nand_1 g03744(n8336, n6703, new_n4121);
not_4  g03745(new_n4121, new_n4122);
nand_1 g03746(n11876, n11222, new_n4123);
not_4  g03747(new_n4123, new_n4124);
nand_1 g03748(n12069, n5645, new_n4125);
not_4  g03749(new_n4125, new_n4126);
nand_1 g03750(new_n4126, new_n4124, new_n4127);
nand_1 g03751(new_n4125, new_n4123, new_n4128);
nand_1 g03752(new_n4128, new_n4127, new_n4129);
not_4  g03753(new_n4129, new_n4130);
nand_1 g03754(new_n4130, new_n4122, new_n4131);
not_4  g03755(new_n4131, new_n4132);
nand_1 g03756(n9640, n8336, new_n4133);
nand_1 g03757(n10928, n6703, new_n4134);
xnor_1 g03758(new_n4134, new_n4133, new_n4135);
not_4  g03759(new_n4135, new_n4136);
nand_1 g03760(new_n4136, new_n4132, new_n4137);
nand_1 g03761(n12391, n5645, new_n4138);
nand_1 g03762(n12069, n1067, new_n4139);
not_4  g03763(new_n4139, new_n4140);
xnor_1 g03764(new_n4140, new_n4138, new_n4141_1);
xnor_1 g03765(new_n4141_1, new_n4127, new_n4142);
nand_1 g03766(n11222, n10898, new_n4143);
nand_1 g03767(n11876, n11153, new_n4144);
xnor_1 g03768(new_n4144, new_n4143, new_n4145);
xnor_1 g03769(new_n4145, new_n4142, new_n4146);
xnor_1 g03770(new_n4136, new_n4131, new_n4147);
nand_1 g03771(new_n4147, new_n4146, new_n4148);
nand_1 g03772(new_n4148, new_n4137, new_n4149);
not_4  g03773(new_n4149, new_n4150);
nand_1 g03774(n10928, n9640, new_n4151);
not_4  g03775(new_n4151, new_n4152);
nand_1 g03776(new_n4152, new_n4121, new_n4153);
nand_1 g03777(n6986, n6703, new_n4154);
nand_1 g03778(n8336, n3022, new_n4155_1);
nand_1 g03779(new_n4155_1, new_n4154, new_n4156);
nand_1 g03780(n6986, n3022, new_n4157);
not_4  g03781(new_n4157, new_n4158);
nand_1 g03782(new_n4158, new_n4122, new_n4159_1);
nand_1 g03783(new_n4159_1, new_n4156, new_n4160);
nand_1 g03784(new_n4160, new_n4153, new_n4161);
not_4  g03785(new_n4161, new_n4162);
not_4  g03786(new_n4156, new_n4163);
nor_1  g03787(new_n4163, new_n4153, new_n4164);
nor_1  g03788(new_n4164, new_n4162, new_n4165);
xnor_1 g03789(new_n4165, new_n4150, new_n4166);
not_4  g03790(new_n4138, new_n4167);
nand_1 g03791(new_n4140, new_n4167, new_n4168);
not_4  g03792(new_n4168, new_n4169);
nand_1 g03793(n12069, n8665, new_n4170);
nand_1 g03794(n12391, n1067, new_n4171);
nand_1 g03795(n7891, n5645, new_n4172);
not_4  g03796(new_n4172, new_n4173);
xnor_1 g03797(new_n4173, new_n4171, new_n4174);
xnor_1 g03798(new_n4174, new_n4170, new_n4175);
not_4  g03799(new_n4175, new_n4176);
xnor_1 g03800(new_n4176, new_n4169, new_n4177);
not_4  g03801(new_n4127, new_n4178);
nor_1  g03802(new_n4141_1, new_n4178, new_n4179);
not_4  g03803(new_n4179, new_n4180);
nand_1 g03804(new_n4145, new_n4142, new_n4181);
nand_1 g03805(new_n4181, new_n4180, new_n4182);
nand_1 g03806(n11153, n10898, new_n4183);
not_4  g03807(new_n4183, new_n4184);
nand_1 g03808(new_n4184, new_n4123, new_n4185);
nand_1 g03809(n11876, n5314, new_n4186);
nand_1 g03810(n11222, n3754, new_n4187_1);
nand_1 g03811(new_n4187_1, new_n4186, new_n4188);
not_4  g03812(new_n4188, new_n4189_1);
nand_1 g03813(new_n4189_1, new_n4185, new_n4190_1);
nand_1 g03814(n5314, n3754, new_n4191);
not_4  g03815(new_n4191, new_n4192);
nand_1 g03816(new_n4192, new_n4124, new_n4193);
nand_1 g03817(new_n4193, new_n4190_1, new_n4194);
nor_1  g03818(new_n4189_1, new_n4185, new_n4195);
nor_1  g03819(new_n4195, new_n4194, new_n4196);
xnor_1 g03820(new_n4196, new_n4182, new_n4197);
xnor_1 g03821(new_n4197, new_n4177, new_n4198);
xnor_1 g03822(new_n4198, new_n4166, new_n4199);
not_4  g03823(new_n4199, new_n4200);
nor_1  g03824(new_n4200, new_n4120, new_n4201);
not_4  g03825(new_n4201, new_n4202);
xnor_1 g03826(new_n4130, new_n4121, new_n4203_1);
nand_1 g03827(new_n4203_1, new_n4087, new_n4204);
nand_1 g03828(n2564, n1798, new_n4205);
nand_1 g03829(n6687, n3932, new_n4206);
xnor_1 g03830(new_n4206, new_n4205, new_n4207);
nand_1 g03831(new_n4207, new_n4204, new_n4208);
xnor_1 g03832(new_n4147, new_n4146, new_n4209);
not_4  g03833(new_n4209, new_n4210);
xnor_1 g03834(new_n4207, new_n4204, new_n4211);
nor_1  g03835(new_n4211, new_n4210, new_n4212);
not_4  g03836(new_n4212, new_n4213);
nand_1 g03837(new_n4213, new_n4208, new_n4214);
not_4  g03838(new_n4214, new_n4215);
xnor_1 g03839(new_n4199, new_n4120, new_n4216);
nand_1 g03840(new_n4216, new_n4215, new_n4217);
nand_1 g03841(new_n4217, new_n4202, new_n4218);
xnor_1 g03842(new_n4218, new_n4117, new_n4219);
nand_1 g03843(new_n4175, new_n4169, new_n4220);
not_4  g03844(new_n4220, new_n4221);
nand_1 g03845(n12069, n11922, new_n4222);
nand_1 g03846(new_n4172, new_n4171, new_n4223);
nand_1 g03847(new_n4174, new_n4170, new_n4224);
nand_1 g03848(new_n4224, new_n4223, new_n4225);
not_4  g03849(new_n4225, new_n4226_1);
xnor_1 g03850(new_n4226_1, new_n4222, new_n4227);
nand_1 g03851(n7160, n5645, new_n4228);
nand_1 g03852(n7891, n1067, new_n4229);
nand_1 g03853(n12391, n8665, new_n4230_1);
not_4  g03854(new_n4230_1, new_n4231);
xnor_1 g03855(new_n4231, new_n4229, new_n4232);
nor_1  g03856(new_n4232, new_n4228, new_n4233);
nand_1 g03857(new_n4232, new_n4228, new_n4234);
not_4  g03858(new_n4234, new_n4235);
nor_1  g03859(new_n4235, new_n4233, new_n4236);
xnor_1 g03860(new_n4236, new_n4227, new_n4237);
xnor_1 g03861(new_n4237, new_n4221, new_n4238);
nand_1 g03862(n11222, n2749, new_n4239);
nand_1 g03863(new_n4193, new_n4183, new_n4240);
nand_1 g03864(new_n4240, new_n4188, new_n4241);
not_4  g03865(new_n4241, new_n4242);
xnor_1 g03866(new_n4242, new_n4239, new_n4243);
nand_1 g03867(n10898, n5314, new_n4244);
nand_1 g03868(n11153, n3754, new_n4245);
nand_1 g03869(n11876, n996, new_n4246);
not_4  g03870(new_n4246, new_n4247);
xnor_1 g03871(new_n4247, new_n4245, new_n4248);
not_4  g03872(new_n4248, new_n4249);
xnor_1 g03873(new_n4249, new_n4244, new_n4250);
xnor_1 g03874(new_n4250, new_n4243, new_n4251);
nand_1 g03875(new_n4194, new_n4184, new_n4252);
xnor_1 g03876(new_n4252, new_n4251, new_n4253);
xnor_1 g03877(new_n4253, new_n4238, new_n4254);
not_4  g03878(new_n4196, new_n4255);
nand_1 g03879(new_n4255, new_n4182, new_n4256);
not_4  g03880(new_n4177, new_n4257);
nand_1 g03881(new_n4197, new_n4257, new_n4258);
nand_1 g03882(new_n4258, new_n4256, new_n4259);
xnor_1 g03883(new_n4259, new_n4254, new_n4260);
not_4  g03884(new_n4260, new_n4261);
nand_1 g03885(n11023, n8336, new_n4262);
nand_1 g03886(new_n4159_1, new_n4151, new_n4263);
nand_1 g03887(new_n4263, new_n4156, new_n4264);
nor_1  g03888(new_n4264, new_n4262, new_n4265);
not_4  g03889(new_n4265, new_n4266);
nand_1 g03890(new_n4264, new_n4262, new_n4267);
nand_1 g03891(new_n4267, new_n4266, new_n4268);
nand_1 g03892(n9640, n6986, new_n4269);
not_4  g03893(new_n4269, new_n4270);
nand_1 g03894(n10928, n3022, new_n4271);
nand_1 g03895(n6703, n2226, new_n4272);
nand_1 g03896(new_n4272, new_n4271, new_n4273);
not_4  g03897(new_n4271, new_n4274);
not_4  g03898(new_n4272, new_n4275);
nand_1 g03899(new_n4275, new_n4274, new_n4276);
nand_1 g03900(new_n4276, new_n4273, new_n4277);
xnor_1 g03901(new_n4277, new_n4270, new_n4278);
xnor_1 g03902(new_n4278, new_n4268, new_n4279);
nand_1 g03903(new_n4162, new_n4152, new_n4280);
xnor_1 g03904(new_n4280, new_n4279, new_n4281);
not_4  g03905(new_n4281, new_n4282);
not_4  g03906(new_n4165, new_n4283);
nand_1 g03907(new_n4283, new_n4150, new_n4284);
nand_1 g03908(new_n4198, new_n4166, new_n4285);
nand_1 g03909(new_n4285, new_n4284, new_n4286);
nor_1  g03910(new_n4286, new_n4282, new_n4287);
not_4  g03911(new_n4287, new_n4288);
nand_1 g03912(new_n4286, new_n4282, new_n4289);
nand_1 g03913(new_n4289, new_n4288, new_n4290);
nand_1 g03914(new_n4290, new_n4261, new_n4291);
not_4  g03915(new_n4290, new_n4292);
nand_1 g03916(new_n4292, new_n4260, new_n4293);
nand_1 g03917(new_n4293, new_n4291, new_n4294);
xnor_1 g03918(new_n4294, new_n4219, n911);
nand_1 g03919(n6687, n3842, new_n4296);
nand_1 g03920(n11917, n6687, new_n4297);
nand_1 g03921(n9956, n4189, new_n4298);
nand_1 g03922(new_n4298, new_n4297, new_n4299);
nand_1 g03923(n9956, n6687, new_n4300_1);
not_4  g03924(new_n4300_1, new_n4301);
nand_1 g03925(n11917, n4189, new_n4302);
not_4  g03926(new_n4302, new_n4303);
nand_1 g03927(new_n4303, new_n4301, new_n4304);
nand_1 g03928(n4921, n2564, new_n4305);
nand_1 g03929(new_n4305, new_n4304, new_n4306);
nand_1 g03930(new_n4306, new_n4299, new_n4307);
nor_1  g03931(new_n4307, new_n4296, new_n4308);
not_4  g03932(new_n4308, new_n4309);
nand_1 g03933(new_n4307, new_n4296, new_n4310);
nand_1 g03934(new_n4310, new_n4309, new_n4311);
nand_1 g03935(n4921, n4189, new_n4312_1);
not_4  g03936(new_n4312_1, new_n4313);
nand_1 g03937(n11917, n2564, new_n4314);
nand_1 g03938(n9956, n6770, new_n4315);
nand_1 g03939(new_n4315, new_n4314, new_n4316);
nor_1  g03940(new_n4315, new_n4314, new_n4317);
not_4  g03941(new_n4317, new_n4318);
nand_1 g03942(new_n4318, new_n4316, new_n4319);
xnor_1 g03943(new_n4319, new_n4313, new_n4320);
xnor_1 g03944(new_n4320, new_n4311, new_n4321);
nand_1 g03945(new_n4304, new_n4299, new_n4322);
not_4  g03946(new_n4322, new_n4323);
nand_1 g03947(n9956, n2564, new_n4324);
not_4  g03948(new_n4324, new_n4325);
nand_1 g03949(n6687, n4921, new_n4326_1);
not_4  g03950(new_n4326_1, new_n4327);
nand_1 g03951(new_n4327, new_n4325, new_n4328);
nor_1  g03952(new_n4328, new_n4323, new_n4329);
nand_1 g03953(new_n4329, new_n4321, new_n4330);
nand_1 g03954(n6687, n2577, new_n4331);
not_4  g03955(new_n4311, new_n4332);
nand_1 g03956(new_n4320, new_n4332, new_n4333_1);
nand_1 g03957(new_n4333_1, new_n4309, new_n4334);
xnor_1 g03958(new_n4334, new_n4331, new_n4335);
nand_1 g03959(n3842, n2564, new_n4336);
nand_1 g03960(new_n4318, new_n4312_1, new_n4337);
nand_1 g03961(new_n4337, new_n4316, new_n4338);
nor_1  g03962(new_n4338, new_n4336, new_n4339);
not_4  g03963(new_n4339, new_n4340);
nand_1 g03964(new_n4338, new_n4336, new_n4341);
nand_1 g03965(new_n4341, new_n4340, new_n4342);
nand_1 g03966(n6770, n4921, new_n4343);
nand_1 g03967(n9956, n9920, new_n4344);
xnor_1 g03968(new_n4344, new_n4303, new_n4345);
xnor_1 g03969(new_n4345, new_n4343, new_n4346);
xnor_1 g03970(new_n4346, new_n4342, new_n4347);
xnor_1 g03971(new_n4347, new_n4335, new_n4348);
not_4  g03972(new_n4348, new_n4349);
xnor_1 g03973(new_n4349, new_n4330, new_n4350);
not_4  g03974(new_n4350, new_n4351);
xnor_1 g03975(new_n4329, new_n4321, new_n4352);
not_4  g03976(new_n4352, new_n4353);
nand_1 g03977(n8595, n8336, new_n4354);
nand_1 g03978(n8336, n6126, new_n4355);
nand_1 g03979(n6986, n3719, new_n4356);
nand_1 g03980(new_n4356, new_n4355, new_n4357);
nand_1 g03981(n8336, n3719, new_n4358);
not_4  g03982(new_n4358, new_n4359);
nand_1 g03983(n6986, n6126, new_n4360);
not_4  g03984(new_n4360, new_n4361);
nand_1 g03985(new_n4361, new_n4359, new_n4362);
nand_1 g03986(n10928, n3602, new_n4363);
nand_1 g03987(new_n4363, new_n4362, new_n4364);
nand_1 g03988(new_n4364, new_n4357, new_n4365);
xnor_1 g03989(new_n4365, new_n4354, new_n4366);
nand_1 g03990(n6986, n3602, new_n4367);
not_4  g03991(new_n4367, new_n4368);
nand_1 g03992(n10928, n6126, new_n4369);
nand_1 g03993(n3719, n2226, new_n4370_1);
nand_1 g03994(new_n4370_1, new_n4369, new_n4371);
nor_1  g03995(new_n4370_1, new_n4369, new_n4372);
not_4  g03996(new_n4372, new_n4373);
nand_1 g03997(new_n4373, new_n4371, new_n4374);
xnor_1 g03998(new_n4374, new_n4368, new_n4375);
not_4  g03999(new_n4375, new_n4376);
nor_1  g04000(new_n4376, new_n4366, new_n4377);
not_4  g04001(new_n4377, new_n4378_1);
nand_1 g04002(new_n4376, new_n4366, new_n4379);
nand_1 g04003(new_n4379, new_n4378_1, new_n4380);
not_4  g04004(new_n4363, new_n4381);
nand_1 g04005(new_n4381, new_n4358, new_n4382);
nand_1 g04006(new_n4362, new_n4357, new_n4383);
nand_1 g04007(new_n4383, new_n4382, new_n4384);
not_4  g04008(new_n4384, new_n4385);
nand_1 g04009(new_n4385, new_n4381, new_n4386);
nand_1 g04010(new_n4386, new_n4380, new_n4387);
not_4  g04011(new_n4380, new_n4388);
not_4  g04012(new_n4386, new_n4389);
nand_1 g04013(new_n4389, new_n4388, new_n4390);
nand_1 g04014(new_n4390, new_n4387, new_n4391);
nand_1 g04015(n12069, n7610, new_n4392);
nand_1 g04016(n12069, n4826, new_n4393);
nand_1 g04017(n12925, n7891, new_n4394);
nand_1 g04018(new_n4394, new_n4393, new_n4395);
nand_1 g04019(n12925, n12069, new_n4396);
not_4  g04020(new_n4396, new_n4397_1);
nand_1 g04021(n7891, n4826, new_n4398);
not_4  g04022(new_n4398, new_n4399);
nand_1 g04023(new_n4399, new_n4397_1, new_n4400);
nand_1 g04024(n12391, n7733, new_n4401);
nand_1 g04025(new_n4401, new_n4400, new_n4402);
nand_1 g04026(new_n4402, new_n4395, new_n4403);
xnor_1 g04027(new_n4403, new_n4392, new_n4404);
nand_1 g04028(n7891, n7733, new_n4405);
nand_1 g04029(n12925, n7160, new_n4406);
nand_1 g04030(n12391, n4826, new_n4407);
not_4  g04031(new_n4407, new_n4408);
xnor_1 g04032(new_n4408, new_n4406, new_n4409);
nor_1  g04033(new_n4409, new_n4405, new_n4410);
nand_1 g04034(new_n4409, new_n4405, new_n4411);
not_4  g04035(new_n4411, new_n4412);
nor_1  g04036(new_n4412, new_n4410, new_n4413);
not_4  g04037(new_n4413, new_n4414);
xnor_1 g04038(new_n4414, new_n4404, new_n4415);
nand_1 g04039(new_n4400, new_n4395, new_n4416);
not_4  g04040(new_n4416, new_n4417);
nand_1 g04041(n12925, n12391, new_n4418);
not_4  g04042(new_n4418, new_n4419);
nand_1 g04043(n12069, n7733, new_n4420);
not_4  g04044(new_n4420, new_n4421);
nand_1 g04045(new_n4421, new_n4419, new_n4422);
nor_1  g04046(new_n4422, new_n4417, new_n4423);
nor_1  g04047(new_n4423, new_n4415, new_n4424);
nand_1 g04048(new_n4423, new_n4415, new_n4425);
not_4  g04049(new_n4425, new_n4426);
nor_1  g04050(new_n4426, new_n4424, new_n4427);
nand_1 g04051(n11222, n217, new_n4428);
nand_1 g04052(n8433, n5314, new_n4429);
nand_1 g04053(n11222, n4086, new_n4430);
nand_1 g04054(new_n4430, new_n4429, new_n4431);
not_4  g04055(new_n4429, new_n4432);
not_4  g04056(new_n4430, new_n4433);
nand_1 g04057(new_n4433, new_n4432, new_n4434);
nand_1 g04058(n11153, n405, new_n4435);
nand_1 g04059(new_n4435, new_n4434, new_n4436_1);
nand_1 g04060(new_n4436_1, new_n4431, new_n4437);
nor_1  g04061(new_n4437, new_n4428, new_n4438);
not_4  g04062(new_n4438, new_n4439);
nand_1 g04063(new_n4437, new_n4428, new_n4440);
nand_1 g04064(new_n4440, new_n4439, new_n4441);
nand_1 g04065(n5314, n405, new_n4442);
not_4  g04066(new_n4442, new_n4443);
nand_1 g04067(n8433, n996, new_n4444);
nand_1 g04068(n11153, n4086, new_n4445);
nand_1 g04069(new_n4445, new_n4444, new_n4446);
not_4  g04070(new_n4444, new_n4447);
not_4  g04071(new_n4445, new_n4448);
nand_1 g04072(new_n4448, new_n4447, new_n4449);
nand_1 g04073(new_n4449, new_n4446, new_n4450);
xnor_1 g04074(new_n4450, new_n4443, new_n4451);
xnor_1 g04075(new_n4451, new_n4441, new_n4452);
not_4  g04076(new_n4435, new_n4453);
not_4  g04077(new_n4431, new_n4454);
nand_1 g04078(n11222, n8433, new_n4455);
nand_1 g04079(new_n4455, new_n4453, new_n4456);
nand_1 g04080(new_n4456, new_n4454, new_n4457);
nand_1 g04081(new_n4457, new_n4434, new_n4458);
nand_1 g04082(new_n4458, new_n4453, new_n4459);
xnor_1 g04083(new_n4459, new_n4452, new_n4460);
not_4  g04084(new_n4460, new_n4461);
xnor_1 g04085(new_n4461, new_n4427, new_n4462);
not_4  g04086(new_n4455, new_n4463);
nand_1 g04087(new_n4463, new_n4397_1, new_n4464);
not_4  g04088(new_n4464, new_n4465);
nand_1 g04089(n11153, n8433, new_n4466);
nand_1 g04090(n11222, n405, new_n4467);
not_4  g04091(new_n4467, new_n4468);
xnor_1 g04092(new_n4468, new_n4466, new_n4469);
nor_1  g04093(new_n4469, new_n4465, new_n4470);
not_4  g04094(new_n4470, new_n4471);
xnor_1 g04095(new_n4469, new_n4464, new_n4472);
nand_1 g04096(new_n4420, new_n4418, new_n4473);
nand_1 g04097(new_n4473, new_n4422, new_n4474);
nand_1 g04098(new_n4474, new_n4472, new_n4475);
nand_1 g04099(new_n4475, new_n4471, new_n4476);
nor_1  g04100(new_n4456, new_n4454, new_n4477);
nor_1  g04101(new_n4477, new_n4458, new_n4478);
not_4  g04102(new_n4478, new_n4479);
nand_1 g04103(new_n4479, new_n4476, new_n4480);
xnor_1 g04104(new_n4478, new_n4476, new_n4481);
nor_1  g04105(new_n4401, new_n4397_1, new_n4482);
not_4  g04106(new_n4482, new_n4483);
nand_1 g04107(new_n4483, new_n4416, new_n4484);
nand_1 g04108(new_n4482, new_n4395, new_n4485);
nand_1 g04109(new_n4485, new_n4484, new_n4486);
nand_1 g04110(new_n4486, new_n4481, new_n4487);
nand_1 g04111(new_n4487, new_n4480, new_n4488);
not_4  g04112(new_n4488, new_n4489);
xnor_1 g04113(new_n4489, new_n4462, new_n4490);
nor_1  g04114(new_n4490, new_n4391, new_n4491);
not_4  g04115(new_n4491, new_n4492);
nand_1 g04116(new_n4490, new_n4391, new_n4493);
nand_1 g04117(new_n4493, new_n4492, new_n4494);
not_4  g04118(new_n4382, new_n4495);
nand_1 g04119(new_n4495, new_n4357, new_n4496);
nand_1 g04120(new_n4496, new_n4384, new_n4497);
not_4  g04121(new_n4486, new_n4498);
xnor_1 g04122(new_n4498, new_n4481, new_n4499_1);
nor_1  g04123(new_n4499_1, new_n4497, new_n4500);
not_4  g04124(new_n4500, new_n4501);
not_4  g04125(new_n4497, new_n4502);
xnor_1 g04126(new_n4499_1, new_n4502, new_n4503);
xnor_1 g04127(new_n4474, new_n4472, new_n4504);
nand_1 g04128(n10928, n3719, new_n4505);
nand_1 g04129(n8336, n3602, new_n4506);
xnor_1 g04130(new_n4506, new_n4505, new_n4507);
not_4  g04131(new_n4507, new_n4508);
nand_1 g04132(new_n4508, new_n4504, new_n4509);
nand_1 g04133(new_n4455, new_n4396, new_n4510);
nand_1 g04134(new_n4510, new_n4464, new_n4511);
not_4  g04135(new_n4511, new_n4512);
nand_1 g04136(new_n4512, new_n4359, new_n4513);
not_4  g04137(new_n4513, new_n4514);
xnor_1 g04138(new_n4507, new_n4504, new_n4515);
nand_1 g04139(new_n4515, new_n4514, new_n4516_1);
nand_1 g04140(new_n4516_1, new_n4509, new_n4517);
nand_1 g04141(new_n4517, new_n4503, new_n4518);
nand_1 g04142(new_n4518, new_n4501, new_n4519);
xnor_1 g04143(new_n4519, new_n4494, new_n4520);
nor_1  g04144(new_n4520, new_n4353, new_n4521);
not_4  g04145(new_n4521, new_n4522);
not_4  g04146(new_n4517, new_n4523);
xnor_1 g04147(new_n4523, new_n4503, new_n4524);
not_4  g04148(new_n4524, new_n4525);
nor_1  g04149(new_n4305, new_n4301, new_n4526);
not_4  g04150(new_n4526, new_n4527);
nand_1 g04151(new_n4527, new_n4322, new_n4528);
nand_1 g04152(new_n4526, new_n4299, new_n4529);
nand_1 g04153(new_n4529, new_n4528, new_n4530);
nand_1 g04154(new_n4530, new_n4525, new_n4531);
xnor_1 g04155(new_n4530, new_n4524, new_n4532);
xnor_1 g04156(new_n4512, new_n4358, new_n4533);
nand_1 g04157(new_n4533, new_n4301, new_n4534);
nand_1 g04158(new_n4326_1, new_n4324, new_n4535);
nand_1 g04159(new_n4535, new_n4328, new_n4536);
nand_1 g04160(new_n4536, new_n4534, new_n4537);
xnor_1 g04161(new_n4515, new_n4513, new_n4538);
xnor_1 g04162(new_n4536, new_n4534, new_n4539);
nor_1  g04163(new_n4539, new_n4538, new_n4540);
not_4  g04164(new_n4540, new_n4541);
nand_1 g04165(new_n4541, new_n4537, new_n4542);
nand_1 g04166(new_n4542, new_n4532, new_n4543);
nand_1 g04167(new_n4543, new_n4531, new_n4544);
xnor_1 g04168(new_n4520, new_n4352, new_n4545);
nand_1 g04169(new_n4545, new_n4544, new_n4546);
nand_1 g04170(new_n4546, new_n4522, new_n4547);
nand_1 g04171(new_n4547, new_n4351, new_n4548);
nor_1  g04172(new_n4547, new_n4351, new_n4549);
not_4  g04173(new_n4549, new_n4550);
nand_1 g04174(new_n4550, new_n4548, new_n4551);
nand_1 g04175(n10439, n8336, new_n4552);
nor_1  g04176(new_n4365, new_n4354, new_n4553_1);
nor_1  g04177(new_n4377, new_n4553_1, new_n4554);
not_4  g04178(new_n4554, new_n4555);
xnor_1 g04179(new_n4555, new_n4552, new_n4556);
nand_1 g04180(n10928, n8595, new_n4557);
nand_1 g04181(new_n4373, new_n4367, new_n4558);
nand_1 g04182(new_n4558, new_n4371, new_n4559);
nor_1  g04183(new_n4559, new_n4557, new_n4560);
not_4  g04184(new_n4560, new_n4561);
nand_1 g04185(new_n4559, new_n4557, new_n4562);
nand_1 g04186(new_n4562, new_n4561, new_n4563);
nand_1 g04187(n3602, n2226, new_n4564);
nand_1 g04188(n3719, n1094, new_n4565);
xnor_1 g04189(new_n4565, new_n4361, new_n4566);
xnor_1 g04190(new_n4566, new_n4564, new_n4567);
xnor_1 g04191(new_n4567, new_n4563, new_n4568);
xnor_1 g04192(new_n4568, new_n4556, new_n4569);
not_4  g04193(new_n4569, new_n4570);
xnor_1 g04194(new_n4570, new_n4390, new_n4571);
not_4  g04195(new_n4571, new_n4572);
not_4  g04196(new_n4452, new_n4573);
nor_1  g04197(new_n4459, new_n4573, new_n4574);
nand_1 g04198(n11222, n6611, new_n4575);
nand_1 g04199(n11153, n217, new_n4576);
nand_1 g04200(n996, n405, new_n4577);
not_4  g04201(new_n4577, new_n4578);
nand_1 g04202(n5314, n4086, new_n4579);
nand_1 g04203(n8433, n5767, new_n4580);
nand_1 g04204(new_n4580, new_n4579, new_n4581);
not_4  g04205(new_n4579, new_n4582);
not_4  g04206(new_n4580, new_n4583);
nand_1 g04207(new_n4583, new_n4582, new_n4584);
nand_1 g04208(new_n4584, new_n4581, new_n4585);
xnor_1 g04209(new_n4585, new_n4578, new_n4586);
xnor_1 g04210(new_n4586, new_n4576, new_n4587);
nand_1 g04211(new_n4449, new_n4442, new_n4588);
nand_1 g04212(new_n4588, new_n4446, new_n4589);
xnor_1 g04213(new_n4589, new_n4587, new_n4590);
xnor_1 g04214(new_n4590, new_n4575, new_n4591);
not_4  g04215(new_n4591, new_n4592);
not_4  g04216(new_n4441, new_n4593);
nand_1 g04217(new_n4451, new_n4593, new_n4594);
nand_1 g04218(new_n4594, new_n4439, new_n4595);
xnor_1 g04219(new_n4595, new_n4592, new_n4596);
xnor_1 g04220(new_n4596, new_n4574, new_n4597);
nand_1 g04221(n12069, n4970, new_n4598);
nand_1 g04222(n12391, n7610, new_n4599);
nand_1 g04223(new_n4407, new_n4406, new_n4600);
nand_1 g04224(new_n4411, new_n4600, new_n4601);
not_4  g04225(new_n4601, new_n4602);
xnor_1 g04226(new_n4602, new_n4599, new_n4603);
nand_1 g04227(n7733, n7160, new_n4604);
nand_1 g04228(n12925, n4828, new_n4605);
xnor_1 g04229(new_n4605, new_n4399, new_n4606);
not_4  g04230(new_n4606, new_n4607);
xnor_1 g04231(new_n4607, new_n4604, new_n4608);
xnor_1 g04232(new_n4608, new_n4603, new_n4609);
xnor_1 g04233(new_n4609, new_n4598, new_n4610);
nor_1  g04234(new_n4403, new_n4392, new_n4611);
nor_1  g04235(new_n4413, new_n4404, new_n4612);
nor_1  g04236(new_n4612, new_n4611, new_n4613);
xnor_1 g04237(new_n4613, new_n4610, new_n4614);
xnor_1 g04238(new_n4614, new_n4425, new_n4615);
nor_1  g04239(new_n4460, new_n4427, new_n4616);
not_4  g04240(new_n4616, new_n4617);
nand_1 g04241(new_n4488, new_n4462, new_n4618);
nand_1 g04242(new_n4618, new_n4617, new_n4619);
xnor_1 g04243(new_n4619, new_n4615, new_n4620);
not_4  g04244(new_n4620, new_n4621);
xnor_1 g04245(new_n4621, new_n4597, new_n4622);
nor_1  g04246(new_n4622, new_n4572, new_n4623);
not_4  g04247(new_n4623, new_n4624);
nand_1 g04248(new_n4622, new_n4572, new_n4625);
nand_1 g04249(new_n4625, new_n4624, new_n4626);
not_4  g04250(new_n4494, new_n4627);
nand_1 g04251(new_n4519, new_n4627, new_n4628);
nand_1 g04252(new_n4628, new_n4492, new_n4629);
xnor_1 g04253(new_n4629, new_n4626, new_n4630);
xnor_1 g04254(new_n4630, new_n4551, n992);
nand_1 g04255(n7265, n6687, new_n4632);
nand_1 g04256(n8336, n7946, new_n4633);
nand_1 g04257(n11222, n9763, new_n4634_1);
not_4  g04258(new_n4634_1, new_n4635);
nand_1 g04259(n12069, n2558, new_n4636);
not_4  g04260(new_n4636, new_n4637);
nand_1 g04261(new_n4637, new_n4635, new_n4638);
nand_1 g04262(new_n4636, new_n4634_1, new_n4639);
nand_1 g04263(new_n4639, new_n4638, new_n4640);
not_4  g04264(new_n4640, new_n4641);
xnor_1 g04265(new_n4641, new_n4633, new_n4642);
xnor_1 g04266(new_n4642, new_n4632, n1020);
xnor_1 g04267(new_n2292, new_n2288, n1136);
xnor_1 g04268(new_n4545, new_n4544, n1138);
nand_1 g04269(n12591, n11757, new_n4646);
nand_1 g04270(n5240, n3932, new_n4647);
not_4  g04271(new_n4647, new_n4648);
nand_1 g04272(n11821, n1798, new_n4649);
not_4  g04273(new_n4649, new_n4650);
nand_1 g04274(new_n4650, new_n4648, new_n4651);
nand_1 g04275(new_n4649, new_n4647, new_n4652);
nand_1 g04276(new_n4652, new_n4651, new_n4653);
not_4  g04277(new_n4653, new_n4654);
xnor_1 g04278(new_n4654, new_n4646, new_n4655);
nand_1 g04279(n5240, n1798, new_n4656);
nand_1 g04280(n12591, n3172, new_n4657);
nand_1 g04281(new_n4657, new_n4656, new_n4658);
not_4  g04282(new_n4656, new_n4659);
not_4  g04283(new_n4657, new_n4660);
nand_1 g04284(new_n4660, new_n4659, new_n4661);
nand_1 g04285(n11757, n3932, new_n4662);
nand_1 g04286(new_n4662, new_n4661, new_n4663);
nand_1 g04287(new_n4663, new_n4658, new_n4664);
xnor_1 g04288(new_n4664, new_n4655, new_n4665);
not_4  g04289(new_n4665, new_n4666);
nand_1 g04290(n7456, n1333, new_n4667);
nand_1 g04291(n11757, n1798, new_n4668);
nand_1 g04292(n12591, n1333, new_n4669);
nand_1 g04293(new_n4669, new_n4668, new_n4670);
not_4  g04294(new_n4668, new_n4671);
not_4  g04295(new_n4669, new_n4672);
nand_1 g04296(new_n4672, new_n4671, new_n4673);
nand_1 g04297(n3932, n3172, new_n4674);
nand_1 g04298(new_n4674, new_n4673, new_n4675);
nand_1 g04299(new_n4675, new_n4670, new_n4676);
nor_1  g04300(new_n4676, new_n4667, new_n4677);
not_4  g04301(new_n4677, new_n4678);
not_4  g04302(new_n4676, new_n4679);
xnor_1 g04303(new_n4679, new_n4667, new_n4680);
not_4  g04304(new_n4662, new_n4681);
nand_1 g04305(new_n4661, new_n4658, new_n4682);
xnor_1 g04306(new_n4682, new_n4681, new_n4683);
nand_1 g04307(new_n4683, new_n4680, new_n4684);
nand_1 g04308(new_n4684, new_n4678, new_n4685);
nand_1 g04309(n11662, n1333, new_n4686_1);
nand_1 g04310(n7456, n3172, new_n4687);
xnor_1 g04311(new_n4687, new_n4686_1, new_n4688);
xnor_1 g04312(new_n4688, new_n4685, new_n4689_1);
not_4  g04313(new_n4689_1, new_n4690);
xnor_1 g04314(new_n4690, new_n4666, new_n4691);
not_4  g04315(new_n4691, new_n4692);
nand_1 g04316(n11662, n7862, new_n4693);
not_4  g04317(new_n4693, new_n4694);
not_4  g04318(new_n4680, new_n4695);
xnor_1 g04319(new_n4683, new_n4695, new_n4696);
nor_1  g04320(new_n4696, new_n4694, new_n4697);
xnor_1 g04321(new_n4696, new_n4694, new_n4698);
nand_1 g04322(n7862, n7456, new_n4699);
not_4  g04323(new_n4699, new_n4700);
nand_1 g04324(n3172, n1798, new_n4701);
not_4  g04325(new_n4701, new_n4702);
nand_1 g04326(n12591, n7862, new_n4703);
not_4  g04327(new_n4703, new_n4704);
nand_1 g04328(new_n4704, new_n4702, new_n4705);
nand_1 g04329(new_n4703, new_n4701, new_n4706);
nand_1 g04330(n3932, n1333, new_n4707);
not_4  g04331(new_n4707, new_n4708);
nand_1 g04332(new_n4708, new_n4706, new_n4709);
nand_1 g04333(new_n4709, new_n4705, new_n4710);
nand_1 g04334(new_n4710, new_n4700, new_n4711);
xnor_1 g04335(new_n4710, new_n4699, new_n4712);
not_4  g04336(new_n4712, new_n4713);
nand_1 g04337(new_n4673, new_n4670, new_n4714);
xnor_1 g04338(new_n4714, new_n4674, new_n4715);
nor_1  g04339(new_n4715, new_n4713, new_n4716);
not_4  g04340(new_n4716, new_n4717);
nand_1 g04341(new_n4717, new_n4711, new_n4718);
nor_1  g04342(new_n4718, new_n4698, new_n4719);
nor_1  g04343(new_n4719, new_n4697, new_n4720);
nand_1 g04344(new_n4720, new_n4692, new_n4721);
not_4  g04345(new_n4646, new_n4722_1);
nand_1 g04346(new_n4654, new_n4722_1, new_n4723);
not_4  g04347(new_n4655, new_n4724);
nor_1  g04348(new_n4664, new_n4724, new_n4725);
not_4  g04349(new_n4725, new_n4726);
nand_1 g04350(new_n4726, new_n4723, new_n4727);
nand_1 g04351(n10327, n1333, new_n4728);
not_4  g04352(new_n4728, new_n4729);
nand_1 g04353(n11662, n3172, new_n4730);
nand_1 g04354(n9583, n7862, new_n4731);
not_4  g04355(new_n4731, new_n4732);
xnor_1 g04356(new_n4732, new_n4730, new_n4733_1);
xnor_1 g04357(new_n4733_1, new_n4729, new_n4734);
xnor_1 g04358(new_n4734, new_n4727, new_n4735);
not_4  g04359(new_n4651, new_n4736);
nand_1 g04360(n11757, n7456, new_n4737);
not_4  g04361(new_n4737, new_n4738);
nand_1 g04362(new_n4738, new_n4736, new_n4739);
nand_1 g04363(new_n4737, new_n4651, new_n4740);
nand_1 g04364(new_n4740, new_n4739, new_n4741);
nand_1 g04365(n11821, n3932, new_n4742);
nand_1 g04366(n12591, n5240, new_n4743);
nand_1 g04367(n9080, n1798, new_n4744);
nand_1 g04368(new_n4744, new_n4743, new_n4745);
not_4  g04369(new_n4743, new_n4746);
not_4  g04370(new_n4744, new_n4747);
nand_1 g04371(new_n4747, new_n4746, new_n4748);
nand_1 g04372(new_n4748, new_n4745, new_n4749);
xnor_1 g04373(new_n4749, new_n4742, new_n4750);
not_4  g04374(new_n4750, new_n4751);
xnor_1 g04375(new_n4751, new_n4741, new_n4752);
xnor_1 g04376(new_n4752, new_n4735, new_n4753);
not_4  g04377(new_n4688, new_n4754);
nand_1 g04378(new_n4754, new_n4685, new_n4755);
nor_1  g04379(new_n4687, new_n4686_1, new_n4756);
nor_1  g04380(new_n4690, new_n4666, new_n4757_1);
xnor_1 g04381(new_n4757_1, new_n4756, new_n4758);
nand_1 g04382(new_n4758, new_n4755, new_n4759);
xnor_1 g04383(new_n4759, new_n4753, new_n4760);
xnor_1 g04384(new_n4760, new_n4721, new_n4761);
nand_1 g04385(n10327, n7862, new_n4762);
not_4  g04386(new_n4762, new_n4763);
xnor_1 g04387(new_n4720, new_n4691, new_n4764);
nand_1 g04388(new_n4764, new_n4763, new_n4765);
xnor_1 g04389(new_n4715, new_n4712, new_n4766);
nand_1 g04390(new_n4706, new_n4705, new_n4767);
not_4  g04391(new_n4767, new_n4768);
nand_1 g04392(n1798, n1333, new_n4769);
not_4  g04393(new_n4769, new_n4770);
nand_1 g04394(n7862, n3932, new_n4771);
not_4  g04395(new_n4771, new_n4772);
nand_1 g04396(new_n4772, new_n4770, new_n4773);
nor_1  g04397(new_n4773, new_n4768, new_n4774);
nand_1 g04398(new_n4774, new_n4766, new_n4775);
not_4  g04399(new_n4775, new_n4776);
xnor_1 g04400(new_n4718, new_n4698, new_n4777);
nand_1 g04401(new_n4777, new_n4776, new_n4778);
not_4  g04402(new_n4778, new_n4779);
xnor_1 g04403(new_n4764, new_n4762, new_n4780);
nand_1 g04404(new_n4780, new_n4779, new_n4781);
nand_1 g04405(new_n4781, new_n4765, new_n4782);
xnor_1 g04406(new_n4782, new_n4761, new_n4783);
nand_1 g04407(n11311, n3022, new_n4784);
not_4  g04408(new_n4784, new_n4785);
nand_1 g04409(n9640, n4187, new_n4786);
nand_1 g04410(n6703, n4203, new_n4787);
not_4  g04411(new_n4787, new_n4788);
xnor_1 g04412(new_n4788, new_n4786, new_n4789);
xnor_1 g04413(new_n4789, new_n4785, new_n4790);
nand_1 g04414(n6703, n4187, new_n4791);
nand_1 g04415(n3022, n2464, new_n4792);
nand_1 g04416(new_n4792, new_n4791, new_n4793);
not_4  g04417(new_n4791, new_n4794);
not_4  g04418(new_n4792, new_n4795);
nand_1 g04419(new_n4795, new_n4794, new_n4796);
nand_1 g04420(n11311, n9640, new_n4797);
nand_1 g04421(new_n4797, new_n4796, new_n4798);
nand_1 g04422(new_n4798, new_n4793, new_n4799);
nor_1  g04423(new_n4799, new_n4790, new_n4800);
not_4  g04424(new_n4800, new_n4801);
nand_1 g04425(new_n4799, new_n4790, new_n4802);
nand_1 g04426(new_n4802, new_n4801, new_n4803);
nand_1 g04427(n10451, n9400, new_n4804);
nand_1 g04428(n11023, n2464, new_n4805_1);
not_4  g04429(new_n4805_1, new_n4806);
xnor_1 g04430(new_n4806, new_n4804, new_n4807);
xnor_1 g04431(new_n4807, new_n4803, new_n4808);
nand_1 g04432(n11023, n9400, new_n4809);
nand_1 g04433(n11311, n6703, new_n4810);
nand_1 g04434(n9400, n3022, new_n4811);
nand_1 g04435(new_n4811, new_n4810, new_n4812);
not_4  g04436(new_n4810, new_n4813);
not_4  g04437(new_n4811, new_n4814);
nand_1 g04438(new_n4814, new_n4813, new_n4815);
nand_1 g04439(n9640, n2464, new_n4816);
nand_1 g04440(new_n4816, new_n4815, new_n4817_1);
nand_1 g04441(new_n4817_1, new_n4812, new_n4818);
nor_1  g04442(new_n4818, new_n4809, new_n4819);
not_4  g04443(new_n4818, new_n4820);
xnor_1 g04444(new_n4820, new_n4809, new_n4821);
not_4  g04445(new_n4821, new_n4822);
nand_1 g04446(new_n4796, new_n4793, new_n4823);
xnor_1 g04447(new_n4823, new_n4797, new_n4824);
nor_1  g04448(new_n4824, new_n4822, new_n4825);
nor_1  g04449(new_n4825, new_n4819, new_n4826_1);
not_4  g04450(new_n4826_1, new_n4827);
xnor_1 g04451(new_n4827, new_n4808, new_n4828_1);
not_4  g04452(new_n4828_1, new_n4829);
nand_1 g04453(n10451, n6877, new_n4830);
not_4  g04454(new_n4830, new_n4831);
xnor_1 g04455(new_n4824, new_n4821, new_n4832);
nand_1 g04456(new_n4832, new_n4831, new_n4833);
nand_1 g04457(n11023, n6877, new_n4834);
nand_1 g04458(n6703, n2464, new_n4835);
nand_1 g04459(n6877, n3022, new_n4836);
nand_1 g04460(new_n4836, new_n4835, new_n4837);
nor_1  g04461(new_n4836, new_n4835, new_n4838);
not_4  g04462(new_n4838, new_n4839);
nand_1 g04463(n9640, n9400, new_n4840);
nand_1 g04464(new_n4840, new_n4839, new_n4841);
nand_1 g04465(new_n4841, new_n4837, new_n4842);
nor_1  g04466(new_n4842, new_n4834, new_n4843);
xnor_1 g04467(new_n4842, new_n4834, new_n4844);
nand_1 g04468(new_n4815, new_n4812, new_n4845);
xnor_1 g04469(new_n4845, new_n4816, new_n4846);
nor_1  g04470(new_n4846, new_n4844, new_n4847);
nor_1  g04471(new_n4847, new_n4843, new_n4848);
not_4  g04472(new_n4848, new_n4849);
xnor_1 g04473(new_n4832, new_n4830, new_n4850);
nand_1 g04474(new_n4850, new_n4849, new_n4851);
nand_1 g04475(new_n4851, new_n4833, new_n4852);
nand_1 g04476(new_n4852, new_n4829, new_n4853);
nand_1 g04477(new_n4789, new_n4785, new_n4854);
nand_1 g04478(new_n4801, new_n4854, new_n4855);
nand_1 g04479(n10278, n9400, new_n4856);
nand_1 g04480(n10451, n2464, new_n4857);
not_4  g04481(new_n4857, new_n4858);
nand_1 g04482(n11423, n6877, new_n4859);
not_4  g04483(new_n4859, new_n4860);
nand_1 g04484(new_n4860, new_n4858, new_n4861);
nand_1 g04485(new_n4859, new_n4857, new_n4862);
nand_1 g04486(new_n4862, new_n4861, new_n4863);
xnor_1 g04487(new_n4863, new_n4856, new_n4864);
xnor_1 g04488(new_n4864, new_n4855, new_n4865);
not_4  g04489(new_n4786, new_n4866);
nand_1 g04490(new_n4788, new_n4866, new_n4867);
not_4  g04491(new_n4867, new_n4868);
nand_1 g04492(n11311, n11023, new_n4869);
not_4  g04493(new_n4869, new_n4870);
nand_1 g04494(new_n4870, new_n4868, new_n4871);
nand_1 g04495(new_n4869, new_n4867, new_n4872);
nand_1 g04496(new_n4872, new_n4871, new_n4873);
nand_1 g04497(n9640, n4203, new_n4874);
nand_1 g04498(n4187, n3022, new_n4875);
nand_1 g04499(n12753, n6703, new_n4876);
nand_1 g04500(new_n4876, new_n4875, new_n4877);
not_4  g04501(new_n4875, new_n4878);
not_4  g04502(new_n4876, new_n4879);
nand_1 g04503(new_n4879, new_n4878, new_n4880);
nand_1 g04504(new_n4880, new_n4877, new_n4881);
xnor_1 g04505(new_n4881, new_n4874, new_n4882);
not_4  g04506(new_n4882, new_n4883);
xnor_1 g04507(new_n4883, new_n4873, new_n4884);
xnor_1 g04508(new_n4884, new_n4865, new_n4885);
not_4  g04509(new_n4803, new_n4886);
nand_1 g04510(new_n4807, new_n4886, new_n4887);
nor_1  g04511(new_n4805_1, new_n4804, new_n4888);
nand_1 g04512(new_n4827, new_n4808, new_n4889);
not_4  g04513(new_n4889, new_n4890);
xnor_1 g04514(new_n4890, new_n4888, new_n4891);
nand_1 g04515(new_n4891, new_n4887, new_n4892);
xnor_1 g04516(new_n4892, new_n4885, new_n4893);
xnor_1 g04517(new_n4893, new_n4853, new_n4894);
nand_1 g04518(n10278, n6877, new_n4895);
not_4  g04519(new_n4895, new_n4896);
xnor_1 g04520(new_n4852, new_n4828_1, new_n4897);
nand_1 g04521(new_n4897, new_n4896, new_n4898);
xnor_1 g04522(new_n4846, new_n4844, new_n4899);
not_4  g04523(new_n4899, new_n4900);
not_4  g04524(new_n4840, new_n4901);
nand_1 g04525(n6877, n6703, new_n4902);
nand_1 g04526(new_n4902, new_n4901, new_n4903_1);
nand_1 g04527(new_n4839, new_n4837, new_n4904);
nand_1 g04528(new_n4904, new_n4903_1, new_n4905);
not_4  g04529(new_n4905, new_n4906);
nand_1 g04530(new_n4906, new_n4901, new_n4907);
not_4  g04531(new_n4907, new_n4908);
nand_1 g04532(new_n4908, new_n4900, new_n4909);
xnor_1 g04533(new_n4850, new_n4848, new_n4910);
not_4  g04534(new_n4910, new_n4911);
nor_1  g04535(new_n4911, new_n4909, new_n4912);
xnor_1 g04536(new_n4897, new_n4895, new_n4913);
nand_1 g04537(new_n4913, new_n4912, new_n4914);
nand_1 g04538(new_n4914, new_n4898, new_n4915);
xnor_1 g04539(new_n4915, new_n4894, new_n4916);
nand_1 g04540(n12826, n4805, new_n4917);
not_4  g04541(new_n4917, new_n4918);
nand_1 g04542(n8665, n137, new_n4919);
nand_1 g04543(n6294, n1067, new_n4920);
nand_1 g04544(n6797, n5645, new_n4921_1);
not_4  g04545(new_n4921_1, new_n4922);
xnor_1 g04546(new_n4922, new_n4920, new_n4923);
xnor_1 g04547(new_n4923, new_n4919, new_n4924);
nand_1 g04548(n6294, n5645, new_n4925);
nand_1 g04549(n8665, n5283, new_n4926);
nand_1 g04550(new_n4926, new_n4925, new_n4927);
nand_1 g04551(n1067, n137, new_n4928_1);
not_4  g04552(new_n4926, new_n4929);
xnor_1 g04553(new_n4929, new_n4925, new_n4930);
nand_1 g04554(new_n4930, new_n4928_1, new_n4931);
nand_1 g04555(new_n4931, new_n4927, new_n4932);
xnor_1 g04556(new_n4932, new_n4924, new_n4933);
nand_1 g04557(n11922, n11478, new_n4934);
nand_1 g04558(n5283, n1067, new_n4935);
nand_1 g04559(n11478, n8665, new_n4936);
nand_1 g04560(new_n4936, new_n4935, new_n4937);
nand_1 g04561(n5645, n137, new_n4938_1);
not_4  g04562(new_n4935, new_n4939);
not_4  g04563(new_n4936, new_n4940);
nor_1  g04564(new_n4940, new_n4939, new_n4941);
nor_1  g04565(new_n4936, new_n4935, new_n4942);
nor_1  g04566(new_n4942, new_n4941, new_n4943);
nand_1 g04567(new_n4943, new_n4938_1, new_n4944);
nand_1 g04568(new_n4944, new_n4937, new_n4945);
nor_1  g04569(new_n4945, new_n4934, new_n4946);
xnor_1 g04570(new_n4930, new_n4928_1, new_n4947);
not_4  g04571(new_n4947, new_n4948);
not_4  g04572(new_n4934, new_n4949);
not_4  g04573(new_n4938_1, new_n4950);
nand_1 g04574(new_n4940, new_n4939, new_n4951);
nand_1 g04575(new_n4951, new_n4937, new_n4952);
nor_1  g04576(new_n4952, new_n4950, new_n4953);
nor_1  g04577(new_n4953, new_n4941, new_n4954);
nand_1 g04578(new_n4954, new_n4949, new_n4955);
nand_1 g04579(new_n4945, new_n4934, new_n4956);
nand_1 g04580(new_n4956, new_n4955, new_n4957);
nor_1  g04581(new_n4957, new_n4948, new_n4958);
nor_1  g04582(new_n4958, new_n4946, new_n4959);
nand_1 g04583(n11478, n2551, new_n4960);
nand_1 g04584(n11922, n5283, new_n4961);
nand_1 g04585(new_n4961, new_n4960, new_n4962);
not_4  g04586(new_n4960, new_n4963);
not_4  g04587(new_n4961, new_n4964);
nand_1 g04588(new_n4964, new_n4963, new_n4965);
nand_1 g04589(new_n4965, new_n4962, new_n4966);
nor_1  g04590(new_n4966, new_n4959, new_n4967);
nor_1  g04591(new_n4954, new_n4949, new_n4968);
nor_1  g04592(new_n4968, new_n4946, new_n4969);
nand_1 g04593(new_n4969, new_n4947, new_n4970_1);
nand_1 g04594(new_n4970_1, new_n4955, new_n4971_1);
not_4  g04595(new_n4966, new_n4972);
nor_1  g04596(new_n4972, new_n4971_1, new_n4973);
nor_1  g04597(new_n4973, new_n4967, new_n4974);
nand_1 g04598(new_n4974, new_n4933, new_n4975);
not_4  g04599(new_n4933, new_n4976);
nand_1 g04600(new_n4972, new_n4971_1, new_n4977);
nand_1 g04601(new_n4966, new_n4959, new_n4978);
nand_1 g04602(new_n4978, new_n4977, new_n4979);
nand_1 g04603(new_n4979, new_n4976, new_n4980);
nand_1 g04604(new_n4980, new_n4975, new_n4981);
nand_1 g04605(n4805, n2551, new_n4982);
not_4  g04606(new_n4982, new_n4983);
nand_1 g04607(n11922, n4805, new_n4984);
not_4  g04608(new_n4984, new_n4985);
nand_1 g04609(n5645, n5283, new_n4986);
not_4  g04610(new_n4986, new_n4987);
nand_1 g04611(n8665, n4805, new_n4988);
not_4  g04612(new_n4988, new_n4989);
nand_1 g04613(new_n4989, new_n4987, new_n4990);
nand_1 g04614(new_n4988, new_n4986, new_n4991);
nand_1 g04615(n11478, n1067, new_n4992);
not_4  g04616(new_n4992, new_n4993);
nand_1 g04617(new_n4993, new_n4991, new_n4994);
nand_1 g04618(new_n4994, new_n4990, new_n4995);
nand_1 g04619(new_n4995, new_n4985, new_n4996);
xnor_1 g04620(new_n4995, new_n4984, new_n4997);
nand_1 g04621(new_n4952, new_n4950, new_n4998);
nand_1 g04622(new_n4998, new_n4944, new_n4999);
nand_1 g04623(new_n4999, new_n4997, new_n5000);
nand_1 g04624(new_n5000, new_n4996, new_n5001);
nor_1  g04625(new_n5001, new_n4983, new_n5002);
not_4  g04626(new_n5002, new_n5003);
nand_1 g04627(new_n4957, new_n4948, new_n5004);
nand_1 g04628(new_n5004, new_n4970_1, new_n5005);
nand_1 g04629(new_n5001, new_n4983, new_n5006);
nand_1 g04630(new_n5006, new_n5003, new_n5007);
not_4  g04631(new_n5007, new_n5008);
nand_1 g04632(new_n5008, new_n5005, new_n5009);
nand_1 g04633(new_n5009, new_n5003, new_n5010);
nor_1  g04634(new_n5010, new_n4981, new_n5011);
nor_1  g04635(new_n4979, new_n4976, new_n5012);
nor_1  g04636(new_n4974, new_n4933, new_n5013);
nor_1  g04637(new_n5013, new_n5012, new_n5014);
not_4  g04638(new_n5010, new_n5015);
nor_1  g04639(new_n5015, new_n5014, new_n5016);
nor_1  g04640(new_n5016, new_n5011, new_n5017);
nand_1 g04641(new_n5017, new_n4918, new_n5018);
not_4  g04642(new_n4997, new_n5019);
xnor_1 g04643(new_n4999, new_n5019, new_n5020);
nand_1 g04644(new_n4991, new_n4990, new_n5021);
not_4  g04645(new_n5021, new_n5022);
nand_1 g04646(n4805, n1067, new_n5023);
not_4  g04647(new_n5023, new_n5024);
nand_1 g04648(n11478, n5645, new_n5025);
not_4  g04649(new_n5025, new_n5026);
nand_1 g04650(new_n5026, new_n5024, new_n5027);
nor_1  g04651(new_n5027, new_n5022, new_n5028);
nand_1 g04652(new_n5028, new_n5020, new_n5029);
xnor_1 g04653(new_n5007, new_n5005, new_n5030_1);
nor_1  g04654(new_n5030_1, new_n5029, new_n5031);
nand_1 g04655(new_n5015, new_n5014, new_n5032);
nand_1 g04656(new_n5010, new_n4981, new_n5033);
nand_1 g04657(new_n5033, new_n5032, new_n5034_1);
nor_1  g04658(new_n5034_1, new_n4917, new_n5035);
nor_1  g04659(new_n5017, new_n4918, new_n5036);
nor_1  g04660(new_n5036, new_n5035, new_n5037);
nand_1 g04661(new_n5037, new_n5031, new_n5038);
nand_1 g04662(new_n5038, new_n5018, new_n5039);
nand_1 g04663(n12826, n11478, new_n5040);
nand_1 g04664(n5283, n2551, new_n5041);
not_4  g04665(new_n5041, new_n5042);
nand_1 g04666(n4805, n4094, new_n5043);
xnor_1 g04667(new_n5043, new_n5042, new_n5044);
xnor_1 g04668(new_n5044, new_n5040, new_n5045);
not_4  g04669(new_n4919, new_n5046);
nand_1 g04670(new_n4923, new_n5046, new_n5047);
not_4  g04671(new_n4932, new_n5048);
nand_1 g04672(new_n5048, new_n4924, new_n5049);
nand_1 g04673(new_n5049, new_n5047, new_n5050);
not_4  g04674(new_n5050, new_n5051);
xnor_1 g04675(new_n5051, new_n5045, new_n5052);
not_4  g04676(new_n4920, new_n5053);
nand_1 g04677(new_n4922, new_n5053, new_n5054);
nand_1 g04678(n11922, n137, new_n5055);
nand_1 g04679(new_n5055, new_n5054, new_n5056);
not_4  g04680(new_n5054, new_n5057);
not_4  g04681(new_n5055, new_n5058);
nand_1 g04682(new_n5058, new_n5057, new_n5059);
nand_1 g04683(new_n5059, new_n5056, new_n5060);
not_4  g04684(new_n5060, new_n5061);
nand_1 g04685(n6797, n1067, new_n5062);
nand_1 g04686(n8665, n6294, new_n5063);
nand_1 g04687(n5645, n3146, new_n5064);
not_4  g04688(new_n5064, new_n5065);
xnor_1 g04689(new_n5065, new_n5063, new_n5066);
xnor_1 g04690(new_n5066, new_n5062, new_n5067);
not_4  g04691(new_n5067, new_n5068);
xnor_1 g04692(new_n5068, new_n5061, new_n5069_1);
xnor_1 g04693(new_n5069_1, new_n5052, new_n5070);
not_4  g04694(new_n5070, new_n5071);
not_4  g04695(new_n4965, new_n5072);
nand_1 g04696(new_n5012, new_n5072, new_n5073);
nand_1 g04697(new_n4975, new_n4965, new_n5074);
nand_1 g04698(new_n5074, new_n5073, new_n5075);
nand_1 g04699(new_n5075, new_n4977, new_n5076);
nand_1 g04700(new_n5076, new_n5071, new_n5077);
nor_1  g04701(new_n4975, new_n4965, new_n5078);
nor_1  g04702(new_n5012, new_n5072, new_n5079);
nor_1  g04703(new_n5079, new_n5078, new_n5080);
nor_1  g04704(new_n5080, new_n4967, new_n5081);
nand_1 g04705(new_n5081, new_n5070, new_n5082);
nand_1 g04706(new_n5082, new_n5077, new_n5083);
nor_1  g04707(new_n5083, new_n5032, new_n5084);
nor_1  g04708(new_n5081, new_n5070, new_n5085);
nor_1  g04709(new_n5076, new_n5071, new_n5086);
nor_1  g04710(new_n5086, new_n5085, new_n5087);
nor_1  g04711(new_n5087, new_n5011, new_n5088);
nor_1  g04712(new_n5088, new_n5084, new_n5089);
nand_1 g04713(new_n5089, new_n5039, new_n5090);
not_4  g04714(new_n5031, new_n5091);
nand_1 g04715(new_n5034_1, new_n4917, new_n5092);
nand_1 g04716(new_n5092, new_n5018, new_n5093);
nor_1  g04717(new_n5093, new_n5091, new_n5094_1);
nor_1  g04718(new_n5094_1, new_n5035, new_n5095);
nand_1 g04719(new_n5087, new_n5011, new_n5096);
nand_1 g04720(new_n5083, new_n5032, new_n5097);
nand_1 g04721(new_n5097, new_n5096, new_n5098);
nand_1 g04722(new_n5098, new_n5095, new_n5099);
nand_1 g04723(new_n5099, new_n5090, new_n5100);
nand_1 g04724(n3992, n2749, new_n5101);
not_4  g04725(new_n5101, new_n5102);
nand_1 g04726(n11876, n6358, new_n5103);
not_4  g04727(new_n5103, new_n5104);
nand_1 g04728(n3992, n3754, new_n5105_1);
not_4  g04729(new_n5105_1, new_n5106);
nor_1  g04730(new_n5106, new_n5104, new_n5107);
nand_1 g04731(n10898, n8384, new_n5108);
not_4  g04732(new_n5108, new_n5109);
nand_1 g04733(new_n5105_1, new_n5103, new_n5110);
nand_1 g04734(new_n5106, new_n5104, new_n5111);
nand_1 g04735(new_n5111, new_n5110, new_n5112);
nor_1  g04736(new_n5112, new_n5109, new_n5113);
nor_1  g04737(new_n5113, new_n5107, new_n5114);
nand_1 g04738(new_n5114, new_n5102, new_n5115);
nor_1  g04739(new_n5105_1, new_n5103, new_n5116);
nor_1  g04740(new_n5116, new_n5107, new_n5117);
nand_1 g04741(new_n5117, new_n5108, new_n5118);
nand_1 g04742(new_n5118, new_n5110, new_n5119);
nor_1  g04743(new_n5119, new_n5101, new_n5120);
nor_1  g04744(new_n5114, new_n5102, new_n5121);
nor_1  g04745(new_n5121, new_n5120, new_n5122);
nand_1 g04746(n10898, n6358, new_n5123);
nand_1 g04747(n11876, n5198, new_n5124);
nand_1 g04748(n8384, n3754, new_n5125);
not_4  g04749(new_n5125, new_n5126);
xnor_1 g04750(new_n5126, new_n5124, new_n5127);
xnor_1 g04751(new_n5127, new_n5123, new_n5128);
nand_1 g04752(new_n5128, new_n5122, new_n5129);
nand_1 g04753(new_n5129, new_n5115, new_n5130);
nand_1 g04754(n8384, n2749, new_n5131);
nand_1 g04755(n3992, n159, new_n5132_1);
nand_1 g04756(new_n5132_1, new_n5131, new_n5133);
not_4  g04757(new_n5131, new_n5134);
not_4  g04758(new_n5132_1, new_n5135);
nand_1 g04759(new_n5135, new_n5134, new_n5136);
nand_1 g04760(new_n5136, new_n5133, new_n5137);
not_4  g04761(new_n5137, new_n5138);
nand_1 g04762(new_n5138, new_n5130, new_n5139);
nand_1 g04763(new_n5119, new_n5101, new_n5140);
nand_1 g04764(new_n5140, new_n5115, new_n5141);
not_4  g04765(new_n5128, new_n5142);
nor_1  g04766(new_n5142, new_n5141, new_n5143);
nor_1  g04767(new_n5143, new_n5120, new_n5144);
nand_1 g04768(new_n5137, new_n5144, new_n5145);
nand_1 g04769(new_n5145, new_n5139, new_n5146);
nand_1 g04770(n6358, n3754, new_n5147);
nand_1 g04771(n10898, n5198, new_n5148);
nand_1 g04772(n11876, n1471, new_n5149);
not_4  g04773(new_n5149, new_n5150);
xnor_1 g04774(new_n5150, new_n5148, new_n5151);
not_4  g04775(new_n5151, new_n5152);
xnor_1 g04776(new_n5152, new_n5147, new_n5153_1);
nand_1 g04777(new_n5125, new_n5124, new_n5154);
nand_1 g04778(new_n5127, new_n5123, new_n5155);
nand_1 g04779(new_n5155, new_n5154, new_n5156);
xnor_1 g04780(new_n5156, new_n5153_1, new_n5157);
nor_1  g04781(new_n5157, new_n5146, new_n5158);
nor_1  g04782(new_n5137, new_n5144, new_n5159);
nor_1  g04783(new_n5138, new_n5130, new_n5160);
nor_1  g04784(new_n5160, new_n5159, new_n5161);
not_4  g04785(new_n5157, new_n5162);
nor_1  g04786(new_n5162, new_n5161, new_n5163);
nor_1  g04787(new_n5163, new_n5158, new_n5164);
nand_1 g04788(n7236, n159, new_n5165);
not_4  g04789(new_n5165, new_n5166);
nand_1 g04790(n7236, n2749, new_n5167);
nand_1 g04791(n11876, n8384, new_n5168);
nand_1 g04792(n7236, n3754, new_n5169);
nand_1 g04793(new_n5169, new_n5168, new_n5170);
nand_1 g04794(n11876, n7236, new_n5171);
not_4  g04795(new_n5171, new_n5172);
nand_1 g04796(new_n5172, new_n5126, new_n5173);
nand_1 g04797(n10898, n3992, new_n5174);
nand_1 g04798(new_n5174, new_n5173, new_n5175);
nand_1 g04799(new_n5175, new_n5170, new_n5176);
nor_1  g04800(new_n5176, new_n5167, new_n5177);
not_4  g04801(new_n5177, new_n5178);
not_4  g04802(new_n5176, new_n5179);
xnor_1 g04803(new_n5179, new_n5167, new_n5180);
xnor_1 g04804(new_n5112, new_n5108, new_n5181);
not_4  g04805(new_n5181, new_n5182);
nand_1 g04806(new_n5182, new_n5180, new_n5183);
nand_1 g04807(new_n5183, new_n5178, new_n5184);
nor_1  g04808(new_n5184, new_n5166, new_n5185);
not_4  g04809(new_n5185, new_n5186);
nand_1 g04810(new_n5142, new_n5141, new_n5187);
nand_1 g04811(new_n5187, new_n5129, new_n5188);
nand_1 g04812(new_n5184, new_n5166, new_n5189);
nand_1 g04813(new_n5189, new_n5186, new_n5190);
not_4  g04814(new_n5190, new_n5191_1);
nand_1 g04815(new_n5191_1, new_n5188, new_n5192);
nand_1 g04816(new_n5192, new_n5186, new_n5193);
not_4  g04817(new_n5193, new_n5194);
nand_1 g04818(new_n5194, new_n5164, new_n5195);
not_4  g04819(new_n5148, new_n5196);
nand_1 g04820(new_n5150, new_n5196, new_n5197);
not_4  g04821(new_n5197, new_n5198_1);
nand_1 g04822(n6358, n2749, new_n5199);
not_4  g04823(new_n5199, new_n5200);
nand_1 g04824(new_n5200, new_n5198_1, new_n5201);
nand_1 g04825(new_n5199, new_n5197, new_n5202);
nand_1 g04826(new_n5202, new_n5201, new_n5203);
not_4  g04827(new_n5203, new_n5204);
nand_1 g04828(n10898, n1471, new_n5205);
nand_1 g04829(n5198, n3754, new_n5206);
nand_1 g04830(n11876, n7646, new_n5207);
not_4  g04831(new_n5207, new_n5208);
xnor_1 g04832(new_n5208, new_n5206, new_n5209);
xnor_1 g04833(new_n5209, new_n5205, new_n5210);
not_4  g04834(new_n5210, new_n5211);
xnor_1 g04835(new_n5211, new_n5204, new_n5212_1);
nand_1 g04836(new_n5152, new_n5147, new_n5213);
not_4  g04837(new_n5153_1, new_n5214);
nand_1 g04838(new_n5156, new_n5214, new_n5215);
nand_1 g04839(new_n5215, new_n5213, new_n5216);
nand_1 g04840(n3992, n1510, new_n5217);
nand_1 g04841(n8384, n159, new_n5218);
nand_1 g04842(n12247, n7236, new_n5219);
not_4  g04843(new_n5219, new_n5220);
xnor_1 g04844(new_n5220, new_n5218, new_n5221);
xnor_1 g04845(new_n5221, new_n5217, new_n5222);
xnor_1 g04846(new_n5222, new_n5216, new_n5223);
xnor_1 g04847(new_n5223, new_n5212_1, new_n5224);
not_4  g04848(new_n5224, new_n5225);
not_4  g04849(new_n5136, new_n5226);
nand_1 g04850(new_n5158, new_n5226, new_n5227);
nand_1 g04851(new_n5162, new_n5161, new_n5228);
nand_1 g04852(new_n5228, new_n5136, new_n5229);
nand_1 g04853(new_n5229, new_n5227, new_n5230);
nand_1 g04854(new_n5230, new_n5139, new_n5231);
nand_1 g04855(new_n5231, new_n5225, new_n5232);
nor_1  g04856(new_n5228, new_n5136, new_n5233);
nor_1  g04857(new_n5158, new_n5226, new_n5234);
nor_1  g04858(new_n5234, new_n5233, new_n5235);
nor_1  g04859(new_n5235, new_n5159, new_n5236);
nand_1 g04860(new_n5236, new_n5224, new_n5237);
nand_1 g04861(new_n5237, new_n5232, new_n5238);
nor_1  g04862(new_n5238, new_n5195, new_n5239);
nand_1 g04863(new_n5157, new_n5146, new_n5240_1);
nand_1 g04864(new_n5240_1, new_n5228, new_n5241);
nor_1  g04865(new_n5193, new_n5241, new_n5242);
nor_1  g04866(new_n5236, new_n5224, new_n5243);
nor_1  g04867(new_n5231, new_n5225, new_n5244);
nor_1  g04868(new_n5244, new_n5243, new_n5245);
nor_1  g04869(new_n5245, new_n5242, new_n5246);
nor_1  g04870(new_n5246, new_n5239, new_n5247);
nand_1 g04871(n7236, n1510, new_n5248);
not_4  g04872(new_n5248, new_n5249);
nor_1  g04873(new_n5194, new_n5164, new_n5250);
nor_1  g04874(new_n5250, new_n5242, new_n5251);
nand_1 g04875(new_n5251, new_n5249, new_n5252);
xnor_1 g04876(new_n5182, new_n5180, new_n5253);
not_4  g04877(new_n5253, new_n5254);
nand_1 g04878(new_n5173, new_n5170, new_n5255);
not_4  g04879(new_n5255, new_n5256);
nand_1 g04880(n11876, n3992, new_n5257_1);
not_4  g04881(new_n5257_1, new_n5258);
nand_1 g04882(n10898, n7236, new_n5259);
not_4  g04883(new_n5259, new_n5260);
nand_1 g04884(new_n5260, new_n5258, new_n5261);
nor_1  g04885(new_n5261, new_n5256, new_n5262);
nand_1 g04886(new_n5262, new_n5254, new_n5263);
xnor_1 g04887(new_n5190, new_n5188, new_n5264);
nor_1  g04888(new_n5264, new_n5263, new_n5265);
nand_1 g04889(new_n5193, new_n5241, new_n5266);
nand_1 g04890(new_n5266, new_n5195, new_n5267);
nor_1  g04891(new_n5267, new_n5248, new_n5268);
nor_1  g04892(new_n5251, new_n5249, new_n5269);
nor_1  g04893(new_n5269, new_n5268, new_n5270);
nand_1 g04894(new_n5270, new_n5265, new_n5271);
nand_1 g04895(new_n5271, new_n5252, new_n5272);
nand_1 g04896(new_n5272, new_n5247, new_n5273);
nand_1 g04897(new_n5245, new_n5242, new_n5274);
nand_1 g04898(new_n5238, new_n5195, new_n5275);
nand_1 g04899(new_n5275, new_n5274, new_n5276);
not_4  g04900(new_n5265, new_n5277);
nand_1 g04901(new_n5267, new_n5248, new_n5278);
nand_1 g04902(new_n5278, new_n5252, new_n5279);
nor_1  g04903(new_n5279, new_n5277, new_n5280);
nor_1  g04904(new_n5280, new_n5268, new_n5281);
nand_1 g04905(new_n5281, new_n5276, new_n5282);
nand_1 g04906(new_n5282, new_n5273, new_n5283_1);
nand_1 g04907(new_n5283_1, new_n5100, new_n5284);
nor_1  g04908(new_n5098, new_n5095, new_n5285);
nor_1  g04909(new_n5089, new_n5039, new_n5286);
nor_1  g04910(new_n5286, new_n5285, new_n5287);
nor_1  g04911(new_n5281, new_n5276, new_n5288);
nor_1  g04912(new_n5272, new_n5247, new_n5289);
nor_1  g04913(new_n5289, new_n5288, new_n5290);
nand_1 g04914(new_n5290, new_n5287, new_n5291);
nand_1 g04915(new_n5291, new_n5284, new_n5292);
nor_1  g04916(new_n5037, new_n5031, new_n5293);
nor_1  g04917(new_n5293, new_n5094_1, new_n5294);
nor_1  g04918(new_n5270, new_n5265, new_n5295);
nor_1  g04919(new_n5295, new_n5280, new_n5296);
nor_1  g04920(new_n5296, new_n5294, new_n5297);
nand_1 g04921(new_n5093, new_n5091, new_n5298);
nand_1 g04922(new_n5298, new_n5038, new_n5299);
nand_1 g04923(new_n5279, new_n5277, new_n5300);
nand_1 g04924(new_n5300, new_n5271, new_n5301);
nand_1 g04925(new_n5301, new_n5299, new_n5302);
nand_1 g04926(new_n5296, new_n5294, new_n5303);
nand_1 g04927(new_n5303, new_n5302, new_n5304);
nand_1 g04928(new_n5264, new_n5263, new_n5305_1);
nand_1 g04929(new_n5305_1, new_n5277, new_n5306);
not_4  g04930(new_n5028, new_n5307);
xnor_1 g04931(new_n5307, new_n5020, new_n5308);
xnor_1 g04932(new_n5262, new_n5253, new_n5309);
nor_1  g04933(new_n5309, new_n5308, new_n5310);
not_4  g04934(new_n5310, new_n5311);
nand_1 g04935(new_n5259, new_n5257_1, new_n5312);
nand_1 g04936(new_n5312, new_n5261, new_n5313);
not_4  g04937(new_n5313, new_n5314_1);
xnor_1 g04938(new_n5026, new_n5023, new_n5315);
nor_1  g04939(new_n5315, new_n5314_1, new_n5316);
not_4  g04940(new_n5316, new_n5317);
nand_1 g04941(n5645, n4805, new_n5318);
not_4  g04942(new_n5318, new_n5319_1);
nand_1 g04943(new_n5319_1, new_n5172, new_n5320_1);
xnor_1 g04944(new_n5315, new_n5313, new_n5321);
nand_1 g04945(new_n5321, new_n5320_1, new_n5322);
nand_1 g04946(new_n5322, new_n5317, new_n5323);
nand_1 g04947(new_n5318, new_n4993, new_n5324);
nor_1  g04948(new_n5324, new_n4991, new_n5325);
not_4  g04949(new_n5325, new_n5326);
nand_1 g04950(new_n5324, new_n5022, new_n5327);
nand_1 g04951(new_n5327, new_n5326, new_n5328);
not_4  g04952(new_n5328, new_n5329);
nand_1 g04953(new_n5329, new_n5323, new_n5330);
xnor_1 g04954(new_n5328, new_n5323, new_n5331_1);
nor_1  g04955(new_n5174, new_n5172, new_n5332);
not_4  g04956(new_n5332, new_n5333);
nand_1 g04957(new_n5333, new_n5255, new_n5334);
nand_1 g04958(new_n5332, new_n5170, new_n5335);
nand_1 g04959(new_n5335, new_n5334, new_n5336);
nand_1 g04960(new_n5336, new_n5331_1, new_n5337);
nand_1 g04961(new_n5337, new_n5330, new_n5338);
not_4  g04962(new_n5309, new_n5339);
xnor_1 g04963(new_n5339, new_n5308, new_n5340);
nand_1 g04964(new_n5340, new_n5338, new_n5341);
nand_1 g04965(new_n5341, new_n5311, new_n5342);
nand_1 g04966(new_n5342, new_n5306, new_n5343);
nand_1 g04967(new_n5030_1, new_n5029, new_n5344);
nand_1 g04968(new_n5344, new_n5091, new_n5345);
xnor_1 g04969(new_n5342, new_n5306, new_n5346);
not_4  g04970(new_n5346, new_n5347);
nand_1 g04971(new_n5347, new_n5345, new_n5348);
nand_1 g04972(new_n5348, new_n5343, new_n5349);
not_4  g04973(new_n5349, new_n5350);
nor_1  g04974(new_n5350, new_n5304, new_n5351);
nor_1  g04975(new_n5351, new_n5297, new_n5352);
nor_1  g04976(new_n5352, new_n5292, new_n5353);
nor_1  g04977(new_n5290, new_n5287, new_n5354);
nor_1  g04978(new_n5283_1, new_n5100, new_n5355);
nor_1  g04979(new_n5355, new_n5354, new_n5356);
nor_1  g04980(new_n5301, new_n5299, new_n5357);
nor_1  g04981(new_n5357, new_n5297, new_n5358);
nand_1 g04982(new_n5349, new_n5358, new_n5359);
nand_1 g04983(new_n5359, new_n5302, new_n5360);
nor_1  g04984(new_n5360, new_n5356, new_n5361);
nor_1  g04985(new_n5361, new_n5353, new_n5362);
nand_1 g04986(new_n5362, new_n4916, new_n5363);
not_4  g04987(new_n4916, new_n5364);
nand_1 g04988(new_n5360, new_n5356, new_n5365);
nand_1 g04989(new_n5352, new_n5292, new_n5366);
nand_1 g04990(new_n5366, new_n5365, new_n5367);
nand_1 g04991(new_n5367, new_n5364, new_n5368);
nand_1 g04992(new_n5368, new_n5363, new_n5369);
xnor_1 g04993(new_n4913, new_n4912, new_n5370);
not_4  g04994(new_n5370, new_n5371);
nand_1 g04995(new_n5350, new_n5304, new_n5372);
nand_1 g04996(new_n5372, new_n5359, new_n5373);
nor_1  g04997(new_n5373, new_n5371, new_n5374);
xnor_1 g04998(new_n4910, new_n4909, new_n5375);
xnor_1 g04999(new_n4907, new_n4900, new_n5376);
xnor_1 g05000(new_n5340, new_n5338, new_n5377);
nand_1 g05001(new_n5377, new_n5376, new_n5378);
not_4  g05002(new_n5376, new_n5379);
xnor_1 g05003(new_n5377, new_n5379, new_n5380);
xnor_1 g05004(new_n5336, new_n5331_1, new_n5381);
not_4  g05005(new_n5381, new_n5382);
not_4  g05006(new_n4903_1, new_n5383);
nand_1 g05007(new_n5383, new_n4837, new_n5384);
nand_1 g05008(new_n5384, new_n4905, new_n5385);
nor_1  g05009(new_n5385, new_n5382, new_n5386);
not_4  g05010(new_n5386, new_n5387);
xnor_1 g05011(new_n5385, new_n5381, new_n5388);
xnor_1 g05012(new_n5321, new_n5320_1, new_n5389);
nand_1 g05013(n9400, n6703, new_n5390);
nand_1 g05014(n9640, n6877, new_n5391);
xnor_1 g05015(new_n5391, new_n5390, new_n5392);
not_4  g05016(new_n5392, new_n5393);
nand_1 g05017(new_n5393, new_n5389, new_n5394);
not_4  g05018(new_n4902, new_n5395);
nand_1 g05019(new_n5318, new_n5171, new_n5396);
nand_1 g05020(new_n5396, new_n5320_1, new_n5397);
not_4  g05021(new_n5397, new_n5398);
nand_1 g05022(new_n5398, new_n5395, new_n5399);
not_4  g05023(new_n5399, new_n5400);
xnor_1 g05024(new_n5392, new_n5389, new_n5401);
nand_1 g05025(new_n5401, new_n5400, new_n5402);
nand_1 g05026(new_n5402, new_n5394, new_n5403);
nand_1 g05027(new_n5403, new_n5388, new_n5404);
nand_1 g05028(new_n5404, new_n5387, new_n5405);
nand_1 g05029(new_n5405, new_n5380, new_n5406);
nand_1 g05030(new_n5406, new_n5378, new_n5407);
nor_1  g05031(new_n5407, new_n5375, new_n5408);
not_4  g05032(new_n5408, new_n5409);
xnor_1 g05033(new_n5347, new_n5345, new_n5410);
not_4  g05034(new_n5410, new_n5411_1);
not_4  g05035(new_n5407, new_n5412);
xnor_1 g05036(new_n5412, new_n5375, new_n5413);
nand_1 g05037(new_n5413, new_n5411_1, new_n5414);
nand_1 g05038(new_n5414, new_n5409, new_n5415);
not_4  g05039(new_n5415, new_n5416);
nor_1  g05040(new_n5349, new_n5358, new_n5417);
nor_1  g05041(new_n5417, new_n5351, new_n5418);
nand_1 g05042(new_n5418, new_n5370, new_n5419);
nand_1 g05043(new_n5373, new_n5371, new_n5420);
nand_1 g05044(new_n5420, new_n5419, new_n5421);
nor_1  g05045(new_n5421, new_n5416, new_n5422);
nor_1  g05046(new_n5422, new_n5374, new_n5423);
nor_1  g05047(new_n5423, new_n5369, new_n5424);
nor_1  g05048(new_n5367, new_n5364, new_n5425);
nor_1  g05049(new_n5362, new_n4916, new_n5426);
nor_1  g05050(new_n5426, new_n5425, new_n5427);
nor_1  g05051(new_n5418, new_n5370, new_n5428);
nor_1  g05052(new_n5428, new_n5374, new_n5429);
nand_1 g05053(new_n5429, new_n5415, new_n5430);
nand_1 g05054(new_n5430, new_n5419, new_n5431);
nor_1  g05055(new_n5431, new_n5427, new_n5432);
nor_1  g05056(new_n5432, new_n5424, new_n5433);
nor_1  g05057(new_n5433, new_n4783, new_n5434);
not_4  g05058(new_n4783, new_n5435_1);
nand_1 g05059(new_n5431, new_n5427, new_n5436);
nand_1 g05060(new_n5423, new_n5369, new_n5437);
nand_1 g05061(new_n5437, new_n5436, new_n5438);
nand_1 g05062(new_n5438, new_n5435_1, new_n5439);
nand_1 g05063(new_n5433, new_n4783, new_n5440);
nand_1 g05064(new_n5440, new_n5439, new_n5441);
xnor_1 g05065(new_n4780, new_n4778, new_n5442);
not_4  g05066(new_n5442, new_n5443);
nor_1  g05067(new_n5429, new_n5415, new_n5444);
nor_1  g05068(new_n5444, new_n5422, new_n5445);
nor_1  g05069(new_n5445, new_n5443, new_n5446);
not_4  g05070(new_n4777, new_n5447);
xnor_1 g05071(new_n5447, new_n4776, new_n5448);
not_4  g05072(new_n5448, new_n5449);
xnor_1 g05073(new_n5413, new_n5410, new_n5450);
nand_1 g05074(new_n5450, new_n5449, new_n5451);
xnor_1 g05075(new_n5450, new_n5448, new_n5452);
not_4  g05076(new_n5452, new_n5453);
xnor_1 g05077(new_n4774, new_n4766, new_n5454);
not_4  g05078(new_n5454, new_n5455);
not_4  g05079(new_n5405, new_n5456);
xnor_1 g05080(new_n5456, new_n5380, new_n5457);
nor_1  g05081(new_n5457, new_n5455, new_n5458);
xnor_1 g05082(new_n5403, new_n5388, new_n5459);
nand_1 g05083(n7862, n1798, new_n5460);
nand_1 g05084(new_n5460, new_n4708, new_n5461);
nand_1 g05085(new_n5461, new_n4767, new_n5462);
not_4  g05086(new_n5461, new_n5463);
nand_1 g05087(new_n5463, new_n4706, new_n5464);
nand_1 g05088(new_n5464, new_n5462, new_n5465);
nand_1 g05089(new_n5465, new_n5459, new_n5466);
xnor_1 g05090(new_n5465, new_n5459, new_n5467);
not_4  g05091(new_n5460, new_n5468);
xnor_1 g05092(new_n5398, new_n4902, new_n5469);
nand_1 g05093(new_n5469, new_n5468, new_n5470);
nand_1 g05094(new_n4771, new_n4769, new_n5471);
nand_1 g05095(new_n5471, new_n4773, new_n5472);
nand_1 g05096(new_n5472, new_n5470, new_n5473);
xnor_1 g05097(new_n5401, new_n5399, new_n5474);
xnor_1 g05098(new_n5472, new_n5470, new_n5475);
nor_1  g05099(new_n5475, new_n5474, new_n5476);
not_4  g05100(new_n5476, new_n5477);
nand_1 g05101(new_n5477, new_n5473, new_n5478);
not_4  g05102(new_n5478, new_n5479);
nor_1  g05103(new_n5479, new_n5467, new_n5480);
not_4  g05104(new_n5480, new_n5481);
nand_1 g05105(new_n5481, new_n5466, new_n5482);
not_4  g05106(new_n5482, new_n5483);
xnor_1 g05107(new_n5457, new_n5455, new_n5484);
nor_1  g05108(new_n5484, new_n5483, new_n5485);
nor_1  g05109(new_n5485, new_n5458, new_n5486);
nor_1  g05110(new_n5486, new_n5453, new_n5487);
not_4  g05111(new_n5487, new_n5488);
nand_1 g05112(new_n5488, new_n5451, new_n5489);
nand_1 g05113(new_n5421, new_n5416, new_n5490);
nand_1 g05114(new_n5490, new_n5430, new_n5491);
nand_1 g05115(new_n5491, new_n5442, new_n5492);
nand_1 g05116(new_n5445, new_n5443, new_n5493);
nand_1 g05117(new_n5493, new_n5492, new_n5494);
nor_1  g05118(new_n5494, new_n5489, new_n5495);
nor_1  g05119(new_n5495, new_n5446, new_n5496);
nor_1  g05120(new_n5496, new_n5441, new_n5497);
nor_1  g05121(new_n5497, new_n5434, new_n5498);
not_4  g05122(new_n4853, new_n5499);
nand_1 g05123(new_n4893, new_n5499, new_n5500);
nand_1 g05124(new_n4915, new_n4894, new_n5501);
nand_1 g05125(new_n5501, new_n5500, new_n5502);
nand_1 g05126(n7862, n753, new_n5503);
not_4  g05127(new_n5045, new_n5504);
nand_1 g05128(new_n5051, new_n5504, new_n5505);
not_4  g05129(new_n5069_1, new_n5506);
nand_1 g05130(new_n5506, new_n5052, new_n5507);
nand_1 g05131(new_n5507, new_n5505, new_n5508);
xnor_1 g05132(new_n5508, new_n5503, new_n5509);
nand_1 g05133(new_n5067, new_n5061, new_n5510);
nand_1 g05134(new_n5510, new_n5059, new_n5511);
nand_1 g05135(n3146, n1067, new_n5512);
nand_1 g05136(n2551, n137, new_n5513);
xnor_1 g05137(new_n5513, new_n5512, new_n5514);
nand_1 g05138(n12826, n5283, new_n5515);
nand_1 g05139(n8665, n6797, new_n5516);
not_4  g05140(new_n5516, new_n5517);
xnor_1 g05141(new_n5517, new_n5515, new_n5518);
xnor_1 g05142(new_n5518, new_n5514, new_n5519);
xnor_1 g05143(new_n5519, new_n5511, new_n5520);
nand_1 g05144(new_n5210, new_n5204, new_n5521);
nand_1 g05145(new_n5521, new_n5201, new_n5522);
nand_1 g05146(new_n5219, new_n5218, new_n5523);
nand_1 g05147(new_n5221, new_n5217, new_n5524);
nand_1 g05148(new_n5524, new_n5523, new_n5525);
nand_1 g05149(n8384, n1510, new_n5526);
nand_1 g05150(n5198, n2749, new_n5527);
not_4  g05151(new_n5527, new_n5528);
xnor_1 g05152(new_n5528, new_n5526, new_n5529);
xnor_1 g05153(new_n5529, new_n5525, new_n5530);
xnor_1 g05154(new_n5530, new_n5522, new_n5531);
xnor_1 g05155(new_n5531, new_n5520, new_n5532);
xnor_1 g05156(new_n5532, new_n5509, new_n5533);
xnor_1 g05157(new_n5533, new_n5502, new_n5534);
nand_1 g05158(new_n4757_1, new_n4756, new_n5535);
not_4  g05159(new_n4753, new_n5536);
nand_1 g05160(new_n4759, new_n5536, new_n5537);
nand_1 g05161(new_n5537, new_n5535, new_n5538);
nand_1 g05162(new_n5077, new_n5073, new_n5539);
xnor_1 g05163(new_n5539, new_n5538, new_n5540);
nand_1 g05164(n12511, n7236, new_n5541);
nand_1 g05165(n6826, n1798, new_n5542);
xnor_1 g05166(new_n5542, new_n5541, new_n5543);
nand_1 g05167(new_n5064, new_n5063, new_n5544);
nand_1 g05168(new_n5066, new_n5062, new_n5545);
nand_1 g05169(new_n5545, new_n5544, new_n5546);
nand_1 g05170(new_n5207, new_n5206, new_n5547);
nand_1 g05171(new_n5209, new_n5205, new_n5548);
nand_1 g05172(new_n5548, new_n5547, new_n5549);
xnor_1 g05173(new_n5549, new_n5546, new_n5550);
xnor_1 g05174(new_n5550, new_n5543, new_n5551);
nand_1 g05175(n6358, n159, new_n5552);
nand_1 g05176(new_n5044, new_n5040, new_n5553);
nand_1 g05177(new_n5553, new_n5042, new_n5554);
nand_1 g05178(n11478, n4094, new_n5555);
nor_1  g05179(new_n5555, new_n5554, new_n5556);
not_4  g05180(new_n5554, new_n5557);
nor_1  g05181(new_n5555, new_n4918, new_n5558);
nor_1  g05182(new_n5558, new_n5557, new_n5559);
nor_1  g05183(new_n5559, new_n5556, new_n5560);
xnor_1 g05184(new_n5560, new_n5552, new_n5561);
xnor_1 g05185(new_n5561, new_n5551, new_n5562);
xnor_1 g05186(new_n5562, new_n5540, new_n5563);
xnor_1 g05187(new_n5563, new_n5534, new_n5564);
nor_1  g05188(new_n5243, new_n5233, new_n5565);
nand_1 g05189(n5645, n4938, new_n5566);
nand_1 g05190(n10898, n7646, new_n5567);
xnor_1 g05191(new_n5567, new_n5566, new_n5568);
xnor_1 g05192(new_n5568, new_n5565, new_n5569);
xnor_1 g05193(new_n5569, new_n5564, new_n5570);
nand_1 g05194(new_n5365, new_n5284, new_n5571);
nand_1 g05195(n11922, n6294, new_n5572);
nand_1 g05196(new_n5090, new_n5096, new_n5573);
xnor_1 g05197(new_n5573, new_n5572, new_n5574);
not_4  g05198(new_n4721, new_n5575);
nand_1 g05199(new_n4760, new_n5575, new_n5576);
nand_1 g05200(new_n4782, new_n4761, new_n5577);
nand_1 g05201(new_n5577, new_n5576, new_n5578);
nand_1 g05202(new_n4890, new_n4888, new_n5579_1);
not_4  g05203(new_n4885, new_n5580);
nand_1 g05204(new_n4892, new_n5580, new_n5581);
nand_1 g05205(new_n5581, new_n5579_1, new_n5582);
not_4  g05206(new_n4855, new_n5583);
nand_1 g05207(new_n4864, new_n5583, new_n5584);
not_4  g05208(new_n4884, new_n5585);
nand_1 g05209(new_n5585, new_n4865, new_n5586);
nand_1 g05210(new_n5586, new_n5584, new_n5587);
not_4  g05211(new_n4874, new_n5588);
nand_1 g05212(new_n4877, new_n5588, new_n5589);
nand_1 g05213(new_n5589, new_n4880, new_n5590);
nand_1 g05214(n4203, n3022, new_n5591);
nand_1 g05215(n11023, n4187, new_n5592);
xnor_1 g05216(new_n5592, new_n5591, new_n5593);
xnor_1 g05217(new_n5593, new_n5590, new_n5594);
nand_1 g05218(n7456, n5240, new_n5595);
nand_1 g05219(n12753, n9640, new_n5596);
not_4  g05220(new_n5596, new_n5597);
xnor_1 g05221(new_n5597, new_n5595, new_n5598);
nand_1 g05222(n9583, n1333, new_n5599);
nand_1 g05223(n12591, n11821, new_n5600);
xnor_1 g05224(new_n5600, new_n5599, new_n5601);
xnor_1 g05225(new_n5601, new_n5598, new_n5602);
xnor_1 g05226(new_n5602, new_n5594, new_n5603);
xnor_1 g05227(new_n5603, new_n5587, new_n5604);
not_4  g05228(new_n4727, new_n5605);
nand_1 g05229(new_n4734, new_n5605, new_n5606);
not_4  g05230(new_n4752, new_n5607);
nand_1 g05231(new_n5607, new_n4735, new_n5608);
nand_1 g05232(new_n5608, new_n5606, new_n5609);
nand_1 g05233(n9080, n3932, new_n5610);
nand_1 g05234(n10174, n6703, new_n5611);
nand_1 g05235(n6877, n2278, new_n5612);
xnor_1 g05236(new_n5612, new_n5611, new_n5613);
xnor_1 g05237(new_n5613, new_n5610, new_n5614);
xnor_1 g05238(new_n5614, new_n5609, new_n5615);
xnor_1 g05239(new_n5615, new_n5604, new_n5616);
xnor_1 g05240(new_n5616, new_n5582, new_n5617);
xnor_1 g05241(new_n5617, new_n5578, new_n5618);
xnor_1 g05242(new_n5618, new_n5574, new_n5619);
xnor_1 g05243(new_n5619, new_n5571, new_n5620);
xnor_1 g05244(new_n5620, new_n5570, new_n5621);
nand_1 g05245(new_n5621, new_n5498, new_n5622);
nor_1  g05246(new_n5438, new_n5435_1, new_n5623);
nor_1  g05247(new_n5623, new_n5434, new_n5624);
not_4  g05248(new_n5489, new_n5625);
nor_1  g05249(new_n5491, new_n5442, new_n5626);
nor_1  g05250(new_n5626, new_n5446, new_n5627);
nand_1 g05251(new_n5627, new_n5625, new_n5628);
nand_1 g05252(new_n5628, new_n5492, new_n5629);
nand_1 g05253(new_n5629, new_n5624, new_n5630);
nand_1 g05254(new_n5630, new_n5439, new_n5631);
not_4  g05255(new_n5621, new_n5632);
nand_1 g05256(new_n5632, new_n5631, new_n5633);
nand_1 g05257(new_n5633, new_n5622, new_n5634);
not_4  g05258(new_n5222, new_n5635);
nand_1 g05259(new_n5635, new_n5216, new_n5636);
not_4  g05260(new_n5212_1, new_n5637);
nand_1 g05261(new_n5223, new_n5637, new_n5638);
nand_1 g05262(new_n5638, new_n5636, new_n5639);
not_4  g05263(new_n4741, new_n5640);
nand_1 g05264(new_n4751, new_n5640, new_n5641_1);
nand_1 g05265(new_n5641_1, new_n4739, new_n5642);
not_4  g05266(new_n4856, new_n5643);
nand_1 g05267(new_n4862, new_n5643, new_n5644);
nand_1 g05268(new_n5644, new_n4861, new_n5645_1);
xnor_1 g05269(new_n5645_1, new_n5642, new_n5646);
nand_1 g05270(new_n4731, new_n4730, new_n5647);
nand_1 g05271(new_n4733_1, new_n4728, new_n5648);
nand_1 g05272(new_n5648, new_n5647, new_n5649);
not_4  g05273(new_n4742, new_n5650);
nand_1 g05274(new_n4745, new_n5650, new_n5651);
nand_1 g05275(new_n5651, new_n4748, new_n5652);
nand_1 g05276(n10278, n2464, new_n5653);
nand_1 g05277(n11757, n11662, new_n5654);
xnor_1 g05278(new_n5654, new_n5653, new_n5655);
nand_1 g05279(n10327, n3172, new_n5656);
nand_1 g05280(n11423, n9400, new_n5657);
xnor_1 g05281(new_n5657, new_n5656, new_n5658);
xnor_1 g05282(new_n5658, new_n5655, new_n5659);
xnor_1 g05283(new_n5659, new_n5652, new_n5660);
xnor_1 g05284(new_n5660, new_n5649, new_n5661);
xnor_1 g05285(new_n5661, new_n5646, new_n5662);
xnor_1 g05286(new_n5662, new_n5639, new_n5663);
nand_1 g05287(n3754, n1471, new_n5664);
nand_1 g05288(n11311, n10451, new_n5665);
xnor_1 g05289(new_n5665, new_n5664, new_n5666);
not_4  g05290(new_n4873, new_n5667);
nand_1 g05291(new_n4883, new_n5667, new_n5668);
nand_1 g05292(new_n5668, new_n4871, new_n5669);
nand_1 g05293(n11876, n4722, new_n5670_1);
nand_1 g05294(n10685, n4805, new_n5671);
nand_1 g05295(n12247, n3992, new_n5672);
xnor_1 g05296(new_n5672, new_n5671, new_n5673);
xnor_1 g05297(new_n5673, new_n5670_1, new_n5674);
xnor_1 g05298(new_n5674, new_n5669, new_n5675);
xnor_1 g05299(new_n5675, new_n5666, new_n5676);
xnor_1 g05300(new_n5676, new_n5663, new_n5677);
nand_1 g05301(new_n5273, new_n5274, new_n5678);
nor_1  g05302(new_n5424, new_n5425, new_n5679);
xnor_1 g05303(new_n5679, new_n5678, new_n5680);
xnor_1 g05304(new_n5680, new_n5677, new_n5681);
nand_1 g05305(new_n5681, new_n5634, new_n5682);
nor_1  g05306(new_n5632, new_n5631, new_n5683);
nor_1  g05307(new_n5621, new_n5498, new_n5684);
nor_1  g05308(new_n5684, new_n5683, new_n5685);
not_4  g05309(new_n5681, new_n5686);
nand_1 g05310(new_n5686, new_n5685, new_n5687);
nand_1 g05311(new_n5687, new_n5682, n1269);
nand_1 g05312(n10223, n4312, new_n5689);
nand_1 g05313(n12705, n7265, new_n5690);
not_4  g05314(new_n5690, new_n5691);
nand_1 g05315(n4312, n2879, new_n5692);
xnor_1 g05316(new_n5691, new_n1103, new_n5693_1);
nand_1 g05317(new_n5693_1, new_n5692, new_n5694_1);
nand_1 g05318(new_n5694_1, new_n5691, new_n5695);
nand_1 g05319(new_n5695, new_n5689, new_n5696);
not_4  g05320(new_n5689, new_n5697);
nand_1 g05321(new_n5695, new_n1113, new_n5698);
nand_1 g05322(new_n5698, new_n5697, new_n5699);
nand_1 g05323(new_n5699, new_n5696, new_n5700);
nand_1 g05324(n12025, n7265, new_n5701);
nand_1 g05325(n12705, n2879, new_n5702);
nand_1 g05326(new_n5702, new_n5701, new_n5703);
not_4  g05327(new_n5701, new_n5704);
not_4  g05328(new_n5702, new_n5705);
nand_1 g05329(new_n5705, new_n5704, new_n5706);
nand_1 g05330(new_n5706, new_n5703, new_n5707);
nand_1 g05331(new_n5707, new_n5700, new_n5708);
nor_1  g05332(new_n5707, new_n5700, new_n5709);
not_4  g05333(new_n5709, new_n5710);
nand_1 g05334(new_n5710, new_n5708, new_n5711);
nand_1 g05335(n9195, n5964, new_n5712);
nand_1 g05336(n4634, n1097, new_n5713);
not_4  g05337(new_n5713, new_n5714);
xnor_1 g05338(new_n5714, new_n5712, new_n5715);
xnor_1 g05339(new_n5715, new_n5711, new_n5716);
nand_1 g05340(n5964, n4634, new_n5717);
nand_1 g05341(new_n1119, new_n1113, new_n5718);
nand_1 g05342(new_n5718, new_n1117, new_n5719);
nor_1  g05343(new_n5719, new_n5717, new_n5720);
not_4  g05344(new_n5720, new_n5721);
xnor_1 g05345(new_n5693_1, new_n5692, new_n5722);
nand_1 g05346(new_n5719, new_n5717, new_n5723);
nand_1 g05347(new_n5723, new_n5721, new_n5724);
not_4  g05348(new_n5724, new_n5725);
nand_1 g05349(new_n5725, new_n5722, new_n5726);
nand_1 g05350(new_n5726, new_n5721, new_n5727);
nand_1 g05351(new_n5727, new_n5716, new_n5728);
not_4  g05352(new_n5728, new_n5729);
nor_1  g05353(new_n5727, new_n5716, new_n5730);
nor_1  g05354(new_n5730, new_n5729, new_n5731);
nand_1 g05355(n9195, n5305, new_n5732);
not_4  g05356(new_n1112, new_n5733);
nand_1 g05357(new_n1121, new_n5733, new_n5734);
nand_1 g05358(new_n5734, new_n1110, new_n5735);
not_4  g05359(new_n5735, new_n5736);
nand_1 g05360(new_n5736, new_n5732, new_n5737);
not_4  g05361(new_n5722, new_n5738);
xnor_1 g05362(new_n5725, new_n5738, new_n5739);
not_4  g05363(new_n5739, new_n5740);
xnor_1 g05364(new_n5735, new_n5732, new_n5741);
nand_1 g05365(new_n5741, new_n5740, new_n5742);
nand_1 g05366(new_n5742, new_n5737, new_n5743);
not_4  g05367(new_n5743, new_n5744);
nand_1 g05368(new_n5744, new_n5731, new_n5745);
nand_1 g05369(new_n5710, new_n5699, new_n5746);
nand_1 g05370(n5964, n2253, new_n5747);
nand_1 g05371(n9195, n1097, new_n5748);
nand_1 g05372(n5305, n3865, new_n5749);
not_4  g05373(new_n5749, new_n5750);
xnor_1 g05374(new_n5750, new_n5748, new_n5751);
not_4  g05375(new_n5751, new_n5752);
xnor_1 g05376(new_n5752, new_n5747, new_n5753);
xnor_1 g05377(new_n5753, new_n5746, new_n5754);
nand_1 g05378(n4634, n4312, new_n5755);
nand_1 g05379(new_n5755, new_n5706, new_n5756);
not_4  g05380(new_n5706, new_n5757);
not_4  g05381(new_n5755, new_n5758);
nand_1 g05382(new_n5758, new_n5757, new_n5759);
nand_1 g05383(new_n5759, new_n5756, new_n5760_1);
not_4  g05384(new_n5760_1, new_n5761);
nand_1 g05385(n12025, n2879, new_n5762);
nand_1 g05386(n11257, n7265, new_n5763);
nand_1 g05387(n12705, n10223, new_n5764);
not_4  g05388(new_n5764, new_n5765);
xnor_1 g05389(new_n5765, new_n5763, new_n5766);
xnor_1 g05390(new_n5766, new_n5762, new_n5767_1);
not_4  g05391(new_n5767_1, new_n5768);
xnor_1 g05392(new_n5768, new_n5761, new_n5769);
xnor_1 g05393(new_n5769, new_n5754, new_n5770);
not_4  g05394(new_n5711, new_n5771);
nand_1 g05395(new_n5715, new_n5771, new_n5772);
nor_1  g05396(new_n5713, new_n5712, new_n5773);
xnor_1 g05397(new_n5729, new_n5773, new_n5774);
nand_1 g05398(new_n5774, new_n5772, new_n5775);
xnor_1 g05399(new_n5775, new_n5770, new_n5776);
xnor_1 g05400(new_n5776, new_n5745, new_n5777);
nand_1 g05401(n5305, n2253, new_n5778);
not_4  g05402(new_n5778, new_n5779);
xnor_1 g05403(new_n5743, new_n5731, new_n5780);
nand_1 g05404(new_n5780, new_n5779, new_n5781);
not_4  g05405(new_n1128, new_n5782);
nand_1 g05406(new_n5782, new_n1122, new_n5783);
xnor_1 g05407(new_n5741, new_n5739, new_n5784);
nor_1  g05408(new_n5784, new_n5783, new_n5785);
xnor_1 g05409(new_n5780, new_n5778, new_n5786);
nand_1 g05410(new_n5786, new_n5785, new_n5787);
nand_1 g05411(new_n5787, new_n5781, new_n5788);
xnor_1 g05412(new_n5788, new_n5777, new_n5789);
xnor_1 g05413(new_n5786, new_n5785, new_n5790);
not_4  g05414(new_n1266, new_n5791);
nand_1 g05415(n12145, n8759, new_n5792);
nor_1  g05416(new_n1245, new_n1243, new_n5793);
nor_1  g05417(new_n1258, new_n5793, new_n5794);
not_4  g05418(new_n5794, new_n5795);
xnor_1 g05419(new_n5795, new_n5792, new_n5796);
nand_1 g05420(n6776, n2522, new_n5797);
nand_1 g05421(new_n1254, new_n1247, new_n5798_1);
nand_1 g05422(new_n5798_1, new_n1251, new_n5799);
not_4  g05423(new_n5799, new_n5800);
xnor_1 g05424(new_n5800, new_n5797, new_n5801);
not_4  g05425(new_n5801, new_n5802);
nand_1 g05426(n7436, n2024, new_n5803);
nand_1 g05427(n12299, n9189, new_n5804);
nand_1 g05428(n8276, n7946, new_n5805);
not_4  g05429(new_n5805, new_n5806);
xnor_1 g05430(new_n5806, new_n5804, new_n5807);
xnor_1 g05431(new_n5807, new_n5803, new_n5808);
xnor_1 g05432(new_n5808, new_n5802, new_n5809);
xnor_1 g05433(new_n5809, new_n5796, new_n5810);
not_4  g05434(new_n5810, new_n5811);
nand_1 g05435(new_n5811, new_n5791, new_n5812);
nand_1 g05436(n12221, n8759, new_n5813);
nor_1  g05437(new_n5799, new_n5797, new_n5814_1);
not_4  g05438(new_n5814_1, new_n5815);
nand_1 g05439(new_n5808, new_n5801, new_n5816);
nand_1 g05440(new_n5816, new_n5815, new_n5817);
nand_1 g05441(n12145, n6776, new_n5818);
nand_1 g05442(n12299, n2522, new_n5819);
not_4  g05443(new_n5819, new_n5820);
xnor_1 g05444(new_n5820, new_n5818, new_n5821);
xnor_1 g05445(new_n5821, new_n5817, new_n5822);
nand_1 g05446(n9189, n7436, new_n5823);
nand_1 g05447(new_n5807, new_n5803, new_n5824);
nand_1 g05448(new_n5824, new_n5806, new_n5825);
nand_1 g05449(new_n5825, new_n5823, new_n5826);
not_4  g05450(new_n5823, new_n5827);
nand_1 g05451(new_n5825, new_n1247, new_n5828);
nand_1 g05452(new_n5828, new_n5827, new_n5829);
nand_1 g05453(new_n5829, new_n5826, new_n5830);
not_4  g05454(new_n5830, new_n5831);
nand_1 g05455(n8276, n2024, new_n5832);
nand_1 g05456(n9241, n7946, new_n5833);
nand_1 g05457(new_n5833, new_n5832, new_n5834);
not_4  g05458(new_n5832, new_n5835);
not_4  g05459(new_n5833, new_n5836);
nand_1 g05460(new_n5836, new_n5835, new_n5837);
nand_1 g05461(new_n5837, new_n5834, new_n5838);
not_4  g05462(new_n5838, new_n5839);
xnor_1 g05463(new_n5839, new_n5831, new_n5840);
xnor_1 g05464(new_n5840, new_n5822, new_n5841);
nor_1  g05465(new_n5794, new_n5792, new_n5842);
not_4  g05466(new_n5842, new_n5843);
nand_1 g05467(new_n5809, new_n5796, new_n5844);
nand_1 g05468(new_n5844, new_n5843, new_n5845);
xnor_1 g05469(new_n5845, new_n5841, new_n5846);
xnor_1 g05470(new_n5846, new_n5813, new_n5847);
xnor_1 g05471(new_n5847, new_n5812, new_n5848);
xnor_1 g05472(new_n5811, new_n1266, new_n5849);
not_4  g05473(new_n1289, new_n5850);
nand_1 g05474(new_n1290, new_n5850, new_n5851);
nand_1 g05475(n6016, n5331, new_n5852);
nand_1 g05476(n8476, n521, new_n5853);
nor_1  g05477(new_n1284, new_n1283, new_n5854);
nor_1  g05478(new_n1281, new_n1280, new_n5855);
nor_1  g05479(new_n5855, new_n5854, new_n5856);
nand_1 g05480(new_n5856, new_n1279, new_n5857_1);
nand_1 g05481(new_n5857_1, new_n1282, new_n5858);
nor_1  g05482(new_n5858, new_n5853, new_n5859);
not_4  g05483(new_n5853, new_n5860_1);
not_4  g05484(new_n1279, new_n5861);
nor_1  g05485(new_n1286, new_n5861, new_n5862);
nor_1  g05486(new_n5862, new_n5854, new_n5863);
nor_1  g05487(new_n5863, new_n5860_1, new_n5864);
nor_1  g05488(new_n5864, new_n5859, new_n5865);
nand_1 g05489(n12648, n2498, new_n5866);
nand_1 g05490(n10545, n2558, new_n5867);
nand_1 g05491(new_n5867, new_n1213, new_n5868);
not_4  g05492(new_n5867, new_n5869);
nand_1 g05493(new_n5869, new_n1214, new_n5870);
nand_1 g05494(new_n5870, new_n5868, new_n5871);
xnor_1 g05495(new_n5871, new_n5866, new_n5872);
not_4  g05496(new_n5872, new_n5873);
nand_1 g05497(new_n5873, new_n5865, new_n5874);
nand_1 g05498(new_n5863, new_n5860_1, new_n5875);
nand_1 g05499(new_n5858, new_n5853, new_n5876);
nand_1 g05500(new_n5876, new_n5875, new_n5877);
nand_1 g05501(new_n5872, new_n5877, new_n5878);
nand_1 g05502(new_n5878, new_n5874, new_n5879);
nor_1  g05503(new_n5879, new_n5852, new_n5880);
not_4  g05504(new_n5852, new_n5881);
nor_1  g05505(new_n5872, new_n5877, new_n5882);
nor_1  g05506(new_n5873, new_n5865, new_n5883);
nor_1  g05507(new_n5883, new_n5882, new_n5884);
nor_1  g05508(new_n5884, new_n5881, new_n5885);
nor_1  g05509(new_n5885, new_n5880, new_n5886);
nor_1  g05510(new_n1276, new_n1274, new_n5887);
not_4  g05511(new_n5887, new_n5888);
nand_1 g05512(new_n1288, new_n1278, new_n5889);
nand_1 g05513(new_n5889, new_n5888, new_n5890);
nand_1 g05514(new_n5890, new_n5886, new_n5891);
nand_1 g05515(new_n5884, new_n5881, new_n5892);
nand_1 g05516(new_n5879, new_n5852, new_n5893);
nand_1 g05517(new_n5893, new_n5892, new_n5894);
not_4  g05518(new_n5890, new_n5895);
nand_1 g05519(new_n5895, new_n5894, new_n5896);
nand_1 g05520(new_n5896, new_n5891, new_n5897);
nor_1  g05521(new_n5897, new_n5851, new_n5898);
not_4  g05522(new_n5851, new_n5899);
nor_1  g05523(new_n5895, new_n5894, new_n5900);
nor_1  g05524(new_n5890, new_n5886, new_n5901);
nor_1  g05525(new_n5901, new_n5900, new_n5902);
nor_1  g05526(new_n5902, new_n5899, new_n5903);
nor_1  g05527(new_n5903, new_n5898, new_n5904);
not_4  g05528(new_n1308, new_n5905);
nand_1 g05529(new_n5905, new_n1307, new_n5906);
nand_1 g05530(n7965, n7270, new_n5907);
nand_1 g05531(n7388, n806, new_n5908);
nor_1  g05532(new_n1302, new_n1301, new_n5909);
nor_1  g05533(new_n1299, new_n1298, new_n5910);
nor_1  g05534(new_n5910, new_n5909, new_n5911);
nand_1 g05535(new_n5911, new_n1297, new_n5912);
nand_1 g05536(new_n5912, new_n1300, new_n5913);
nor_1  g05537(new_n5913, new_n5908, new_n5914);
not_4  g05538(new_n5908, new_n5915);
not_4  g05539(new_n1297, new_n5916);
nor_1  g05540(new_n1304, new_n5916, new_n5917);
nor_1  g05541(new_n5917, new_n5909, new_n5918);
nor_1  g05542(new_n5918, new_n5915, new_n5919);
nor_1  g05543(new_n5919, new_n5914, new_n5920);
nand_1 g05544(n9111, n2393, new_n5921);
nand_1 g05545(n9763, n5860, new_n5922);
nand_1 g05546(new_n5922, new_n1191, new_n5923);
not_4  g05547(new_n5922, new_n5924);
nand_1 g05548(new_n5924, new_n1192, new_n5925);
nand_1 g05549(new_n5925, new_n5923, new_n5926);
xnor_1 g05550(new_n5926, new_n5921, new_n5927);
not_4  g05551(new_n5927, new_n5928);
nand_1 g05552(new_n5928, new_n5920, new_n5929);
nand_1 g05553(new_n5918, new_n5915, new_n5930);
nand_1 g05554(new_n5913, new_n5908, new_n5931);
nand_1 g05555(new_n5931, new_n5930, new_n5932);
nand_1 g05556(new_n5927, new_n5932, new_n5933);
nand_1 g05557(new_n5933, new_n5929, new_n5934_1);
nor_1  g05558(new_n5934_1, new_n5907, new_n5935);
not_4  g05559(new_n5907, new_n5936);
nor_1  g05560(new_n5927, new_n5932, new_n5937);
nor_1  g05561(new_n5928, new_n5920, new_n5938);
nor_1  g05562(new_n5938, new_n5937, new_n5939);
nor_1  g05563(new_n5939, new_n5936, new_n5940);
nor_1  g05564(new_n5940, new_n5935, new_n5941);
not_4  g05565(new_n1292, new_n5942);
nand_1 g05566(new_n1294, new_n5942, new_n5943);
nor_1  g05567(new_n1305, new_n1296, new_n5944);
not_4  g05568(new_n5944, new_n5945);
nand_1 g05569(new_n5945, new_n5943, new_n5946);
nand_1 g05570(new_n5946, new_n5941, new_n5947);
nand_1 g05571(new_n5939, new_n5936, new_n5948);
nand_1 g05572(new_n5934_1, new_n5907, new_n5949);
nand_1 g05573(new_n5949, new_n5948, new_n5950);
not_4  g05574(new_n5946, new_n5951);
nand_1 g05575(new_n5951, new_n5950, new_n5952);
nand_1 g05576(new_n5952, new_n5947, new_n5953);
nor_1  g05577(new_n5953, new_n5906, new_n5954);
not_4  g05578(new_n5906, new_n5955);
nor_1  g05579(new_n5951, new_n5950, new_n5956);
nor_1  g05580(new_n5946, new_n5941, new_n5957);
nor_1  g05581(new_n5957, new_n5956, new_n5958);
nor_1  g05582(new_n5958, new_n5955, new_n5959);
nor_1  g05583(new_n5959, new_n5954, new_n5960);
nand_1 g05584(new_n5960, new_n5904, new_n5961);
nand_1 g05585(new_n5902, new_n5899, new_n5962);
nand_1 g05586(new_n5897, new_n5851, new_n5963);
nand_1 g05587(new_n5963, new_n5962, new_n5964_1);
nand_1 g05588(new_n5958, new_n5955, new_n5965);
nand_1 g05589(new_n5953, new_n5906, new_n5966);
nand_1 g05590(new_n5966, new_n5965, new_n5967);
nand_1 g05591(new_n5967, new_n5964_1, new_n5968);
nand_1 g05592(new_n5968, new_n5961, new_n5969);
nand_1 g05593(new_n1322, new_n1312, new_n5970);
not_4  g05594(new_n5970, new_n5971);
nand_1 g05595(new_n5971, new_n5969, new_n5972);
nor_1  g05596(new_n5967, new_n5964_1, new_n5973);
nor_1  g05597(new_n5960, new_n5904, new_n5974);
nor_1  g05598(new_n5974, new_n5973, new_n5975);
nand_1 g05599(new_n5970, new_n5975, new_n5976);
nand_1 g05600(new_n5976, new_n5972, new_n5977);
nand_1 g05601(new_n5977, new_n5849, new_n5978);
nor_1  g05602(new_n1271, new_n1267, new_n5979);
not_4  g05603(new_n5979, new_n5980);
nand_1 g05604(new_n1323, new_n1273, new_n5981);
nand_1 g05605(new_n5981, new_n5980, new_n5982);
not_4  g05606(new_n5849, new_n5983);
nor_1  g05607(new_n5970, new_n5975, new_n5984);
nor_1  g05608(new_n5971, new_n5969, new_n5985);
nor_1  g05609(new_n5985, new_n5984, new_n5986);
nor_1  g05610(new_n5986, new_n5983, new_n5987);
nor_1  g05611(new_n5977, new_n5849, new_n5988);
nor_1  g05612(new_n5988, new_n5987, new_n5989);
nand_1 g05613(new_n5989, new_n5982, new_n5990);
nand_1 g05614(new_n5990, new_n5978, new_n5991);
nor_1  g05615(new_n5991, new_n5848, new_n5992);
not_4  g05616(new_n5848, new_n5993);
not_4  g05617(new_n5982, new_n5994);
nand_1 g05618(new_n5986, new_n5983, new_n5995);
nand_1 g05619(new_n5995, new_n5978, new_n5996);
nor_1  g05620(new_n5996, new_n5994, new_n5997);
nor_1  g05621(new_n5997, new_n5987, new_n5998);
nor_1  g05622(new_n5998, new_n5993, new_n5999);
nor_1  g05623(new_n5999, new_n5992, new_n6000);
nand_1 g05624(n5798, n5331, new_n6001);
nand_1 g05625(n12648, n5579, new_n6002);
nand_1 g05626(n10545, n2498, new_n6003);
nand_1 g05627(n7690, n2558, new_n6004);
not_4  g05628(new_n6004, new_n6005);
xnor_1 g05629(new_n6005, new_n6003, new_n6006);
not_4  g05630(new_n6006, new_n6007);
xnor_1 g05631(new_n6007, new_n6002, new_n6008);
nand_1 g05632(new_n5870, new_n5866, new_n6009);
nand_1 g05633(new_n6009, new_n5868, new_n6010);
xnor_1 g05634(new_n6010, new_n6008, new_n6011);
nand_1 g05635(n8476, n6016, new_n6012);
nand_1 g05636(n2530, n521, new_n6013);
not_4  g05637(new_n6013, new_n6014);
xnor_1 g05638(new_n6014, new_n6012, new_n6015);
xnor_1 g05639(new_n6015, new_n6011, new_n6016_1);
nor_1  g05640(new_n5882, new_n5859, new_n6017);
xnor_1 g05641(new_n6017, new_n6016_1, new_n6018);
nor_1  g05642(new_n5900, new_n5880, new_n6019);
xnor_1 g05643(new_n6019, new_n6018, new_n6020);
xnor_1 g05644(new_n6020, new_n6001, new_n6021);
xnor_1 g05645(new_n6021, new_n5962, new_n6022);
nand_1 g05646(n7965, n5153, new_n6023);
nand_1 g05647(n3342, n2393, new_n6024);
nand_1 g05648(n9763, n3986, new_n6025);
nand_1 g05649(n9111, n5860, new_n6026);
not_4  g05650(new_n6026, new_n6027);
xnor_1 g05651(new_n6027, new_n6025, new_n6028);
xnor_1 g05652(new_n6028, new_n6024, new_n6029);
nand_1 g05653(new_n5925, new_n5921, new_n6030);
nand_1 g05654(new_n6030, new_n5923, new_n6031);
xnor_1 g05655(new_n6031, new_n6029, new_n6032);
nand_1 g05656(n7388, n7270, new_n6033);
nand_1 g05657(n11892, n806, new_n6034);
nand_1 g05658(new_n6034, new_n6033, new_n6035);
not_4  g05659(new_n6033, new_n6036);
not_4  g05660(new_n6034, new_n6037);
nand_1 g05661(new_n6037, new_n6036, new_n6038_1);
nand_1 g05662(new_n6038_1, new_n6035, new_n6039);
not_4  g05663(new_n6039, new_n6040);
nand_1 g05664(new_n6040, new_n6032, new_n6041);
not_4  g05665(new_n6031, new_n6042);
xnor_1 g05666(new_n6042, new_n6029, new_n6043);
nand_1 g05667(new_n6039, new_n6043, new_n6044);
nand_1 g05668(new_n6044, new_n6041, new_n6045);
nor_1  g05669(new_n5937, new_n5914, new_n6046);
not_4  g05670(new_n6046, new_n6047);
xnor_1 g05671(new_n6047, new_n6045, new_n6048);
nor_1  g05672(new_n5956, new_n5935, new_n6049);
xnor_1 g05673(new_n6049, new_n6048, new_n6050);
xnor_1 g05674(new_n6050, new_n6023, new_n6051);
xnor_1 g05675(new_n6051, new_n5954, new_n6052);
xnor_1 g05676(new_n6052, new_n6022, new_n6053);
nand_1 g05677(new_n5976, new_n5968, new_n6054);
xnor_1 g05678(new_n6054, new_n6053, new_n6055);
nand_1 g05679(new_n6055, new_n6000, new_n6056);
nand_1 g05680(new_n5998, new_n5993, new_n6057);
nand_1 g05681(new_n5991, new_n5848, new_n6058);
nand_1 g05682(new_n6058, new_n6057, new_n6059);
not_4  g05683(new_n6055, new_n6060);
nand_1 g05684(new_n6060, new_n6059, new_n6061);
nand_1 g05685(new_n6061, new_n6056, new_n6062);
nand_1 g05686(new_n6062, new_n5790, new_n6063);
not_4  g05687(new_n5790, new_n6064);
nor_1  g05688(new_n6060, new_n6059, new_n6065);
nor_1  g05689(new_n6055, new_n6000, new_n6066);
nor_1  g05690(new_n6066, new_n6065, new_n6067);
nor_1  g05691(new_n6067, new_n6064, new_n6068);
nor_1  g05692(new_n6062, new_n5790, new_n6069);
nor_1  g05693(new_n6069, new_n6068, new_n6070);
xnor_1 g05694(new_n5784, new_n5783, new_n6071);
not_4  g05695(new_n6071, new_n6072);
xnor_1 g05696(new_n5996, new_n5982, new_n6073);
nor_1  g05697(new_n6073, new_n6072, new_n6074);
nand_1 g05698(new_n1240, new_n1129, new_n6075);
nor_1  g05699(new_n1324, new_n1241, new_n6076);
not_4  g05700(new_n6076, new_n6077);
nand_1 g05701(new_n6077, new_n6075, new_n6078);
not_4  g05702(new_n6074, new_n6079);
nand_1 g05703(new_n6073, new_n6072, new_n6080);
nand_1 g05704(new_n6080, new_n6079, new_n6081);
nor_1  g05705(new_n6081, new_n6078, new_n6082);
nor_1  g05706(new_n6082, new_n6074, new_n6083);
not_4  g05707(new_n6083, new_n6084);
nand_1 g05708(new_n6084, new_n6070, new_n6085);
nand_1 g05709(new_n6085, new_n6063, new_n6086);
nor_1  g05710(new_n6086, new_n5789, new_n6087);
not_4  g05711(new_n5789, new_n6088);
nand_1 g05712(new_n6067, new_n6064, new_n6089_1);
nand_1 g05713(new_n6089_1, new_n6063, new_n6090);
nor_1  g05714(new_n6083, new_n6090, new_n6091);
nor_1  g05715(new_n6091, new_n6068, new_n6092);
nor_1  g05716(new_n6092, new_n6088, new_n6093);
nor_1  g05717(new_n6093, new_n6087, new_n6094);
not_4  g05718(new_n5813, new_n6095);
nand_1 g05719(new_n5846, new_n6095, new_n6096);
not_4  g05720(new_n5812, new_n6097);
nand_1 g05721(new_n5847, new_n6097, new_n6098);
nand_1 g05722(new_n6098, new_n6096, new_n6099);
not_4  g05723(new_n5841, new_n6100);
nand_1 g05724(new_n5845, new_n6100, new_n6101);
nand_1 g05725(new_n5839, new_n5831, new_n6102);
nand_1 g05726(new_n6102, new_n5829, new_n6103);
nand_1 g05727(n12221, n6776, new_n6104);
nand_1 g05728(n12299, n12145, new_n6105);
nand_1 g05729(n10217, n8759, new_n6106);
not_4  g05730(new_n6106, new_n6107);
xnor_1 g05731(new_n6107, new_n6105, new_n6108);
not_4  g05732(new_n6108, new_n6109);
xnor_1 g05733(new_n6109, new_n6104, new_n6110);
not_4  g05734(new_n6110, new_n6111);
xnor_1 g05735(new_n6111, new_n6103, new_n6112);
not_4  g05736(new_n5837, new_n6113);
nand_1 g05737(n7436, n2522, new_n6114);
not_4  g05738(new_n6114, new_n6115);
nand_1 g05739(new_n6115, new_n6113, new_n6116);
nand_1 g05740(new_n6114, new_n5837, new_n6117);
nand_1 g05741(new_n6117, new_n6116, new_n6118);
not_4  g05742(new_n6118, new_n6119);
nand_1 g05743(n9241, n2024, new_n6120);
not_4  g05744(new_n6120, new_n6121);
nand_1 g05745(n10510, n7946, new_n6122);
nand_1 g05746(n9189, n8276, new_n6123);
nand_1 g05747(new_n6123, new_n6122, new_n6124);
not_4  g05748(new_n6122, new_n6125);
not_4  g05749(new_n6123, new_n6126_1);
nand_1 g05750(new_n6126_1, new_n6125, new_n6127);
nand_1 g05751(new_n6127, new_n6124, new_n6128);
xnor_1 g05752(new_n6128, new_n6121, new_n6129);
not_4  g05753(new_n6129, new_n6130);
xnor_1 g05754(new_n6130, new_n6119, new_n6131);
not_4  g05755(new_n6131, new_n6132);
xnor_1 g05756(new_n6132, new_n6112, new_n6133);
nand_1 g05757(new_n5821, new_n5817, new_n6134);
nor_1  g05758(new_n5819, new_n5818, new_n6135);
nor_1  g05759(new_n5840, new_n5822, new_n6136);
xnor_1 g05760(new_n6136, new_n6135, new_n6137);
nand_1 g05761(new_n6137, new_n6134, new_n6138);
xnor_1 g05762(new_n6138, new_n6133, new_n6139);
xnor_1 g05763(new_n6139, new_n6101, new_n6140);
xnor_1 g05764(new_n6140, new_n6099, new_n6141);
nand_1 g05765(new_n6056, new_n6058, new_n6142);
xnor_1 g05766(new_n6142, new_n6141, new_n6143);
not_4  g05767(new_n6143, new_n6144);
not_4  g05768(new_n6019, new_n6145);
nand_1 g05769(new_n6145, new_n6018, new_n6146);
nand_1 g05770(n8476, n5798, new_n6147);
nand_1 g05771(n6016, n2530, new_n6148);
not_4  g05772(new_n6148, new_n6149);
nand_1 g05773(n5331, n2347, new_n6150);
xnor_1 g05774(new_n6150, new_n6149, new_n6151);
xnor_1 g05775(new_n6151, new_n6147, new_n6152);
nor_1  g05776(new_n6007, new_n6002, new_n6153);
nor_1  g05777(new_n6010, new_n6008, new_n6154);
nor_1  g05778(new_n6154, new_n6153, new_n6155);
xnor_1 g05779(new_n6155, new_n6152, new_n6156);
not_4  g05780(new_n6003, new_n6157);
nand_1 g05781(new_n6005, new_n6157, new_n6158);
nand_1 g05782(n12648, n521, new_n6159);
xnor_1 g05783(new_n6159, new_n6158, new_n6160);
nand_1 g05784(n7690, n2498, new_n6161);
not_4  g05785(new_n6161, new_n6162);
nand_1 g05786(n10545, n5579, new_n6163);
nand_1 g05787(n3616, n2558, new_n6164);
not_4  g05788(new_n6164, new_n6165);
xnor_1 g05789(new_n6165, new_n6163, new_n6166);
xnor_1 g05790(new_n6166, new_n6162, new_n6167);
xnor_1 g05791(new_n6167, new_n6160, new_n6168);
xnor_1 g05792(new_n6168, new_n6156, new_n6169);
not_4  g05793(new_n6169, new_n6170);
not_4  g05794(new_n6011, new_n6171);
nand_1 g05795(new_n6015, new_n6171, new_n6172);
nor_1  g05796(new_n6013, new_n6012, new_n6173);
not_4  g05797(new_n6016_1, new_n6174);
nor_1  g05798(new_n6017, new_n6174, new_n6175);
xnor_1 g05799(new_n6175, new_n6173, new_n6176);
nand_1 g05800(new_n6176, new_n6172, new_n6177);
xnor_1 g05801(new_n6177, new_n6170, new_n6178);
xnor_1 g05802(new_n6178, new_n6146, new_n6179);
not_4  g05803(new_n6001, new_n6180);
nand_1 g05804(new_n6020, new_n6180, new_n6181);
nand_1 g05805(new_n6021, new_n5898, new_n6182);
nand_1 g05806(new_n6182, new_n6181, new_n6183);
xnor_1 g05807(new_n6183, new_n6179, new_n6184);
not_4  g05808(new_n6048, new_n6185);
nor_1  g05809(new_n6049, new_n6185, new_n6186);
not_4  g05810(new_n6024, new_n6187);
nand_1 g05811(new_n6028, new_n6187, new_n6188);
nand_1 g05812(new_n6042, new_n6029, new_n6189);
nand_1 g05813(new_n6189, new_n6188, new_n6190);
nand_1 g05814(n7388, n5153, new_n6191);
not_4  g05815(new_n6191, new_n6192_1);
nand_1 g05816(n11892, n7270, new_n6193);
nand_1 g05817(n7965, n2507, new_n6194);
not_4  g05818(new_n6194, new_n6195);
xnor_1 g05819(new_n6195, new_n6193, new_n6196);
xnor_1 g05820(new_n6196, new_n6192_1, new_n6197);
xnor_1 g05821(new_n6197, new_n6190, new_n6198);
not_4  g05822(new_n6025, new_n6199);
nand_1 g05823(new_n6027, new_n6199, new_n6200);
not_4  g05824(new_n6200, new_n6201);
nand_1 g05825(n2393, n806, new_n6202);
not_4  g05826(new_n6202, new_n6203);
nand_1 g05827(new_n6203, new_n6201, new_n6204);
nand_1 g05828(new_n6202, new_n6200, new_n6205);
nand_1 g05829(new_n6205, new_n6204, new_n6206);
not_4  g05830(new_n6206, new_n6207);
nand_1 g05831(n9111, n3986, new_n6208);
nand_1 g05832(n5860, n3342, new_n6209);
nand_1 g05833(n9763, n5857, new_n6210);
not_4  g05834(new_n6210, new_n6211);
xnor_1 g05835(new_n6211, new_n6209, new_n6212);
xnor_1 g05836(new_n6212, new_n6208, new_n6213);
not_4  g05837(new_n6213, new_n6214);
xnor_1 g05838(new_n6214, new_n6207, new_n6215);
xnor_1 g05839(new_n6215, new_n6198, new_n6216);
not_4  g05840(new_n6216, new_n6217);
not_4  g05841(new_n6041, new_n6218);
nor_1  g05842(new_n6046, new_n6045, new_n6219);
xnor_1 g05843(new_n6219, new_n6038_1, new_n6220);
nor_1  g05844(new_n6220, new_n6218, new_n6221);
xnor_1 g05845(new_n6221, new_n6217, new_n6222);
not_4  g05846(new_n6222, new_n6223);
xnor_1 g05847(new_n6223, new_n6186, new_n6224);
not_4  g05848(new_n6023, new_n6225);
nor_1  g05849(new_n6050, new_n6225, new_n6226);
not_4  g05850(new_n6226, new_n6227);
nand_1 g05851(new_n6051, new_n5965, new_n6228);
nand_1 g05852(new_n6228, new_n6227, new_n6229);
xnor_1 g05853(new_n6229, new_n6224, new_n6230);
xnor_1 g05854(new_n6230, new_n6184, new_n6231);
not_4  g05855(new_n6022, new_n6232);
nand_1 g05856(new_n6052, new_n6232, new_n6233);
nand_1 g05857(new_n6054, new_n6053, new_n6234);
nand_1 g05858(new_n6234, new_n6233, new_n6235);
xnor_1 g05859(new_n6235, new_n6231, new_n6236);
xnor_1 g05860(new_n6236, new_n6144, new_n6237);
not_4  g05861(new_n6237, new_n6238);
nand_1 g05862(new_n6238, new_n6094, new_n6239);
nand_1 g05863(new_n6092, new_n6088, new_n6240);
nand_1 g05864(new_n6086, new_n5789, new_n6241);
nand_1 g05865(new_n6241, new_n6240, new_n6242);
nand_1 g05866(new_n6237, new_n6242, new_n6243);
nand_1 g05867(new_n6243, new_n6239, n1523);
nand_1 g05868(n6687, n4634, new_n6245);
not_4  g05869(new_n4632, new_n6246);
nand_1 g05870(n10223, n4189, new_n6247);
not_4  g05871(new_n6247, new_n6248);
nand_1 g05872(new_n6248, new_n6246, new_n6249);
nand_1 g05873(n10223, n6687, new_n6250);
nand_1 g05874(n7265, n4189, new_n6251);
nand_1 g05875(new_n6251, new_n6250, new_n6252);
nand_1 g05876(n2879, n2564, new_n6253);
not_4  g05877(new_n6253, new_n6254_1);
nand_1 g05878(new_n6254_1, new_n6252, new_n6255);
nand_1 g05879(new_n6255, new_n6249, new_n6256);
xnor_1 g05880(new_n6256, new_n6245, new_n6257);
nand_1 g05881(n4189, n2879, new_n6258);
nand_1 g05882(n10223, n2564, new_n6259);
nand_1 g05883(n7265, n6770, new_n6260);
xnor_1 g05884(new_n6260, new_n6259, new_n6261);
xnor_1 g05885(new_n6261, new_n6258, new_n6262);
xnor_1 g05886(new_n6262, new_n6257, new_n6263);
nand_1 g05887(new_n6252, new_n6249, new_n6264);
not_4  g05888(new_n6264, new_n6265);
nand_1 g05889(n7265, n2564, new_n6266);
not_4  g05890(new_n6266, new_n6267);
nand_1 g05891(n6687, n2879, new_n6268);
not_4  g05892(new_n6268, new_n6269);
nand_1 g05893(new_n6269, new_n6267, new_n6270);
nor_1  g05894(new_n6270, new_n6265, new_n6271);
nand_1 g05895(new_n6271, new_n6263, new_n6272);
nand_1 g05896(n9195, n6687, new_n6273_1);
nand_1 g05897(n4634, n2564, new_n6274);
nand_1 g05898(n6770, n2879, new_n6275);
nand_1 g05899(n9920, n7265, new_n6276);
nand_1 g05900(new_n6276, new_n6247, new_n6277);
not_4  g05901(new_n6276, new_n6278);
nand_1 g05902(new_n6278, new_n6248, new_n6279);
nand_1 g05903(new_n6279, new_n6277, new_n6280);
xnor_1 g05904(new_n6280, new_n6275, new_n6281);
not_4  g05905(new_n6281, new_n6282);
xnor_1 g05906(new_n6282, new_n6274, new_n6283);
nand_1 g05907(new_n6260, new_n6259, new_n6284);
not_4  g05908(new_n6261, new_n6285);
nand_1 g05909(new_n6285, new_n6258, new_n6286);
nand_1 g05910(new_n6286, new_n6284, new_n6287);
xnor_1 g05911(new_n6287, new_n6283, new_n6288);
xnor_1 g05912(new_n6288, new_n6273_1, new_n6289);
not_4  g05913(new_n6245, new_n6290);
nand_1 g05914(new_n6256, new_n6290, new_n6291);
not_4  g05915(new_n6257, new_n6292);
nor_1  g05916(new_n6262, new_n6292, new_n6293);
not_4  g05917(new_n6293, new_n6294_1);
nand_1 g05918(new_n6294_1, new_n6291, new_n6295);
xnor_1 g05919(new_n6295, new_n6289, new_n6296);
not_4  g05920(new_n6296, new_n6297);
xnor_1 g05921(new_n6297, new_n6272, new_n6298);
nand_1 g05922(n8336, n2522, new_n6299);
nand_1 g05923(n9189, n8336, new_n6300);
nand_1 g05924(n7946, n6986, new_n6301);
nand_1 g05925(new_n6301, new_n6300, new_n6302);
not_4  g05926(new_n4633, new_n6303);
nand_1 g05927(n9189, n6986, new_n6304);
not_4  g05928(new_n6304, new_n6305);
nand_1 g05929(new_n6305, new_n6303, new_n6306);
nand_1 g05930(n10928, n2024, new_n6307);
nand_1 g05931(new_n6307, new_n6306, new_n6308);
nand_1 g05932(new_n6308, new_n6302, new_n6309);
not_4  g05933(new_n6309, new_n6310);
xnor_1 g05934(new_n6310, new_n6299, new_n6311);
nand_1 g05935(n6986, n2024, new_n6312);
not_4  g05936(new_n6312, new_n6313);
nand_1 g05937(n10928, n9189, new_n6314);
nand_1 g05938(n7946, n2226, new_n6315);
nand_1 g05939(new_n6315, new_n6314, new_n6316);
not_4  g05940(new_n6314, new_n6317);
not_4  g05941(new_n6315, new_n6318);
nand_1 g05942(new_n6318, new_n6317, new_n6319);
nand_1 g05943(new_n6319, new_n6316, new_n6320);
xnor_1 g05944(new_n6320, new_n6313, new_n6321);
xnor_1 g05945(new_n6321, new_n6311, new_n6322);
not_4  g05946(new_n6322, new_n6323);
not_4  g05947(new_n6307, new_n6324);
nand_1 g05948(new_n6324, new_n4633, new_n6325);
nand_1 g05949(new_n6306, new_n6302, new_n6326);
nand_1 g05950(new_n6326, new_n6325, new_n6327);
not_4  g05951(new_n6327, new_n6328);
nand_1 g05952(new_n6328, new_n6324, new_n6329);
not_4  g05953(new_n6329, new_n6330);
nand_1 g05954(new_n6330, new_n6323, new_n6331);
nand_1 g05955(n12145, n8336, new_n6332);
nand_1 g05956(n10928, n2522, new_n6333);
nand_1 g05957(new_n6319, new_n6312, new_n6334);
nand_1 g05958(new_n6334, new_n6316, new_n6335);
not_4  g05959(new_n6335, new_n6336);
xnor_1 g05960(new_n6336, new_n6333, new_n6337);
nand_1 g05961(n2226, n2024, new_n6338);
nand_1 g05962(n7946, n1094, new_n6339);
nand_1 g05963(new_n6339, new_n6304, new_n6340);
not_4  g05964(new_n6339, new_n6341);
nand_1 g05965(new_n6341, new_n6305, new_n6342);
nand_1 g05966(new_n6342, new_n6340, new_n6343);
xnor_1 g05967(new_n6343, new_n6338, new_n6344);
xnor_1 g05968(new_n6344, new_n6337, new_n6345);
xnor_1 g05969(new_n6345, new_n6332, new_n6346);
nor_1  g05970(new_n6309, new_n6299, new_n6347);
not_4  g05971(new_n6347, new_n6348);
nand_1 g05972(new_n6321, new_n6311, new_n6349);
nand_1 g05973(new_n6349, new_n6348, new_n6350);
xnor_1 g05974(new_n6350, new_n6346, new_n6351);
not_4  g05975(new_n6351, new_n6352);
xnor_1 g05976(new_n6352, new_n6331, new_n6353);
xnor_1 g05977(new_n6329, new_n6323, new_n6354);
not_4  g05978(new_n6354, new_n6355);
nand_1 g05979(n12069, n521, new_n6356);
nand_1 g05980(n7891, n5579, new_n6357);
not_4  g05981(new_n6357, new_n6358_1);
nand_1 g05982(new_n6358_1, new_n4637, new_n6359_1);
nand_1 g05983(n12069, n5579, new_n6360);
nand_1 g05984(n7891, n2558, new_n6361);
nand_1 g05985(new_n6361, new_n6360, new_n6362);
nand_1 g05986(n12391, n2498, new_n6363);
not_4  g05987(new_n6363, new_n6364);
nand_1 g05988(new_n6364, new_n6362, new_n6365);
nand_1 g05989(new_n6365, new_n6359_1, new_n6366);
xnor_1 g05990(new_n6366, new_n6356, new_n6367);
nand_1 g05991(n7891, n2498, new_n6368);
not_4  g05992(new_n6368, new_n6369);
nand_1 g05993(n12391, n5579, new_n6370);
nand_1 g05994(n7160, n2558, new_n6371);
nand_1 g05995(new_n6371, new_n6370, new_n6372);
not_4  g05996(new_n6370, new_n6373);
not_4  g05997(new_n6371, new_n6374);
nand_1 g05998(new_n6374, new_n6373, new_n6375);
nand_1 g05999(new_n6375, new_n6372, new_n6376);
xnor_1 g06000(new_n6376, new_n6369, new_n6377);
not_4  g06001(new_n6377, new_n6378);
xnor_1 g06002(new_n6378, new_n6367, new_n6379);
nand_1 g06003(new_n6362, new_n6359_1, new_n6380);
not_4  g06004(new_n6380, new_n6381);
nand_1 g06005(n12391, n2558, new_n6382);
not_4  g06006(new_n6382, new_n6383);
nand_1 g06007(n12069, n2498, new_n6384);
not_4  g06008(new_n6384, new_n6385);
nand_1 g06009(new_n6385, new_n6383, new_n6386);
nor_1  g06010(new_n6386, new_n6381, new_n6387);
nor_1  g06011(new_n6387, new_n6379, new_n6388);
nand_1 g06012(new_n6387, new_n6379, new_n6389);
not_4  g06013(new_n6389, new_n6390);
nor_1  g06014(new_n6390, new_n6388, new_n6391);
nand_1 g06015(n11222, n806, new_n6392);
nand_1 g06016(n11222, n3342, new_n6393);
nand_1 g06017(n9763, n5314, new_n6394);
nand_1 g06018(new_n6394, new_n6393, new_n6395);
nand_1 g06019(n5314, n3342, new_n6396);
not_4  g06020(new_n6396, new_n6397);
nand_1 g06021(new_n6397, new_n4635, new_n6398);
nand_1 g06022(n11153, n9111, new_n6399);
nand_1 g06023(new_n6399, new_n6398, new_n6400);
nand_1 g06024(new_n6400, new_n6395, new_n6401);
nor_1  g06025(new_n6401, new_n6392, new_n6402);
not_4  g06026(new_n6402, new_n6403);
nand_1 g06027(new_n6401, new_n6392, new_n6404);
nand_1 g06028(new_n6404, new_n6403, new_n6405);
nand_1 g06029(n9111, n5314, new_n6406);
not_4  g06030(new_n6406, new_n6407);
nand_1 g06031(n11153, n3342, new_n6408);
nand_1 g06032(n9763, n996, new_n6409);
nand_1 g06033(new_n6409, new_n6408, new_n6410);
not_4  g06034(new_n6408, new_n6411);
not_4  g06035(new_n6409, new_n6412);
nand_1 g06036(new_n6412, new_n6411, new_n6413);
nand_1 g06037(new_n6413, new_n6410, new_n6414);
xnor_1 g06038(new_n6414, new_n6407, new_n6415);
xnor_1 g06039(new_n6415, new_n6405, new_n6416);
not_4  g06040(new_n6399, new_n6417);
not_4  g06041(new_n6395, new_n6418);
nand_1 g06042(new_n6417, new_n4634_1, new_n6419);
nand_1 g06043(new_n6419, new_n6418, new_n6420);
nand_1 g06044(new_n6420, new_n6398, new_n6421);
nand_1 g06045(new_n6421, new_n6417, new_n6422);
xnor_1 g06046(new_n6422, new_n6416, new_n6423);
not_4  g06047(new_n6423, new_n6424);
xnor_1 g06048(new_n6424, new_n6391, new_n6425);
nor_1  g06049(new_n6419, new_n6418, new_n6426);
nor_1  g06050(new_n6426, new_n6421, new_n6427);
not_4  g06051(new_n6427, new_n6428);
not_4  g06052(new_n4638, new_n6429_1);
xnor_1 g06053(new_n6385, new_n6382, new_n6430);
nor_1  g06054(new_n6430, new_n6429_1, new_n6431_1);
not_4  g06055(new_n6431_1, new_n6432);
xnor_1 g06056(new_n6430, new_n4638, new_n6433);
nand_1 g06057(n11153, n9763, new_n6434);
nand_1 g06058(n11222, n9111, new_n6435);
xnor_1 g06059(new_n6435, new_n6434, new_n6436);
nand_1 g06060(new_n6436, new_n6433, new_n6437);
nand_1 g06061(new_n6437, new_n6432, new_n6438);
nand_1 g06062(new_n6438, new_n6428, new_n6439);
xnor_1 g06063(new_n6438, new_n6427, new_n6440);
nand_1 g06064(new_n6364, new_n4636, new_n6441_1);
nand_1 g06065(new_n6441_1, new_n6380, new_n6442);
not_4  g06066(new_n6441_1, new_n6443);
nand_1 g06067(new_n6443, new_n6362, new_n6444);
nand_1 g06068(new_n6444, new_n6442, new_n6445_1);
nand_1 g06069(new_n6445_1, new_n6440, new_n6446);
nand_1 g06070(new_n6446, new_n6439, new_n6447);
nor_1  g06071(new_n6447, new_n6425, new_n6448);
nand_1 g06072(new_n6447, new_n6425, new_n6449);
not_4  g06073(new_n6449, new_n6450);
nor_1  g06074(new_n6450, new_n6448, new_n6451);
nor_1  g06075(new_n6451, new_n6355, new_n6452);
not_4  g06076(new_n6452, new_n6453);
xnor_1 g06077(new_n6451, new_n6354, new_n6454);
not_4  g06078(new_n6325, new_n6455);
nand_1 g06079(new_n6455, new_n6302, new_n6456);
nand_1 g06080(new_n6456, new_n6327, new_n6457);
xnor_1 g06081(new_n6445_1, new_n6440, new_n6458);
not_4  g06082(new_n6458, new_n6459);
nor_1  g06083(new_n6459, new_n6457, new_n6460);
not_4  g06084(new_n6460, new_n6461);
xnor_1 g06085(new_n6458, new_n6457, new_n6462);
xnor_1 g06086(new_n6436, new_n6433, new_n6463);
nand_1 g06087(n10928, n7946, new_n6464);
nand_1 g06088(n8336, n2024, new_n6465);
xnor_1 g06089(new_n6465, new_n6464, new_n6466);
not_4  g06090(new_n6466, new_n6467);
nand_1 g06091(new_n6467, new_n6463, new_n6468);
nand_1 g06092(new_n4641, new_n6303, new_n6469);
not_4  g06093(new_n6469, new_n6470);
xnor_1 g06094(new_n6466, new_n6463, new_n6471);
nand_1 g06095(new_n6471, new_n6470, new_n6472);
nand_1 g06096(new_n6472, new_n6468, new_n6473);
nand_1 g06097(new_n6473, new_n6462, new_n6474);
nand_1 g06098(new_n6474, new_n6461, new_n6475);
nand_1 g06099(new_n6475, new_n6454, new_n6476);
nand_1 g06100(new_n6476, new_n6453, new_n6477);
not_4  g06101(new_n6477, new_n6478);
xnor_1 g06102(new_n6478, new_n6353, new_n6479);
nand_1 g06103(n12069, n6016, new_n6480);
nand_1 g06104(n12391, n521, new_n6481);
nand_1 g06105(new_n6375, new_n6368, new_n6482);
nand_1 g06106(new_n6482, new_n6372, new_n6483);
not_4  g06107(new_n6483, new_n6484);
xnor_1 g06108(new_n6484, new_n6481, new_n6485);
nand_1 g06109(n7160, n2498, new_n6486);
not_4  g06110(new_n6486, new_n6487);
nand_1 g06111(n4828, n2558, new_n6488);
not_4  g06112(new_n6488, new_n6489);
xnor_1 g06113(new_n6489, new_n6357, new_n6490);
xnor_1 g06114(new_n6490, new_n6487, new_n6491);
xnor_1 g06115(new_n6491, new_n6485, new_n6492);
xnor_1 g06116(new_n6492, new_n6480, new_n6493);
not_4  g06117(new_n6356, new_n6494);
nand_1 g06118(new_n6366, new_n6494, new_n6495);
nand_1 g06119(new_n6377, new_n6367, new_n6496);
nand_1 g06120(new_n6496, new_n6495, new_n6497);
nor_1  g06121(new_n6497, new_n6493, new_n6498);
nand_1 g06122(new_n6497, new_n6493, new_n6499);
not_4  g06123(new_n6499, new_n6500);
nor_1  g06124(new_n6500, new_n6498, new_n6501);
xnor_1 g06125(new_n6501, new_n6389, new_n6502);
not_4  g06126(new_n6416, new_n6503);
nor_1  g06127(new_n6422, new_n6503, new_n6504);
nand_1 g06128(n11222, n7270, new_n6505);
nand_1 g06129(n11153, n806, new_n6506);
nand_1 g06130(new_n6413, new_n6406, new_n6507);
nand_1 g06131(new_n6507, new_n6410, new_n6508);
nor_1  g06132(new_n6508, new_n6506, new_n6509);
not_4  g06133(new_n6509, new_n6510);
nand_1 g06134(new_n6508, new_n6506, new_n6511);
nand_1 g06135(new_n6511, new_n6510, new_n6512);
nand_1 g06136(n9111, n996, new_n6513);
not_4  g06137(new_n6513, new_n6514);
nand_1 g06138(n9763, n5767, new_n6515);
nand_1 g06139(new_n6515, new_n6396, new_n6516);
nor_1  g06140(new_n6515, new_n6396, new_n6517);
not_4  g06141(new_n6517, new_n6518);
nand_1 g06142(new_n6518, new_n6516, new_n6519);
xnor_1 g06143(new_n6519, new_n6514, new_n6520);
xnor_1 g06144(new_n6520, new_n6512, new_n6521);
xnor_1 g06145(new_n6521, new_n6505, new_n6522);
not_4  g06146(new_n6522, new_n6523);
not_4  g06147(new_n6405, new_n6524);
nand_1 g06148(new_n6415, new_n6524, new_n6525);
nand_1 g06149(new_n6525, new_n6403, new_n6526);
xnor_1 g06150(new_n6526, new_n6523, new_n6527);
nand_1 g06151(new_n6527, new_n6504, new_n6528);
not_4  g06152(new_n6528, new_n6529);
nor_1  g06153(new_n6527, new_n6504, new_n6530);
nor_1  g06154(new_n6530, new_n6529, new_n6531);
nand_1 g06155(new_n6531, new_n6502, new_n6532);
nor_1  g06156(new_n6531, new_n6502, new_n6533);
not_4  g06157(new_n6533, new_n6534);
nand_1 g06158(new_n6534, new_n6532, new_n6535);
not_4  g06159(new_n6535, new_n6536);
nor_1  g06160(new_n6423, new_n6391, new_n6537);
nor_1  g06161(new_n6450, new_n6537, new_n6538);
not_4  g06162(new_n6538, new_n6539);
nand_1 g06163(new_n6539, new_n6536, new_n6540);
nand_1 g06164(new_n6538, new_n6535, new_n6541);
nand_1 g06165(new_n6541, new_n6540, new_n6542);
not_4  g06166(new_n6542, new_n6543);
xnor_1 g06167(new_n6543, new_n6479, new_n6544);
nor_1  g06168(new_n6544, new_n6298, new_n6545);
not_4  g06169(new_n6545, new_n6546);
nand_1 g06170(new_n6544, new_n6298, new_n6547);
nand_1 g06171(new_n6547, new_n6546, new_n6548);
xnor_1 g06172(new_n6271, new_n6263, new_n6549);
xnor_1 g06173(new_n6475, new_n6454, new_n6550);
nand_1 g06174(new_n6550, new_n6549, new_n6551);
xnor_1 g06175(new_n6473, new_n6462, new_n6552);
nand_1 g06176(new_n6254_1, new_n4632, new_n6553);
nand_1 g06177(new_n6553, new_n6264, new_n6554);
not_4  g06178(new_n6553, new_n6555);
nand_1 g06179(new_n6555, new_n6252, new_n6556);
nand_1 g06180(new_n6556, new_n6554, new_n6557);
nand_1 g06181(new_n6557, new_n6552, new_n6558);
xnor_1 g06182(new_n6557, new_n6552, new_n6559);
nand_1 g06183(new_n4642, new_n6246, new_n6560);
nand_1 g06184(new_n6268, new_n6266, new_n6561);
nand_1 g06185(new_n6561, new_n6270, new_n6562);
nand_1 g06186(new_n6562, new_n6560, new_n6563);
xnor_1 g06187(new_n6471, new_n6469, new_n6564);
xnor_1 g06188(new_n6562, new_n6560, new_n6565);
nor_1  g06189(new_n6565, new_n6564, new_n6566);
not_4  g06190(new_n6566, new_n6567);
nand_1 g06191(new_n6567, new_n6563, new_n6568);
not_4  g06192(new_n6568, new_n6569);
nor_1  g06193(new_n6569, new_n6559, new_n6570);
not_4  g06194(new_n6570, new_n6571);
nand_1 g06195(new_n6571, new_n6558, new_n6572);
not_4  g06196(new_n6572, new_n6573);
xnor_1 g06197(new_n6550, new_n6549, new_n6574);
nor_1  g06198(new_n6574, new_n6573, new_n6575);
not_4  g06199(new_n6575, new_n6576);
nand_1 g06200(new_n6576, new_n6551, new_n6577);
not_4  g06201(new_n6577, new_n6578_1);
nand_1 g06202(new_n6578_1, new_n6548, new_n6579);
nor_1  g06203(new_n6578_1, new_n6548, new_n6580);
not_4  g06204(new_n6580, new_n6581);
nand_1 g06205(new_n6581, new_n6579, n1658);
nand_1 g06206(n7862, n4634, new_n6583);
nand_1 g06207(n10223, n7862, new_n6584);
nand_1 g06208(n7265, n3172, new_n6585);
nand_1 g06209(new_n6585, new_n6584, new_n6586);
nand_1 g06210(n7862, n7265, new_n6587);
not_4  g06211(new_n6587, new_n6588);
nand_1 g06212(n10223, n3172, new_n6589);
not_4  g06213(new_n6589, new_n6590);
nand_1 g06214(new_n6590, new_n6588, new_n6591);
nand_1 g06215(n2879, n1333, new_n6592);
nand_1 g06216(new_n6592, new_n6591, new_n6593);
nand_1 g06217(new_n6593, new_n6586, new_n6594);
nor_1  g06218(new_n6594, new_n6583, new_n6595);
not_4  g06219(new_n6595, new_n6596);
nand_1 g06220(new_n6594, new_n6583, new_n6597);
nand_1 g06221(new_n6597, new_n6596, new_n6598);
nand_1 g06222(n3172, n2879, new_n6599);
not_4  g06223(new_n6599, new_n6600);
nand_1 g06224(n10223, n1333, new_n6601);
nand_1 g06225(n11757, n7265, new_n6602);
nand_1 g06226(new_n6602, new_n6601, new_n6603);
nor_1  g06227(new_n6602, new_n6601, new_n6604_1);
not_4  g06228(new_n6604_1, new_n6605);
nand_1 g06229(new_n6605, new_n6603, new_n6606);
xnor_1 g06230(new_n6606, new_n6600, new_n6607);
xnor_1 g06231(new_n6607, new_n6598, new_n6608);
not_4  g06232(new_n6592, new_n6609);
not_4  g06233(new_n6586, new_n6610);
nand_1 g06234(new_n6609, new_n6587, new_n6611_1);
nand_1 g06235(new_n6611_1, new_n6610, new_n6612);
nand_1 g06236(new_n6612, new_n6591, new_n6613);
nand_1 g06237(new_n6613, new_n6609, new_n6614);
xnor_1 g06238(new_n6614, new_n6608, new_n6615);
nand_1 g06239(n6877, n2522, new_n6616);
nand_1 g06240(n2464, n2024, new_n6617);
not_4  g06241(new_n6617, new_n6618);
nand_1 g06242(n9400, n9189, new_n6619);
nand_1 g06243(n11311, n7946, new_n6620);
not_4  g06244(new_n6620, new_n6621);
xnor_1 g06245(new_n6621, new_n6619, new_n6622);
xnor_1 g06246(new_n6622, new_n6618, new_n6623);
nor_1  g06247(new_n6623, new_n6616, new_n6624);
not_4  g06248(new_n6624, new_n6625);
nand_1 g06249(new_n6623, new_n6616, new_n6626);
nand_1 g06250(new_n6626, new_n6625, new_n6627);
nand_1 g06251(n9189, n6877, new_n6628);
nand_1 g06252(n7946, n2464, new_n6629);
nand_1 g06253(new_n6629, new_n6628, new_n6630);
nand_1 g06254(n7946, n6877, new_n6631);
not_4  g06255(new_n6631, new_n6632);
nand_1 g06256(n9189, n2464, new_n6633);
not_4  g06257(new_n6633, new_n6634);
nand_1 g06258(new_n6634, new_n6632, new_n6635);
nand_1 g06259(n9400, n2024, new_n6636);
nand_1 g06260(new_n6636, new_n6635, new_n6637);
nand_1 g06261(new_n6637, new_n6630, new_n6638);
nor_1  g06262(new_n6638, new_n6627, new_n6639);
not_4  g06263(new_n6639, new_n6640);
nand_1 g06264(new_n6638, new_n6627, new_n6641);
nand_1 g06265(new_n6641, new_n6640, new_n6642);
not_4  g06266(new_n6636, new_n6643);
nand_1 g06267(new_n6643, new_n6631, new_n6644);
nand_1 g06268(new_n6635, new_n6630, new_n6645_1);
nand_1 g06269(new_n6645_1, new_n6644, new_n6646);
not_4  g06270(new_n6646, new_n6647);
nand_1 g06271(new_n6647, new_n6643, new_n6648);
nand_1 g06272(new_n6648, new_n6642, new_n6649);
not_4  g06273(new_n6642, new_n6650);
not_4  g06274(new_n6648, new_n6651);
nand_1 g06275(new_n6651, new_n6650, new_n6652);
nand_1 g06276(new_n6652, new_n6649, new_n6653);
not_4  g06277(new_n6653, new_n6654);
not_4  g06278(new_n6644, new_n6655);
nand_1 g06279(new_n6655, new_n6630, new_n6656);
nand_1 g06280(new_n6656, new_n6646, new_n6657);
nand_1 g06281(n4805, n2558, new_n6658);
nand_1 g06282(n9763, n7236, new_n6659);
not_4  g06283(new_n6659, new_n6660);
xnor_1 g06284(new_n6660, new_n6658, new_n6661);
nand_1 g06285(new_n6661, new_n6632, new_n6662);
not_4  g06286(new_n6662, new_n6663);
nand_1 g06287(n9400, n7946, new_n6664);
nand_1 g06288(n6877, n2024, new_n6665);
not_4  g06289(new_n6665, new_n6666);
xnor_1 g06290(new_n6666, new_n6664, new_n6667);
nand_1 g06291(new_n6667, new_n6663, new_n6668);
not_4  g06292(new_n6668, new_n6669);
nor_1  g06293(new_n6659, new_n6658, new_n6670);
nand_1 g06294(n9111, n7236, new_n6671);
nand_1 g06295(n9763, n3992, new_n6672);
nand_1 g06296(new_n6672, new_n6671, new_n6673);
not_4  g06297(new_n6671, new_n6674);
not_4  g06298(new_n6672, new_n6675);
nand_1 g06299(new_n6675, new_n6674, new_n6676);
nand_1 g06300(new_n6676, new_n6673, new_n6677);
xnor_1 g06301(new_n6677, new_n6670, new_n6678);
not_4  g06302(new_n6678, new_n6679);
nand_1 g06303(n4805, n2498, new_n6680);
nand_1 g06304(n11478, n2558, new_n6681);
xnor_1 g06305(new_n6681, new_n6680, new_n6682);
xnor_1 g06306(new_n6682, new_n6679, new_n6683);
xnor_1 g06307(new_n6667, new_n6662, new_n6684);
not_4  g06308(new_n6684, new_n6685);
nor_1  g06309(new_n6685, new_n6683, new_n6686);
nor_1  g06310(new_n6686, new_n6669, new_n6687_1);
nand_1 g06311(new_n6687_1, new_n6657, new_n6688);
not_4  g06312(new_n6670, new_n6689_1);
nand_1 g06313(new_n6677, new_n6689_1, new_n6690);
nand_1 g06314(new_n6682, new_n6678, new_n6691);
nand_1 g06315(new_n6691, new_n6690, new_n6692);
nand_1 g06316(n11478, n2498, new_n6693);
not_4  g06317(new_n6693, new_n6694);
nand_1 g06318(new_n6694, new_n6658, new_n6695);
nand_1 g06319(n5283, n2558, new_n6696);
nand_1 g06320(n5579, n4805, new_n6697);
nand_1 g06321(new_n6697, new_n6696, new_n6698);
not_4  g06322(new_n6696, new_n6699);
not_4  g06323(new_n6697, new_n6700);
nand_1 g06324(new_n6700, new_n6699, new_n6701);
nand_1 g06325(new_n6701, new_n6698, new_n6702);
nand_1 g06326(new_n6702, new_n6695, new_n6703_1);
not_4  g06327(new_n6698, new_n6704);
nor_1  g06328(new_n6704, new_n6695, new_n6705);
not_4  g06329(new_n6705, new_n6706);
nand_1 g06330(new_n6706, new_n6703_1, new_n6707);
xnor_1 g06331(new_n6707, new_n6692, new_n6708);
not_4  g06332(new_n6708, new_n6709);
nand_1 g06333(n9111, n3992, new_n6710);
not_4  g06334(new_n6710, new_n6711);
nand_1 g06335(new_n6711, new_n6659, new_n6712);
not_4  g06336(new_n6712, new_n6713);
nand_1 g06337(n9763, n8384, new_n6714);
nand_1 g06338(n7236, n3342, new_n6715);
nand_1 g06339(new_n6715, new_n6714, new_n6716);
not_4  g06340(new_n6716, new_n6717);
nand_1 g06341(new_n6717, new_n6713, new_n6718);
not_4  g06342(new_n6714, new_n6719);
not_4  g06343(new_n6715, new_n6720);
nand_1 g06344(new_n6720, new_n6719, new_n6721);
nand_1 g06345(new_n6721, new_n6716, new_n6722);
not_4  g06346(new_n6722, new_n6723);
nand_1 g06347(new_n6723, new_n6712, new_n6724);
nand_1 g06348(new_n6724, new_n6718, new_n6725);
xnor_1 g06349(new_n6725, new_n6709, new_n6726);
not_4  g06350(new_n6726, new_n6727);
xnor_1 g06351(new_n6687_1, new_n6657, new_n6728);
nor_1  g06352(new_n6728, new_n6727, new_n6729);
not_4  g06353(new_n6729, new_n6730);
nand_1 g06354(new_n6730, new_n6688, new_n6731);
xnor_1 g06355(new_n6731, new_n6654, new_n6732);
not_4  g06356(new_n6732, new_n6733);
nand_1 g06357(n4805, n521, new_n6734);
nand_1 g06358(new_n6701, new_n6693, new_n6735);
nand_1 g06359(new_n6735, new_n6698, new_n6736);
xnor_1 g06360(new_n6736, new_n6734, new_n6737);
nand_1 g06361(n5283, n2498, new_n6738);
nand_1 g06362(n2558, n137, new_n6739);
nand_1 g06363(n11478, n5579, new_n6740);
nand_1 g06364(new_n6740, new_n6739, new_n6741);
not_4  g06365(new_n6739, new_n6742_1);
not_4  g06366(new_n6740, new_n6743);
nand_1 g06367(new_n6743, new_n6742_1, new_n6744);
nand_1 g06368(new_n6744, new_n6741, new_n6745);
xnor_1 g06369(new_n6745, new_n6738, new_n6746);
not_4  g06370(new_n6746, new_n6747);
xnor_1 g06371(new_n6747, new_n6737, new_n6748);
nor_1  g06372(new_n6703_1, new_n6693, new_n6749);
xnor_1 g06373(new_n6749, new_n6748, new_n6750);
nand_1 g06374(n7236, n806, new_n6751);
nand_1 g06375(new_n6716, new_n6711, new_n6752);
nand_1 g06376(new_n6752, new_n6721, new_n6753);
xnor_1 g06377(new_n6753, new_n6751, new_n6754);
nand_1 g06378(n9111, n8384, new_n6755);
not_4  g06379(new_n6755, new_n6756);
nand_1 g06380(n9763, n6358, new_n6757);
nand_1 g06381(n3992, n3342, new_n6758);
nand_1 g06382(new_n6758, new_n6757, new_n6759);
not_4  g06383(new_n6757, new_n6760);
not_4  g06384(new_n6758, new_n6761);
nand_1 g06385(new_n6761, new_n6760, new_n6762);
nand_1 g06386(new_n6762, new_n6759, new_n6763);
xnor_1 g06387(new_n6763, new_n6756, new_n6764);
xnor_1 g06388(new_n6764, new_n6754, new_n6765);
nor_1  g06389(new_n6723, new_n6676, new_n6766);
xnor_1 g06390(new_n6766, new_n6765, new_n6767);
xnor_1 g06391(new_n6767, new_n6750, new_n6768);
nand_1 g06392(new_n6707, new_n6692, new_n6769);
not_4  g06393(new_n6725, new_n6770_1);
nand_1 g06394(new_n6770_1, new_n6709, new_n6771);
nand_1 g06395(new_n6771, new_n6769, new_n6772);
xnor_1 g06396(new_n6772, new_n6768, new_n6773);
xnor_1 g06397(new_n6773, new_n6733, new_n6774);
nand_1 g06398(new_n6774, new_n6615, new_n6775);
nor_1  g06399(new_n6774, new_n6615, new_n6776_1);
not_4  g06400(new_n6776_1, new_n6777);
nand_1 g06401(new_n6777, new_n6775, new_n6778);
nor_1  g06402(new_n6611_1, new_n6610, new_n6779);
nor_1  g06403(new_n6779, new_n6613, new_n6780);
nand_1 g06404(new_n6728, new_n6727, new_n6781);
nand_1 g06405(new_n6781, new_n6730, new_n6782);
nand_1 g06406(new_n6782, new_n6780, new_n6783);
xnor_1 g06407(new_n6661, new_n6631, new_n6784);
nand_1 g06408(new_n6784, new_n6588, new_n6785);
nand_1 g06409(n7265, n1333, new_n6786);
nand_1 g06410(n7862, n2879, new_n6787);
xnor_1 g06411(new_n6787, new_n6786, new_n6788);
nand_1 g06412(new_n6788, new_n6785, new_n6789);
xnor_1 g06413(new_n6684, new_n6683, new_n6790);
xnor_1 g06414(new_n6788, new_n6785, new_n6791);
nor_1  g06415(new_n6791, new_n6790, new_n6792);
not_4  g06416(new_n6792, new_n6793);
nand_1 g06417(new_n6793, new_n6789, new_n6794);
xnor_1 g06418(new_n6782, new_n6780, new_n6795);
nor_1  g06419(new_n6795, new_n6794, new_n6796);
not_4  g06420(new_n6796, new_n6797_1);
nand_1 g06421(new_n6797_1, new_n6783, new_n6798);
xnor_1 g06422(new_n6798, new_n6778, n1847);
nand_1 g06423(n5305, n1798, new_n6800);
not_4  g06424(new_n6800, new_n6801);
nand_1 g06425(n8759, n6703, new_n6802);
nand_1 g06426(n5645, n5331, new_n6803);
not_4  g06427(new_n6803, new_n6804);
nand_1 g06428(n11876, n7965, new_n6805);
not_4  g06429(new_n6805, new_n6806_1);
nand_1 g06430(new_n6806_1, new_n6804, new_n6807);
nand_1 g06431(new_n6805, new_n6803, new_n6808);
nand_1 g06432(new_n6808, new_n6807, new_n6809_1);
not_4  g06433(new_n6809_1, new_n6810);
xnor_1 g06434(new_n6810, new_n6802, new_n6811);
nand_1 g06435(new_n6811, new_n6801, new_n6812);
not_4  g06436(new_n6812, new_n6813);
nand_1 g06437(n5305, n3932, new_n6814);
nand_1 g06438(n5964, n1798, new_n6815);
nand_1 g06439(new_n6815, new_n6814, new_n6816);
not_4  g06440(new_n6814, new_n6817);
not_4  g06441(new_n6815, new_n6818);
nand_1 g06442(new_n6818, new_n6817, new_n6819);
nand_1 g06443(new_n6819, new_n6816, new_n6820);
xnor_1 g06444(new_n6820, new_n6813, new_n6821);
not_4  g06445(new_n6802, new_n6822_1);
nand_1 g06446(new_n6810, new_n6822_1, new_n6823);
nand_1 g06447(n9640, n8759, new_n6824);
nand_1 g06448(n6776, n6703, new_n6825);
xnor_1 g06449(new_n6825, new_n6824, new_n6826_1);
not_4  g06450(new_n6826_1, new_n6827);
xnor_1 g06451(new_n6827, new_n6823, new_n6828);
nand_1 g06452(n10898, n7965, new_n6829);
nand_1 g06453(n11876, n7388, new_n6830);
xnor_1 g06454(new_n6830, new_n6829, new_n6831);
not_4  g06455(new_n6831, new_n6832);
xnor_1 g06456(new_n6832, new_n6807, new_n6833);
not_4  g06457(new_n6833, new_n6834);
nand_1 g06458(n5331, n1067, new_n6835);
nand_1 g06459(n8476, n5645, new_n6836);
nand_1 g06460(new_n6836, new_n6835, new_n6837);
not_4  g06461(new_n6835, new_n6838);
not_4  g06462(new_n6836, new_n6839);
nand_1 g06463(new_n6839, new_n6838, new_n6840);
nand_1 g06464(new_n6840, new_n6837, new_n6841);
nand_1 g06465(new_n6841, new_n6834, new_n6842);
not_4  g06466(new_n6841, new_n6843);
nand_1 g06467(new_n6843, new_n6833, new_n6844);
nand_1 g06468(new_n6844, new_n6842, new_n6845);
xnor_1 g06469(new_n6845, new_n6828, new_n6846);
not_4  g06470(new_n6846, new_n6847);
xnor_1 g06471(new_n6847, new_n6821, n2096);
not_4  g06472(new_n3923, new_n6849);
xnor_1 g06473(new_n3926, new_n6849, n2131);
nand_1 g06474(n7456, n2564, new_n6851);
not_4  g06475(new_n6851, new_n6852);
nand_1 g06476(new_n4100, new_n4095, new_n6853);
nand_1 g06477(new_n6853, new_n4098, new_n6854);
not_4  g06478(new_n6854, new_n6855);
nand_1 g06479(new_n6855, new_n6852, new_n6856);
xnor_1 g06480(new_n6854, new_n6852, new_n6857);
nand_1 g06481(n6770, n3932, new_n6858);
nand_1 g06482(n9920, n1798, new_n6859);
nand_1 g06483(new_n6859, new_n4088_1, new_n6860_1);
not_4  g06484(new_n6860_1, new_n6861);
nor_1  g06485(new_n6859, new_n4088_1, new_n6862);
nor_1  g06486(new_n6862, new_n6861, new_n6863);
xnor_1 g06487(new_n6863, new_n6858, new_n6864);
nand_1 g06488(new_n6864, new_n6857, new_n6865);
nand_1 g06489(new_n6865, new_n6856, new_n6866);
nand_1 g06490(n11662, n2564, new_n6867);
nand_1 g06491(n7456, n4189, new_n6868);
not_4  g06492(new_n6868, new_n6869);
xnor_1 g06493(new_n6869, new_n6867, new_n6870);
xnor_1 g06494(new_n6870, new_n6866, new_n6871);
not_4  g06495(new_n6871, new_n6872);
nand_1 g06496(n12591, n6770, new_n6873);
nand_1 g06497(n3627, n1798, new_n6874);
nand_1 g06498(n9920, n3932, new_n6875);
not_4  g06499(new_n6875, new_n6876);
xnor_1 g06500(new_n6876, new_n6874, new_n6877_1);
xnor_1 g06501(new_n6877_1, new_n6873, new_n6878);
not_4  g06502(new_n6878, new_n6879);
not_4  g06503(new_n6858, new_n6880);
nor_1  g06504(new_n6862, new_n6880, new_n6881);
nor_1  g06505(new_n6881, new_n6861, new_n6882);
not_4  g06506(new_n6882, new_n6883);
xnor_1 g06507(new_n6883, new_n6879, new_n6884);
xnor_1 g06508(new_n6884, new_n6872, new_n6885);
nand_1 g06509(n11662, n6687, new_n6886);
nor_1  g06510(new_n4093, new_n4082, new_n6887);
nor_1  g06511(new_n4103, new_n6887, new_n6888);
nand_1 g06512(new_n6888, new_n6886, new_n6889);
xnor_1 g06513(new_n6864, new_n6857, new_n6890);
not_4  g06514(new_n6888, new_n6891);
xnor_1 g06515(new_n6891, new_n6886, new_n6892);
nand_1 g06516(new_n6892, new_n6890, new_n6893);
nand_1 g06517(new_n6893, new_n6889, new_n6894);
not_4  g06518(new_n6894, new_n6895);
nand_1 g06519(new_n6895, new_n6885, new_n6896);
not_4  g06520(new_n6873, new_n6897);
nand_1 g06521(new_n6877_1, new_n6897, new_n6898);
nand_1 g06522(new_n6882, new_n6878, new_n6899);
nand_1 g06523(new_n6899, new_n6898, new_n6900);
nand_1 g06524(n10327, n2564, new_n6901);
nand_1 g06525(n11662, n4189, new_n6902);
nand_1 g06526(n9583, n6687, new_n6903);
not_4  g06527(new_n6903, new_n6904);
xnor_1 g06528(new_n6904, new_n6902, new_n6905);
xnor_1 g06529(new_n6905, new_n6901, new_n6906);
not_4  g06530(new_n6906, new_n6907);
xnor_1 g06531(new_n6907, new_n6900, new_n6908);
not_4  g06532(new_n6874, new_n6909);
nand_1 g06533(new_n6876, new_n6909, new_n6910);
nand_1 g06534(n7456, n6770, new_n6911);
xnor_1 g06535(new_n6911, new_n6910, new_n6912);
nand_1 g06536(n3932, n3627, new_n6913);
nand_1 g06537(n12591, n9920, new_n6914);
nand_1 g06538(n4516, n1798, new_n6915);
nand_1 g06539(new_n6915, new_n6914, new_n6916);
not_4  g06540(new_n6914, new_n6917);
not_4  g06541(new_n6915, new_n6918);
nand_1 g06542(new_n6918, new_n6917, new_n6919);
nand_1 g06543(new_n6919, new_n6916, new_n6920);
xnor_1 g06544(new_n6920, new_n6913, new_n6921);
not_4  g06545(new_n6921, new_n6922);
xnor_1 g06546(new_n6922, new_n6912, new_n6923);
xnor_1 g06547(new_n6923, new_n6908, new_n6924);
nand_1 g06548(new_n6870, new_n6866, new_n6925);
nor_1  g06549(new_n6868, new_n6867, new_n6926);
nor_1  g06550(new_n6884, new_n6871, new_n6927);
xnor_1 g06551(new_n6927, new_n6926, new_n6928);
nand_1 g06552(new_n6928, new_n6925, new_n6929);
xnor_1 g06553(new_n6929, new_n6924, new_n6930);
xnor_1 g06554(new_n6930, new_n6896, new_n6931);
nand_1 g06555(n10327, n6687, new_n6932);
not_4  g06556(new_n6932, new_n6933);
xnor_1 g06557(new_n6894, new_n6885, new_n6934);
nand_1 g06558(new_n6934, new_n6933, new_n6935);
not_4  g06559(new_n4115, new_n6936);
xnor_1 g06560(new_n6892, new_n6890, new_n6937);
nand_1 g06561(new_n6937, new_n6936, new_n6938);
not_4  g06562(new_n6938, new_n6939);
xnor_1 g06563(new_n6934, new_n6932, new_n6940);
nand_1 g06564(new_n6940, new_n6939, new_n6941);
nand_1 g06565(new_n6941, new_n6935, new_n6942);
xnor_1 g06566(new_n6942, new_n6931, new_n6943);
not_4  g06567(new_n6943, new_n6944);
nand_1 g06568(n3022, n2226, new_n6945);
nand_1 g06569(n9640, n1094, new_n6946);
nand_1 g06570(n10678, n6703, new_n6947);
not_4  g06571(new_n6947, new_n6948);
xnor_1 g06572(new_n6948, new_n6946, new_n6949);
xnor_1 g06573(new_n6949, new_n6945, new_n6950);
nand_1 g06574(n6703, n1094, new_n6951);
nand_1 g06575(new_n6951, new_n4157, new_n6952);
nor_1  g06576(new_n6951, new_n4157, new_n6953);
not_4  g06577(new_n6953, new_n6954);
nand_1 g06578(n9640, n2226, new_n6955);
nand_1 g06579(new_n6955, new_n6954, new_n6956);
nand_1 g06580(new_n6956, new_n6952, new_n6957);
xnor_1 g06581(new_n6957, new_n6950, new_n6958);
not_4  g06582(new_n6958, new_n6959);
nand_1 g06583(n10928, n10451, new_n6960);
nand_1 g06584(n11023, n6986, new_n6961);
not_4  g06585(new_n6961, new_n6962);
xnor_1 g06586(new_n6962, new_n6960, new_n6963);
xnor_1 g06587(new_n6963, new_n6959, new_n6964);
nand_1 g06588(n11023, n10928, new_n6965);
nand_1 g06589(new_n4276, new_n4269, new_n6966);
nand_1 g06590(new_n6966, new_n4273, new_n6967);
nor_1  g06591(new_n6967, new_n6965, new_n6968);
not_4  g06592(new_n6967, new_n6969);
xnor_1 g06593(new_n6969, new_n6965, new_n6970);
not_4  g06594(new_n6970, new_n6971);
nand_1 g06595(new_n6954, new_n6952, new_n6972);
xnor_1 g06596(new_n6972, new_n6955, new_n6973);
nor_1  g06597(new_n6973, new_n6971, new_n6974);
nor_1  g06598(new_n6974, new_n6968, new_n6975);
not_4  g06599(new_n6975, new_n6976);
xnor_1 g06600(new_n6976, new_n6964, new_n6977);
not_4  g06601(new_n6977, new_n6978);
nand_1 g06602(n10451, n8336, new_n6979);
not_4  g06603(new_n6979, new_n6980);
xnor_1 g06604(new_n6973, new_n6970, new_n6981);
nand_1 g06605(new_n6981, new_n6980, new_n6982);
not_4  g06606(new_n4268, new_n6983);
nand_1 g06607(new_n4278, new_n6983, new_n6984);
nand_1 g06608(new_n6984, new_n4266, new_n6985);
xnor_1 g06609(new_n6981, new_n6979, new_n6986_1);
nand_1 g06610(new_n6986_1, new_n6985, new_n6987);
nand_1 g06611(new_n6987, new_n6982, new_n6988);
nand_1 g06612(new_n6988, new_n6978, new_n6989);
not_4  g06613(new_n6945, new_n6990);
nand_1 g06614(new_n6949, new_n6990, new_n6991);
not_4  g06615(new_n6950, new_n6992);
nor_1  g06616(new_n6957, new_n6992, new_n6993);
not_4  g06617(new_n6993, new_n6994);
nand_1 g06618(new_n6994, new_n6991, new_n6995);
nand_1 g06619(n10928, n10278, new_n6996);
nand_1 g06620(n10451, n6986, new_n6997);
not_4  g06621(new_n6997, new_n6998);
nand_1 g06622(n11423, n8336, new_n6999);
not_4  g06623(new_n6999, new_n7000);
xnor_1 g06624(new_n7000, new_n6998, new_n7001);
xnor_1 g06625(new_n7001, new_n6996, new_n7002);
xnor_1 g06626(new_n7002, new_n6995, new_n7003);
not_4  g06627(new_n7003, new_n7004);
not_4  g06628(new_n6946, new_n7005);
nand_1 g06629(new_n6948, new_n7005, new_n7006);
nand_1 g06630(n11023, n2226, new_n7007);
not_4  g06631(new_n7007, new_n7008);
xnor_1 g06632(new_n7008, new_n7006, new_n7009);
nand_1 g06633(n10678, n9640, new_n7010);
nand_1 g06634(n3022, n1094, new_n7011);
nand_1 g06635(n7320, n6703, new_n7012);
not_4  g06636(new_n7012, new_n7013);
xnor_1 g06637(new_n7013, new_n7011, new_n7014);
xnor_1 g06638(new_n7014, new_n7010, new_n7015);
xnor_1 g06639(new_n7015, new_n7009, new_n7016);
xnor_1 g06640(new_n7016, new_n7004, new_n7017);
nand_1 g06641(new_n6963, new_n6958, new_n7018);
nor_1  g06642(new_n6961, new_n6960, new_n7019);
nand_1 g06643(new_n6976, new_n6964, new_n7020);
not_4  g06644(new_n7020, new_n7021);
xnor_1 g06645(new_n7021, new_n7019, new_n7022);
nand_1 g06646(new_n7022, new_n7018, new_n7023);
xnor_1 g06647(new_n7023, new_n7017, new_n7024);
xnor_1 g06648(new_n7024, new_n6989, new_n7025);
nand_1 g06649(n10278, n8336, new_n7026);
not_4  g06650(new_n7026, new_n7027);
xnor_1 g06651(new_n6988, new_n6977, new_n7028);
nor_1  g06652(new_n7028, new_n7027, new_n7029);
not_4  g06653(new_n7029, new_n7030);
not_4  g06654(new_n4280, new_n7031);
nand_1 g06655(new_n7031, new_n4279, new_n7032);
xnor_1 g06656(new_n6986_1, new_n6985, new_n7033);
nor_1  g06657(new_n7033, new_n7032, new_n7034);
not_4  g06658(new_n7034, new_n7035);
xnor_1 g06659(new_n7028, new_n7026, new_n7036);
nand_1 g06660(new_n7036, new_n7035, new_n7037);
nand_1 g06661(new_n7037, new_n7030, new_n7038);
xnor_1 g06662(new_n7038, new_n7025, new_n7039);
not_4  g06663(new_n7039, new_n7040);
nand_1 g06664(n8665, n7160, new_n7041);
nand_1 g06665(n4828, n1067, new_n7042);
nand_1 g06666(n5645, n2515, new_n7043);
not_4  g06667(new_n7043, new_n7044);
xnor_1 g06668(new_n7044, new_n7042, new_n7045);
xnor_1 g06669(new_n7045, new_n7041, new_n7046);
not_4  g06670(new_n7046, new_n7047);
nand_1 g06671(n5645, n4828, new_n7048);
nand_1 g06672(n8665, n7891, new_n7049);
nand_1 g06673(new_n7049, new_n7048, new_n7050);
nand_1 g06674(n7160, n1067, new_n7051);
xnor_1 g06675(new_n7049, new_n7048, new_n7052);
not_4  g06676(new_n7052, new_n7053);
nand_1 g06677(new_n7053, new_n7051, new_n7054);
nand_1 g06678(new_n7054, new_n7050, new_n7055);
xnor_1 g06679(new_n7055, new_n7047, new_n7056);
nand_1 g06680(n12391, n2551, new_n7057);
nand_1 g06681(n11922, n7891, new_n7058);
nand_1 g06682(new_n7058, new_n7057, new_n7059);
not_4  g06683(new_n7057, new_n7060);
not_4  g06684(new_n7058, new_n7061);
nand_1 g06685(new_n7061, new_n7060, new_n7062);
nand_1 g06686(new_n7062, new_n7059, new_n7063);
not_4  g06687(new_n7063, new_n7064);
xnor_1 g06688(new_n7064, new_n7056, new_n7065);
nand_1 g06689(n12391, n11922, new_n7066);
nand_1 g06690(new_n4230_1, new_n4229, new_n7067);
nand_1 g06691(new_n4234, new_n7067, new_n7068);
nor_1  g06692(new_n7068, new_n7066, new_n7069);
not_4  g06693(new_n7069, new_n7070);
xnor_1 g06694(new_n7053, new_n7051, new_n7071);
not_4  g06695(new_n7068, new_n7072);
xnor_1 g06696(new_n7072, new_n7066, new_n7073);
nand_1 g06697(new_n7073, new_n7071, new_n7074);
nand_1 g06698(new_n7074, new_n7070, new_n7075);
xnor_1 g06699(new_n7075, new_n7065, new_n7076);
not_4  g06700(new_n7076, new_n7077);
nand_1 g06701(n12069, n2551, new_n7078);
not_4  g06702(new_n7078, new_n7079);
xnor_1 g06703(new_n7073, new_n7071, new_n7080);
not_4  g06704(new_n7080, new_n7081);
nand_1 g06705(new_n7081, new_n7079, new_n7082);
nand_1 g06706(new_n7080, new_n7078, new_n7083);
nor_1  g06707(new_n4225, new_n4222, new_n7084);
not_4  g06708(new_n7084, new_n7085);
not_4  g06709(new_n4236, new_n7086);
nand_1 g06710(new_n7086, new_n4227, new_n7087);
nand_1 g06711(new_n7087, new_n7085, new_n7088);
nand_1 g06712(new_n7088, new_n7083, new_n7089);
nand_1 g06713(new_n7089, new_n7082, new_n7090);
nand_1 g06714(new_n7090, new_n7077, new_n7091);
not_4  g06715(new_n7041, new_n7092);
nand_1 g06716(new_n7045, new_n7092, new_n7093);
not_4  g06717(new_n7093, new_n7094);
not_4  g06718(new_n7055, new_n7095);
nand_1 g06719(new_n7095, new_n7046, new_n7096);
not_4  g06720(new_n7096, new_n7097);
nor_1  g06721(new_n7097, new_n7094, new_n7098);
nand_1 g06722(n12826, n12391, new_n7099);
not_4  g06723(new_n7099, new_n7100);
nand_1 g06724(n7891, n2551, new_n7101);
nand_1 g06725(n12069, n4094, new_n7102);
not_4  g06726(new_n7102, new_n7103);
xnor_1 g06727(new_n7103, new_n7101, new_n7104);
xnor_1 g06728(new_n7104, new_n7100, new_n7105);
not_4  g06729(new_n7105, new_n7106);
xnor_1 g06730(new_n7106, new_n7098, new_n7107);
not_4  g06731(new_n7042, new_n7108);
nand_1 g06732(new_n7044, new_n7108, new_n7109);
nand_1 g06733(n11922, n7160, new_n7110);
nand_1 g06734(new_n7110, new_n7109, new_n7111);
not_4  g06735(new_n7109, new_n7112);
not_4  g06736(new_n7110, new_n7113);
nand_1 g06737(new_n7113, new_n7112, new_n7114);
nand_1 g06738(new_n7114, new_n7111, new_n7115);
nand_1 g06739(n2515, n1067, new_n7116);
nand_1 g06740(n8665, n4828, new_n7117);
nand_1 g06741(n5645, n1199, new_n7118);
nand_1 g06742(new_n7118, new_n7117, new_n7119);
not_4  g06743(new_n7117, new_n7120);
not_4  g06744(new_n7118, new_n7121);
nand_1 g06745(new_n7121, new_n7120, new_n7122);
nand_1 g06746(new_n7122, new_n7119, new_n7123);
xnor_1 g06747(new_n7123, new_n7116, new_n7124);
not_4  g06748(new_n7124, new_n7125);
xnor_1 g06749(new_n7125, new_n7115, new_n7126);
not_4  g06750(new_n7126, new_n7127);
xnor_1 g06751(new_n7127, new_n7107, new_n7128);
not_4  g06752(new_n7056, new_n7129);
nand_1 g06753(new_n7064, new_n7129, new_n7130);
nand_1 g06754(new_n7075, new_n7065, new_n7131);
xnor_1 g06755(new_n7131, new_n7062, new_n7132);
nand_1 g06756(new_n7132, new_n7130, new_n7133);
not_4  g06757(new_n7133, new_n7134);
xnor_1 g06758(new_n7134, new_n7128, new_n7135);
xnor_1 g06759(new_n7135, new_n7091, new_n7136);
nand_1 g06760(n12826, n12069, new_n7137);
xnor_1 g06761(new_n7090, new_n7076, new_n7138);
not_4  g06762(new_n7138, new_n7139);
nand_1 g06763(new_n7139, new_n7137, new_n7140);
nand_1 g06764(new_n4237, new_n4221, new_n7141);
not_4  g06765(new_n7088, new_n7142);
nand_1 g06766(new_n7083, new_n7082, new_n7143);
xnor_1 g06767(new_n7143, new_n7142, new_n7144);
nor_1  g06768(new_n7144, new_n7141, new_n7145);
not_4  g06769(new_n7145, new_n7146);
xnor_1 g06770(new_n7138, new_n7137, new_n7147);
nand_1 g06771(new_n7147, new_n7146, new_n7148);
nand_1 g06772(new_n7148, new_n7140, new_n7149);
xnor_1 g06773(new_n7149, new_n7136, new_n7150);
nand_1 g06774(n3754, n996, new_n7151);
nand_1 g06775(n10898, n5767, new_n7152);
nand_1 g06776(n11876, n5319, new_n7153);
not_4  g06777(new_n7153, new_n7154);
xnor_1 g06778(new_n7154, new_n7152, new_n7155);
xnor_1 g06779(new_n7155, new_n7151, new_n7156);
nand_1 g06780(n10898, n996, new_n7157);
nand_1 g06781(new_n7157, new_n4191, new_n7158);
nand_1 g06782(n11876, n5767, new_n7159_1);
not_4  g06783(new_n7157, new_n7160_1);
xnor_1 g06784(new_n7160_1, new_n4191, new_n7161);
nand_1 g06785(new_n7161, new_n7159_1, new_n7162);
nand_1 g06786(new_n7162, new_n7158, new_n7163);
not_4  g06787(new_n7163, new_n7164);
xnor_1 g06788(new_n7164, new_n7156, new_n7165);
nand_1 g06789(n11153, n159, new_n7166);
nand_1 g06790(n5314, n2749, new_n7167);
not_4  g06791(new_n7167, new_n7168);
xnor_1 g06792(new_n7168, new_n7166, new_n7169);
xnor_1 g06793(new_n7169, new_n7165, new_n7170);
nand_1 g06794(n11153, n2749, new_n7171);
nand_1 g06795(new_n4246, new_n4245, new_n7172);
nand_1 g06796(new_n4248, new_n4244, new_n7173);
nand_1 g06797(new_n7173, new_n7172, new_n7174);
nor_1  g06798(new_n7174, new_n7171, new_n7175);
not_4  g06799(new_n7175, new_n7176);
not_4  g06800(new_n7174, new_n7177);
xnor_1 g06801(new_n7177, new_n7171, new_n7178);
not_4  g06802(new_n7161, new_n7179);
xnor_1 g06803(new_n7179, new_n7159_1, new_n7180);
not_4  g06804(new_n7180, new_n7181);
nand_1 g06805(new_n7181, new_n7178, new_n7182);
nand_1 g06806(new_n7182, new_n7176, new_n7183);
xnor_1 g06807(new_n7183, new_n7170, new_n7184);
not_4  g06808(new_n7184, new_n7185);
nand_1 g06809(n11222, n159, new_n7186);
not_4  g06810(new_n7186, new_n7187);
xnor_1 g06811(new_n7181, new_n7178, new_n7188);
not_4  g06812(new_n7188, new_n7189);
nand_1 g06813(new_n7189, new_n7187, new_n7190);
nand_1 g06814(new_n7188, new_n7186, new_n7191);
nor_1  g06815(new_n4241, new_n4239, new_n7192);
not_4  g06816(new_n4243, new_n7193_1);
nor_1  g06817(new_n4250, new_n7193_1, new_n7194);
nor_1  g06818(new_n7194, new_n7192, new_n7195);
not_4  g06819(new_n7195, new_n7196);
nand_1 g06820(new_n7196, new_n7191, new_n7197);
nand_1 g06821(new_n7197, new_n7190, new_n7198);
nand_1 g06822(new_n7198, new_n7185, new_n7199);
not_4  g06823(new_n7165, new_n7200);
nand_1 g06824(new_n7169, new_n7200, new_n7201);
nor_1  g06825(new_n7167, new_n7166, new_n7202);
nand_1 g06826(new_n7183, new_n7170, new_n7203);
not_4  g06827(new_n7203, new_n7204);
xnor_1 g06828(new_n7204, new_n7202, new_n7205);
nand_1 g06829(new_n7205, new_n7201, new_n7206);
not_4  g06830(new_n7151, new_n7207);
nand_1 g06831(new_n7155, new_n7207, new_n7208);
nand_1 g06832(new_n7164, new_n7156, new_n7209);
nand_1 g06833(new_n7209, new_n7208, new_n7210);
nand_1 g06834(n11153, n1510, new_n7211);
nand_1 g06835(n5314, n159, new_n7212);
nand_1 g06836(n12247, n11222, new_n7213);
not_4  g06837(new_n7213, new_n7214);
xnor_1 g06838(new_n7214, new_n7212, new_n7215);
xnor_1 g06839(new_n7215, new_n7211, new_n7216);
xnor_1 g06840(new_n7216, new_n7210, new_n7217);
not_4  g06841(new_n7152, new_n7218);
nand_1 g06842(new_n7154, new_n7218, new_n7219);
nand_1 g06843(n2749, n996, new_n7220);
not_4  g06844(new_n7220, new_n7221);
xnor_1 g06845(new_n7221, new_n7219, new_n7222);
nand_1 g06846(n10898, n5319, new_n7223);
nand_1 g06847(n11876, n9457, new_n7224);
nand_1 g06848(n5767, n3754, new_n7225);
not_4  g06849(new_n7225, new_n7226);
xnor_1 g06850(new_n7226, new_n7224, new_n7227);
xnor_1 g06851(new_n7227, new_n7223, new_n7228);
not_4  g06852(new_n7228, new_n7229);
xnor_1 g06853(new_n7229, new_n7222, new_n7230);
xnor_1 g06854(new_n7230, new_n7217, new_n7231);
not_4  g06855(new_n7231, new_n7232);
xnor_1 g06856(new_n7232, new_n7206, new_n7233);
xnor_1 g06857(new_n7233, new_n7199, new_n7234);
nand_1 g06858(n11222, n1510, new_n7235);
not_4  g06859(new_n7235, new_n7236_1);
xnor_1 g06860(new_n7198, new_n7184, new_n7237);
nor_1  g06861(new_n7237, new_n7236_1, new_n7238);
not_4  g06862(new_n4251, new_n7239);
nor_1  g06863(new_n4252, new_n7239, new_n7240);
nand_1 g06864(new_n7191, new_n7190, new_n7241);
xnor_1 g06865(new_n7241, new_n7196, new_n7242);
nand_1 g06866(new_n7242, new_n7240, new_n7243);
not_4  g06867(new_n7243, new_n7244);
not_4  g06868(new_n7238, new_n7245);
nand_1 g06869(new_n7237, new_n7236_1, new_n7246);
nand_1 g06870(new_n7246, new_n7245, new_n7247);
nor_1  g06871(new_n7247, new_n7244, new_n7248);
nor_1  g06872(new_n7248, new_n7238, new_n7249);
xnor_1 g06873(new_n7249, new_n7234, new_n7250);
not_4  g06874(new_n7250, new_n7251);
xnor_1 g06875(new_n7247, new_n7244, new_n7252);
xnor_1 g06876(new_n7147, new_n7145, new_n7253);
not_4  g06877(new_n7253, new_n7254);
nand_1 g06878(new_n7254, new_n7252, new_n7255);
xnor_1 g06879(new_n7247, new_n7243, new_n7256);
nand_1 g06880(new_n7253, new_n7256, new_n7257);
nand_1 g06881(new_n7144, new_n7141, new_n7258);
nand_1 g06882(new_n7258, new_n7146, new_n7259);
not_4  g06883(new_n4238, new_n7260);
nor_1  g06884(new_n4253, new_n7260, new_n7261);
not_4  g06885(new_n7261, new_n7262);
nand_1 g06886(new_n4259, new_n4254, new_n7263);
nand_1 g06887(new_n7263, new_n7262, new_n7264);
nand_1 g06888(new_n7264, new_n7259, new_n7265_1);
xnor_1 g06889(new_n7242, new_n7240, new_n7266);
xnor_1 g06890(new_n7264, new_n7259, new_n7267);
not_4  g06891(new_n7267, new_n7268);
nand_1 g06892(new_n7268, new_n7266, new_n7269);
nand_1 g06893(new_n7269, new_n7265_1, new_n7270_1);
not_4  g06894(new_n7270_1, new_n7271);
nand_1 g06895(new_n7271, new_n7257, new_n7272);
nand_1 g06896(new_n7272, new_n7255, new_n7273);
nand_1 g06897(new_n7273, new_n7251, new_n7274);
not_4  g06898(new_n7255, new_n7275);
nor_1  g06899(new_n7254, new_n7252, new_n7276);
nor_1  g06900(new_n7270_1, new_n7276, new_n7277);
nor_1  g06901(new_n7277, new_n7275, new_n7278);
nand_1 g06902(new_n7278, new_n7250, new_n7279);
nand_1 g06903(new_n7279, new_n7274, new_n7280);
not_4  g06904(new_n7280, new_n7281);
xnor_1 g06905(new_n7281, new_n7150, new_n7282);
nor_1  g06906(new_n7282, new_n7040, new_n7283);
not_4  g06907(new_n7283, new_n7284);
nand_1 g06908(new_n7282, new_n7040, new_n7285);
nand_1 g06909(new_n7285, new_n7284, new_n7286);
xnor_1 g06910(new_n7036, new_n7034, new_n7287);
not_4  g06911(new_n7287, new_n7288);
nand_1 g06912(new_n7033, new_n7032, new_n7289);
nand_1 g06913(new_n7289, new_n7035, new_n7290);
xnor_1 g06914(new_n7267, new_n7266, new_n7291);
nor_1  g06915(new_n7291, new_n7290, new_n7292);
not_4  g06916(new_n7292, new_n7293);
nand_1 g06917(new_n4293, new_n4288, new_n7294_1);
nand_1 g06918(new_n7291, new_n7290, new_n7295);
nand_1 g06919(new_n7295, new_n7293, new_n7296);
not_4  g06920(new_n7296, new_n7297);
nand_1 g06921(new_n7297, new_n7294_1, new_n7298);
nand_1 g06922(new_n7298, new_n7293, new_n7299);
nand_1 g06923(new_n7299, new_n7288, new_n7300);
not_4  g06924(new_n7299, new_n7301);
xnor_1 g06925(new_n7301, new_n7288, new_n7302);
nand_1 g06926(new_n7257, new_n7255, new_n7303);
not_4  g06927(new_n7303, new_n7304);
xnor_1 g06928(new_n7304, new_n7270_1, new_n7305);
nand_1 g06929(new_n7305, new_n7302, new_n7306);
nand_1 g06930(new_n7306, new_n7300, new_n7307);
not_4  g06931(new_n7307, new_n7308);
nor_1  g06932(new_n7308, new_n7286, new_n7309);
not_4  g06933(new_n7309, new_n7310);
nand_1 g06934(new_n7308, new_n7286, new_n7311);
nand_1 g06935(new_n7311, new_n7310, new_n7312);
not_4  g06936(new_n7312, new_n7313);
nand_1 g06937(new_n7313, new_n6944, new_n7314);
nand_1 g06938(new_n7312, new_n6943, new_n7315);
nand_1 g06939(new_n7315, new_n7314, new_n7316);
xnor_1 g06940(new_n6940, new_n6938, new_n7317);
xnor_1 g06941(new_n7305, new_n7302, new_n7318);
not_4  g06942(new_n7318, new_n7319);
nand_1 g06943(new_n7319, new_n7317, new_n7320_1);
not_4  g06944(new_n7317, new_n7321);
nand_1 g06945(new_n7318, new_n7321, new_n7322);
xnor_1 g06946(new_n6937, new_n4115, new_n7323);
xnor_1 g06947(new_n7296, new_n7294_1, new_n7324);
nor_1  g06948(new_n7324, new_n7323, new_n7325);
not_4  g06949(new_n4117, new_n7326);
nand_1 g06950(new_n4218, new_n7326, new_n7327);
not_4  g06951(new_n4294, new_n7328);
nand_1 g06952(new_n7328, new_n4219, new_n7329);
nand_1 g06953(new_n7329, new_n7327, new_n7330);
xnor_1 g06954(new_n7324, new_n7323, new_n7331);
nor_1  g06955(new_n7331, new_n7330, new_n7332);
nor_1  g06956(new_n7332, new_n7325, new_n7333);
nand_1 g06957(new_n7333, new_n7322, new_n7334);
nand_1 g06958(new_n7334, new_n7320_1, new_n7335);
xnor_1 g06959(new_n7335, new_n7316, n2301);
xnor_1 g06960(new_n4216, new_n4214, n2316);
nand_1 g06961(n4634, n1333, new_n7338);
nand_1 g06962(new_n6605, new_n6599, new_n7339);
nand_1 g06963(new_n7339, new_n6603, new_n7340);
nor_1  g06964(new_n7340, new_n7338, new_n7341);
not_4  g06965(new_n7341, new_n7342);
nand_1 g06966(new_n7340, new_n7338, new_n7343);
nand_1 g06967(new_n7343, new_n7342, new_n7344);
not_4  g06968(new_n7344, new_n7345);
nand_1 g06969(n11757, n2879, new_n7346);
nand_1 g06970(n7265, n5240, new_n7347);
nand_1 g06971(new_n7347, new_n6589, new_n7348);
not_4  g06972(new_n7347, new_n7349);
nand_1 g06973(new_n7349, new_n6590, new_n7350);
nand_1 g06974(new_n7350, new_n7348, new_n7351);
xnor_1 g06975(new_n7351, new_n7346, new_n7352);
not_4  g06976(new_n7352, new_n7353);
nand_1 g06977(new_n7353, new_n7345, new_n7354_1);
nand_1 g06978(new_n7354_1, new_n7342, new_n7355);
nand_1 g06979(n4634, n3172, new_n7356);
nand_1 g06980(n9195, n1333, new_n7357);
not_4  g06981(new_n7357, new_n7358);
xnor_1 g06982(new_n7358, new_n7356, new_n7359);
xnor_1 g06983(new_n7359, new_n7355, new_n7360);
nand_1 g06984(n11757, n10223, new_n7361);
nand_1 g06985(n5240, n2879, new_n7362);
nand_1 g06986(n11821, n7265, new_n7363);
nand_1 g06987(new_n7363, new_n7362, new_n7364);
not_4  g06988(new_n7362, new_n7365);
not_4  g06989(new_n7363, new_n7366);
nand_1 g06990(new_n7366, new_n7365, new_n7367);
nand_1 g06991(new_n7367, new_n7364, new_n7368);
xnor_1 g06992(new_n7368, new_n7361, new_n7369);
nand_1 g06993(new_n7350, new_n7346, new_n7370);
nand_1 g06994(new_n7370, new_n7348, new_n7371);
xnor_1 g06995(new_n7371, new_n7369, new_n7372);
xnor_1 g06996(new_n7372, new_n7360, new_n7373);
not_4  g06997(new_n7373, new_n7374);
nand_1 g06998(n9195, n7862, new_n7375);
not_4  g06999(new_n7375, new_n7376);
nand_1 g07000(new_n7352, new_n7344, new_n7377);
nand_1 g07001(new_n7377, new_n7354_1, new_n7378);
not_4  g07002(new_n7378, new_n7379);
nand_1 g07003(new_n7379, new_n7376, new_n7380);
not_4  g07004(new_n6598, new_n7381);
nand_1 g07005(new_n6607, new_n7381, new_n7382);
nand_1 g07006(new_n7382, new_n6596, new_n7383);
xnor_1 g07007(new_n7379, new_n7375, new_n7384);
nand_1 g07008(new_n7384, new_n7383, new_n7385);
nand_1 g07009(new_n7385, new_n7380, new_n7386);
nand_1 g07010(new_n7386, new_n7374, new_n7387);
nand_1 g07011(new_n7368, new_n7361, new_n7388_1);
not_4  g07012(new_n7369, new_n7389);
nand_1 g07013(new_n7371, new_n7389, new_n7390);
nand_1 g07014(new_n7390, new_n7388_1, new_n7391);
nand_1 g07015(n2253, n1333, new_n7392);
nand_1 g07016(n9195, n3172, new_n7393);
not_4  g07017(new_n7393, new_n7394);
nand_1 g07018(n7862, n3865, new_n7395);
not_4  g07019(new_n7395, new_n7396);
nand_1 g07020(new_n7396, new_n7394, new_n7397);
nand_1 g07021(new_n7395, new_n7393, new_n7398);
nand_1 g07022(new_n7398, new_n7397, new_n7399);
xnor_1 g07023(new_n7399, new_n7392, new_n7400);
xnor_1 g07024(new_n7400, new_n7391, new_n7401);
nand_1 g07025(n11757, n4634, new_n7402);
xnor_1 g07026(new_n7402, new_n7367, new_n7403);
nand_1 g07027(n11821, n2879, new_n7404);
not_4  g07028(new_n7404, new_n7405);
nand_1 g07029(n10223, n5240, new_n7406);
nand_1 g07030(n9080, n7265, new_n7407);
not_4  g07031(new_n7407, new_n7408);
xnor_1 g07032(new_n7408, new_n7406, new_n7409);
xnor_1 g07033(new_n7409, new_n7405, new_n7410);
xnor_1 g07034(new_n7410, new_n7403, new_n7411);
xnor_1 g07035(new_n7411, new_n7401, new_n7412);
nand_1 g07036(new_n7359, new_n7355, new_n7413);
nor_1  g07037(new_n7357, new_n7356, new_n7414);
nor_1  g07038(new_n7372, new_n7360, new_n7415);
xnor_1 g07039(new_n7415, new_n7414, new_n7416);
nand_1 g07040(new_n7416, new_n7413, new_n7417);
xnor_1 g07041(new_n7417, new_n7412, new_n7418);
xnor_1 g07042(new_n7418, new_n7387, new_n7419);
nand_1 g07043(n7862, n2253, new_n7420);
not_4  g07044(new_n7420, new_n7421);
xnor_1 g07045(new_n7386, new_n7373, new_n7422);
nand_1 g07046(new_n7422, new_n7421, new_n7423);
not_4  g07047(new_n6608, new_n7424);
nor_1  g07048(new_n6614, new_n7424, new_n7425);
xnor_1 g07049(new_n7384, new_n7383, new_n7426);
not_4  g07050(new_n7426, new_n7427);
nand_1 g07051(new_n7427, new_n7425, new_n7428);
not_4  g07052(new_n7428, new_n7429);
xnor_1 g07053(new_n7422, new_n7420, new_n7430);
nand_1 g07054(new_n7430, new_n7429, new_n7431);
nand_1 g07055(new_n7431, new_n7423, new_n7432);
xnor_1 g07056(new_n7432, new_n7419, new_n7433);
xnor_1 g07057(new_n7430, new_n7428, new_n7434);
xnor_1 g07058(new_n7426, new_n7425, new_n7435);
nand_1 g07059(n12145, n6877, new_n7436_1);
nand_1 g07060(n9400, n2522, new_n7437);
nand_1 g07061(n11311, n2024, new_n7438);
not_4  g07062(new_n7438, new_n7439);
nand_1 g07063(n7946, n4187, new_n7440);
nand_1 g07064(new_n7440, new_n6633, new_n7441);
not_4  g07065(new_n7440, new_n7442);
nand_1 g07066(new_n7442, new_n6634, new_n7443);
nand_1 g07067(new_n7443, new_n7441, new_n7444);
xnor_1 g07068(new_n7444, new_n7439, new_n7445);
not_4  g07069(new_n7445, new_n7446);
xnor_1 g07070(new_n7446, new_n7437, new_n7447);
nand_1 g07071(new_n6620, new_n6619, new_n7448);
nand_1 g07072(new_n6622, new_n6617, new_n7449);
nand_1 g07073(new_n7449, new_n7448, new_n7450);
xnor_1 g07074(new_n7450, new_n7447, new_n7451);
nor_1  g07075(new_n7451, new_n7436_1, new_n7452);
not_4  g07076(new_n7452, new_n7453);
nand_1 g07077(new_n7451, new_n7436_1, new_n7454);
nand_1 g07078(new_n7454, new_n7453, new_n7455);
not_4  g07079(new_n7455, new_n7456_1);
nand_1 g07080(new_n6640, new_n6625, new_n7457);
nand_1 g07081(new_n7457, new_n7456_1, new_n7458);
not_4  g07082(new_n7457, new_n7459);
nand_1 g07083(new_n7459, new_n7455, new_n7460);
nand_1 g07084(new_n7460, new_n7458, new_n7461);
not_4  g07085(new_n7461, new_n7462);
xnor_1 g07086(new_n7462, new_n6652, new_n7463);
not_4  g07087(new_n6731, new_n7464);
nand_1 g07088(new_n7464, new_n6654, new_n7465);
nand_1 g07089(new_n6773, new_n6732, new_n7466);
nand_1 g07090(new_n7466, new_n7465, new_n7467);
xnor_1 g07091(new_n7467, new_n7463, new_n7468);
nand_1 g07092(new_n6749, new_n6748, new_n7469);
nand_1 g07093(n11478, n521, new_n7470);
nand_1 g07094(new_n6744, new_n6738, new_n7471);
nand_1 g07095(new_n7471, new_n6741, new_n7472);
not_4  g07096(new_n7472, new_n7473);
xnor_1 g07097(new_n7473, new_n7470, new_n7474);
nand_1 g07098(n2498, n137, new_n7475);
not_4  g07099(new_n7475, new_n7476);
nand_1 g07100(n5579, n5283, new_n7477);
nand_1 g07101(n6294, n2558, new_n7478);
nand_1 g07102(new_n7478, new_n7477, new_n7479);
not_4  g07103(new_n7477, new_n7480);
not_4  g07104(new_n7478, new_n7481);
nand_1 g07105(new_n7481, new_n7480, new_n7482);
nand_1 g07106(new_n7482, new_n7479, new_n7483);
xnor_1 g07107(new_n7483, new_n7476, new_n7484);
xnor_1 g07108(new_n7484, new_n7474, new_n7485);
not_4  g07109(new_n7485, new_n7486);
nand_1 g07110(n6016, n4805, new_n7487);
nor_1  g07111(new_n6736, new_n6734, new_n7488);
nor_1  g07112(new_n6746, new_n6737, new_n7489);
nor_1  g07113(new_n7489, new_n7488, new_n7490);
not_4  g07114(new_n7490, new_n7491);
xnor_1 g07115(new_n7491, new_n7487, new_n7492);
xnor_1 g07116(new_n7492, new_n7486, new_n7493);
nor_1  g07117(new_n7493, new_n7469, new_n7494);
not_4  g07118(new_n7494, new_n7495);
nand_1 g07119(new_n7493, new_n7469, new_n7496);
nand_1 g07120(new_n7496, new_n7495, new_n7497);
not_4  g07121(new_n6765, new_n7498);
nand_1 g07122(new_n6766, new_n7498, new_n7499);
nand_1 g07123(n7270, n7236, new_n7500_1);
not_4  g07124(new_n7500_1, new_n7501);
not_4  g07125(new_n6751, new_n7502);
nand_1 g07126(new_n6753, new_n7502, new_n7503);
nand_1 g07127(new_n6764, new_n6754, new_n7504);
nand_1 g07128(new_n7504, new_n7503, new_n7505);
xnor_1 g07129(new_n7505, new_n7501, new_n7506);
nand_1 g07130(n3992, n806, new_n7507);
nand_1 g07131(new_n6762, new_n6755, new_n7508);
nand_1 g07132(new_n7508, new_n6759, new_n7509);
not_4  g07133(new_n7509, new_n7510);
xnor_1 g07134(new_n7510, new_n7507, new_n7511);
nand_1 g07135(n9111, n6358, new_n7512);
not_4  g07136(new_n7512, new_n7513);
nand_1 g07137(n8384, n3342, new_n7514);
nand_1 g07138(n9763, n5198, new_n7515);
xnor_1 g07139(new_n7515, new_n7514, new_n7516);
xnor_1 g07140(new_n7516, new_n7513, new_n7517);
xnor_1 g07141(new_n7517, new_n7511, new_n7518);
xnor_1 g07142(new_n7518, new_n7506, new_n7519);
not_4  g07143(new_n7519, new_n7520);
xnor_1 g07144(new_n7520, new_n7499, new_n7521);
xnor_1 g07145(new_n7521, new_n7497, new_n7522);
not_4  g07146(new_n6767, new_n7523_1);
nand_1 g07147(new_n7523_1, new_n6750, new_n7524);
nand_1 g07148(new_n6772, new_n6768, new_n7525);
nand_1 g07149(new_n7525, new_n7524, new_n7526);
xnor_1 g07150(new_n7526, new_n7522, new_n7527);
xnor_1 g07151(new_n7527, new_n7468, new_n7528);
nor_1  g07152(new_n7528, new_n7435, new_n7529);
not_4  g07153(new_n7529, new_n7530);
nand_1 g07154(new_n7528, new_n7435, new_n7531);
nand_1 g07155(new_n7531, new_n7530, new_n7532);
not_4  g07156(new_n6798, new_n7533);
nand_1 g07157(new_n7533, new_n6775, new_n7534);
nand_1 g07158(new_n7534, new_n6777, new_n7535);
not_4  g07159(new_n7535, new_n7536);
nor_1  g07160(new_n7536, new_n7532, new_n7537);
nor_1  g07161(new_n7537, new_n7529, new_n7538);
nor_1  g07162(new_n7538, new_n7434, new_n7539);
not_4  g07163(new_n7539, new_n7540);
nor_1  g07164(new_n7467, new_n7463, new_n7541);
nor_1  g07165(new_n7527, new_n7468, new_n7542);
nor_1  g07166(new_n7542, new_n7541, new_n7543);
not_4  g07167(new_n6652, new_n7544);
nand_1 g07168(new_n7462, new_n7544, new_n7545);
nand_1 g07169(n12221, n6877, new_n7546_1);
nand_1 g07170(new_n7458, new_n7453, new_n7547);
nand_1 g07171(new_n7446, new_n7437, new_n7548);
not_4  g07172(new_n7447, new_n7549);
nand_1 g07173(new_n7450, new_n7549, new_n7550);
nand_1 g07174(new_n7550, new_n7548, new_n7551);
nand_1 g07175(n11311, n9189, new_n7552);
nand_1 g07176(n7946, n4203, new_n7553);
nand_1 g07177(n4187, n2024, new_n7554);
nand_1 g07178(new_n7554, new_n7553, new_n7555);
not_4  g07179(new_n7553, new_n7556);
not_4  g07180(new_n7554, new_n7557);
nand_1 g07181(new_n7557, new_n7556, new_n7558);
nand_1 g07182(new_n7558, new_n7555, new_n7559);
xnor_1 g07183(new_n7559, new_n7552, new_n7560);
nand_1 g07184(new_n7443, new_n7438, new_n7561);
nand_1 g07185(new_n7561, new_n7441, new_n7562);
xnor_1 g07186(new_n7562, new_n7560, new_n7563);
nand_1 g07187(n12145, n9400, new_n7564);
nand_1 g07188(n2522, n2464, new_n7565);
nand_1 g07189(new_n7565, new_n7564, new_n7566);
not_4  g07190(new_n7564, new_n7567);
not_4  g07191(new_n7565, new_n7568_1);
nand_1 g07192(new_n7568_1, new_n7567, new_n7569);
nand_1 g07193(new_n7569, new_n7566, new_n7570);
nand_1 g07194(new_n7570, new_n7563, new_n7571);
nor_1  g07195(new_n7570, new_n7563, new_n7572);
not_4  g07196(new_n7572, new_n7573);
nand_1 g07197(new_n7573, new_n7571, new_n7574);
xnor_1 g07198(new_n7574, new_n7551, new_n7575);
xnor_1 g07199(new_n7575, new_n7547, new_n7576);
xnor_1 g07200(new_n7576, new_n7546_1, new_n7577);
xnor_1 g07201(new_n7577, new_n7545, new_n7578);
not_4  g07202(new_n7578, new_n7579);
xnor_1 g07203(new_n7579, new_n7543, new_n7580);
nor_1  g07204(new_n7519, new_n7499, new_n7581);
not_4  g07205(new_n7581, new_n7582);
nand_1 g07206(n7236, n5153, new_n7583);
not_4  g07207(new_n7583, new_n7584);
nand_1 g07208(n6358, n3342, new_n7585);
nand_1 g07209(n9111, n5198, new_n7586);
nand_1 g07210(n9763, n1471, new_n7587);
not_4  g07211(new_n7587, new_n7588);
xnor_1 g07212(new_n7588, new_n7586, new_n7589);
xnor_1 g07213(new_n7589, new_n7585, new_n7590);
nand_1 g07214(new_n7515, new_n7514, new_n7591);
not_4  g07215(new_n7591, new_n7592);
nor_1  g07216(new_n7516, new_n7513, new_n7593);
nor_1  g07217(new_n7593, new_n7592, new_n7594);
nand_1 g07218(new_n7594, new_n7590, new_n7595);
not_4  g07219(new_n7595, new_n7596);
nor_1  g07220(new_n7594, new_n7590, new_n7597);
nor_1  g07221(new_n7597, new_n7596, new_n7598);
nand_1 g07222(n7270, n3992, new_n7599);
nand_1 g07223(n8384, n806, new_n7600);
nand_1 g07224(new_n7600, new_n7599, new_n7601);
not_4  g07225(new_n7599, new_n7602);
not_4  g07226(new_n7600, new_n7603);
nand_1 g07227(new_n7603, new_n7602, new_n7604);
nand_1 g07228(new_n7604, new_n7601, new_n7605);
xnor_1 g07229(new_n7605, new_n7598, new_n7606);
nor_1  g07230(new_n7509, new_n7507, new_n7607);
not_4  g07231(new_n7607, new_n7608);
nand_1 g07232(new_n7517, new_n7511, new_n7609);
nand_1 g07233(new_n7609, new_n7608, new_n7610_1);
not_4  g07234(new_n7610_1, new_n7611);
xnor_1 g07235(new_n7611, new_n7606, new_n7612);
nor_1  g07236(new_n7505, new_n7501, new_n7613);
not_4  g07237(new_n7518, new_n7614);
nor_1  g07238(new_n7614, new_n7506, new_n7615);
nor_1  g07239(new_n7615, new_n7613, new_n7616);
nand_1 g07240(new_n7616, new_n7612, new_n7617);
not_4  g07241(new_n7617, new_n7618);
nor_1  g07242(new_n7616, new_n7612, new_n7619);
nor_1  g07243(new_n7619, new_n7618, new_n7620);
nand_1 g07244(new_n7620, new_n7584, new_n7621);
not_4  g07245(new_n7620, new_n7622);
nand_1 g07246(new_n7622, new_n7583, new_n7623);
nand_1 g07247(new_n7623, new_n7621, new_n7624);
xnor_1 g07248(new_n7624, new_n7582, new_n7625);
not_4  g07249(new_n7625, new_n7626);
nand_1 g07250(n5798, n4805, new_n7627);
nand_1 g07251(n5579, n137, new_n7628);
nand_1 g07252(n6797, n2558, new_n7629);
nand_1 g07253(n6294, n2498, new_n7630);
not_4  g07254(new_n7630, new_n7631);
xnor_1 g07255(new_n7631, new_n7629, new_n7632);
not_4  g07256(new_n7632, new_n7633);
xnor_1 g07257(new_n7633, new_n7628, new_n7634);
nand_1 g07258(new_n7482, new_n7475, new_n7635);
nand_1 g07259(new_n7635, new_n7479, new_n7636);
xnor_1 g07260(new_n7636, new_n7634, new_n7637);
nand_1 g07261(n11478, n6016, new_n7638);
nand_1 g07262(n5283, n521, new_n7639);
not_4  g07263(new_n7639, new_n7640);
xnor_1 g07264(new_n7640, new_n7638, new_n7641);
xnor_1 g07265(new_n7641, new_n7637, new_n7642);
nor_1  g07266(new_n7472, new_n7470, new_n7643);
not_4  g07267(new_n7643, new_n7644);
nand_1 g07268(new_n7484, new_n7474, new_n7645);
nand_1 g07269(new_n7645, new_n7644, new_n7646_1);
xnor_1 g07270(new_n7646_1, new_n7642, new_n7647);
nand_1 g07271(new_n7490, new_n7487, new_n7648);
nand_1 g07272(new_n7492, new_n7485, new_n7649);
nand_1 g07273(new_n7649, new_n7648, new_n7650);
nor_1  g07274(new_n7650, new_n7647, new_n7651);
not_4  g07275(new_n7651, new_n7652);
nand_1 g07276(new_n7650, new_n7647, new_n7653);
nand_1 g07277(new_n7653, new_n7652, new_n7654);
nand_1 g07278(new_n7654, new_n7627, new_n7655);
not_4  g07279(new_n7627, new_n7656);
not_4  g07280(new_n7654, new_n7657);
nand_1 g07281(new_n7657, new_n7656, new_n7658);
nand_1 g07282(new_n7658, new_n7655, new_n7659);
xnor_1 g07283(new_n7659, new_n7495, new_n7660);
xnor_1 g07284(new_n7660, new_n7626, new_n7661);
not_4  g07285(new_n7521, new_n7662);
nand_1 g07286(new_n7662, new_n7497, new_n7663);
nand_1 g07287(new_n7526, new_n7522, new_n7664);
nand_1 g07288(new_n7664, new_n7663, new_n7665);
xnor_1 g07289(new_n7665, new_n7661, new_n7666);
xnor_1 g07290(new_n7666, new_n7580, new_n7667);
not_4  g07291(new_n7667, new_n7668);
nand_1 g07292(new_n7538, new_n7434, new_n7669);
nand_1 g07293(new_n7669, new_n7540, new_n7670);
nor_1  g07294(new_n7670, new_n7668, new_n7671);
not_4  g07295(new_n7671, new_n7672);
nand_1 g07296(new_n7672, new_n7540, new_n7673);
nand_1 g07297(new_n7673, new_n7433, new_n7674);
not_4  g07298(new_n7674, new_n7675);
nor_1  g07299(new_n7673, new_n7433, new_n7676_1);
nor_1  g07300(new_n7676_1, new_n7675, new_n7677);
not_4  g07301(new_n7575, new_n7678);
nand_1 g07302(new_n7678, new_n7547, new_n7679);
nand_1 g07303(new_n7559, new_n7552, new_n7680);
not_4  g07304(new_n7560, new_n7681);
nand_1 g07305(new_n7562, new_n7681, new_n7682);
nand_1 g07306(new_n7682, new_n7680, new_n7683);
nand_1 g07307(n12221, n9400, new_n7684);
nand_1 g07308(n12145, n2464, new_n7685);
nand_1 g07309(n10217, n6877, new_n7686);
not_4  g07310(new_n7686, new_n7687);
xnor_1 g07311(new_n7687, new_n7685, new_n7688);
xnor_1 g07312(new_n7688, new_n7684, new_n7689);
xnor_1 g07313(new_n7689, new_n7683, new_n7690_1);
nand_1 g07314(n11311, n2522, new_n7691);
nand_1 g07315(new_n7691, new_n7558, new_n7692);
not_4  g07316(new_n7558, new_n7693);
not_4  g07317(new_n7691, new_n7694);
nand_1 g07318(new_n7694, new_n7693, new_n7695);
nand_1 g07319(new_n7695, new_n7692, new_n7696);
nand_1 g07320(n4203, n2024, new_n7697);
nand_1 g07321(n9189, n4187, new_n7698);
nand_1 g07322(n12753, n7946, new_n7699);
nand_1 g07323(new_n7699, new_n7698, new_n7700);
not_4  g07324(new_n7698, new_n7701);
not_4  g07325(new_n7699, new_n7702);
nand_1 g07326(new_n7702, new_n7701, new_n7703);
nand_1 g07327(new_n7703, new_n7700, new_n7704);
xnor_1 g07328(new_n7704, new_n7697, new_n7705);
not_4  g07329(new_n7705, new_n7706);
xnor_1 g07330(new_n7706, new_n7696, new_n7707);
not_4  g07331(new_n7707, new_n7708);
xnor_1 g07332(new_n7708, new_n7690_1, new_n7709);
not_4  g07333(new_n7571, new_n7710);
nor_1  g07334(new_n7710, new_n7551, new_n7711);
xnor_1 g07335(new_n7711, new_n7569, new_n7712);
nor_1  g07336(new_n7712, new_n7572, new_n7713);
xnor_1 g07337(new_n7713, new_n7709, new_n7714);
xnor_1 g07338(new_n7714, new_n7679, new_n7715);
not_4  g07339(new_n7546_1, new_n7716);
nand_1 g07340(new_n7576, new_n7716, new_n7717);
not_4  g07341(new_n7545, new_n7718);
nand_1 g07342(new_n7577, new_n7718, new_n7719);
nand_1 g07343(new_n7719, new_n7717, new_n7720);
xnor_1 g07344(new_n7720, new_n7715, new_n7721);
nand_1 g07345(n4805, n2347, new_n7722);
nand_1 g07346(n6016, n5283, new_n7723);
nand_1 g07347(n11478, n5798, new_n7724);
not_4  g07348(new_n7724, new_n7725);
xnor_1 g07349(new_n7725, new_n7723, new_n7726);
xnor_1 g07350(new_n7726, new_n7722, new_n7727);
nor_1  g07351(new_n7633, new_n7628, new_n7728);
nor_1  g07352(new_n7636, new_n7634, new_n7729);
nor_1  g07353(new_n7729, new_n7728, new_n7730_1);
xnor_1 g07354(new_n7730_1, new_n7727, new_n7731);
not_4  g07355(new_n7629, new_n7732);
nand_1 g07356(new_n7631, new_n7732, new_n7733_1);
not_4  g07357(new_n7733_1, new_n7734);
nand_1 g07358(n521, n137, new_n7735);
not_4  g07359(new_n7735, new_n7736);
nand_1 g07360(new_n7736, new_n7734, new_n7737);
nand_1 g07361(new_n7735, new_n7733_1, new_n7738);
nand_1 g07362(new_n7738, new_n7737, new_n7739);
not_4  g07363(new_n7739, new_n7740);
nand_1 g07364(n6797, n2498, new_n7741);
nand_1 g07365(n6294, n5579, new_n7742);
nand_1 g07366(n3146, n2558, new_n7743);
not_4  g07367(new_n7743, new_n7744);
xnor_1 g07368(new_n7744, new_n7742, new_n7745);
xnor_1 g07369(new_n7745, new_n7741, new_n7746);
not_4  g07370(new_n7746, new_n7747);
xnor_1 g07371(new_n7747, new_n7740, new_n7748);
xnor_1 g07372(new_n7748, new_n7731, new_n7749);
not_4  g07373(new_n7637, new_n7750);
nand_1 g07374(new_n7641, new_n7750, new_n7751);
nor_1  g07375(new_n7639, new_n7638, new_n7752);
nand_1 g07376(new_n7646_1, new_n7642, new_n7753);
not_4  g07377(new_n7753, new_n7754);
xnor_1 g07378(new_n7754, new_n7752, new_n7755);
nand_1 g07379(new_n7755, new_n7751, new_n7756);
xnor_1 g07380(new_n7756, new_n7749, new_n7757);
xnor_1 g07381(new_n7757, new_n7652, new_n7758);
not_4  g07382(new_n7758, new_n7759);
nand_1 g07383(new_n7655, new_n7494, new_n7760);
nand_1 g07384(new_n7760, new_n7658, new_n7761);
xnor_1 g07385(new_n7761, new_n7759, new_n7762);
not_4  g07386(new_n7762, new_n7763);
not_4  g07387(new_n7605, new_n7764);
nand_1 g07388(new_n7764, new_n7598, new_n7765);
nand_1 g07389(new_n7610_1, new_n7606, new_n7766);
xnor_1 g07390(new_n7766, new_n7604, new_n7767);
nand_1 g07391(new_n7767, new_n7765, new_n7768);
not_4  g07392(new_n7586, new_n7769);
nand_1 g07393(new_n7588, new_n7769, new_n7770);
not_4  g07394(new_n7770, new_n7771);
nand_1 g07395(n6358, n806, new_n7772);
not_4  g07396(new_n7772, new_n7773);
nand_1 g07397(new_n7773, new_n7771, new_n7774);
nand_1 g07398(new_n7772, new_n7770, new_n7775);
nand_1 g07399(new_n7775, new_n7774, new_n7776);
nand_1 g07400(n9111, n1471, new_n7777);
nand_1 g07401(n5198, n3342, new_n7778);
nand_1 g07402(n9763, n7646, new_n7779);
nand_1 g07403(new_n7779, new_n7778, new_n7780);
not_4  g07404(new_n7778, new_n7781);
not_4  g07405(new_n7779, new_n7782);
nand_1 g07406(new_n7782, new_n7781, new_n7783);
nand_1 g07407(new_n7783, new_n7780, new_n7784);
xnor_1 g07408(new_n7784, new_n7777, new_n7785);
not_4  g07409(new_n7785, new_n7786);
xnor_1 g07410(new_n7786, new_n7776, new_n7787);
not_4  g07411(new_n7585, new_n7788);
nand_1 g07412(new_n7589, new_n7788, new_n7789);
nand_1 g07413(new_n7595, new_n7789, new_n7790);
nand_1 g07414(n5153, n3992, new_n7791);
not_4  g07415(new_n7791, new_n7792);
nand_1 g07416(n8384, n7270, new_n7793);
nand_1 g07417(n7236, n2507, new_n7794);
not_4  g07418(new_n7794, new_n7795);
xnor_1 g07419(new_n7795, new_n7793, new_n7796);
xnor_1 g07420(new_n7796, new_n7792, new_n7797);
xnor_1 g07421(new_n7797, new_n7790, new_n7798);
xnor_1 g07422(new_n7798, new_n7787, new_n7799);
xnor_1 g07423(new_n7799, new_n7768, new_n7800);
xnor_1 g07424(new_n7800, new_n7617, new_n7801);
nand_1 g07425(new_n7621, new_n7582, new_n7802);
nand_1 g07426(new_n7802, new_n7623, new_n7803);
xnor_1 g07427(new_n7803, new_n7801, new_n7804);
not_4  g07428(new_n7804, new_n7805);
xnor_1 g07429(new_n7805, new_n7763, new_n7806);
nand_1 g07430(new_n7660, new_n7625, new_n7807);
nand_1 g07431(new_n7665, new_n7661, new_n7808);
nand_1 g07432(new_n7808, new_n7807, new_n7809);
xnor_1 g07433(new_n7809, new_n7806, new_n7810);
not_4  g07434(new_n7810, new_n7811);
xnor_1 g07435(new_n7811, new_n7721, new_n7812);
nand_1 g07436(new_n7578, new_n7543, new_n7813);
nand_1 g07437(new_n7666, new_n7580, new_n7814);
nand_1 g07438(new_n7814, new_n7813, new_n7815);
xnor_1 g07439(new_n7815, new_n7812, new_n7816);
nand_1 g07440(new_n7816, new_n7677, new_n7817);
nand_1 g07441(new_n7817, new_n7674, new_n7818);
not_4  g07442(new_n7721, new_n7819);
nand_1 g07443(new_n7811, new_n7819, new_n7820);
nand_1 g07444(new_n7815, new_n7812, new_n7821);
nand_1 g07445(new_n7821, new_n7820, new_n7822);
nand_1 g07446(n4805, n1576, new_n7823_1);
nand_1 g07447(new_n7754, new_n7752, new_n7824);
not_4  g07448(new_n7749, new_n7825);
nand_1 g07449(new_n7756, new_n7825, new_n7826);
nand_1 g07450(new_n7826, new_n7824, new_n7827);
xnor_1 g07451(new_n7827, new_n7823_1, new_n7828);
xnor_1 g07452(new_n7828, new_n7822, new_n7829);
not_4  g07453(new_n7679, new_n7830);
nand_1 g07454(new_n7714, new_n7830, new_n7831);
nand_1 g07455(new_n7720, new_n7715, new_n7832);
nand_1 g07456(new_n7832, new_n7831, new_n7833);
nand_1 g07457(new_n7800, new_n7618, new_n7834);
not_4  g07458(new_n7803, new_n7835);
nand_1 g07459(new_n7835, new_n7801, new_n7836);
nand_1 g07460(new_n7836, new_n7834, new_n7837);
not_4  g07461(new_n7689, new_n7838);
nand_1 g07462(new_n7838, new_n7683, new_n7839);
nand_1 g07463(new_n7708, new_n7690_1, new_n7840);
nand_1 g07464(new_n7840, new_n7839, new_n7841);
nand_1 g07465(n9189, n4203, new_n7842);
nand_1 g07466(n4187, n2522, new_n7843);
xnor_1 g07467(new_n7843, new_n7842, new_n7844);
nand_1 g07468(n9763, n4722, new_n7845);
nand_1 g07469(n10217, n9400, new_n7846);
xnor_1 g07470(new_n7846, new_n7845, new_n7847);
xnor_1 g07471(new_n7847, new_n7844, new_n7848);
nand_1 g07472(n9111, n7646, new_n7849);
nand_1 g07473(n12221, n2464, new_n7850);
nand_1 g07474(n12145, n11311, new_n7851);
xnor_1 g07475(new_n7851, new_n7850, new_n7852);
xnor_1 g07476(new_n7852, new_n7849, new_n7853);
xnor_1 g07477(new_n7853, new_n7848, new_n7854);
xnor_1 g07478(new_n7854, new_n7841, new_n7855);
xnor_1 g07479(new_n7855, new_n7837, new_n7856);
xnor_1 g07480(new_n7856, new_n7833, new_n7857);
not_4  g07481(new_n7569, new_n7858);
nand_1 g07482(new_n7711, new_n7858, new_n7859);
not_4  g07483(new_n7713, new_n7860);
nand_1 g07484(new_n7860, new_n7709, new_n7861);
nand_1 g07485(new_n7861, new_n7859, new_n7862_1);
nor_1  g07486(new_n7766, new_n7604, new_n7863);
not_4  g07487(new_n7768, new_n7864);
nor_1  g07488(new_n7799, new_n7864, new_n7865);
nor_1  g07489(new_n7865, new_n7863, new_n7866);
xnor_1 g07490(new_n7866, new_n7862_1, new_n7867);
nand_1 g07491(n11821, n10223, new_n7868);
nand_1 g07492(n9080, n2879, new_n7869);
xnor_1 g07493(new_n7869, new_n7868, new_n7870);
nand_1 g07494(n11757, n9195, new_n7871);
nand_1 g07495(n7862, n2512, new_n7872);
xnor_1 g07496(new_n7872, new_n7871, new_n7873);
xnor_1 g07497(new_n7873, new_n7870, new_n7874);
not_4  g07498(new_n7392, new_n7875);
nand_1 g07499(new_n7398, new_n7875, new_n7876);
nand_1 g07500(new_n7876, new_n7397, new_n7877);
xnor_1 g07501(new_n7877, new_n7874, new_n7878);
nand_1 g07502(n12753, n2024, new_n7879);
not_4  g07503(new_n7879, new_n7880);
nand_1 g07504(n3865, n1333, new_n7881);
nand_1 g07505(n5240, n4634, new_n7882);
xnor_1 g07506(new_n7882, new_n7881, new_n7883);
xnor_1 g07507(new_n7883, new_n7880, new_n7884);
xnor_1 g07508(new_n7884, new_n7878, new_n7885);
xnor_1 g07509(new_n7885, new_n7867, new_n7886);
nand_1 g07510(new_n7415, new_n7414, new_n7887);
not_4  g07511(new_n7412, new_n7888);
nand_1 g07512(new_n7417, new_n7888, new_n7889);
nand_1 g07513(new_n7889, new_n7887, new_n7890);
nand_1 g07514(new_n7400, new_n7391, new_n7891_1);
not_4  g07515(new_n7401, new_n7892);
nand_1 g07516(new_n7411, new_n7892, new_n7893);
nand_1 g07517(new_n7893, new_n7891_1, new_n7894);
not_4  g07518(new_n7696, new_n7895);
nand_1 g07519(new_n7706, new_n7895, new_n7896);
nand_1 g07520(new_n7896, new_n7695, new_n7897);
nand_1 g07521(n8384, n5153, new_n7898);
nand_1 g07522(n7270, n6358, new_n7899);
xnor_1 g07523(new_n7899, new_n7898, new_n7900);
not_4  g07524(new_n7697, new_n7901);
nand_1 g07525(new_n7700, new_n7901, new_n7902);
nand_1 g07526(new_n7902, new_n7703, new_n7903);
xnor_1 g07527(new_n7903, new_n7900, new_n7904);
xnor_1 g07528(new_n7904, new_n7897, new_n7905);
xnor_1 g07529(new_n7905, new_n7894, new_n7906);
nand_1 g07530(n5198, n806, new_n7907);
nand_1 g07531(n3992, n2507, new_n7908);
xnor_1 g07532(new_n7908, new_n7907, new_n7909);
nand_1 g07533(n7823, n6877, new_n7910);
nand_1 g07534(n3342, n1471, new_n7911);
xnor_1 g07535(new_n7911, new_n7910, new_n7912);
xnor_1 g07536(new_n7912, new_n7909, new_n7913);
not_4  g07537(new_n7777, new_n7914);
nand_1 g07538(new_n7780, new_n7914, new_n7915);
nand_1 g07539(new_n7915, new_n7783, new_n7916);
xnor_1 g07540(new_n7916, new_n7913, new_n7917);
xnor_1 g07541(new_n7917, new_n7906, new_n7918);
not_4  g07542(new_n7790, new_n7919);
nand_1 g07543(new_n7797, new_n7919, new_n7920);
not_4  g07544(new_n7787, new_n7921);
nand_1 g07545(new_n7798, new_n7921, new_n7922);
nand_1 g07546(new_n7922, new_n7920, new_n7923);
nand_1 g07547(new_n7686, new_n7685, new_n7924);
nand_1 g07548(new_n7688, new_n7684, new_n7925);
nand_1 g07549(new_n7925, new_n7924, new_n7926);
nand_1 g07550(n7236, n6431, new_n7927);
nand_1 g07551(n10174, n7946, new_n7928);
not_4  g07552(new_n7928, new_n7929);
xnor_1 g07553(new_n7929, new_n7927, new_n7930);
xnor_1 g07554(new_n7930, new_n7926, new_n7931);
xnor_1 g07555(new_n7931, new_n7923, new_n7932);
xnor_1 g07556(new_n7932, new_n7918, new_n7933);
xnor_1 g07557(new_n7933, new_n7890, new_n7934);
xnor_1 g07558(new_n7934, new_n7886, new_n7935);
xnor_1 g07559(new_n7935, new_n7857, new_n7936);
nand_1 g07560(new_n7805, new_n7763, new_n7937);
not_4  g07561(new_n7806, new_n7938);
nand_1 g07562(new_n7809, new_n7938, new_n7939);
nand_1 g07563(new_n7939, new_n7937, new_n7940);
not_4  g07564(new_n7387, new_n7941);
nand_1 g07565(new_n7418, new_n7941, new_n7942);
nand_1 g07566(new_n7432, new_n7419, new_n7943);
nand_1 g07567(new_n7943, new_n7942, new_n7944);
nand_1 g07568(new_n7757, new_n7651, new_n7945);
nand_1 g07569(new_n7761, new_n7758, new_n7946_1);
nand_1 g07570(new_n7946_1, new_n7945, new_n7947);
not_4  g07571(new_n7776, new_n7948);
nand_1 g07572(new_n7786, new_n7948, new_n7949);
nand_1 g07573(new_n7949, new_n7774, new_n7950);
nand_1 g07574(new_n7746, new_n7740, new_n7951);
nand_1 g07575(new_n7951, new_n7737, new_n7952);
xnor_1 g07576(new_n7952, new_n7950, new_n7953);
nand_1 g07577(new_n7402, new_n7367, new_n7954);
not_4  g07578(new_n7403, new_n7955);
nand_1 g07579(new_n7410, new_n7955, new_n7956);
nand_1 g07580(new_n7956, new_n7954, new_n7957);
nand_1 g07581(n3172, n2253, new_n7958);
nand_1 g07582(n6797, n5579, new_n7959);
nand_1 g07583(n5798, n5283, new_n7960);
xnor_1 g07584(new_n7960, new_n7959, new_n7961);
xnor_1 g07585(new_n7961, new_n7958, new_n7962);
xnor_1 g07586(new_n7962, new_n7957, new_n7963);
nand_1 g07587(new_n7724, new_n7723, new_n7964);
nand_1 g07588(new_n7726, new_n7722, new_n7965_1);
nand_1 g07589(new_n7965_1, new_n7964, new_n7966_1);
nand_1 g07590(new_n7743, new_n7742, new_n7967);
nand_1 g07591(new_n7745, new_n7741, new_n7968);
nand_1 g07592(new_n7968, new_n7967, new_n7969);
xnor_1 g07593(new_n7969, new_n7966_1, new_n7970);
nand_1 g07594(n11478, n2347, new_n7971);
nand_1 g07595(n3146, n2498, new_n7972);
xnor_1 g07596(new_n7972, new_n7971, new_n7973);
xnor_1 g07597(new_n7973, new_n7970, new_n7974);
xnor_1 g07598(new_n7974, new_n7963, new_n7975);
xnor_1 g07599(new_n7975, new_n7953, new_n7976);
not_4  g07600(new_n7727, new_n7977);
nand_1 g07601(new_n7730_1, new_n7977, new_n7978);
not_4  g07602(new_n7748, new_n7979);
nand_1 g07603(new_n7979, new_n7731, new_n7980);
nand_1 g07604(new_n7980, new_n7978, new_n7981_1);
nand_1 g07605(new_n7407, new_n7406, new_n7982);
nand_1 g07606(new_n7409, new_n7404, new_n7983);
nand_1 g07607(new_n7983, new_n7982, new_n7984);
nand_1 g07608(n6016, n137, new_n7985);
not_4  g07609(new_n7985, new_n7986);
nand_1 g07610(n7265, n6826, new_n7987);
nand_1 g07611(n6294, n521, new_n7988);
xnor_1 g07612(new_n7988, new_n7987, new_n7989);
xnor_1 g07613(new_n7989, new_n7986, new_n7990);
xnor_1 g07614(new_n7990, new_n7984, new_n7991);
nand_1 g07615(n4938, n2558, new_n7992);
nand_1 g07616(new_n7794, new_n7793, new_n7993);
nand_1 g07617(new_n7796, new_n7791, new_n7994);
nand_1 g07618(new_n7994, new_n7993, new_n7995);
xnor_1 g07619(new_n7995, new_n7992, new_n7996);
xnor_1 g07620(new_n7996, new_n7991, new_n7997);
xnor_1 g07621(new_n7997, new_n7981_1, new_n7998);
xnor_1 g07622(new_n7998, new_n7976, new_n7999);
xnor_1 g07623(new_n7999, new_n7947, new_n8000);
xnor_1 g07624(new_n8000, new_n7944, new_n8001);
xnor_1 g07625(new_n8001, new_n7940, new_n8002);
xnor_1 g07626(new_n8002, new_n7936, new_n8003);
xnor_1 g07627(new_n8003, new_n7829, new_n8004);
xnor_1 g07628(new_n8004, new_n7818, n2383);
nand_1 g07629(new_n6569, new_n6559, new_n8006);
nand_1 g07630(new_n8006, new_n6571, n2425);
xnor_1 g07631(new_n3175, new_n3122, n2431);
xnor_1 g07632(new_n2283, new_n2282, n2434);
nand_1 g07633(new_n5475, new_n5474, new_n8010);
nand_1 g07634(new_n8010, new_n5477, n2581);
nand_1 g07635(new_n7322, new_n7320_1, new_n8012);
xnor_1 g07636(new_n8012, new_n7333, n2624);
nand_1 g07637(n11917, n6770, new_n8014);
not_4  g07638(new_n8014, new_n8015);
nand_1 g07639(n9920, n4921, new_n8016);
nand_1 g07640(n9956, n3627, new_n8017);
not_4  g07641(new_n8017, new_n8018);
xnor_1 g07642(new_n8018, new_n8016, new_n8019);
nor_1  g07643(new_n8019, new_n8015, new_n8020);
not_4  g07644(new_n8020, new_n8021);
nand_1 g07645(new_n8019, new_n8015, new_n8022);
nand_1 g07646(new_n8022, new_n8021, new_n8023);
nand_1 g07647(new_n4344, new_n4302, new_n8024);
nand_1 g07648(new_n4345, new_n4343, new_n8025);
nand_1 g07649(new_n8025, new_n8024, new_n8026);
xnor_1 g07650(new_n8026, new_n8023, new_n8027);
nand_1 g07651(n2577, n2564, new_n8028_1);
nand_1 g07652(n4189, n3842, new_n8029);
not_4  g07653(new_n8029, new_n8030);
xnor_1 g07654(new_n8030, new_n8028_1, new_n8031);
xnor_1 g07655(new_n8031, new_n8027, new_n8032);
not_4  g07656(new_n4342, new_n8033);
nand_1 g07657(new_n4346, new_n8033, new_n8034);
nand_1 g07658(new_n8034, new_n4340, new_n8035);
xnor_1 g07659(new_n8035, new_n8032, new_n8036);
not_4  g07660(new_n8036, new_n8037);
not_4  g07661(new_n4331, new_n8038);
nand_1 g07662(new_n4334, new_n8038, new_n8039);
nand_1 g07663(new_n4347, new_n4335, new_n8040);
nand_1 g07664(new_n8040, new_n8039, new_n8041);
nand_1 g07665(new_n8041, new_n8037, new_n8042);
not_4  g07666(new_n8016, new_n8043);
nand_1 g07667(new_n8018, new_n8043, new_n8044);
nand_1 g07668(n6770, n3842, new_n8045);
not_4  g07669(new_n8045, new_n8046);
xnor_1 g07670(new_n8046, new_n8044, new_n8047);
not_4  g07671(new_n8047, new_n8048);
nand_1 g07672(n4921, n3627, new_n8049);
nand_1 g07673(n11917, n9920, new_n8050);
nand_1 g07674(n9956, n4516, new_n8051);
not_4  g07675(new_n8051, new_n8052);
xnor_1 g07676(new_n8052, new_n8050, new_n8053);
xnor_1 g07677(new_n8053, new_n8049, new_n8054);
not_4  g07678(new_n8054, new_n8055);
xnor_1 g07679(new_n8055, new_n8048, new_n8056);
not_4  g07680(new_n8023, new_n8057);
nand_1 g07681(new_n8026, new_n8057, new_n8058);
nand_1 g07682(new_n8058, new_n8021, new_n8059);
nand_1 g07683(n9637, n2564, new_n8060);
nand_1 g07684(n4189, n2577, new_n8061);
nand_1 g07685(n6687, n1835, new_n8062);
not_4  g07686(new_n8062, new_n8063);
xnor_1 g07687(new_n8063, new_n8061, new_n8064);
xnor_1 g07688(new_n8064, new_n8060, new_n8065_1);
xnor_1 g07689(new_n8065_1, new_n8059, new_n8066);
xnor_1 g07690(new_n8066, new_n8056, new_n8067);
not_4  g07691(new_n8067, new_n8068);
not_4  g07692(new_n8027, new_n8069);
nand_1 g07693(new_n8031, new_n8069, new_n8070);
nor_1  g07694(new_n8029, new_n8028_1, new_n8071);
nand_1 g07695(new_n8035, new_n8032, new_n8072);
not_4  g07696(new_n8072, new_n8073);
xnor_1 g07697(new_n8073, new_n8071, new_n8074);
nand_1 g07698(new_n8074, new_n8070, new_n8075);
xnor_1 g07699(new_n8075, new_n8068, new_n8076);
xnor_1 g07700(new_n8076, new_n8042, new_n8077);
nand_1 g07701(n9637, n6687, new_n8078);
not_4  g07702(new_n8078, new_n8079);
xnor_1 g07703(new_n8041, new_n8036, new_n8080);
nand_1 g07704(new_n8080, new_n8079, new_n8081);
not_4  g07705(new_n4330, new_n8082);
nand_1 g07706(new_n4349, new_n8082, new_n8083);
not_4  g07707(new_n8083, new_n8084);
xnor_1 g07708(new_n8080, new_n8078, new_n8085);
nand_1 g07709(new_n8085, new_n8084, new_n8086);
nand_1 g07710(new_n8086, new_n8081, new_n8087);
xnor_1 g07711(new_n8087, new_n8077, new_n8088);
nand_1 g07712(n6126, n2226, new_n8089);
nand_1 g07713(n3602, n1094, new_n8090);
nand_1 g07714(n10678, n3719, new_n8091);
not_4  g07715(new_n8091, new_n8092);
xnor_1 g07716(new_n8092, new_n8090, new_n8093);
not_4  g07717(new_n8093, new_n8094);
xnor_1 g07718(new_n8094, new_n8089, new_n8095);
nand_1 g07719(new_n4565, new_n4360, new_n8096);
nand_1 g07720(new_n4566, new_n4564, new_n8097);
nand_1 g07721(new_n8097, new_n8096, new_n8098);
xnor_1 g07722(new_n8098, new_n8095, new_n8099);
not_4  g07723(new_n8099, new_n8100_1);
nand_1 g07724(n10928, n10439, new_n8101);
nand_1 g07725(n8595, n6986, new_n8102);
nand_1 g07726(new_n8102, new_n8101, new_n8103);
not_4  g07727(new_n8101, new_n8104);
not_4  g07728(new_n8102, new_n8105);
nand_1 g07729(new_n8105, new_n8104, new_n8106);
nand_1 g07730(new_n8106, new_n8103, new_n8107);
xnor_1 g07731(new_n8107, new_n8100_1, new_n8108);
not_4  g07732(new_n4563, new_n8109);
nand_1 g07733(new_n4567, new_n8109, new_n8110);
nand_1 g07734(new_n8110, new_n4561, new_n8111);
xnor_1 g07735(new_n8111, new_n8108, new_n8112);
not_4  g07736(new_n8112, new_n8113);
nor_1  g07737(new_n4554, new_n4552, new_n8114);
not_4  g07738(new_n8114, new_n8115);
nand_1 g07739(new_n4568, new_n4556, new_n8116);
nand_1 g07740(new_n8116, new_n8115, new_n8117);
nand_1 g07741(new_n8117, new_n8113, new_n8118);
nand_1 g07742(new_n8094, new_n8089, new_n8119);
not_4  g07743(new_n8095, new_n8120);
nand_1 g07744(new_n8098, new_n8120, new_n8121);
nand_1 g07745(new_n8121, new_n8119, new_n8122);
nand_1 g07746(n10928, n8065, new_n8123);
nand_1 g07747(n10439, n6986, new_n8124);
nand_1 g07748(n10391, n8336, new_n8125);
not_4  g07749(new_n8125, new_n8126);
xnor_1 g07750(new_n8126, new_n8124, new_n8127);
xnor_1 g07751(new_n8127, new_n8123, new_n8128);
xnor_1 g07752(new_n8128, new_n8122, new_n8129);
not_4  g07753(new_n8090, new_n8130);
nand_1 g07754(new_n8092, new_n8130, new_n8131);
nand_1 g07755(n8595, n2226, new_n8132);
nand_1 g07756(new_n8132, new_n8131, new_n8133);
not_4  g07757(new_n8131, new_n8134);
not_4  g07758(new_n8132, new_n8135);
nand_1 g07759(new_n8135, new_n8134, new_n8136);
nand_1 g07760(new_n8136, new_n8133, new_n8137);
not_4  g07761(new_n8137, new_n8138_1);
nand_1 g07762(n10678, n3602, new_n8139);
nand_1 g07763(n6126, n1094, new_n8140);
nand_1 g07764(n7320, n3719, new_n8141);
not_4  g07765(new_n8141, new_n8142);
xnor_1 g07766(new_n8142, new_n8140, new_n8143);
xnor_1 g07767(new_n8143, new_n8139, new_n8144);
not_4  g07768(new_n8144, new_n8145);
xnor_1 g07769(new_n8145, new_n8138_1, new_n8146);
xnor_1 g07770(new_n8146, new_n8129, new_n8147);
not_4  g07771(new_n8147, new_n8148);
not_4  g07772(new_n8107, new_n8149);
nand_1 g07773(new_n8149, new_n8100_1, new_n8150);
not_4  g07774(new_n8150, new_n8151);
nand_1 g07775(new_n8111, new_n8108, new_n8152);
not_4  g07776(new_n8152, new_n8153);
xnor_1 g07777(new_n8153, new_n8106, new_n8154);
nor_1  g07778(new_n8154, new_n8151, new_n8155);
xnor_1 g07779(new_n8155, new_n8148, new_n8156);
not_4  g07780(new_n8156, new_n8157);
xnor_1 g07781(new_n8157, new_n8118, new_n8158);
nand_1 g07782(n8336, n8065, new_n8159);
not_4  g07783(new_n8159, new_n8160);
xnor_1 g07784(new_n8117, new_n8112, new_n8161);
nor_1  g07785(new_n8161, new_n8160, new_n8162);
not_4  g07786(new_n8162, new_n8163);
not_4  g07787(new_n4390, new_n8164);
nand_1 g07788(new_n4570, new_n8164, new_n8165);
nand_1 g07789(new_n8161, new_n8160, new_n8166);
nand_1 g07790(new_n8166, new_n8163, new_n8167);
not_4  g07791(new_n8167, new_n8168);
nand_1 g07792(new_n8168, new_n8165, new_n8169);
nand_1 g07793(new_n8169, new_n8163, new_n8170);
xnor_1 g07794(new_n8170, new_n8158, new_n8171);
nand_1 g07795(n7160, n4826, new_n8172);
not_4  g07796(new_n8172, new_n8173);
nand_1 g07797(n7733, n4828, new_n8174);
nand_1 g07798(n12925, n2515, new_n8175);
not_4  g07799(new_n8175, new_n8176);
xnor_1 g07800(new_n8176, new_n8174, new_n8177);
xnor_1 g07801(new_n8177, new_n8173, new_n8178);
nand_1 g07802(new_n4605, new_n4398, new_n8179);
nand_1 g07803(new_n4606, new_n4604, new_n8180);
nand_1 g07804(new_n8180, new_n8179, new_n8181);
nor_1  g07805(new_n8181, new_n8178, new_n8182);
not_4  g07806(new_n8182, new_n8183);
nand_1 g07807(new_n8181, new_n8178, new_n8184);
nand_1 g07808(new_n8184, new_n8183, new_n8185);
nand_1 g07809(n12391, n4970, new_n8186);
nand_1 g07810(n7891, n7610, new_n8187);
not_4  g07811(new_n8187, new_n8188);
xnor_1 g07812(new_n8188, new_n8186, new_n8189);
xnor_1 g07813(new_n8189, new_n8185, new_n8190);
nor_1  g07814(new_n4601, new_n4599, new_n8191);
not_4  g07815(new_n4603, new_n8192);
nor_1  g07816(new_n4608, new_n8192, new_n8193);
nor_1  g07817(new_n8193, new_n8191, new_n8194);
xnor_1 g07818(new_n8194, new_n8190, new_n8195);
not_4  g07819(new_n4598, new_n8196);
nand_1 g07820(new_n4609, new_n8196, new_n8197);
not_4  g07821(new_n4613, new_n8198);
nand_1 g07822(new_n8198, new_n4610, new_n8199);
nand_1 g07823(new_n8199, new_n8197, new_n8200);
nand_1 g07824(new_n8200, new_n8195, new_n8201);
nand_1 g07825(new_n8177, new_n8173, new_n8202_1);
nand_1 g07826(new_n8183, new_n8202_1, new_n8203);
nand_1 g07827(n12391, n503, new_n8204);
nand_1 g07828(n7891, n4970, new_n8205);
nand_1 g07829(n12069, n10965, new_n8206);
not_4  g07830(new_n8206, new_n8207);
xnor_1 g07831(new_n8207, new_n8205, new_n8208);
xnor_1 g07832(new_n8208, new_n8204, new_n8209);
not_4  g07833(new_n8209, new_n8210);
xnor_1 g07834(new_n8210, new_n8203, new_n8211);
not_4  g07835(new_n8174, new_n8212);
nand_1 g07836(new_n8176, new_n8212, new_n8213);
not_4  g07837(new_n8213, new_n8214);
nand_1 g07838(n7610, n7160, new_n8215);
not_4  g07839(new_n8215, new_n8216);
nand_1 g07840(new_n8216, new_n8214, new_n8217);
nand_1 g07841(new_n8215, new_n8213, new_n8218);
nand_1 g07842(new_n8218, new_n8217, new_n8219);
nand_1 g07843(n7733, n2515, new_n8220);
nand_1 g07844(n4828, n4826, new_n8221);
nand_1 g07845(n12925, n1199, new_n8222);
not_4  g07846(new_n8222, new_n8223);
xnor_1 g07847(new_n8223, new_n8221, new_n8224);
xnor_1 g07848(new_n8224, new_n8220, new_n8225);
xnor_1 g07849(new_n8225, new_n8219, new_n8226);
xnor_1 g07850(new_n8226, new_n8211, new_n8227);
not_4  g07851(new_n8185, new_n8228);
nand_1 g07852(new_n8189, new_n8228, new_n8229);
nor_1  g07853(new_n8187, new_n8186, new_n8230);
not_4  g07854(new_n8194, new_n8231);
nand_1 g07855(new_n8231, new_n8190, new_n8232);
not_4  g07856(new_n8232, new_n8233);
xnor_1 g07857(new_n8233, new_n8230, new_n8234);
nand_1 g07858(new_n8234, new_n8229, new_n8235);
xnor_1 g07859(new_n8235, new_n8227, new_n8236_1);
xnor_1 g07860(new_n8236_1, new_n8201, new_n8237);
nand_1 g07861(n12069, n503, new_n8238);
not_4  g07862(new_n8238, new_n8239);
not_4  g07863(new_n8201, new_n8240);
nor_1  g07864(new_n8200, new_n8195, new_n8241);
nor_1  g07865(new_n8241, new_n8240, new_n8242);
nand_1 g07866(new_n8242, new_n8239, new_n8243);
nand_1 g07867(new_n4614, new_n4426, new_n8244);
xnor_1 g07868(new_n8242, new_n8238, new_n8245);
not_4  g07869(new_n8245, new_n8246);
nor_1  g07870(new_n8246, new_n8244, new_n8247);
not_4  g07871(new_n8247, new_n8248);
nand_1 g07872(new_n8248, new_n8243, new_n8249);
not_4  g07873(new_n8249, new_n8250);
xnor_1 g07874(new_n8250, new_n8237, new_n8251);
not_4  g07875(new_n8251, new_n8252);
nand_1 g07876(n11222, n6359, new_n8253);
not_4  g07877(new_n8253, new_n8254);
nand_1 g07878(n4086, n996, new_n8255);
not_4  g07879(new_n8255, new_n8256);
nand_1 g07880(n5767, n405, new_n8257);
nand_1 g07881(n8433, n5319, new_n8258);
not_4  g07882(new_n8258, new_n8259);
xnor_1 g07883(new_n8259, new_n8257, new_n8260);
xnor_1 g07884(new_n8260, new_n8256, new_n8261);
nand_1 g07885(new_n4584, new_n4577, new_n8262);
nand_1 g07886(new_n8262, new_n4581, new_n8263);
nor_1  g07887(new_n8263, new_n8261, new_n8264);
not_4  g07888(new_n8264, new_n8265);
nand_1 g07889(new_n8263, new_n8261, new_n8266);
nand_1 g07890(new_n8266, new_n8265, new_n8267);
nand_1 g07891(n11153, n6611, new_n8268);
nand_1 g07892(n5314, n217, new_n8269);
nand_1 g07893(new_n8269, new_n8268, new_n8270);
not_4  g07894(new_n8268, new_n8271);
not_4  g07895(new_n8269, new_n8272);
nand_1 g07896(new_n8272, new_n8271, new_n8273);
nand_1 g07897(new_n8273, new_n8270, new_n8274);
not_4  g07898(new_n8274, new_n8275);
xnor_1 g07899(new_n8275, new_n8267, new_n8276_1);
not_4  g07900(new_n4576, new_n8277);
nand_1 g07901(new_n4586, new_n8277, new_n8278);
not_4  g07902(new_n4589, new_n8279);
nand_1 g07903(new_n8279, new_n4587, new_n8280);
nand_1 g07904(new_n8280, new_n8278, new_n8281);
xnor_1 g07905(new_n8281, new_n8276_1, new_n8282);
not_4  g07906(new_n4575, new_n8283);
nand_1 g07907(new_n4590, new_n8283, new_n8284);
nand_1 g07908(new_n4595, new_n4591, new_n8285);
nand_1 g07909(new_n8285, new_n8284, new_n8286);
xnor_1 g07910(new_n8286, new_n8282, new_n8287);
nand_1 g07911(new_n8287, new_n8254, new_n8288);
not_4  g07912(new_n8288, new_n8289);
nand_1 g07913(new_n4596, new_n4574, new_n8290);
not_4  g07914(new_n8282, new_n8291);
xnor_1 g07915(new_n8286, new_n8291, new_n8292);
nand_1 g07916(new_n8292, new_n8253, new_n8293);
nand_1 g07917(new_n8293, new_n8288, new_n8294);
nor_1  g07918(new_n8294, new_n8290, new_n8295);
nor_1  g07919(new_n8295, new_n8289, new_n8296);
nand_1 g07920(new_n8286, new_n8291, new_n8297);
not_4  g07921(new_n8257, new_n8298);
nand_1 g07922(new_n8259, new_n8298, new_n8299);
not_4  g07923(new_n8299, new_n8300);
nand_1 g07924(n996, n217, new_n8301);
not_4  g07925(new_n8301, new_n8302);
nand_1 g07926(new_n8302, new_n8300, new_n8303_1);
nand_1 g07927(new_n8301, new_n8299, new_n8304);
nand_1 g07928(new_n8304, new_n8303_1, new_n8305);
not_4  g07929(new_n8305, new_n8306);
nand_1 g07930(n5319, n405, new_n8307);
nand_1 g07931(n5767, n4086, new_n8308);
nand_1 g07932(n9457, n8433, new_n8309);
not_4  g07933(new_n8309, new_n8310);
xnor_1 g07934(new_n8310, new_n8308, new_n8311);
not_4  g07935(new_n8311, new_n8312);
xnor_1 g07936(new_n8312, new_n8307, new_n8313);
not_4  g07937(new_n8313, new_n8314);
nand_1 g07938(new_n8314, new_n8306, new_n8315);
nand_1 g07939(new_n8313, new_n8305, new_n8316);
nand_1 g07940(new_n8316, new_n8315, new_n8317);
nand_1 g07941(n11153, n6359, new_n8318);
nand_1 g07942(n6611, n5314, new_n8319);
not_4  g07943(new_n8319, new_n8320);
nand_1 g07944(n11296, n11222, new_n8321);
xnor_1 g07945(new_n8321, new_n8320, new_n8322);
xnor_1 g07946(new_n8322, new_n8318, new_n8323);
not_4  g07947(new_n8323, new_n8324);
nand_1 g07948(new_n8260, new_n8256, new_n8325);
nand_1 g07949(new_n8265, new_n8325, new_n8326);
xnor_1 g07950(new_n8326, new_n8324, new_n8327);
xnor_1 g07951(new_n8327, new_n8317, new_n8328);
not_4  g07952(new_n8267, new_n8329);
nand_1 g07953(new_n8275, new_n8329, new_n8330);
nand_1 g07954(new_n8281, new_n8276_1, new_n8331);
nor_1  g07955(new_n8331, new_n8273, new_n8332);
not_4  g07956(new_n8332, new_n8333);
nand_1 g07957(new_n8331, new_n8273, new_n8334);
nand_1 g07958(new_n8334, new_n8333, new_n8335);
nand_1 g07959(new_n8335, new_n8330, new_n8336_1);
nand_1 g07960(new_n8336_1, new_n8328, new_n8337);
not_4  g07961(new_n8337, new_n8338);
nor_1  g07962(new_n8336_1, new_n8328, new_n8339);
nor_1  g07963(new_n8339, new_n8338, new_n8340);
xnor_1 g07964(new_n8340, new_n8297, new_n8341);
not_4  g07965(new_n8341, new_n8342);
xnor_1 g07966(new_n8342, new_n8296, new_n8343);
nand_1 g07967(new_n8343, new_n8252, new_n8344);
xnor_1 g07968(new_n8341, new_n8296, new_n8345);
nand_1 g07969(new_n8345, new_n8251, new_n8346);
nand_1 g07970(new_n8346, new_n8344, new_n8347);
xnor_1 g07971(new_n8245, new_n8244, new_n8348);
not_4  g07972(new_n8290, new_n8349);
xnor_1 g07973(new_n8294, new_n8349, new_n8350);
nor_1  g07974(new_n8350, new_n8348, new_n8351);
not_4  g07975(new_n4615, new_n8352);
nand_1 g07976(new_n4619, new_n8352, new_n8353);
nand_1 g07977(new_n4620, new_n4597, new_n8354);
nand_1 g07978(new_n8354, new_n8353, new_n8355);
not_4  g07979(new_n8355, new_n8356);
not_4  g07980(new_n8348, new_n8357);
xnor_1 g07981(new_n8294, new_n8290, new_n8358);
nand_1 g07982(new_n8358, new_n8357, new_n8359);
nand_1 g07983(new_n8350, new_n8348, new_n8360);
nand_1 g07984(new_n8360, new_n8359, new_n8361);
nor_1  g07985(new_n8361, new_n8356, new_n8362);
nor_1  g07986(new_n8362, new_n8351, new_n8363);
nor_1  g07987(new_n8363, new_n8347, new_n8364);
nor_1  g07988(new_n8345, new_n8251, new_n8365);
nor_1  g07989(new_n8343, new_n8252, new_n8366);
nor_1  g07990(new_n8366, new_n8365, new_n8367);
nor_1  g07991(new_n8358, new_n8357, new_n8368);
nor_1  g07992(new_n8368, new_n8351, new_n8369);
nand_1 g07993(new_n8369, new_n8355, new_n8370);
nand_1 g07994(new_n8370, new_n8359, new_n8371);
nor_1  g07995(new_n8371, new_n8367, new_n8372);
nor_1  g07996(new_n8372, new_n8364, new_n8373);
nand_1 g07997(new_n8373, new_n8171, new_n8374);
not_4  g07998(new_n8171, new_n8375);
nand_1 g07999(new_n8371, new_n8367, new_n8376);
nand_1 g08000(new_n8363, new_n8347, new_n8377);
nand_1 g08001(new_n8377, new_n8376, new_n8378);
nand_1 g08002(new_n8378, new_n8375, new_n8379);
nand_1 g08003(new_n8379, new_n8374, new_n8380);
not_4  g08004(new_n8165, new_n8381);
nand_1 g08005(new_n8167, new_n8381, new_n8382);
nand_1 g08006(new_n8382, new_n8169, new_n8383);
nand_1 g08007(new_n8361, new_n8356, new_n8384_1);
nand_1 g08008(new_n8384_1, new_n8370, new_n8385);
nor_1  g08009(new_n8385, new_n8383, new_n8386);
not_4  g08010(new_n8383, new_n8387);
nor_1  g08011(new_n8369, new_n8355, new_n8388);
nor_1  g08012(new_n8388, new_n8362, new_n8389);
nand_1 g08013(new_n8389, new_n8387, new_n8390);
nand_1 g08014(new_n8385, new_n8383, new_n8391);
nand_1 g08015(new_n8391, new_n8390, new_n8392);
not_4  g08016(new_n4626, new_n8393);
nand_1 g08017(new_n4629, new_n8393, new_n8394);
nand_1 g08018(new_n8394, new_n4624, new_n8395);
nor_1  g08019(new_n8395, new_n8392, new_n8396);
nor_1  g08020(new_n8396, new_n8386, new_n8397);
nor_1  g08021(new_n8397, new_n8380, new_n8398_1);
nor_1  g08022(new_n8378, new_n8375, new_n8399);
nor_1  g08023(new_n8373, new_n8171, new_n8400);
nor_1  g08024(new_n8400, new_n8399, new_n8401);
nor_1  g08025(new_n8389, new_n8387, new_n8402);
nor_1  g08026(new_n8402, new_n8386, new_n8403);
not_4  g08027(new_n8395, new_n8404);
nand_1 g08028(new_n8404, new_n8403, new_n8405);
nand_1 g08029(new_n8405, new_n8390, new_n8406);
nor_1  g08030(new_n8406, new_n8401, new_n8407);
nor_1  g08031(new_n8407, new_n8398_1, new_n8408);
nor_1  g08032(new_n8408, new_n8088, new_n8409);
xnor_1 g08033(new_n8085, new_n8083, new_n8410);
not_4  g08034(new_n4551, new_n8411);
nand_1 g08035(new_n4630, new_n8411, new_n8412);
nand_1 g08036(new_n8412, new_n4550, new_n8413);
nor_1  g08037(new_n8413, new_n8410, new_n8414);
not_4  g08038(new_n8414, new_n8415);
nand_1 g08039(new_n8395, new_n8392, new_n8416);
nand_1 g08040(new_n8416, new_n8405, new_n8417);
nand_1 g08041(new_n8413, new_n8410, new_n8418);
nand_1 g08042(new_n8418, new_n8415, new_n8419);
nor_1  g08043(new_n8419, new_n8417, new_n8420);
not_4  g08044(new_n8420, new_n8421);
nand_1 g08045(new_n8421, new_n8415, new_n8422);
not_4  g08046(new_n8088, new_n8423);
nand_1 g08047(new_n8406, new_n8401, new_n8424);
nand_1 g08048(new_n8397, new_n8380, new_n8425);
nand_1 g08049(new_n8425, new_n8424, new_n8426);
nand_1 g08050(new_n8426, new_n8423, new_n8427);
nand_1 g08051(new_n8408, new_n8088, new_n8428);
nand_1 g08052(new_n8428, new_n8427, new_n8429);
nor_1  g08053(new_n8429, new_n8422, new_n8430);
nor_1  g08054(new_n8430, new_n8409, new_n8431);
nand_1 g08055(new_n8233, new_n8230, new_n8432);
not_4  g08056(new_n8227, new_n8433_1);
nand_1 g08057(new_n8235, new_n8433_1, new_n8434);
nand_1 g08058(new_n8434, new_n8432, new_n8435);
not_4  g08059(new_n8219, new_n8436);
nand_1 g08060(new_n8225, new_n8436, new_n8437);
nand_1 g08061(new_n8437, new_n8217, new_n8438);
nand_1 g08062(new_n8062, new_n8061, new_n8439);
nand_1 g08063(new_n8064, new_n8060, new_n8440);
nand_1 g08064(new_n8440, new_n8439, new_n8441);
nand_1 g08065(n6770, n2577, new_n8442);
xnor_1 g08066(new_n8442, new_n8441, new_n8443);
nand_1 g08067(n9637, n4189, new_n8444);
nand_1 g08068(n11917, n3627, new_n8445);
xnor_1 g08069(new_n8445, new_n8444, new_n8446);
xnor_1 g08070(new_n8446, new_n8443, new_n8447);
not_4  g08071(new_n8447, new_n8448);
nand_1 g08072(new_n8206, new_n8205, new_n8449);
nand_1 g08073(new_n8208, new_n8204, new_n8450);
nand_1 g08074(new_n8450, new_n8449, new_n8451);
nand_1 g08075(new_n8045, new_n8044, new_n8452);
nand_1 g08076(new_n8055, new_n8047, new_n8453);
nand_1 g08077(new_n8453, new_n8452, new_n8454);
xnor_1 g08078(new_n8454, new_n8451, new_n8455);
xnor_1 g08079(new_n8455, new_n8448, new_n8456);
xnor_1 g08080(new_n8456, new_n8438, new_n8457);
nor_1  g08081(new_n8209, new_n8203, new_n8458);
not_4  g08082(new_n8211, new_n8459);
nor_1  g08083(new_n8226, new_n8459, new_n8460);
nor_1  g08084(new_n8460, new_n8458, new_n8461);
nand_1 g08085(new_n8141, new_n8140, new_n8462);
nand_1 g08086(new_n8143, new_n8139, new_n8463);
nand_1 g08087(new_n8463, new_n8462, new_n8464);
nand_1 g08088(n7523, n3719, new_n8465);
nand_1 g08089(n11222, n1357, new_n8466);
xnor_1 g08090(new_n8466, new_n8465, new_n8467);
nand_1 g08091(n8336, n4190, new_n8468);
nand_1 g08092(n7320, n3602, new_n8469);
xnor_1 g08093(new_n8469, new_n8468, new_n8470);
xnor_1 g08094(new_n8470, new_n8467, new_n8471);
xnor_1 g08095(new_n8471, new_n8464, new_n8472);
xnor_1 g08096(new_n8472, new_n8461, new_n8473);
xnor_1 g08097(new_n8473, new_n8457, new_n8474);
nand_1 g08098(new_n8073, new_n8071, new_n8475);
nand_1 g08099(new_n8075, new_n8067, new_n8476_1);
nand_1 g08100(new_n8476_1, new_n8475, new_n8477);
nor_1  g08101(new_n8152, new_n8106, new_n8478);
nor_1  g08102(new_n8155, new_n8147, new_n8479);
nor_1  g08103(new_n8479, new_n8478, new_n8480);
xnor_1 g08104(new_n8480, new_n8477, new_n8481);
xnor_1 g08105(new_n8481, new_n8474, new_n8482);
xnor_1 g08106(new_n8482, new_n8435, new_n8483);
nor_1  g08107(new_n8157, new_n8118, new_n8484);
nor_1  g08108(new_n8170, new_n8158, new_n8485);
nor_1  g08109(new_n8485, new_n8484, new_n8486);
nand_1 g08110(new_n8125, new_n8124, new_n8487);
nand_1 g08111(new_n8127, new_n8123, new_n8488);
nand_1 g08112(new_n8488, new_n8487, new_n8489);
nand_1 g08113(n5319, n4086, new_n8490);
nand_1 g08114(n10928, n10391, new_n8491);
xnor_1 g08115(new_n8491, new_n8490, new_n8492);
xnor_1 g08116(new_n8492, new_n8489, new_n8493);
xnor_1 g08117(new_n8493, new_n8486, new_n8494);
xnor_1 g08118(new_n8494, new_n8483, new_n8495);
nand_1 g08119(new_n8236_1, new_n8240, new_n8496);
nand_1 g08120(new_n8249, new_n8237, new_n8497);
nand_1 g08121(new_n8497, new_n8496, new_n8498);
not_4  g08122(new_n8340, new_n8499);
nor_1  g08123(new_n8499, new_n8297, new_n8500);
nor_1  g08124(new_n8342, new_n8296, new_n8501);
nor_1  g08125(new_n8501, new_n8500, new_n8502);
xnor_1 g08126(new_n8502, new_n8498, new_n8503);
xnor_1 g08127(new_n8503, new_n8495, new_n8504);
nand_1 g08128(n4826, n2515, new_n8505);
nand_1 g08129(n12925, n6578, new_n8506);
xnor_1 g08130(new_n8506, new_n8505, new_n8507);
nand_1 g08131(n6359, n5314, new_n8508);
nand_1 g08132(n12069, n7546, new_n8509);
xnor_1 g08133(new_n8509, new_n8508, new_n8510);
xnor_1 g08134(new_n8510, new_n8507, new_n8511);
nand_1 g08135(new_n8309, new_n8308, new_n8512);
nand_1 g08136(new_n8311, new_n8307, new_n8513);
nand_1 g08137(new_n8513, new_n8512, new_n8514);
nand_1 g08138(new_n8322, new_n8318, new_n8515);
nand_1 g08139(new_n8515, new_n8320, new_n8516);
not_4  g08140(new_n8516, new_n8517);
nand_1 g08141(n11296, n11153, new_n8518);
not_4  g08142(new_n8518, new_n8519);
nand_1 g08143(new_n8519, new_n8517, new_n8520);
nand_1 g08144(new_n8519, new_n8253, new_n8521);
nand_1 g08145(new_n8521, new_n8516, new_n8522);
nand_1 g08146(new_n8522, new_n8520, new_n8523);
xnor_1 g08147(new_n8523, new_n8514, new_n8524);
xnor_1 g08148(new_n8524, new_n8511, new_n8525);
xnor_1 g08149(new_n8525, new_n8504, new_n8526);
not_4  g08150(new_n8526, new_n8527);
nor_1  g08151(new_n8398_1, new_n8399, new_n8528);
nand_1 g08152(new_n8376, new_n8344, new_n8529);
not_4  g08153(new_n8042, new_n8530);
nand_1 g08154(new_n8076, new_n8530, new_n8531);
nand_1 g08155(new_n8087, new_n8077, new_n8532);
nand_1 g08156(new_n8532, new_n8531, new_n8533);
nand_1 g08157(new_n8337, new_n8333, new_n8534);
not_4  g08158(new_n8059, new_n8535);
nand_1 g08159(new_n8065_1, new_n8535, new_n8536);
not_4  g08160(new_n8056, new_n8537);
nand_1 g08161(new_n8066, new_n8537, new_n8538);
nand_1 g08162(new_n8538, new_n8536, new_n8539);
not_4  g08163(new_n8128, new_n8540);
nand_1 g08164(new_n8540, new_n8122, new_n8541);
not_4  g08165(new_n8146, new_n8542);
nand_1 g08166(new_n8542, new_n8129, new_n8543);
nand_1 g08167(new_n8543, new_n8541, new_n8544);
xnor_1 g08168(new_n8544, new_n8539, new_n8545);
nand_1 g08169(new_n8315, new_n8303_1, new_n8546);
nand_1 g08170(n8595, n1094, new_n8547);
nand_1 g08171(n2564, n1835, new_n8548);
not_4  g08172(new_n8548, new_n8549);
xnor_1 g08173(new_n8549, new_n8547, new_n8550);
xnor_1 g08174(new_n8550, new_n8546, new_n8551);
nand_1 g08175(new_n8222, new_n8221, new_n8552);
nand_1 g08176(new_n8224, new_n8220, new_n8553);
nand_1 g08177(new_n8553, new_n8552, new_n8554);
nand_1 g08178(n12391, n10965, new_n8555);
not_4  g08179(new_n8555, new_n8556);
nand_1 g08180(n7891, n503, new_n8557);
nand_1 g08181(n9457, n405, new_n8558);
xnor_1 g08182(new_n8558, new_n8557, new_n8559);
xnor_1 g08183(new_n8559, new_n8556, new_n8560);
xnor_1 g08184(new_n8560, new_n8554, new_n8561);
nand_1 g08185(n8065, n6986, new_n8562);
nand_1 g08186(n10439, n2226, new_n8563);
xnor_1 g08187(new_n8563, new_n8562, new_n8564);
xnor_1 g08188(new_n8564, new_n8561, new_n8565);
xnor_1 g08189(new_n8565, new_n8551, new_n8566);
nand_1 g08190(new_n8051, new_n8050, new_n8567);
nand_1 g08191(new_n8053, new_n8049, new_n8568);
nand_1 g08192(new_n8568, new_n8567, new_n8569);
nand_1 g08193(n11536, n6687, new_n8570);
nand_1 g08194(n6611, n996, new_n8571);
xnor_1 g08195(new_n8571, new_n8570, new_n8572);
nand_1 g08196(n4921, n4516, new_n8573);
nand_1 g08197(n9920, n3842, new_n8574);
xnor_1 g08198(new_n8574, new_n8573, new_n8575);
xnor_1 g08199(new_n8575, new_n8572, new_n8576);
xnor_1 g08200(new_n8576, new_n8569, new_n8577);
nand_1 g08201(n9956, n2087, new_n8578);
nand_1 g08202(n7733, n1199, new_n8579);
nand_1 g08203(n5767, n217, new_n8580);
xnor_1 g08204(new_n8580, new_n8579, new_n8581);
nand_1 g08205(n7160, n4970, new_n8582);
nand_1 g08206(n7610, n4828, new_n8583);
xnor_1 g08207(new_n8583, new_n8582, new_n8584);
xnor_1 g08208(new_n8584, new_n8581, new_n8585);
xnor_1 g08209(new_n8585, new_n8578, new_n8586);
xnor_1 g08210(new_n8586, new_n8577, new_n8587);
nand_1 g08211(new_n8144, new_n8138_1, new_n8588);
nand_1 g08212(new_n8588, new_n8136, new_n8589);
nand_1 g08213(n8433, n4817, new_n8590);
nand_1 g08214(n10678, n6126, new_n8591);
xnor_1 g08215(new_n8591, new_n8590, new_n8592);
xnor_1 g08216(new_n8592, new_n8589, new_n8593);
xnor_1 g08217(new_n8593, new_n8587, new_n8594);
xnor_1 g08218(new_n8594, new_n8566, new_n8595_1);
xnor_1 g08219(new_n8595_1, new_n8545, new_n8596);
xnor_1 g08220(new_n8596, new_n8534, new_n8597);
xnor_1 g08221(new_n8597, new_n8533, new_n8598);
not_4  g08222(new_n8598, new_n8599);
nor_1  g08223(new_n8599, new_n8529, new_n8600);
nor_1  g08224(new_n8364, new_n8365, new_n8601);
nor_1  g08225(new_n8598, new_n8601, new_n8602);
nor_1  g08226(new_n8602, new_n8600, new_n8603);
not_4  g08227(new_n8326, new_n8604);
nand_1 g08228(new_n8604, new_n8324, new_n8605);
nand_1 g08229(new_n8327, new_n8317, new_n8606);
nand_1 g08230(new_n8606, new_n8605, new_n8607);
not_4  g08231(new_n8607, new_n8608);
nand_1 g08232(new_n8608, new_n8603, new_n8609);
nand_1 g08233(new_n8598, new_n8601, new_n8610);
nand_1 g08234(new_n8599, new_n8529, new_n8611);
nand_1 g08235(new_n8611, new_n8610, new_n8612);
nand_1 g08236(new_n8607, new_n8612, new_n8613);
nand_1 g08237(new_n8613, new_n8609, new_n8614);
nand_1 g08238(new_n8614, new_n8528, new_n8615);
nand_1 g08239(new_n8424, new_n8374, new_n8616);
nor_1  g08240(new_n8607, new_n8612, new_n8617);
nor_1  g08241(new_n8608, new_n8603, new_n8618);
nor_1  g08242(new_n8618, new_n8617, new_n8619);
nand_1 g08243(new_n8619, new_n8616, new_n8620);
nand_1 g08244(new_n8620, new_n8615, new_n8621);
nor_1  g08245(new_n8621, new_n8527, new_n8622);
nor_1  g08246(new_n8619, new_n8616, new_n8623);
nor_1  g08247(new_n8614, new_n8528, new_n8624);
nor_1  g08248(new_n8624, new_n8623, new_n8625);
nor_1  g08249(new_n8625, new_n8526, new_n8626);
nor_1  g08250(new_n8626, new_n8622, new_n8627);
nand_1 g08251(new_n8627, new_n8431, new_n8628);
not_4  g08252(new_n8422, new_n8629);
nor_1  g08253(new_n8426, new_n8423, new_n8630);
nor_1  g08254(new_n8630, new_n8409, new_n8631);
nand_1 g08255(new_n8631, new_n8629, new_n8632);
nand_1 g08256(new_n8632, new_n8427, new_n8633);
nand_1 g08257(new_n8625, new_n8526, new_n8634);
nand_1 g08258(new_n8621, new_n8527, new_n8635);
nand_1 g08259(new_n8635, new_n8634, new_n8636);
nand_1 g08260(new_n8636, new_n8633, new_n8637);
nand_1 g08261(new_n8637, new_n8628, n2679);
not_4  g08262(new_n6272, new_n8639);
nand_1 g08263(new_n6297, new_n8639, new_n8640);
not_4  g08264(new_n8640, new_n8641);
nand_1 g08265(n6687, n2253, new_n8642);
not_4  g08266(new_n8642, new_n8643);
nand_1 g08267(n10223, n6770, new_n8644);
nand_1 g08268(n9920, n2879, new_n8645);
nand_1 g08269(n7265, n3627, new_n8646);
not_4  g08270(new_n8646, new_n8647);
xnor_1 g08271(new_n8647, new_n8645, new_n8648);
xnor_1 g08272(new_n8648, new_n8644, new_n8649);
not_4  g08273(new_n6277, new_n8650);
not_4  g08274(new_n6275, new_n8651);
nor_1  g08275(new_n6280, new_n8651, new_n8652);
nor_1  g08276(new_n8652, new_n8650, new_n8653);
xnor_1 g08277(new_n8653, new_n8649, new_n8654);
nand_1 g08278(n9195, n2564, new_n8655);
nand_1 g08279(n4634, n4189, new_n8656);
not_4  g08280(new_n8656, new_n8657);
xnor_1 g08281(new_n8657, new_n8655, new_n8658);
xnor_1 g08282(new_n8658, new_n8654, new_n8659);
nor_1  g08283(new_n6281, new_n6274, new_n8660);
not_4  g08284(new_n8660, new_n8661);
not_4  g08285(new_n6287, new_n8662);
nand_1 g08286(new_n8662, new_n6283, new_n8663);
nand_1 g08287(new_n8663, new_n8661, new_n8664);
xnor_1 g08288(new_n8664, new_n8659, new_n8665_1);
not_4  g08289(new_n6273_1, new_n8666);
nand_1 g08290(new_n6288, new_n8666, new_n8667);
nand_1 g08291(new_n6295, new_n6289, new_n8668);
nand_1 g08292(new_n8668, new_n8667, new_n8669);
xnor_1 g08293(new_n8669, new_n8665_1, new_n8670);
nand_1 g08294(new_n8670, new_n8643, new_n8671);
nor_1  g08295(new_n8670, new_n8643, new_n8672);
not_4  g08296(new_n8672, new_n8673);
nand_1 g08297(new_n8673, new_n8671, new_n8674);
nand_1 g08298(new_n8674, new_n8641, new_n8675);
not_4  g08299(new_n8674, new_n8676);
nand_1 g08300(new_n8676, new_n8640, new_n8677);
nand_1 g08301(new_n8677, new_n8675, new_n8678);
nand_1 g08302(new_n6581, new_n6546, new_n8679);
xnor_1 g08303(new_n8679, new_n8678, new_n8680);
not_4  g08304(new_n6331, new_n8681);
nand_1 g08305(new_n6352, new_n8681, new_n8682);
nand_1 g08306(n12221, n8336, new_n8683);
nand_1 g08307(n9189, n2226, new_n8684);
nand_1 g08308(n2024, n1094, new_n8685);
nand_1 g08309(n10678, n7946, new_n8686);
not_4  g08310(new_n8686, new_n8687);
xnor_1 g08311(new_n8687, new_n8685, new_n8688);
xnor_1 g08312(new_n8688, new_n8684, new_n8689);
not_4  g08313(new_n6340, new_n8690);
not_4  g08314(new_n6338, new_n8691);
nor_1  g08315(new_n6343, new_n8691, new_n8692);
nor_1  g08316(new_n8692, new_n8690, new_n8693);
nand_1 g08317(new_n8693, new_n8689, new_n8694);
not_4  g08318(new_n8694, new_n8695);
nor_1  g08319(new_n8693, new_n8689, new_n8696);
nor_1  g08320(new_n8696, new_n8695, new_n8697);
nand_1 g08321(n12145, n10928, new_n8698);
nand_1 g08322(n6986, n2522, new_n8699);
xnor_1 g08323(new_n8699, new_n8698, new_n8700);
xnor_1 g08324(new_n8700, new_n8697, new_n8701);
nor_1  g08325(new_n6335, new_n6333, new_n8702);
not_4  g08326(new_n6337, new_n8703);
nor_1  g08327(new_n6344, new_n8703, new_n8704);
nor_1  g08328(new_n8704, new_n8702, new_n8705);
not_4  g08329(new_n8705, new_n8706);
xnor_1 g08330(new_n8706, new_n8701, new_n8707);
not_4  g08331(new_n6332, new_n8708);
nand_1 g08332(new_n6345, new_n8708, new_n8709);
nand_1 g08333(new_n6350, new_n6346, new_n8710);
nand_1 g08334(new_n8710, new_n8709, new_n8711);
xnor_1 g08335(new_n8711, new_n8707, new_n8712);
xnor_1 g08336(new_n8712, new_n8683, new_n8713);
xnor_1 g08337(new_n8713, new_n8682, new_n8714);
nand_1 g08338(new_n6477, new_n6353, new_n8715);
nand_1 g08339(new_n6542, new_n6479, new_n8716);
nand_1 g08340(new_n8716, new_n8715, new_n8717_1);
xnor_1 g08341(new_n8717_1, new_n8714, new_n8718);
nand_1 g08342(new_n6501, new_n6390, new_n8719);
not_4  g08343(new_n8719, new_n8720);
nand_1 g08344(n12069, n5798, new_n8721);
not_4  g08345(new_n8721, new_n8722);
nand_1 g08346(n7160, n5579, new_n8723);
nand_1 g08347(new_n6490, new_n6486, new_n8724);
nand_1 g08348(new_n8724, new_n6489, new_n8725);
nand_1 g08349(new_n8725, new_n8723, new_n8726);
not_4  g08350(new_n8723, new_n8727);
nand_1 g08351(new_n8725, new_n6368, new_n8728);
nand_1 g08352(new_n8728, new_n8727, new_n8729);
nand_1 g08353(new_n8729, new_n8726, new_n8730);
nand_1 g08354(n4828, n2498, new_n8731);
nand_1 g08355(n2558, n2515, new_n8732);
nand_1 g08356(new_n8732, new_n8731, new_n8733);
not_4  g08357(new_n8731, new_n8734);
not_4  g08358(new_n8732, new_n8735);
nand_1 g08359(new_n8735, new_n8734, new_n8736);
nand_1 g08360(new_n8736, new_n8733, new_n8737);
nand_1 g08361(new_n8737, new_n8730, new_n8738);
not_4  g08362(new_n8726, new_n8739);
xnor_1 g08363(new_n6489, new_n6358_1, new_n8740);
nor_1  g08364(new_n8740, new_n6487, new_n8741);
nor_1  g08365(new_n8741, new_n6488, new_n8742);
nor_1  g08366(new_n8742, new_n6369, new_n8743);
nor_1  g08367(new_n8743, new_n8723, new_n8744);
nor_1  g08368(new_n8744, new_n8739, new_n8745);
not_4  g08369(new_n8737, new_n8746);
nand_1 g08370(new_n8746, new_n8745, new_n8747);
nand_1 g08371(new_n8747, new_n8738, new_n8748);
not_4  g08372(new_n8748, new_n8749);
nand_1 g08373(n12391, n6016, new_n8750);
nand_1 g08374(n7891, n521, new_n8751);
nand_1 g08375(new_n8751, new_n8750, new_n8752);
not_4  g08376(new_n8750, new_n8753);
not_4  g08377(new_n8751, new_n8754);
nand_1 g08378(new_n8754, new_n8753, new_n8755);
nand_1 g08379(new_n8755, new_n8752, new_n8756);
xnor_1 g08380(new_n8756, new_n8749, new_n8757);
not_4  g08381(new_n8757, new_n8758);
nor_1  g08382(new_n6483, new_n6481, new_n8759_1);
not_4  g08383(new_n6485, new_n8760);
nor_1  g08384(new_n6491, new_n8760, new_n8761);
nor_1  g08385(new_n8761, new_n8759_1, new_n8762);
nor_1  g08386(new_n8762, new_n8758, new_n8763);
not_4  g08387(new_n8763, new_n8764);
nand_1 g08388(new_n8762, new_n8758, new_n8765);
nand_1 g08389(new_n8765, new_n8764, new_n8766);
not_4  g08390(new_n6480, new_n8767);
nand_1 g08391(new_n6492, new_n8767, new_n8768);
nand_1 g08392(new_n6499, new_n8768, new_n8769);
not_4  g08393(new_n8769, new_n8770);
nor_1  g08394(new_n8770, new_n8766, new_n8771);
not_4  g08395(new_n8771, new_n8772);
nand_1 g08396(new_n8770, new_n8766, new_n8773);
nand_1 g08397(new_n8773, new_n8772, new_n8774);
not_4  g08398(new_n8774, new_n8775);
nand_1 g08399(new_n8775, new_n8722, new_n8776);
nand_1 g08400(new_n8774, new_n8721, new_n8777);
nand_1 g08401(new_n8777, new_n8776, new_n8778);
not_4  g08402(new_n8778, new_n8779);
nand_1 g08403(new_n8779, new_n8720, new_n8780);
nand_1 g08404(new_n8778, new_n8719, new_n8781);
nand_1 g08405(new_n8781, new_n8780, new_n8782);
not_4  g08406(new_n8782, new_n8783);
nand_1 g08407(n11222, n5153, new_n8784);
nand_1 g08408(n3342, n996, new_n8785);
nand_1 g08409(n9111, n5767, new_n8786);
nand_1 g08410(n9763, n5319, new_n8787);
not_4  g08411(new_n8787, new_n8788);
xnor_1 g08412(new_n8788, new_n8786, new_n8789);
xnor_1 g08413(new_n8789, new_n8785, new_n8790);
nand_1 g08414(new_n6518, new_n6513, new_n8791);
nand_1 g08415(new_n8791, new_n6516, new_n8792);
xnor_1 g08416(new_n8792, new_n8790, new_n8793);
not_4  g08417(new_n8793, new_n8794);
nand_1 g08418(n11153, n7270, new_n8795);
nand_1 g08419(n5314, n806, new_n8796);
not_4  g08420(new_n8796, new_n8797);
xnor_1 g08421(new_n8797, new_n8795, new_n8798);
xnor_1 g08422(new_n8798, new_n8794, new_n8799);
not_4  g08423(new_n6512, new_n8800);
nand_1 g08424(new_n6520, new_n8800, new_n8801);
nand_1 g08425(new_n8801, new_n6510, new_n8802);
xnor_1 g08426(new_n8802, new_n8799, new_n8803);
not_4  g08427(new_n6505, new_n8804);
nand_1 g08428(new_n6521, new_n8804, new_n8805);
nand_1 g08429(new_n6526, new_n6522, new_n8806);
nand_1 g08430(new_n8806, new_n8805, new_n8807);
xnor_1 g08431(new_n8807, new_n8803, new_n8808);
xnor_1 g08432(new_n8808, new_n8784, new_n8809);
xnor_1 g08433(new_n8809, new_n6529, new_n8810);
not_4  g08434(new_n8810, new_n8811);
nand_1 g08435(new_n8811, new_n8783, new_n8812);
nand_1 g08436(new_n8810, new_n8782, new_n8813);
nand_1 g08437(new_n8813, new_n8812, new_n8814);
nand_1 g08438(new_n6540, new_n6534, new_n8815);
nor_1  g08439(new_n8815, new_n8814, new_n8816);
not_4  g08440(new_n8816, new_n8817);
nand_1 g08441(new_n8815, new_n8814, new_n8818);
nand_1 g08442(new_n8818, new_n8817, new_n8819_1);
nor_1  g08443(new_n8819_1, new_n8718, new_n8820);
not_4  g08444(new_n8820, new_n8821);
nand_1 g08445(new_n8819_1, new_n8718, new_n8822);
nand_1 g08446(new_n8822, new_n8821, new_n8823);
xnor_1 g08447(new_n8823, new_n8680, n2708);
nand_1 g08448(new_n933, new_n932, new_n8825);
nand_1 g08449(new_n8825, new_n935, n2818);
nand_1 g08450(new_n2285, new_n2253_1, new_n8827);
nand_1 g08451(new_n8827, new_n2287, n2902);
nand_1 g08452(n11407, n5305, new_n8829);
nand_1 g08453(n12709, n8759, new_n8830);
nand_1 g08454(n12489, n5331, new_n8831);
not_4  g08455(new_n8831, new_n8832);
nand_1 g08456(n10990, n7965, new_n8833);
not_4  g08457(new_n8833, new_n8834);
nand_1 g08458(new_n8834, new_n8832, new_n8835);
nand_1 g08459(new_n8833, new_n8831, new_n8836);
nand_1 g08460(new_n8836, new_n8835, new_n8837);
not_4  g08461(new_n8837, new_n8838);
xnor_1 g08462(new_n8838, new_n8830, new_n8839);
xnor_1 g08463(new_n8839, new_n8829, n3071);
nand_1 g08464(new_n3165, new_n3164, new_n8841);
nand_1 g08465(new_n8841, new_n3167, n3124);
not_4  g08466(new_n8829, new_n8843);
nand_1 g08467(new_n8839, new_n8843, new_n8844);
nand_1 g08468(n11407, n5964, new_n8845);
nand_1 g08469(n5305, n5212, new_n8846);
xnor_1 g08470(new_n8846, new_n8845, new_n8847);
nand_1 g08471(new_n8847, new_n8844, new_n8848);
not_4  g08472(new_n8830, new_n8849);
nand_1 g08473(new_n8838, new_n8849, new_n8850);
nand_1 g08474(n11728, n8759, new_n8851);
nand_1 g08475(n12709, n6776, new_n8852);
xnor_1 g08476(new_n8852, new_n8851, new_n8853);
not_4  g08477(new_n8853, new_n8854);
xnor_1 g08478(new_n8854, new_n8850, new_n8855);
not_4  g08479(new_n8855, new_n8856);
nand_1 g08480(n7159, n5331, new_n8857);
nand_1 g08481(n12489, n8476, new_n8858);
xnor_1 g08482(new_n8858, new_n8857, new_n8859);
xnor_1 g08483(new_n8859, new_n8835, new_n8860);
nand_1 g08484(n7965, n5760, new_n8861);
nand_1 g08485(n10990, n7388, new_n8862);
xnor_1 g08486(new_n8862, new_n8861, new_n8863);
xnor_1 g08487(new_n8863, new_n8860, new_n8864);
nor_1  g08488(new_n8864, new_n8856, new_n8865);
not_4  g08489(new_n8865, new_n8866);
nand_1 g08490(new_n8864, new_n8856, new_n8867);
nand_1 g08491(new_n8867, new_n8866, new_n8868);
not_4  g08492(new_n8868, new_n8869);
xnor_1 g08493(new_n8847, new_n8844, new_n8870);
nor_1  g08494(new_n8870, new_n8869, new_n8871);
not_4  g08495(new_n8871, new_n8872);
nand_1 g08496(new_n8872, new_n8848, new_n8873);
nand_1 g08497(n5964, n5212, new_n8874);
not_4  g08498(new_n8874, new_n8875);
nand_1 g08499(new_n8875, new_n8829, new_n8876);
nand_1 g08500(n11407, n1097, new_n8877);
nand_1 g08501(n11877, n5305, new_n8878);
nand_1 g08502(new_n8878, new_n8877, new_n8879);
nor_1  g08503(new_n8878, new_n8877, new_n8880);
not_4  g08504(new_n8880, new_n8881);
nand_1 g08505(new_n8881, new_n8879, new_n8882);
nand_1 g08506(new_n8882, new_n8876, new_n8883);
not_4  g08507(new_n8883, new_n8884);
not_4  g08508(new_n8879, new_n8885);
nor_1  g08509(new_n8885, new_n8876, new_n8886);
nor_1  g08510(new_n8886, new_n8884, new_n8887);
not_4  g08511(new_n8887, new_n8888);
xnor_1 g08512(new_n8888, new_n8873, new_n8889);
not_4  g08513(new_n8889, new_n8890);
not_4  g08514(new_n8850, new_n8891);
nand_1 g08515(new_n8854, new_n8891, new_n8892);
nand_1 g08516(new_n8866, new_n8892, new_n8893);
nand_1 g08517(n11728, n6776, new_n8894);
not_4  g08518(new_n8894, new_n8895);
nand_1 g08519(new_n8895, new_n8830, new_n8896);
nand_1 g08520(n12709, n12299, new_n8897);
nand_1 g08521(n8759, n6429, new_n8898);
nand_1 g08522(new_n8898, new_n8897, new_n8899);
nor_1  g08523(new_n8898, new_n8897, new_n8900);
not_4  g08524(new_n8900, new_n8901);
nand_1 g08525(new_n8901, new_n8899, new_n8902);
nand_1 g08526(new_n8902, new_n8896, new_n8903);
not_4  g08527(new_n8903, new_n8904);
not_4  g08528(new_n8899, new_n8905);
nor_1  g08529(new_n8905, new_n8896, new_n8906);
nor_1  g08530(new_n8906, new_n8904, new_n8907);
xnor_1 g08531(new_n8907, new_n8893, new_n8908);
not_4  g08532(new_n8908, new_n8909);
nand_1 g08533(n8476, n7159, new_n8910);
not_4  g08534(new_n8910, new_n8911);
nand_1 g08535(new_n8911, new_n8831, new_n8912);
nand_1 g08536(n12489, n2530, new_n8913);
nand_1 g08537(n12777, n5331, new_n8914);
nand_1 g08538(new_n8914, new_n8913, new_n8915);
nand_1 g08539(n12777, n2530, new_n8916);
not_4  g08540(new_n8916, new_n8917);
nand_1 g08541(new_n8917, new_n8832, new_n8918);
nand_1 g08542(new_n8918, new_n8915, new_n8919);
nand_1 g08543(new_n8919, new_n8912, new_n8920);
not_4  g08544(new_n8920, new_n8921);
not_4  g08545(new_n8915, new_n8922);
nor_1  g08546(new_n8922, new_n8912, new_n8923);
nor_1  g08547(new_n8923, new_n8921, new_n8924);
nand_1 g08548(n7388, n5760, new_n8925);
not_4  g08549(new_n8925, new_n8926);
nand_1 g08550(new_n8926, new_n8833, new_n8927);
nand_1 g08551(n11892, n10990, new_n8928);
nand_1 g08552(n7965, n1478, new_n8929);
nand_1 g08553(new_n8929, new_n8928, new_n8930);
not_4  g08554(new_n8928, new_n8931);
not_4  g08555(new_n8929, new_n8932);
nand_1 g08556(new_n8932, new_n8931, new_n8933);
nand_1 g08557(new_n8933, new_n8930, new_n8934);
nand_1 g08558(new_n8934, new_n8927, new_n8935);
not_4  g08559(new_n8935, new_n8936);
not_4  g08560(new_n8930, new_n8937);
nor_1  g08561(new_n8937, new_n8927, new_n8938);
nor_1  g08562(new_n8938, new_n8936, new_n8939);
xnor_1 g08563(new_n8939, new_n8924, new_n8940);
nand_1 g08564(new_n8859, new_n8835, new_n8941);
not_4  g08565(new_n8860, new_n8942);
nand_1 g08566(new_n8863, new_n8942, new_n8943);
nand_1 g08567(new_n8943, new_n8941, new_n8944);
nor_1  g08568(new_n8944, new_n8940, new_n8945);
not_4  g08569(new_n8945, new_n8946);
nand_1 g08570(new_n8944, new_n8940, new_n8947);
nand_1 g08571(new_n8947, new_n8946, new_n8948);
not_4  g08572(new_n8948, new_n8949);
nand_1 g08573(new_n8949, new_n8909, new_n8950);
nand_1 g08574(new_n8948, new_n8908, new_n8951);
nand_1 g08575(new_n8951, new_n8950, new_n8952);
xnor_1 g08576(new_n8952, new_n8890, n3214);
xnor_1 g08577(new_n6081, new_n6078, n3230);
xnor_1 g08578(new_n5496, new_n5624, n3272);
nand_1 g08579(n5964, n4370, new_n8956);
nand_1 g08580(n11407, n4312, new_n8957);
nand_1 g08581(n11877, n5964, new_n8958);
nand_1 g08582(new_n8958, new_n8957, new_n8959);
nor_1  g08583(new_n8958, new_n8957, new_n8960);
not_4  g08584(new_n8960, new_n8961);
nand_1 g08585(n5212, n1097, new_n8962);
nand_1 g08586(new_n8962, new_n8961, new_n8963);
nand_1 g08587(new_n8963, new_n8959, new_n8964);
nor_1  g08588(new_n8964, new_n8956, new_n8965);
not_4  g08589(new_n8965, new_n8966);
nand_1 g08590(new_n8964, new_n8956, new_n8967);
nand_1 g08591(new_n8967, new_n8966, new_n8968);
not_4  g08592(new_n8968, new_n8969);
nand_1 g08593(n5212, n4312, new_n8970);
nand_1 g08594(n11877, n1097, new_n8971);
nand_1 g08595(n12705, n11407, new_n8972);
nand_1 g08596(new_n8972, new_n8971, new_n8973);
not_4  g08597(new_n8971, new_n8974);
not_4  g08598(new_n8972, new_n8975);
nand_1 g08599(new_n8975, new_n8974, new_n8976);
nand_1 g08600(new_n8976, new_n8973, new_n8977);
xnor_1 g08601(new_n8977, new_n8970, new_n8978);
not_4  g08602(new_n8978, new_n8979);
nand_1 g08603(new_n8979, new_n8969, new_n8980);
nand_1 g08604(new_n8980, new_n8966, new_n8981);
nand_1 g08605(n5964, n5320, new_n8982);
not_4  g08606(new_n8982, new_n8983);
nand_1 g08607(n4370, n1097, new_n8984);
not_4  g08608(new_n8984, new_n8985);
nand_1 g08609(new_n8985, new_n8983, new_n8986);
nand_1 g08610(new_n8984, new_n8982, new_n8987);
nand_1 g08611(new_n8987, new_n8986, new_n8988);
xnor_1 g08612(new_n8988, new_n8981, new_n8989);
nand_1 g08613(n11877, n4312, new_n8990);
nand_1 g08614(n12705, n5212, new_n8991);
nand_1 g08615(n12025, n11407, new_n8992);
not_4  g08616(new_n8992, new_n8993);
xnor_1 g08617(new_n8993, new_n8991, new_n8994);
xnor_1 g08618(new_n8994, new_n8990, new_n8995);
nand_1 g08619(new_n8976, new_n8970, new_n8996);
nand_1 g08620(new_n8996, new_n8973, new_n8997);
xnor_1 g08621(new_n8997, new_n8995, new_n8998);
xnor_1 g08622(new_n8998, new_n8989, new_n8999);
nand_1 g08623(n5320, n5305, new_n9000);
nand_1 g08624(new_n8978, new_n8968, new_n9001);
nand_1 g08625(new_n9001, new_n8980, new_n9002);
nand_1 g08626(new_n9002, new_n9000, new_n9003);
xnor_1 g08627(new_n9002, new_n9000, new_n9004);
not_4  g08628(new_n9004, new_n9005);
nand_1 g08629(n5305, n4370, new_n9006);
nand_1 g08630(new_n8881, new_n8874, new_n9007);
nand_1 g08631(new_n9007, new_n8879, new_n9008);
nor_1  g08632(new_n9008, new_n9006, new_n9009);
xnor_1 g08633(new_n9008, new_n9006, new_n9010);
nand_1 g08634(new_n8961, new_n8959, new_n9011);
xnor_1 g08635(new_n9011, new_n8962, new_n9012);
nor_1  g08636(new_n9012, new_n9010, new_n9013);
nor_1  g08637(new_n9013, new_n9009, new_n9014);
nand_1 g08638(new_n9014, new_n9005, new_n9015);
nand_1 g08639(new_n9015, new_n9003, new_n9016);
nor_1  g08640(new_n9016, new_n8999, new_n9017);
not_4  g08641(new_n8994, new_n9018);
nand_1 g08642(new_n9018, new_n8990, new_n9019);
nand_1 g08643(new_n8997, new_n8995, new_n9020);
nand_1 g08644(new_n9020, new_n9019, new_n9021);
nand_1 g08645(n12000, n5964, new_n9022);
nand_1 g08646(n5320, n1097, new_n9023);
nand_1 g08647(n9725, n5305, new_n9024);
not_4  g08648(new_n9024, new_n9025);
xnor_1 g08649(new_n9025, new_n9023, new_n9026);
xnor_1 g08650(new_n9026, new_n9022, new_n9027);
xnor_1 g08651(new_n9027, new_n9021, new_n9028);
not_4  g08652(new_n9028, new_n9029);
not_4  g08653(new_n8991, new_n9030);
nand_1 g08654(new_n8993, new_n9030, new_n9031);
nand_1 g08655(n4370, n4312, new_n9032);
xnor_1 g08656(new_n9032, new_n9031, new_n9033);
nand_1 g08657(n12025, n5212, new_n9034);
not_4  g08658(new_n9034, new_n9035);
nand_1 g08659(n12705, n11877, new_n9036);
nand_1 g08660(n11407, n11257, new_n9037);
not_4  g08661(new_n9037, new_n9038);
xnor_1 g08662(new_n9038, new_n9036, new_n9039);
xnor_1 g08663(new_n9039, new_n9035, new_n9040);
xnor_1 g08664(new_n9040, new_n9033, new_n9041);
xnor_1 g08665(new_n9041, new_n9029, new_n9042);
not_4  g08666(new_n8988, new_n9043);
nand_1 g08667(new_n9043, new_n8981, new_n9044);
nand_1 g08668(new_n8998, new_n8989, new_n9045);
xnor_1 g08669(new_n9045, new_n8986, new_n9046);
nand_1 g08670(new_n9046, new_n9044, new_n9047);
xnor_1 g08671(new_n9047, new_n9042, new_n9048);
xnor_1 g08672(new_n9048, new_n9017, new_n9049);
nand_1 g08673(n12000, n5305, new_n9050);
not_4  g08674(new_n9050, new_n9051);
not_4  g08675(new_n8999, new_n9052);
xnor_1 g08676(new_n9016, new_n9052, new_n9053);
nand_1 g08677(new_n9053, new_n9051, new_n9054);
xnor_1 g08678(new_n9012, new_n9010, new_n9055);
not_4  g08679(new_n9055, new_n9056);
nand_1 g08680(new_n8884, new_n8875, new_n9057);
not_4  g08681(new_n9057, new_n9058);
nand_1 g08682(new_n9058, new_n9056, new_n9059);
xnor_1 g08683(new_n9014, new_n9004, new_n9060);
nor_1  g08684(new_n9060, new_n9059, new_n9061);
xnor_1 g08685(new_n9053, new_n9050, new_n9062);
nand_1 g08686(new_n9062, new_n9061, new_n9063);
nand_1 g08687(new_n9063, new_n9054, new_n9064);
xnor_1 g08688(new_n9064, new_n9049, new_n9065);
not_4  g08689(new_n9065, new_n9066);
nand_1 g08690(n8759, n8717, new_n9067);
not_4  g08691(new_n9067, new_n9068);
nand_1 g08692(n7436, n6429, new_n9069);
not_4  g08693(new_n9069, new_n9070);
nand_1 g08694(n12709, n9241, new_n9071);
nand_1 g08695(n11728, n8276, new_n9072);
not_4  g08696(new_n9072, new_n9073);
xnor_1 g08697(new_n9073, new_n9071, new_n9074);
nor_1  g08698(new_n9074, new_n9070, new_n9075);
not_4  g08699(new_n9075, new_n9076);
nand_1 g08700(new_n9074, new_n9070, new_n9077);
nand_1 g08701(new_n9077, new_n9076, new_n9078);
nand_1 g08702(n12299, n6429, new_n9079);
nand_1 g08703(n12709, n8276, new_n9080_1);
nand_1 g08704(new_n9080_1, new_n9079, new_n9081);
not_4  g08705(new_n9079, new_n9082);
not_4  g08706(new_n9080_1, new_n9083);
nand_1 g08707(new_n9083, new_n9082, new_n9084);
nand_1 g08708(n11728, n7436, new_n9085);
nand_1 g08709(new_n9085, new_n9084, new_n9086);
nand_1 g08710(new_n9086, new_n9081, new_n9087);
xnor_1 g08711(new_n9087, new_n9078, new_n9088);
nand_1 g08712(n6776, n2433, new_n9089);
nand_1 g08713(n12299, n8819, new_n9090);
not_4  g08714(new_n9090, new_n9091);
xnor_1 g08715(new_n9091, new_n9089, new_n9092);
xnor_1 g08716(new_n9092, new_n9088, new_n9093);
nand_1 g08717(n8819, n6776, new_n9094);
nand_1 g08718(n12709, n7436, new_n9095);
nand_1 g08719(n6776, n6429, new_n9096);
nand_1 g08720(new_n9096, new_n9095, new_n9097);
not_4  g08721(new_n9095, new_n9098);
not_4  g08722(new_n9096, new_n9099);
nand_1 g08723(new_n9099, new_n9098, new_n9100);
nand_1 g08724(n12299, n11728, new_n9101);
nand_1 g08725(new_n9101, new_n9100, new_n9102);
nand_1 g08726(new_n9102, new_n9097, new_n9103);
nor_1  g08727(new_n9103, new_n9094, new_n9104);
not_4  g08728(new_n9103, new_n9105);
xnor_1 g08729(new_n9105, new_n9094, new_n9106);
not_4  g08730(new_n9106, new_n9107);
nand_1 g08731(new_n9084, new_n9081, new_n9108);
xnor_1 g08732(new_n9108, new_n9085, new_n9109);
nor_1  g08733(new_n9109, new_n9107, new_n9110);
nor_1  g08734(new_n9110, new_n9104, new_n9111_1);
xnor_1 g08735(new_n9111_1, new_n9093, new_n9112);
nand_1 g08736(n8759, n2433, new_n9113);
not_4  g08737(new_n9113, new_n9114);
xnor_1 g08738(new_n9109, new_n9106, new_n9115);
nor_1  g08739(new_n9115, new_n9114, new_n9116);
not_4  g08740(new_n9116, new_n9117);
xnor_1 g08741(new_n9115, new_n9113, new_n9118);
nand_1 g08742(n8819, n8759, new_n9119);
nand_1 g08743(new_n8901, new_n8894, new_n9120);
nand_1 g08744(new_n9120, new_n8899, new_n9121);
nor_1  g08745(new_n9121, new_n9119, new_n9122);
xnor_1 g08746(new_n9121, new_n9119, new_n9123);
nand_1 g08747(new_n9100, new_n9097, new_n9124);
xnor_1 g08748(new_n9124, new_n9101, new_n9125);
nor_1  g08749(new_n9125, new_n9123, new_n9126);
nor_1  g08750(new_n9126, new_n9122, new_n9127);
nand_1 g08751(new_n9127, new_n9118, new_n9128);
nand_1 g08752(new_n9128, new_n9117, new_n9129);
xnor_1 g08753(new_n9129, new_n9112, new_n9130);
nand_1 g08754(new_n9130, new_n9068, new_n9131);
xnor_1 g08755(new_n9125, new_n9123, new_n9132);
not_4  g08756(new_n9132, new_n9133);
nand_1 g08757(new_n8904, new_n8895, new_n9134);
not_4  g08758(new_n9134, new_n9135);
nand_1 g08759(new_n9135, new_n9133, new_n9136);
not_4  g08760(new_n9136, new_n9137_1);
xnor_1 g08761(new_n9127, new_n9118, new_n9138);
nand_1 g08762(new_n9138, new_n9137_1, new_n9139);
not_4  g08763(new_n9139, new_n9140);
xnor_1 g08764(new_n9130, new_n9067, new_n9141);
nand_1 g08765(new_n9141, new_n9140, new_n9142);
nand_1 g08766(new_n9142, new_n9131, new_n9143);
not_4  g08767(new_n9129, new_n9144);
nand_1 g08768(new_n9144, new_n9112, new_n9145);
not_4  g08769(new_n9078, new_n9146);
nand_1 g08770(new_n9087, new_n9146, new_n9147);
nand_1 g08771(new_n9147, new_n9076, new_n9148);
not_4  g08772(new_n9148, new_n9149);
nand_1 g08773(n8717, n6776, new_n9150);
nand_1 g08774(n12299, n2433, new_n9151);
not_4  g08775(new_n9151, new_n9152);
nand_1 g08776(n8759, n7730, new_n9153);
not_4  g08777(new_n9153, new_n9154);
nand_1 g08778(new_n9154, new_n9152, new_n9155);
nand_1 g08779(new_n9153, new_n9151, new_n9156);
nand_1 g08780(new_n9156, new_n9155, new_n9157);
xnor_1 g08781(new_n9157, new_n9150, new_n9158);
xnor_1 g08782(new_n9158, new_n9149, new_n9159);
not_4  g08783(new_n9071, new_n9160);
nand_1 g08784(new_n9073, new_n9160, new_n9161);
nand_1 g08785(n8819, n7436, new_n9162);
not_4  g08786(new_n9162, new_n9163);
xnor_1 g08787(new_n9163, new_n9161, new_n9164);
nand_1 g08788(n11728, n9241, new_n9165);
nand_1 g08789(n8276, n6429, new_n9166);
nand_1 g08790(n12709, n10510, new_n9167);
not_4  g08791(new_n9167, new_n9168);
xnor_1 g08792(new_n9168, new_n9166, new_n9169);
xnor_1 g08793(new_n9169, new_n9165, new_n9170);
not_4  g08794(new_n9170, new_n9171);
xnor_1 g08795(new_n9171, new_n9164, new_n9172);
xnor_1 g08796(new_n9172, new_n9159, new_n9173);
not_4  g08797(new_n9088, new_n9174);
nand_1 g08798(new_n9092, new_n9174, new_n9175);
nor_1  g08799(new_n9090, new_n9089, new_n9176);
not_4  g08800(new_n9111_1, new_n9177);
nand_1 g08801(new_n9177, new_n9093, new_n9178);
not_4  g08802(new_n9178, new_n9179);
xnor_1 g08803(new_n9179, new_n9176, new_n9180);
nand_1 g08804(new_n9180, new_n9175, new_n9181);
xnor_1 g08805(new_n9181, new_n9173, new_n9182);
xnor_1 g08806(new_n9182, new_n9145, new_n9183);
xnor_1 g08807(new_n9183, new_n9143, new_n9184);
nand_1 g08808(n2393, n1478, new_n9185);
nand_1 g08809(n5860, n5760, new_n9186);
nand_1 g08810(n10990, n3986, new_n9187);
not_4  g08811(new_n9187, new_n9188);
xnor_1 g08812(new_n9188, new_n9186, new_n9189_1);
not_4  g08813(new_n9189_1, new_n9190);
xnor_1 g08814(new_n9190, new_n9185, new_n9191);
nand_1 g08815(n11892, n1478, new_n9192);
nand_1 g08816(n10990, n5860, new_n9193);
nand_1 g08817(new_n9193, new_n9192, new_n9194);
not_4  g08818(new_n9192, new_n9195_1);
not_4  g08819(new_n9193, new_n9196);
nand_1 g08820(new_n9196, new_n9195_1, new_n9197);
nand_1 g08821(n5760, n2393, new_n9198);
nand_1 g08822(new_n9198, new_n9197, new_n9199);
nand_1 g08823(new_n9199, new_n9194, new_n9200);
xnor_1 g08824(new_n9200, new_n9191, new_n9201);
nand_1 g08825(n12947, n7388, new_n9202);
nand_1 g08826(n11892, n11791, new_n9203);
not_4  g08827(new_n9203, new_n9204);
xnor_1 g08828(new_n9204, new_n9202, new_n9205);
xnor_1 g08829(new_n9205, new_n9201, new_n9206);
nand_1 g08830(n11791, n7388, new_n9207);
nand_1 g08831(n10990, n2393, new_n9208);
nand_1 g08832(n7388, n1478, new_n9209);
nand_1 g08833(new_n9209, new_n9208, new_n9210);
not_4  g08834(new_n9208, new_n9211);
not_4  g08835(new_n9209, new_n9212);
nand_1 g08836(new_n9212, new_n9211, new_n9213);
nand_1 g08837(n11892, n5760, new_n9214);
nand_1 g08838(new_n9214, new_n9213, new_n9215);
nand_1 g08839(new_n9215, new_n9210, new_n9216);
nor_1  g08840(new_n9216, new_n9207, new_n9217);
not_4  g08841(new_n9217, new_n9218);
not_4  g08842(new_n9216, new_n9219);
xnor_1 g08843(new_n9219, new_n9207, new_n9220);
not_4  g08844(new_n9198, new_n9221);
nand_1 g08845(new_n9197, new_n9194, new_n9222);
xnor_1 g08846(new_n9222, new_n9221, new_n9223);
nand_1 g08847(new_n9223, new_n9220, new_n9224);
nand_1 g08848(new_n9224, new_n9218, new_n9225);
xnor_1 g08849(new_n9225, new_n9206, new_n9226);
nand_1 g08850(n12947, n7965, new_n9227);
nand_1 g08851(n11791, n7965, new_n9228);
nand_1 g08852(new_n8933, new_n8925, new_n9229);
nand_1 g08853(new_n9229, new_n8930, new_n9230);
nor_1  g08854(new_n9230, new_n9228, new_n9231);
xnor_1 g08855(new_n9230, new_n9228, new_n9232);
nand_1 g08856(new_n9213, new_n9210, new_n9233);
xnor_1 g08857(new_n9233, new_n9214, new_n9234);
nor_1  g08858(new_n9234, new_n9232, new_n9235);
nor_1  g08859(new_n9235, new_n9231, new_n9236);
nand_1 g08860(new_n9236, new_n9227, new_n9237);
xnor_1 g08861(new_n9223, new_n9220, new_n9238);
not_4  g08862(new_n9236, new_n9239);
xnor_1 g08863(new_n9239, new_n9227, new_n9240);
nand_1 g08864(new_n9240, new_n9238, new_n9241_1);
nand_1 g08865(new_n9241_1, new_n9237, new_n9242);
nor_1  g08866(new_n9242, new_n9226, new_n9243);
not_4  g08867(new_n9186, new_n9244);
nand_1 g08868(new_n9188, new_n9244, new_n9245);
nand_1 g08869(n11791, n2393, new_n9246);
xnor_1 g08870(new_n9246, new_n9245, new_n9247);
nand_1 g08871(n5760, n3986, new_n9248);
nand_1 g08872(n5860, n1478, new_n9249);
nand_1 g08873(n10990, n5857, new_n9250);
nand_1 g08874(new_n9250, new_n9249, new_n9251);
not_4  g08875(new_n9249, new_n9252);
not_4  g08876(new_n9250, new_n9253);
nand_1 g08877(new_n9253, new_n9252, new_n9254);
nand_1 g08878(new_n9254, new_n9251, new_n9255);
xnor_1 g08879(new_n9255, new_n9248, new_n9256);
not_4  g08880(new_n9256, new_n9257);
xnor_1 g08881(new_n9257, new_n9247, new_n9258);
nand_1 g08882(n7388, n6441, new_n9259);
nand_1 g08883(n12947, n11892, new_n9260);
not_4  g08884(new_n9260, new_n9261);
nand_1 g08885(n11999, n7965, new_n9262);
xnor_1 g08886(new_n9262, new_n9261, new_n9263);
xnor_1 g08887(new_n9263, new_n9259, new_n9264);
nor_1  g08888(new_n9190, new_n9185, new_n9265);
nor_1  g08889(new_n9200, new_n9191, new_n9266);
nor_1  g08890(new_n9266, new_n9265, new_n9267);
xnor_1 g08891(new_n9267, new_n9264, new_n9268);
xnor_1 g08892(new_n9268, new_n9258, new_n9269);
not_4  g08893(new_n9201, new_n9270);
nand_1 g08894(new_n9205, new_n9270, new_n9271);
nor_1  g08895(new_n9203, new_n9202, new_n9272);
nand_1 g08896(new_n9225, new_n9206, new_n9273);
not_4  g08897(new_n9273, new_n9274);
xnor_1 g08898(new_n9274, new_n9272, new_n9275);
nand_1 g08899(new_n9275, new_n9271, new_n9276);
xnor_1 g08900(new_n9276, new_n9269, new_n9277);
xnor_1 g08901(new_n9277, new_n9243, new_n9278);
nand_1 g08902(n7965, n6441, new_n9279);
not_4  g08903(new_n9279, new_n9280);
xnor_1 g08904(new_n9242, new_n9226, new_n9281);
not_4  g08905(new_n9281, new_n9282);
nand_1 g08906(new_n9282, new_n9280, new_n9283);
nand_1 g08907(new_n9281, new_n9279, new_n9284);
xnor_1 g08908(new_n9234, new_n9232, new_n9285);
not_4  g08909(new_n9285, new_n9286);
nand_1 g08910(new_n8936, new_n8926, new_n9287);
not_4  g08911(new_n9287, new_n9288);
nand_1 g08912(new_n9288, new_n9286, new_n9289);
not_4  g08913(new_n9238, new_n9290);
xnor_1 g08914(new_n9240, new_n9290, new_n9291);
nor_1  g08915(new_n9291, new_n9289, new_n9292);
nand_1 g08916(new_n9292, new_n9284, new_n9293);
nand_1 g08917(new_n9293, new_n9283, new_n9294);
xnor_1 g08918(new_n9294, new_n9278, new_n9295);
not_4  g08919(new_n9295, new_n9296);
nand_1 g08920(n12777, n12648, new_n9297);
nand_1 g08921(n10545, n7159, new_n9298);
nand_1 g08922(n12489, n7690, new_n9299);
not_4  g08923(new_n9299, new_n9300);
xnor_1 g08924(new_n9300, new_n9298, new_n9301);
not_4  g08925(new_n9301, new_n9302);
xnor_1 g08926(new_n9302, new_n9297, new_n9303);
nand_1 g08927(n12489, n10545, new_n9304);
nand_1 g08928(new_n9304, new_n8916, new_n9305);
not_4  g08929(new_n9304, new_n9306);
nand_1 g08930(new_n9306, new_n8917, new_n9307);
nand_1 g08931(n12648, n7159, new_n9308);
nand_1 g08932(new_n9308, new_n9307, new_n9309);
nand_1 g08933(new_n9309, new_n9305, new_n9310);
xnor_1 g08934(new_n9310, new_n9303, new_n9311);
nand_1 g08935(n6254, n2530, new_n9312);
nand_1 g08936(n11967, n8476, new_n9313);
not_4  g08937(new_n9313, new_n9314);
xnor_1 g08938(new_n9314, new_n9312, new_n9315);
xnor_1 g08939(new_n9315, new_n9311, new_n9316);
nand_1 g08940(n8476, n6254, new_n9317);
nand_1 g08941(n12648, n12489, new_n9318);
nand_1 g08942(n12777, n8476, new_n9319);
nand_1 g08943(new_n9319, new_n9318, new_n9320);
not_4  g08944(new_n9318, new_n9321);
not_4  g08945(new_n9319, new_n9322);
nand_1 g08946(new_n9322, new_n9321, new_n9323);
nand_1 g08947(n7159, n2530, new_n9324);
nand_1 g08948(new_n9324, new_n9323, new_n9325);
nand_1 g08949(new_n9325, new_n9320, new_n9326);
nor_1  g08950(new_n9326, new_n9317, new_n9327);
not_4  g08951(new_n9327, new_n9328);
not_4  g08952(new_n9326, new_n9329);
xnor_1 g08953(new_n9329, new_n9317, new_n9330);
not_4  g08954(new_n9308, new_n9331);
nand_1 g08955(new_n9307, new_n9305, new_n9332);
xnor_1 g08956(new_n9332, new_n9331, new_n9333);
nand_1 g08957(new_n9333, new_n9330, new_n9334);
nand_1 g08958(new_n9334, new_n9328, new_n9335);
xnor_1 g08959(new_n9335, new_n9316, new_n9336);
nand_1 g08960(n11967, n5331, new_n9337);
not_4  g08961(new_n9337, new_n9338);
not_4  g08962(new_n9330, new_n9339);
xnor_1 g08963(new_n9333, new_n9339, new_n9340);
nor_1  g08964(new_n9340, new_n9338, new_n9341);
not_4  g08965(new_n9341, new_n9342);
xnor_1 g08966(new_n9340, new_n9337, new_n9343);
nand_1 g08967(n6254, n5331, new_n9344);
nand_1 g08968(new_n8918, new_n8910, new_n9345);
nand_1 g08969(new_n9345, new_n8915, new_n9346);
nor_1  g08970(new_n9346, new_n9344, new_n9347);
xnor_1 g08971(new_n9346, new_n9344, new_n9348);
nand_1 g08972(new_n9323, new_n9320, new_n9349);
xnor_1 g08973(new_n9349, new_n9324, new_n9350);
nor_1  g08974(new_n9350, new_n9348, new_n9351);
nor_1  g08975(new_n9351, new_n9347, new_n9352);
nand_1 g08976(new_n9352, new_n9343, new_n9353);
nand_1 g08977(new_n9353, new_n9342, new_n9354);
nor_1  g08978(new_n9354, new_n9336, new_n9355);
nand_1 g08979(n5331, n1353, new_n9356);
nand_1 g08980(n11967, n2530, new_n9357);
nand_1 g08981(n8476, n447, new_n9358);
not_4  g08982(new_n9358, new_n9359);
xnor_1 g08983(new_n9359, new_n9357, new_n9360);
xnor_1 g08984(new_n9360, new_n9356, new_n9361);
nor_1  g08985(new_n9302, new_n9297, new_n9362);
nor_1  g08986(new_n9310, new_n9303, new_n9363);
nor_1  g08987(new_n9363, new_n9362, new_n9364);
xnor_1 g08988(new_n9364, new_n9361, new_n9365);
not_4  g08989(new_n9298, new_n9366);
nand_1 g08990(new_n9300, new_n9366, new_n9367);
not_4  g08991(new_n9367, new_n9368);
nand_1 g08992(n12648, n6254, new_n9369);
not_4  g08993(new_n9369, new_n9370);
nand_1 g08994(new_n9370, new_n9368, new_n9371);
nand_1 g08995(new_n9369, new_n9367, new_n9372);
nand_1 g08996(new_n9372, new_n9371, new_n9373);
not_4  g08997(new_n9373, new_n9374);
nand_1 g08998(n7690, n7159, new_n9375);
nand_1 g08999(n12777, n10545, new_n9376);
nand_1 g09000(n12489, n3616, new_n9377);
not_4  g09001(new_n9377, new_n9378);
xnor_1 g09002(new_n9378, new_n9376, new_n9379);
xnor_1 g09003(new_n9379, new_n9375, new_n9380);
not_4  g09004(new_n9380, new_n9381);
xnor_1 g09005(new_n9381, new_n9374, new_n9382);
xnor_1 g09006(new_n9382, new_n9365, new_n9383);
not_4  g09007(new_n9311, new_n9384);
nand_1 g09008(new_n9315, new_n9384, new_n9385);
nor_1  g09009(new_n9313, new_n9312, new_n9386);
nand_1 g09010(new_n9335, new_n9316, new_n9387_1);
not_4  g09011(new_n9387_1, new_n9388);
xnor_1 g09012(new_n9388, new_n9386, new_n9389);
nand_1 g09013(new_n9389, new_n9385, new_n9390);
xnor_1 g09014(new_n9390, new_n9383, new_n9391);
xnor_1 g09015(new_n9391, new_n9355, new_n9392);
nand_1 g09016(n5331, n447, new_n9393);
not_4  g09017(new_n9393, new_n9394);
xnor_1 g09018(new_n9354, new_n9336, new_n9395);
not_4  g09019(new_n9395, new_n9396);
nand_1 g09020(new_n9396, new_n9394, new_n9397);
nand_1 g09021(new_n9395, new_n9393, new_n9398);
xnor_1 g09022(new_n9350, new_n9348, new_n9399);
not_4  g09023(new_n9399, new_n9400_1);
nand_1 g09024(new_n8921, new_n8911, new_n9401);
not_4  g09025(new_n9401, new_n9402);
nand_1 g09026(new_n9402, new_n9400_1, new_n9403);
not_4  g09027(new_n9352, new_n9404);
xnor_1 g09028(new_n9404, new_n9343, new_n9405);
nor_1  g09029(new_n9405, new_n9403, new_n9406);
nand_1 g09030(new_n9406, new_n9398, new_n9407);
nand_1 g09031(new_n9407, new_n9397, new_n9408);
xnor_1 g09032(new_n9408, new_n9392, new_n9409);
not_4  g09033(new_n9409, new_n9410);
xnor_1 g09034(new_n9410, new_n9296, new_n9411);
not_4  g09035(new_n9292, new_n9412);
nand_1 g09036(new_n9284, new_n9283, new_n9413);
xnor_1 g09037(new_n9413, new_n9412, new_n9414);
nand_1 g09038(new_n9398, new_n9397, new_n9415);
xnor_1 g09039(new_n9415, new_n9406, new_n9416);
not_4  g09040(new_n9416, new_n9417);
nand_1 g09041(new_n9417, new_n9414, new_n9418);
xnor_1 g09042(new_n9405, new_n9403, new_n9419);
not_4  g09043(new_n9291, new_n9420);
xnor_1 g09044(new_n9420, new_n9289, new_n9421);
not_4  g09045(new_n9421, new_n9422);
nand_1 g09046(new_n9422, new_n9419, new_n9423);
xnor_1 g09047(new_n9421, new_n9419, new_n9424);
xnor_1 g09048(new_n9401, new_n9400_1, new_n9425);
xnor_1 g09049(new_n9287, new_n9286, new_n9426);
nand_1 g09050(new_n9426, new_n9425, new_n9427);
nand_1 g09051(new_n8939, new_n8924, new_n9428);
nand_1 g09052(new_n8946, new_n9428, new_n9429);
xnor_1 g09053(new_n9426, new_n9425, new_n9430);
not_4  g09054(new_n9430, new_n9431);
nand_1 g09055(new_n9431, new_n9429, new_n9432);
nand_1 g09056(new_n9432, new_n9427, new_n9433);
not_4  g09057(new_n9433, new_n9434);
nand_1 g09058(new_n9434, new_n9424, new_n9435);
nand_1 g09059(new_n9435, new_n9423, new_n9436);
xnor_1 g09060(new_n9416, new_n9414, new_n9437);
nand_1 g09061(new_n9437, new_n9436, new_n9438);
nand_1 g09062(new_n9438, new_n9418, new_n9439);
xnor_1 g09063(new_n9439, new_n9411, new_n9440);
xnor_1 g09064(new_n9440, new_n9184, new_n9441);
xnor_1 g09065(new_n9141, new_n9139, new_n9442);
not_4  g09066(new_n9442, new_n9443);
not_4  g09067(new_n9437, new_n9444);
xnor_1 g09068(new_n9444, new_n9436, new_n9445);
nand_1 g09069(new_n9445, new_n9443, new_n9446);
xnor_1 g09070(new_n9445, new_n9442, new_n9447);
xnor_1 g09071(new_n9138, new_n9136, new_n9448);
not_4  g09072(new_n9448, new_n9449);
xnor_1 g09073(new_n9433, new_n9424, new_n9450);
nor_1  g09074(new_n9450, new_n9449, new_n9451);
not_4  g09075(new_n9451, new_n9452);
xnor_1 g09076(new_n9134, new_n9133, new_n9453);
xnor_1 g09077(new_n9430, new_n9429, new_n9454);
nand_1 g09078(new_n9454, new_n9453, new_n9455);
xnor_1 g09079(new_n9454, new_n9453, new_n9456);
not_4  g09080(new_n9456, new_n9457_1);
nand_1 g09081(new_n8907, new_n8893, new_n9458);
nand_1 g09082(new_n8950, new_n9458, new_n9459);
nand_1 g09083(new_n9459, new_n9457_1, new_n9460);
nand_1 g09084(new_n9460, new_n9455, new_n9461);
nand_1 g09085(new_n9450, new_n9449, new_n9462);
nand_1 g09086(new_n9462, new_n9452, new_n9463);
not_4  g09087(new_n9463, new_n9464);
nand_1 g09088(new_n9464, new_n9461, new_n9465);
nand_1 g09089(new_n9465, new_n9452, new_n9466);
not_4  g09090(new_n9466, new_n9467);
nand_1 g09091(new_n9467, new_n9447, new_n9468);
nand_1 g09092(new_n9468, new_n9446, new_n9469);
xnor_1 g09093(new_n9469, new_n9441, new_n9470);
nor_1  g09094(new_n9470, new_n9066, new_n9471);
xnor_1 g09095(new_n9470, new_n9065, new_n9472);
not_4  g09096(new_n9472, new_n9473);
xnor_1 g09097(new_n9062, new_n9061, new_n9474);
xnor_1 g09098(new_n9466, new_n9447, new_n9475);
nand_1 g09099(new_n9475, new_n9474, new_n9476);
not_4  g09100(new_n9474, new_n9477);
xnor_1 g09101(new_n9475, new_n9477, new_n9478);
xnor_1 g09102(new_n9060, new_n9059, new_n9479);
not_4  g09103(new_n9479, new_n9480);
xnor_1 g09104(new_n9463, new_n9461, new_n9481);
nor_1  g09105(new_n9481, new_n9480, new_n9482);
xnor_1 g09106(new_n9481, new_n9480, new_n9483);
xnor_1 g09107(new_n9057, new_n9056, new_n9484);
xnor_1 g09108(new_n9459, new_n9456, new_n9485);
nor_1  g09109(new_n9485, new_n9484, new_n9486);
nor_1  g09110(new_n8888, new_n8873, new_n9487);
nor_1  g09111(new_n8952, new_n8889, new_n9488);
nor_1  g09112(new_n9488, new_n9487, new_n9489);
not_4  g09113(new_n9489, new_n9490);
xnor_1 g09114(new_n9485, new_n9484, new_n9491);
nor_1  g09115(new_n9491, new_n9490, new_n9492);
nor_1  g09116(new_n9492, new_n9486, new_n9493);
nor_1  g09117(new_n9493, new_n9483, new_n9494);
nor_1  g09118(new_n9494, new_n9482, new_n9495);
not_4  g09119(new_n9495, new_n9496);
nand_1 g09120(new_n9496, new_n9478, new_n9497);
nand_1 g09121(new_n9497, new_n9476, new_n9498);
nor_1  g09122(new_n9498, new_n9473, new_n9499);
nor_1  g09123(new_n9499, new_n9471, new_n9500);
nand_1 g09124(new_n9440, new_n9184, new_n9501);
not_4  g09125(new_n9441, new_n9502);
nand_1 g09126(new_n9469, new_n9502, new_n9503);
nand_1 g09127(new_n9503, new_n9501, new_n9504);
nand_1 g09128(new_n9048, new_n9017, new_n9505);
not_4  g09129(new_n9049, new_n9506);
nand_1 g09130(new_n9064, new_n9506, new_n9507);
nand_1 g09131(new_n9507, new_n9505, new_n9508);
nand_1 g09132(new_n9037, new_n9036, new_n9509);
nand_1 g09133(new_n9039, new_n9034, new_n9510);
nand_1 g09134(new_n9510, new_n9509, new_n9511);
nand_1 g09135(new_n9024, new_n9023, new_n9512);
nand_1 g09136(new_n9026, new_n9022, new_n9513);
nand_1 g09137(new_n9513, new_n9512, new_n9514);
nand_1 g09138(n9725, n5964, new_n9515);
xnor_1 g09139(new_n9515, new_n9514, new_n9516);
xnor_1 g09140(new_n9516, new_n9511, new_n9517);
xnor_1 g09141(new_n9517, new_n9508, new_n9518);
not_4  g09142(new_n9145, new_n9519);
nand_1 g09143(new_n9182, new_n9519, new_n9520);
nand_1 g09144(new_n9183, new_n9143, new_n9521);
nand_1 g09145(new_n9521, new_n9520, new_n9522);
nand_1 g09146(new_n9391, new_n9355, new_n9523);
not_4  g09147(new_n9392, new_n9524);
nand_1 g09148(new_n9408, new_n9524, new_n9525);
nand_1 g09149(new_n9525, new_n9523, new_n9526);
xnor_1 g09150(new_n9526, new_n9522, new_n9527);
nand_1 g09151(new_n9277, new_n9243, new_n9528);
not_4  g09152(new_n9278, new_n9529);
nand_1 g09153(new_n9294, new_n9529, new_n9530);
nand_1 g09154(new_n9530, new_n9528, new_n9531);
not_4  g09155(new_n9361, new_n9532);
nand_1 g09156(new_n9364, new_n9532, new_n9533);
not_4  g09157(new_n9382, new_n9534);
nand_1 g09158(new_n9534, new_n9365, new_n9535);
nand_1 g09159(new_n9535, new_n9533, new_n9536);
not_4  g09160(new_n9150, new_n9537);
nand_1 g09161(new_n9156, new_n9537, new_n9538);
nand_1 g09162(new_n9538, new_n9155, new_n9539);
nand_1 g09163(n3986, n1478, new_n9540);
nand_1 g09164(n9241, n6429, new_n9541);
nand_1 g09165(n10022, n7965, new_n9542);
xnor_1 g09166(new_n9542, new_n9541, new_n9543);
xnor_1 g09167(new_n9543, new_n9540, new_n9544);
xnor_1 g09168(new_n9544, new_n9539, new_n9545);
xnor_1 g09169(new_n9545, new_n9536, new_n9546);
nand_1 g09170(new_n9377, new_n9376, new_n9547);
nand_1 g09171(new_n9379, new_n9375, new_n9548);
nand_1 g09172(new_n9548, new_n9547, new_n9549);
nand_1 g09173(new_n9263, new_n9259, new_n9550);
nand_1 g09174(new_n9550, new_n9261, new_n9551);
not_4  g09175(new_n9551, new_n9552);
nand_1 g09176(n11999, n7388, new_n9553);
not_4  g09177(new_n9553, new_n9554);
nand_1 g09178(new_n9554, new_n9552, new_n9555);
nand_1 g09179(new_n9554, new_n9279, new_n9556);
nand_1 g09180(new_n9556, new_n9551, new_n9557);
nand_1 g09181(new_n9557, new_n9555, new_n9558);
xnor_1 g09182(new_n9558, new_n9549, new_n9559);
nand_1 g09183(new_n9380, new_n9374, new_n9560);
nand_1 g09184(new_n9560, new_n9371, new_n9561);
not_4  g09185(new_n9248, new_n9562);
nand_1 g09186(new_n9251, new_n9562, new_n9563);
nand_1 g09187(new_n9563, new_n9254, new_n9564);
nand_1 g09188(n2530, n447, new_n9565);
nand_1 g09189(n12777, n7690, new_n9566);
nand_1 g09190(n8476, n1353, new_n9567);
xnor_1 g09191(new_n9567, new_n9566, new_n9568);
xnor_1 g09192(new_n9568, new_n9565, new_n9569);
xnor_1 g09193(new_n9569, new_n9564, new_n9570);
xnor_1 g09194(new_n9570, new_n9561, new_n9571_1);
xnor_1 g09195(new_n9571_1, new_n9559, new_n9572);
nand_1 g09196(n8759, n1198, new_n9573);
nand_1 g09197(n11728, n10510, new_n9574);
xnor_1 g09198(new_n9574, new_n9573, new_n9575);
nand_1 g09199(n12489, n4499, new_n9576);
nand_1 g09200(n10545, n6254, new_n9577);
xnor_1 g09201(new_n9577, new_n9576, new_n9578_1);
nand_1 g09202(n5331, n4436, new_n9579);
nand_1 g09203(n12947, n2393, new_n9580);
xnor_1 g09204(new_n9580, new_n9579, new_n9581);
xnor_1 g09205(new_n9581, new_n9578_1, new_n9582);
xnor_1 g09206(new_n9582, new_n9575, new_n9583_1);
nand_1 g09207(n12648, n11967, new_n9584);
not_4  g09208(new_n9584, new_n9585);
nand_1 g09209(n7159, n3616, new_n9586);
nand_1 g09210(n12709, n10644, new_n9587);
xnor_1 g09211(new_n9587, new_n9586, new_n9588);
xnor_1 g09212(new_n9588, new_n9585, new_n9589);
nand_1 g09213(n8819, n8276, new_n9590);
nand_1 g09214(n7730, n6776, new_n9591);
xnor_1 g09215(new_n9591, new_n9590, new_n9592);
xnor_1 g09216(new_n9592, new_n9589, new_n9593);
xnor_1 g09217(new_n9593, new_n9583_1, new_n9594);
xnor_1 g09218(new_n9594, new_n9572, new_n9595);
xnor_1 g09219(new_n9595, new_n9546, new_n9596);
nand_1 g09220(new_n9274, new_n9272, new_n9597);
not_4  g09221(new_n9269, new_n9598);
nand_1 g09222(new_n9276, new_n9598, new_n9599);
nand_1 g09223(new_n9599, new_n9597, new_n9600);
nand_1 g09224(n12705, n4370, new_n9601);
not_4  g09225(new_n9027, new_n9602);
nand_1 g09226(new_n9602, new_n9021, new_n9603);
nand_1 g09227(new_n9041, new_n9028, new_n9604);
nand_1 g09228(new_n9604, new_n9603, new_n9605);
not_4  g09229(new_n9264, new_n9606);
nand_1 g09230(new_n9267, new_n9606, new_n9607);
not_4  g09231(new_n9258, new_n9608);
nand_1 g09232(new_n9268, new_n9608, new_n9609);
nand_1 g09233(new_n9609, new_n9607, new_n9610);
xnor_1 g09234(new_n9610, new_n9605, new_n9611);
xnor_1 g09235(new_n9611, new_n9601, new_n9612);
xnor_1 g09236(new_n9612, new_n9600, new_n9613);
xnor_1 g09237(new_n9613, new_n9596, new_n9614);
xnor_1 g09238(new_n9614, new_n9531, new_n9615);
xnor_1 g09239(new_n9615, new_n9527, new_n9616);
xnor_1 g09240(new_n9616, new_n9518, new_n9617);
nand_1 g09241(new_n9410, new_n9296, new_n9618);
not_4  g09242(new_n9411, new_n9619);
nand_1 g09243(new_n9439, new_n9619, new_n9620);
nand_1 g09244(new_n9620, new_n9618, new_n9621);
nand_1 g09245(new_n9179, new_n9176, new_n9622);
not_4  g09246(new_n9173, new_n9623);
nand_1 g09247(new_n9181, new_n9623, new_n9624);
nand_1 g09248(new_n9624, new_n9622, new_n9625);
nand_1 g09249(n11407, n10547, new_n9626);
nand_1 g09250(n5320, n4312, new_n9627);
xnor_1 g09251(new_n9627, new_n9626, new_n9628);
nand_1 g09252(n12299, n8717, new_n9629);
nand_1 g09253(n5857, n5760, new_n9630);
xnor_1 g09254(new_n9630, new_n9629, new_n9631);
nand_1 g09255(n12025, n11877, new_n9632);
nand_1 g09256(n12000, n1097, new_n9633);
xnor_1 g09257(new_n9633, new_n9632, new_n9634);
xnor_1 g09258(new_n9634, new_n9631, new_n9635);
xnor_1 g09259(new_n9635, new_n9628, new_n9636);
nand_1 g09260(new_n9167, new_n9166, new_n9637_1);
nand_1 g09261(new_n9169, new_n9165, new_n9638);
nand_1 g09262(new_n9638, new_n9637_1, new_n9639);
nand_1 g09263(n10990, n45, new_n9640_1);
xnor_1 g09264(new_n9640_1, new_n9639, new_n9641);
xnor_1 g09265(new_n9641, new_n9636, new_n9642);
not_4  g09266(new_n9161, new_n9643);
nand_1 g09267(new_n9163, new_n9643, new_n9644);
nand_1 g09268(new_n9170, new_n9164, new_n9645);
nand_1 g09269(new_n9645, new_n9644, new_n9646);
nand_1 g09270(n7436, n2433, new_n9647);
xnor_1 g09271(new_n9647, new_n9646, new_n9648);
xnor_1 g09272(new_n9648, new_n9642, new_n9649);
nand_1 g09273(new_n9358, new_n9357, new_n9650);
nand_1 g09274(new_n9360, new_n9356, new_n9651);
nand_1 g09275(new_n9651, new_n9650, new_n9652);
not_4  g09276(new_n9158, new_n9653);
nor_1  g09277(new_n9653, new_n9149, new_n9654);
not_4  g09278(new_n9159, new_n9655);
nor_1  g09279(new_n9172, new_n9655, new_n9656);
nor_1  g09280(new_n9656, new_n9654, new_n9657);
xnor_1 g09281(new_n9657, new_n9652, new_n9658);
xnor_1 g09282(new_n9658, new_n9649, new_n9659);
xnor_1 g09283(new_n9659, new_n9625, new_n9660);
nand_1 g09284(new_n9388, new_n9386, new_n9661);
not_4  g09285(new_n9383, new_n9662);
nand_1 g09286(new_n9390, new_n9662, new_n9663);
nand_1 g09287(new_n9663, new_n9661, new_n9664);
nor_1  g09288(new_n9246, new_n9245, new_n9665);
nor_1  g09289(new_n9256, new_n9247, new_n9666);
nor_1  g09290(new_n9666, new_n9665, new_n9667);
nand_1 g09291(n11892, n6441, new_n9668);
nand_1 g09292(n11791, n5860, new_n9669);
xnor_1 g09293(new_n9669, new_n9668, new_n9670);
nand_1 g09294(n11257, n5212, new_n9671);
nand_1 g09295(n6604, n5305, new_n9672);
xnor_1 g09296(new_n9672, new_n9671, new_n9673);
xnor_1 g09297(new_n9673, new_n9670, new_n9674);
xnor_1 g09298(new_n9674, new_n9667, new_n9675);
xnor_1 g09299(new_n9675, new_n9664, new_n9676);
xnor_1 g09300(new_n9676, new_n9660, new_n9677);
nand_1 g09301(new_n9032, new_n9031, new_n9678);
not_4  g09302(new_n9033, new_n9679);
nand_1 g09303(new_n9040, new_n9679, new_n9680);
nand_1 g09304(new_n9680, new_n9678, new_n9681);
nor_1  g09305(new_n9045, new_n8986, new_n9682);
not_4  g09306(new_n9047, new_n9683);
nor_1  g09307(new_n9683, new_n9042, new_n9684);
nor_1  g09308(new_n9684, new_n9682, new_n9685);
xnor_1 g09309(new_n9685, new_n9681, new_n9686);
xnor_1 g09310(new_n9686, new_n9677, new_n9687);
xnor_1 g09311(new_n9687, new_n9621, new_n9688);
xnor_1 g09312(new_n9688, new_n9617, new_n9689);
xnor_1 g09313(new_n9689, new_n9504, new_n9690);
xnor_1 g09314(new_n9690, new_n9500, n3287);
xnor_1 g09315(new_n9496, new_n9478, n3339);
xnor_1 g09316(new_n4211, new_n4210, n3456);
nand_1 g09317(n6687, n4005, new_n9694);
not_4  g09318(new_n9694, new_n9695);
nand_1 g09319(n12720, n6770, new_n9696);
nand_1 g09320(n9920, n2509, new_n9697);
nand_1 g09321(n6038, n3627, new_n9698);
nand_1 g09322(new_n9698, new_n9697, new_n9699);
not_4  g09323(new_n9697, new_n9700);
not_4  g09324(new_n9698, new_n9701);
nand_1 g09325(new_n9701, new_n9700, new_n9702);
nand_1 g09326(new_n9702, new_n9699, new_n9703);
xnor_1 g09327(new_n9703, new_n9696, new_n9704);
nand_1 g09328(n9920, n6038, new_n9705);
nand_1 g09329(n12720, n4189, new_n9706_1);
nand_1 g09330(new_n9706_1, new_n9705, new_n9707);
nand_1 g09331(n6770, n2509, new_n9708);
not_4  g09332(new_n9706_1, new_n9709);
xnor_1 g09333(new_n9709, new_n9705, new_n9710);
nand_1 g09334(new_n9710, new_n9708, new_n9711);
nand_1 g09335(new_n9711, new_n9707, new_n9712);
xnor_1 g09336(new_n9712, new_n9704, new_n9713);
not_4  g09337(new_n9713, new_n9714);
nand_1 g09338(n2564, n2508, new_n9715);
not_4  g09339(new_n9715, new_n9716);
nand_1 g09340(n6770, n6038, new_n9717);
nand_1 g09341(n4189, n2509, new_n9718);
nand_1 g09342(new_n9718, new_n9717, new_n9719);
not_4  g09343(new_n9719, new_n9720);
nand_1 g09344(n12720, n2564, new_n9721);
not_4  g09345(new_n9721, new_n9722);
xnor_1 g09346(new_n9718, new_n9717, new_n9723);
nor_1  g09347(new_n9723, new_n9722, new_n9724);
nor_1  g09348(new_n9724, new_n9720, new_n9725_1);
nand_1 g09349(new_n9725_1, new_n9716, new_n9726);
xnor_1 g09350(new_n9710, new_n9708, new_n9727);
xnor_1 g09351(new_n9725_1, new_n9715, new_n9728);
nand_1 g09352(new_n9728, new_n9727, new_n9729);
nand_1 g09353(new_n9729, new_n9726, new_n9730);
nand_1 g09354(n2585, n2564, new_n9731);
nand_1 g09355(n4189, n2508, new_n9732);
xnor_1 g09356(new_n9732, new_n9731, new_n9733);
not_4  g09357(new_n9733, new_n9734);
xnor_1 g09358(new_n9734, new_n9730, new_n9735);
xnor_1 g09359(new_n9735, new_n9714, new_n9736);
nand_1 g09360(n6687, n2585, new_n9737);
not_4  g09361(new_n9737, new_n9738);
nand_1 g09362(n6687, n2508, new_n9739);
not_4  g09363(new_n9739, new_n9740);
not_4  g09364(new_n377, new_n9741);
nand_1 g09365(new_n9709, new_n9741, new_n9742);
nand_1 g09366(n6038, n4189, new_n9743);
nand_1 g09367(n12720, n6687, new_n9744);
nand_1 g09368(new_n9744, new_n9743, new_n9745);
nand_1 g09369(n2564, n2509, new_n9746);
not_4  g09370(new_n9746, new_n9747);
nand_1 g09371(new_n9747, new_n9745, new_n9748);
nand_1 g09372(new_n9748, new_n9742, new_n9749);
nand_1 g09373(new_n9749, new_n9740, new_n9750);
xnor_1 g09374(new_n9749, new_n9739, new_n9751);
xnor_1 g09375(new_n9723, new_n9722, new_n9752);
nand_1 g09376(new_n9752, new_n9751, new_n9753);
nand_1 g09377(new_n9753, new_n9750, new_n9754);
nor_1  g09378(new_n9754, new_n9738, new_n9755);
not_4  g09379(new_n9727, new_n9756_1);
xnor_1 g09380(new_n9728, new_n9756_1, new_n9757);
xnor_1 g09381(new_n9754, new_n9738, new_n9758);
nor_1  g09382(new_n9758, new_n9757, new_n9759);
nor_1  g09383(new_n9759, new_n9755, new_n9760);
nand_1 g09384(new_n9760, new_n9736, new_n9761);
not_4  g09385(new_n9761, new_n9762);
nor_1  g09386(new_n9760, new_n9736, new_n9763_1);
nor_1  g09387(new_n9763_1, new_n9762, new_n9764);
nand_1 g09388(new_n9764, new_n9695, new_n9765);
not_4  g09389(new_n9765, new_n9766);
xnor_1 g09390(new_n9752, new_n9751, new_n9767_1);
not_4  g09391(new_n9767_1, new_n9768);
nand_1 g09392(new_n9745, new_n9742, new_n9769);
not_4  g09393(new_n9769, new_n9770);
nand_1 g09394(n6687, n2509, new_n9771);
not_4  g09395(new_n9771, new_n9772);
nand_1 g09396(n6038, n2564, new_n9773);
not_4  g09397(new_n9773, new_n9774);
nand_1 g09398(new_n9774, new_n9772, new_n9775);
nor_1  g09399(new_n9775, new_n9770, new_n9776);
nand_1 g09400(new_n9776, new_n9768, new_n9777);
not_4  g09401(new_n9777, new_n9778);
xnor_1 g09402(new_n9758, new_n9757, new_n9779);
nand_1 g09403(new_n9779, new_n9778, new_n9780);
xnor_1 g09404(new_n9764, new_n9695, new_n9781);
nor_1  g09405(new_n9781, new_n9780, new_n9782);
nor_1  g09406(new_n9782, new_n9766, new_n9783);
not_4  g09407(new_n9783, new_n9784);
nand_1 g09408(new_n9703, new_n9696, new_n9785);
not_4  g09409(new_n9704, new_n9786);
nand_1 g09410(new_n9712, new_n9786, new_n9787);
nand_1 g09411(new_n9787, new_n9785, new_n9788);
nand_1 g09412(n4005, n2564, new_n9789);
nand_1 g09413(n4189, n2585, new_n9790);
nand_1 g09414(n12706, n6687, new_n9791);
xnor_1 g09415(new_n9791, new_n9790, new_n9792);
xnor_1 g09416(new_n9792, new_n9789, new_n9793);
xnor_1 g09417(new_n9793, new_n9788, new_n9794);
nand_1 g09418(n6770, n2508, new_n9795);
xnor_1 g09419(new_n9795, new_n9702, new_n9796);
nand_1 g09420(n3627, n2509, new_n9797);
nand_1 g09421(n12720, n9920, new_n9798);
not_4  g09422(new_n9798, new_n9799);
nand_1 g09423(n6038, n4516, new_n9800);
not_4  g09424(new_n9800, new_n9801);
nand_1 g09425(new_n9801, new_n9799, new_n9802);
nand_1 g09426(new_n9800, new_n9798, new_n9803);
nand_1 g09427(new_n9803, new_n9802, new_n9804);
xnor_1 g09428(new_n9804, new_n9797, new_n9805);
xnor_1 g09429(new_n9805, new_n9796, new_n9806);
xnor_1 g09430(new_n9806, new_n9794, new_n9807);
nand_1 g09431(new_n9734, new_n9730, new_n9808);
nor_1  g09432(new_n9732, new_n9731, new_n9809);
nor_1  g09433(new_n9735, new_n9713, new_n9810);
xnor_1 g09434(new_n9810, new_n9809, new_n9811);
nand_1 g09435(new_n9811, new_n9808, new_n9812);
xnor_1 g09436(new_n9812, new_n9807, new_n9813);
nand_1 g09437(new_n9813, new_n9762, new_n9814);
not_4  g09438(new_n9807, new_n9815);
xnor_1 g09439(new_n9812, new_n9815, new_n9816);
nand_1 g09440(new_n9816, new_n9761, new_n9817);
nand_1 g09441(new_n9817, new_n9814, new_n9818);
xnor_1 g09442(new_n9818, new_n9784, new_n9819);
not_4  g09443(new_n9819, new_n9820_1);
nand_1 g09444(n8336, n5105, new_n9821);
nand_1 g09445(n10928, n7500, new_n9822);
not_4  g09446(new_n9822, new_n9823);
nand_1 g09447(n8336, n1209, new_n9824);
nand_1 g09448(n7354, n6986, new_n9825);
nand_1 g09449(new_n9825, new_n9824, new_n9826);
nand_1 g09450(new_n9826, new_n9823, new_n9827);
nor_1  g09451(new_n9825, new_n9824, new_n9828);
not_4  g09452(new_n9828, new_n9829);
nand_1 g09453(new_n9829, new_n9827, new_n9830);
xnor_1 g09454(new_n9830, new_n9821, new_n9831);
nand_1 g09455(n7500, n6986, new_n9832);
not_4  g09456(new_n9832, new_n9833);
nand_1 g09457(n7354, n2226, new_n9834);
nand_1 g09458(n10928, n1209, new_n9835);
nand_1 g09459(new_n9835, new_n9834, new_n9836);
nor_1  g09460(new_n9835, new_n9834, new_n9837);
not_4  g09461(new_n9837, new_n9838);
nand_1 g09462(new_n9838, new_n9836, new_n9839);
xnor_1 g09463(new_n9839, new_n9833, new_n9840);
xnor_1 g09464(new_n9840, new_n9831, new_n9841);
not_4  g09465(new_n9841, new_n9842);
nand_1 g09466(new_n9829, new_n9826, new_n9843);
not_4  g09467(new_n9843, new_n9844);
nand_1 g09468(n10928, n7354, new_n9845);
not_4  g09469(new_n9845, new_n9846);
nand_1 g09470(n8336, n7500, new_n9847);
not_4  g09471(new_n9847, new_n9848);
nand_1 g09472(new_n9848, new_n9846, new_n9849);
nor_1  g09473(new_n9849, new_n9844, new_n9850);
nand_1 g09474(new_n9850, new_n9842, new_n9851);
not_4  g09475(new_n9851, new_n9852);
nand_1 g09476(n8336, n4141, new_n9853);
not_4  g09477(new_n9853, new_n9854);
not_4  g09478(new_n9821, new_n9855);
nand_1 g09479(new_n9830, new_n9855, new_n9856);
nand_1 g09480(new_n9840, new_n9831, new_n9857);
nand_1 g09481(new_n9857, new_n9856, new_n9858);
nor_1  g09482(new_n9858, new_n9854, new_n9859);
not_4  g09483(new_n9859, new_n9860);
nand_1 g09484(new_n9858, new_n9854, new_n9861);
nand_1 g09485(new_n9861, new_n9860, new_n9862);
not_4  g09486(new_n9862, new_n9863);
nand_1 g09487(n10928, n5105, new_n9864);
nand_1 g09488(new_n9838, new_n9832, new_n9865);
nand_1 g09489(new_n9865, new_n9836, new_n9866);
nor_1  g09490(new_n9866, new_n9864, new_n9867);
not_4  g09491(new_n9867, new_n9868);
nand_1 g09492(new_n9866, new_n9864, new_n9869);
nand_1 g09493(new_n9869, new_n9868, new_n9870);
not_4  g09494(new_n9870, new_n9871);
nand_1 g09495(n6986, n1209, new_n9872);
nand_1 g09496(n7354, n1094, new_n9873);
nand_1 g09497(n7500, n2226, new_n9874);
not_4  g09498(new_n9874, new_n9875);
xnor_1 g09499(new_n9875, new_n9873, new_n9876);
xnor_1 g09500(new_n9876, new_n9872, new_n9877);
nand_1 g09501(new_n9877, new_n9871, new_n9878);
not_4  g09502(new_n9877, new_n9879);
nand_1 g09503(new_n9879, new_n9870, new_n9880);
nand_1 g09504(new_n9880, new_n9878, new_n9881);
nand_1 g09505(new_n9881, new_n9863, new_n9882);
not_4  g09506(new_n9881, new_n9883);
nand_1 g09507(new_n9883, new_n9862, new_n9884);
nand_1 g09508(new_n9884, new_n9882, new_n9885);
nand_1 g09509(new_n9885, new_n9852, new_n9886);
nand_1 g09510(n8336, n4928, new_n9887);
nand_1 g09511(n2226, n1209, new_n9888);
nand_1 g09512(new_n9874, new_n9873, new_n9889);
nand_1 g09513(new_n9876, new_n9872, new_n9890);
nand_1 g09514(new_n9890, new_n9889, new_n9891);
not_4  g09515(new_n9891, new_n9892);
xnor_1 g09516(new_n9892, new_n9888, new_n9893);
nand_1 g09517(n7500, n1094, new_n9894);
nand_1 g09518(n10678, n7354, new_n9895);
nand_1 g09519(new_n9895, new_n9894, new_n9896);
not_4  g09520(new_n9894, new_n9897);
not_4  g09521(new_n9895, new_n9898);
nand_1 g09522(new_n9898, new_n9897, new_n9899);
nand_1 g09523(new_n9899, new_n9896, new_n9900);
xnor_1 g09524(new_n9900, new_n9893, new_n9901);
nand_1 g09525(n10928, n4141, new_n9902);
nand_1 g09526(n6986, n5105, new_n9903);
not_4  g09527(new_n9903, new_n9904);
xnor_1 g09528(new_n9904, new_n9902, new_n9905);
xnor_1 g09529(new_n9905, new_n9901, new_n9906);
nand_1 g09530(new_n9878, new_n9868, new_n9907);
xnor_1 g09531(new_n9907, new_n9906, new_n9908);
nand_1 g09532(new_n9882, new_n9860, new_n9909);
not_4  g09533(new_n9909, new_n9910);
xnor_1 g09534(new_n9910, new_n9908, new_n9911);
xnor_1 g09535(new_n9911, new_n9887, new_n9912);
xnor_1 g09536(new_n9912, new_n9886, new_n9913);
nand_1 g09537(n11222, n7294, new_n9914);
nand_1 g09538(n11222, n1980, new_n9915);
not_4  g09539(new_n9915, new_n9916);
nand_1 g09540(n8028, n5314, new_n9917);
not_4  g09541(new_n9917, new_n9918);
nand_1 g09542(new_n9918, new_n9916, new_n9919);
nand_1 g09543(new_n9917, new_n9915, new_n9920_1);
nand_1 g09544(n11153, n10848, new_n9921);
not_4  g09545(new_n9921, new_n9922);
nand_1 g09546(new_n9922, new_n9920_1, new_n9923);
nand_1 g09547(new_n9923, new_n9919, new_n9924);
xnor_1 g09548(new_n9924, new_n9914, new_n9925);
nand_1 g09549(n10848, n5314, new_n9926);
not_4  g09550(new_n9926, new_n9927);
nand_1 g09551(n8028, n996, new_n9928);
not_4  g09552(new_n9928, new_n9929);
nand_1 g09553(n11153, n1980, new_n9930);
not_4  g09554(new_n9930, new_n9931);
nand_1 g09555(new_n9931, new_n9929, new_n9932);
nand_1 g09556(new_n9930, new_n9928, new_n9933);
nand_1 g09557(new_n9933, new_n9932, new_n9934);
xnor_1 g09558(new_n9934, new_n9927, new_n9935);
nand_1 g09559(new_n9935, new_n9925, new_n9936);
not_4  g09560(new_n9936, new_n9937);
nor_1  g09561(new_n9935, new_n9925, new_n9938_1);
nor_1  g09562(new_n9938_1, new_n9937, new_n9939);
nand_1 g09563(new_n9920_1, new_n9919, new_n9940);
not_4  g09564(new_n9940, new_n9941);
nand_1 g09565(n11153, n8028, new_n9942);
not_4  g09566(new_n9942, new_n9943);
nand_1 g09567(n11222, n10848, new_n9944);
not_4  g09568(new_n9944, new_n9945);
nand_1 g09569(new_n9945, new_n9943, new_n9946);
nor_1  g09570(new_n9946, new_n9941, new_n9947);
nand_1 g09571(new_n9947, new_n9939, new_n9948);
not_4  g09572(new_n9914, new_n9949);
nand_1 g09573(new_n9924, new_n9949, new_n9950);
nand_1 g09574(new_n9936, new_n9950, new_n9951);
not_4  g09575(new_n9951, new_n9952);
nand_1 g09576(n12704, n11222, new_n9953);
not_4  g09577(new_n9953, new_n9954);
nand_1 g09578(n11153, n7294, new_n9955);
nand_1 g09579(new_n9932, new_n9926, new_n9956_1);
nand_1 g09580(new_n9956_1, new_n9933, new_n9957);
not_4  g09581(new_n9957, new_n9958);
xnor_1 g09582(new_n9958, new_n9955, new_n9959);
nand_1 g09583(n10848, n996, new_n9960);
not_4  g09584(new_n9960, new_n9961);
nand_1 g09585(n5314, n1980, new_n9962);
not_4  g09586(new_n9962, new_n9963);
nand_1 g09587(n8028, n5767, new_n9964);
not_4  g09588(new_n9964, new_n9965);
nand_1 g09589(new_n9965, new_n9963, new_n9966);
nand_1 g09590(new_n9964, new_n9962, new_n9967);
nand_1 g09591(new_n9967, new_n9966, new_n9968);
xnor_1 g09592(new_n9968, new_n9961, new_n9969);
nand_1 g09593(new_n9969, new_n9959, new_n9970);
not_4  g09594(new_n9970, new_n9971);
nor_1  g09595(new_n9969, new_n9959, new_n9972);
nor_1  g09596(new_n9972, new_n9971, new_n9973);
nor_1  g09597(new_n9973, new_n9954, new_n9974);
not_4  g09598(new_n9974, new_n9975);
nand_1 g09599(new_n9973, new_n9954, new_n9976);
nand_1 g09600(new_n9976, new_n9975, new_n9977);
xnor_1 g09601(new_n9977, new_n9952, new_n9978);
nor_1  g09602(new_n9978, new_n9948, new_n9979);
nand_1 g09603(n11222, n5814, new_n9980);
nand_1 g09604(n1980, n996, new_n9981);
not_4  g09605(new_n9981, new_n9982);
nand_1 g09606(n8028, n5319, new_n9983);
nand_1 g09607(n10848, n5767, new_n9984);
not_4  g09608(new_n9984, new_n9985);
xnor_1 g09609(new_n9985, new_n9983, new_n9986);
xnor_1 g09610(new_n9986, new_n9982, new_n9987);
nand_1 g09611(new_n9966, new_n9960, new_n9988);
nand_1 g09612(new_n9988, new_n9967, new_n9989);
nor_1  g09613(new_n9989, new_n9987, new_n9990);
not_4  g09614(new_n9990, new_n9991);
nand_1 g09615(new_n9989, new_n9987, new_n9992);
nand_1 g09616(new_n9992, new_n9991, new_n9993);
nand_1 g09617(n12704, n11153, new_n9994);
nand_1 g09618(n7294, n5314, new_n9995);
not_4  g09619(new_n9995, new_n9996);
xnor_1 g09620(new_n9996, new_n9994, new_n9997);
xnor_1 g09621(new_n9997, new_n9993, new_n9998);
nor_1  g09622(new_n9957, new_n9955, new_n9999);
nor_1  g09623(new_n9971, new_n9999, new_n10000);
xnor_1 g09624(new_n10000, new_n9998, new_n10001);
nor_1  g09625(new_n9977, new_n9951, new_n10002);
nor_1  g09626(new_n10002, new_n9974, new_n10003);
nand_1 g09627(new_n10003, new_n10001, new_n10004);
not_4  g09628(new_n10000, new_n10005);
xnor_1 g09629(new_n10005, new_n9998, new_n10006);
not_4  g09630(new_n10003, new_n10007);
nand_1 g09631(new_n10007, new_n10006, new_n10008);
nand_1 g09632(new_n10008, new_n10004, new_n10009);
not_4  g09633(new_n10009, new_n10010);
xnor_1 g09634(new_n10010, new_n9980, new_n10011);
xnor_1 g09635(new_n10011, new_n9979, new_n10012);
nand_1 g09636(n12069, n2802, new_n10013);
nand_1 g09637(n7891, n1564, new_n10014);
nand_1 g09638(n12069, n533, new_n10015);
nand_1 g09639(new_n10015, new_n10014, new_n10016);
nand_1 g09640(n12391, n1512, new_n10017);
not_4  g09641(new_n10017, new_n10018);
nand_1 g09642(new_n10018, new_n10016, new_n10019);
not_4  g09643(new_n10014, new_n10020);
not_4  g09644(new_n10015, new_n10021);
nand_1 g09645(new_n10021, new_n10020, new_n10022_1);
nand_1 g09646(new_n10022_1, new_n10019, new_n10023);
xnor_1 g09647(new_n10023, new_n10013, new_n10024);
nand_1 g09648(n7891, n1512, new_n10025);
nand_1 g09649(n7160, n1564, new_n10026);
nand_1 g09650(n12391, n533, new_n10027);
nand_1 g09651(new_n10027, new_n10026, new_n10028);
not_4  g09652(new_n10026, new_n10029);
not_4  g09653(new_n10027, new_n10030);
nand_1 g09654(new_n10030, new_n10029, new_n10031);
nand_1 g09655(new_n10031, new_n10028, new_n10032);
xnor_1 g09656(new_n10032, new_n10025, new_n10033);
xnor_1 g09657(new_n10033, new_n10024, new_n10034);
nand_1 g09658(new_n10022_1, new_n10016, new_n10035);
not_4  g09659(new_n10035, new_n10036);
nand_1 g09660(n12391, n1564, new_n10037);
not_4  g09661(new_n10037, new_n10038);
nand_1 g09662(n12069, n1512, new_n10039);
not_4  g09663(new_n10039, new_n10040);
nand_1 g09664(new_n10040, new_n10038, new_n10041);
nor_1  g09665(new_n10041, new_n10036, new_n10042);
nand_1 g09666(new_n10042, new_n10034, new_n10043);
not_4  g09667(new_n10043, new_n10044);
nand_1 g09668(n12069, n6806, new_n10045);
not_4  g09669(new_n10045, new_n10046);
nand_1 g09670(n12391, n2802, new_n10047);
not_4  g09671(new_n10047, new_n10048);
nor_1  g09672(new_n10030, new_n10029, new_n10049);
not_4  g09673(new_n10025, new_n10050);
nor_1  g09674(new_n10032, new_n10050, new_n10051);
nor_1  g09675(new_n10051, new_n10049, new_n10052);
nand_1 g09676(new_n10052, new_n10048, new_n10053);
nor_1  g09677(new_n10027, new_n10026, new_n10054);
nor_1  g09678(new_n10054, new_n10049, new_n10055);
nand_1 g09679(new_n10055, new_n10025, new_n10056);
nand_1 g09680(new_n10056, new_n10028, new_n10057);
nand_1 g09681(new_n10057, new_n10047, new_n10058);
nand_1 g09682(new_n10058, new_n10053, new_n10059);
nand_1 g09683(n7891, n533, new_n10060);
nand_1 g09684(n4828, n1564, new_n10061);
nand_1 g09685(n7160, n1512, new_n10062);
not_4  g09686(new_n10062, new_n10063);
xnor_1 g09687(new_n10063, new_n10061, new_n10064);
xnor_1 g09688(new_n10064, new_n10060, new_n10065);
not_4  g09689(new_n10065, new_n10066);
nor_1  g09690(new_n10066, new_n10059, new_n10067);
nor_1  g09691(new_n10057, new_n10047, new_n10068);
nor_1  g09692(new_n10052, new_n10048, new_n10069);
nor_1  g09693(new_n10069, new_n10068, new_n10070);
nor_1  g09694(new_n10065, new_n10070, new_n10071);
nor_1  g09695(new_n10071, new_n10067, new_n10072);
nor_1  g09696(new_n10072, new_n10046, new_n10073);
nand_1 g09697(new_n10065, new_n10070, new_n10074);
nand_1 g09698(new_n10066, new_n10059, new_n10075);
nand_1 g09699(new_n10075, new_n10074, new_n10076);
nor_1  g09700(new_n10076, new_n10045, new_n10077);
nor_1  g09701(new_n10077, new_n10073, new_n10078);
not_4  g09702(new_n10013, new_n10079);
nand_1 g09703(new_n10023, new_n10079, new_n10080);
not_4  g09704(new_n10033, new_n10081);
nand_1 g09705(new_n10081, new_n10024, new_n10082);
nand_1 g09706(new_n10082, new_n10080, new_n10083);
not_4  g09707(new_n10083, new_n10084);
nand_1 g09708(new_n10084, new_n10078, new_n10085);
nand_1 g09709(new_n10076, new_n10045, new_n10086);
nand_1 g09710(new_n10072, new_n10046, new_n10087);
nand_1 g09711(new_n10087, new_n10086, new_n10088);
nand_1 g09712(new_n10083, new_n10088, new_n10089);
nand_1 g09713(new_n10089, new_n10085, new_n10090);
nand_1 g09714(new_n10090, new_n10044, new_n10091);
not_4  g09715(new_n10091, new_n10092);
nand_1 g09716(n12069, n5069, new_n10093);
nand_1 g09717(n7160, n533, new_n10094);
not_4  g09718(new_n10094, new_n10095);
nand_1 g09719(n2515, n1564, new_n10096);
nand_1 g09720(n4828, n1512, new_n10097);
not_4  g09721(new_n10097, new_n10098);
xnor_1 g09722(new_n10098, new_n10096, new_n10099);
xnor_1 g09723(new_n10099, new_n10095, new_n10100);
nand_1 g09724(new_n10062, new_n10061, new_n10101);
nand_1 g09725(new_n10064, new_n10060, new_n10102);
nand_1 g09726(new_n10102, new_n10101, new_n10103);
nor_1  g09727(new_n10103, new_n10100, new_n10104);
not_4  g09728(new_n10104, new_n10105);
nand_1 g09729(new_n10103, new_n10100, new_n10106);
nand_1 g09730(new_n10106, new_n10105, new_n10107);
nand_1 g09731(n7891, n2802, new_n10108);
nand_1 g09732(n12391, n6806, new_n10109);
not_4  g09733(new_n10109, new_n10110);
xnor_1 g09734(new_n10110, new_n10108, new_n10111);
xnor_1 g09735(new_n10111, new_n10107, new_n10112);
nand_1 g09736(new_n10074, new_n10053, new_n10113);
xnor_1 g09737(new_n10113, new_n10112, new_n10114);
not_4  g09738(new_n10114, new_n10115);
nor_1  g09739(new_n10083, new_n10088, new_n10116);
nor_1  g09740(new_n10116, new_n10073, new_n10117);
nand_1 g09741(new_n10117, new_n10115, new_n10118);
nand_1 g09742(new_n10085, new_n10086, new_n10119);
nand_1 g09743(new_n10119, new_n10114, new_n10120);
nand_1 g09744(new_n10120, new_n10118, new_n10121);
nand_1 g09745(new_n10121, new_n10093, new_n10122);
not_4  g09746(new_n10093, new_n10123);
nor_1  g09747(new_n10119, new_n10114, new_n10124);
nor_1  g09748(new_n10117, new_n10115, new_n10125);
nor_1  g09749(new_n10125, new_n10124, new_n10126);
nand_1 g09750(new_n10126, new_n10123, new_n10127);
nand_1 g09751(new_n10127, new_n10122, new_n10128);
nor_1  g09752(new_n10128, new_n10092, new_n10129);
nor_1  g09753(new_n10126, new_n10123, new_n10130);
nor_1  g09754(new_n10121, new_n10093, new_n10131);
nor_1  g09755(new_n10131, new_n10130, new_n10132);
nor_1  g09756(new_n10132, new_n10091, new_n10133);
nor_1  g09757(new_n10133, new_n10129, new_n10134);
nand_1 g09758(new_n10134, new_n10012, new_n10135);
not_4  g09759(new_n10012, new_n10136);
nand_1 g09760(new_n10132, new_n10091, new_n10137);
nand_1 g09761(new_n10128, new_n10092, new_n10138);
nand_1 g09762(new_n10138, new_n10137, new_n10139);
nand_1 g09763(new_n10139, new_n10136, new_n10140);
nand_1 g09764(new_n10140, new_n10135, new_n10141);
not_4  g09765(new_n9978, new_n10142);
xnor_1 g09766(new_n10142, new_n9948, new_n10143);
not_4  g09767(new_n10143, new_n10144);
xnor_1 g09768(new_n10042, new_n10034, new_n10145);
xnor_1 g09769(new_n9947, new_n9939, new_n10146);
nand_1 g09770(new_n10146, new_n10145, new_n10147);
nand_1 g09771(new_n10018, new_n381_1, new_n10148);
nand_1 g09772(new_n10148, new_n10035, new_n10149);
nor_1  g09773(new_n10019, new_n382, new_n10150);
not_4  g09774(new_n10150, new_n10151);
nand_1 g09775(new_n10151, new_n10149, new_n10152);
nand_1 g09776(new_n9922, new_n379, new_n10153);
nand_1 g09777(new_n10153, new_n9940, new_n10154);
not_4  g09778(new_n10153, new_n10155);
nand_1 g09779(new_n10155, new_n9920_1, new_n10156);
nand_1 g09780(new_n10156, new_n10154, new_n10157);
nor_1  g09781(new_n10157, new_n10152, new_n10158);
nand_1 g09782(new_n9944, new_n9942, new_n10159);
nand_1 g09783(new_n10159, new_n9946, new_n10160);
nand_1 g09784(new_n10160, new_n383, new_n10161);
xnor_1 g09785(new_n10160, new_n383, new_n10162);
not_4  g09786(new_n10162, new_n10163);
nand_1 g09787(new_n10039, new_n10037, new_n10164);
nand_1 g09788(new_n10164, new_n10041, new_n10165);
nand_1 g09789(new_n10165, new_n10163, new_n10166);
nand_1 g09790(new_n10166, new_n10161, new_n10167);
xnor_1 g09791(new_n10157, new_n10152, new_n10168);
nor_1  g09792(new_n10168, new_n10167, new_n10169);
nor_1  g09793(new_n10169, new_n10158, new_n10170);
not_4  g09794(new_n10145, new_n10171);
xnor_1 g09795(new_n10146, new_n10171, new_n10172);
nand_1 g09796(new_n10172, new_n10170, new_n10173);
nand_1 g09797(new_n10173, new_n10147, new_n10174_1);
nand_1 g09798(new_n10174_1, new_n10144, new_n10175);
xnor_1 g09799(new_n10090, new_n10043, new_n10176);
not_4  g09800(new_n10176, new_n10177);
xnor_1 g09801(new_n10174_1, new_n10143, new_n10178);
nand_1 g09802(new_n10178, new_n10177, new_n10179);
nand_1 g09803(new_n10179, new_n10175, new_n10180);
xnor_1 g09804(new_n10180, new_n10141, new_n10181);
nor_1  g09805(new_n10181, new_n9913, new_n10182);
not_4  g09806(new_n10182, new_n10183);
not_4  g09807(new_n10181, new_n10184);
xnor_1 g09808(new_n10184, new_n9913, new_n10185);
xnor_1 g09809(new_n9885, new_n9851, new_n10186);
not_4  g09810(new_n10186, new_n10187);
xnor_1 g09811(new_n10178, new_n10176, new_n10188);
nor_1  g09812(new_n10188, new_n10187, new_n10189);
xnor_1 g09813(new_n10188, new_n10187, new_n10190);
xnor_1 g09814(new_n9850, new_n9841, new_n10191);
not_4  g09815(new_n10191, new_n10192);
not_4  g09816(new_n10172, new_n10193);
xnor_1 g09817(new_n10193, new_n10170, new_n10194);
nor_1  g09818(new_n10194, new_n10192, new_n10195);
not_4  g09819(new_n10195, new_n10196);
xnor_1 g09820(new_n10194, new_n10191, new_n10197);
xnor_1 g09821(new_n10168, new_n10167, new_n10198);
nand_1 g09822(new_n9823, new_n378, new_n10199);
nor_1  g09823(new_n10199, new_n9826, new_n10200);
not_4  g09824(new_n10200, new_n10201);
nand_1 g09825(new_n10199, new_n9844, new_n10202);
nand_1 g09826(new_n10202, new_n10201, new_n10203);
not_4  g09827(new_n10203, new_n10204);
nand_1 g09828(new_n10204, new_n10198, new_n10205);
xnor_1 g09829(new_n10203, new_n10198, new_n10206);
xnor_1 g09830(new_n10165, new_n10162, new_n10207);
not_4  g09831(new_n10207, new_n10208);
nand_1 g09832(new_n9847, new_n9845, new_n10209);
nand_1 g09833(new_n10209, new_n9849, new_n10210);
not_4  g09834(new_n10210, new_n10211);
nand_1 g09835(new_n10211, new_n10208, new_n10212);
not_4  g09836(new_n378, new_n10213);
nand_1 g09837(new_n386, new_n10213, new_n10214);
not_4  g09838(new_n10214, new_n10215);
xnor_1 g09839(new_n10210, new_n10208, new_n10216);
nand_1 g09840(new_n10216, new_n10215, new_n10217_1);
nand_1 g09841(new_n10217_1, new_n10212, new_n10218);
not_4  g09842(new_n10218, new_n10219);
nand_1 g09843(new_n10219, new_n10206, new_n10220);
nand_1 g09844(new_n10220, new_n10205, new_n10221);
not_4  g09845(new_n10221, new_n10222);
nand_1 g09846(new_n10222, new_n10197, new_n10223_1);
nand_1 g09847(new_n10223_1, new_n10196, new_n10224);
not_4  g09848(new_n10224, new_n10225);
nor_1  g09849(new_n10225, new_n10190, new_n10226);
nor_1  g09850(new_n10226, new_n10189, new_n10227);
not_4  g09851(new_n10227, new_n10228);
nand_1 g09852(new_n10228, new_n10185, new_n10229);
nand_1 g09853(new_n10229, new_n10183, new_n10230);
nand_1 g09854(new_n9910, new_n9908, new_n10231);
nor_1  g09855(new_n9891, new_n9888, new_n10232);
not_4  g09856(new_n10232, new_n10233);
not_4  g09857(new_n9900, new_n10234);
nand_1 g09858(new_n10234, new_n9893, new_n10235);
nand_1 g09859(new_n10235, new_n10233, new_n10236);
not_4  g09860(new_n10236, new_n10237);
nand_1 g09861(n10928, n4928, new_n10238);
nand_1 g09862(n6986, n4141, new_n10239);
nand_1 g09863(n8336, n8236, new_n10240);
not_4  g09864(new_n10240, new_n10241);
xnor_1 g09865(new_n10241, new_n10239, new_n10242);
xnor_1 g09866(new_n10242, new_n10238, new_n10243);
xnor_1 g09867(new_n10243, new_n10237, new_n10244);
not_4  g09868(new_n9899, new_n10245);
nand_1 g09869(n5105, n2226, new_n10246);
not_4  g09870(new_n10246, new_n10247);
nand_1 g09871(new_n10247, new_n10245, new_n10248);
nand_1 g09872(new_n10246, new_n9899, new_n10249);
nand_1 g09873(new_n10249, new_n10248, new_n10250);
nand_1 g09874(n10678, n7500, new_n10251);
nand_1 g09875(n7354, n7320, new_n10252);
nand_1 g09876(n1209, n1094, new_n10253);
not_4  g09877(new_n10253, new_n10254);
xnor_1 g09878(new_n10254, new_n10252, new_n10255);
xnor_1 g09879(new_n10255, new_n10251, new_n10256);
xnor_1 g09880(new_n10256, new_n10250, new_n10257);
xnor_1 g09881(new_n10257, new_n10244, new_n10258);
nand_1 g09882(new_n9905, new_n9901, new_n10259);
nor_1  g09883(new_n9903, new_n9902, new_n10260);
not_4  g09884(new_n9906, new_n10261);
nand_1 g09885(new_n9907, new_n10261, new_n10262);
not_4  g09886(new_n10262, new_n10263);
xnor_1 g09887(new_n10263, new_n10260, new_n10264);
nand_1 g09888(new_n10264, new_n10259, new_n10265);
xnor_1 g09889(new_n10265, new_n10258, new_n10266);
xnor_1 g09890(new_n10266, new_n10231, new_n10267);
nand_1 g09891(new_n9911, new_n9887, new_n10268);
not_4  g09892(new_n9912, new_n10269);
nand_1 g09893(new_n10269, new_n9886, new_n10270);
nand_1 g09894(new_n10270, new_n10268, new_n10271);
xnor_1 g09895(new_n10271, new_n10267, new_n10272);
not_4  g09896(new_n10272, new_n10273);
nand_1 g09897(new_n9986, new_n9982, new_n10274);
nand_1 g09898(new_n9991, new_n10274, new_n10275);
nand_1 g09899(n11153, n5814, new_n10276);
not_4  g09900(new_n10276, new_n10277);
nand_1 g09901(n12704, n5314, new_n10278_1);
nand_1 g09902(n11222, n4903, new_n10279);
not_4  g09903(new_n10279, new_n10280);
xnor_1 g09904(new_n10280, new_n10278_1, new_n10281);
xnor_1 g09905(new_n10281, new_n10277, new_n10282);
xnor_1 g09906(new_n10282, new_n10275, new_n10283);
not_4  g09907(new_n9983, new_n10284);
nand_1 g09908(new_n9985, new_n10284, new_n10285);
not_4  g09909(new_n10285, new_n10286);
nand_1 g09910(n7294, n996, new_n10287);
not_4  g09911(new_n10287, new_n10288);
nand_1 g09912(new_n10288, new_n10286, new_n10289);
nand_1 g09913(new_n10287, new_n10285, new_n10290);
nand_1 g09914(new_n10290, new_n10289, new_n10291);
not_4  g09915(new_n10291, new_n10292);
nand_1 g09916(n10848, n5319, new_n10293);
nand_1 g09917(n5767, n1980, new_n10294);
nand_1 g09918(n9457, n8028, new_n10295);
not_4  g09919(new_n10295, new_n10296);
xnor_1 g09920(new_n10296, new_n10294, new_n10297);
xnor_1 g09921(new_n10297, new_n10293, new_n10298);
not_4  g09922(new_n10298, new_n10299);
xnor_1 g09923(new_n10299, new_n10292, new_n10300);
xnor_1 g09924(new_n10300, new_n10283, new_n10301);
not_4  g09925(new_n9993, new_n10302);
nand_1 g09926(new_n9997, new_n10302, new_n10303);
nor_1  g09927(new_n9995, new_n9994, new_n10304);
nand_1 g09928(new_n10005, new_n9998, new_n10305);
not_4  g09929(new_n10305, new_n10306);
xnor_1 g09930(new_n10306, new_n10304, new_n10307);
nand_1 g09931(new_n10307, new_n10303, new_n10308);
xnor_1 g09932(new_n10308, new_n10301, new_n10309);
xnor_1 g09933(new_n10309, new_n10004, new_n10310);
not_4  g09934(new_n9980, new_n10311);
nand_1 g09935(new_n10010, new_n10311, new_n10312);
nand_1 g09936(new_n10011, new_n9979, new_n10313);
nand_1 g09937(new_n10313, new_n10312, new_n10314);
xnor_1 g09938(new_n10314, new_n10310, new_n10315);
not_4  g09939(new_n10315, new_n10316);
not_4  g09940(new_n10107, new_n10317);
nand_1 g09941(new_n10111, new_n10317, new_n10318);
nor_1  g09942(new_n10109, new_n10108, new_n10319);
nand_1 g09943(new_n10113, new_n10112, new_n10320);
not_4  g09944(new_n10320, new_n10321);
xnor_1 g09945(new_n10321, new_n10319, new_n10322);
nand_1 g09946(new_n10322, new_n10318, new_n10323);
not_4  g09947(new_n10096, new_n10324);
nand_1 g09948(new_n10098, new_n10324, new_n10325);
not_4  g09949(new_n10325, new_n10326);
nand_1 g09950(n7160, n2802, new_n10327_1);
not_4  g09951(new_n10327_1, new_n10328);
nand_1 g09952(new_n10328, new_n10326, new_n10329);
nand_1 g09953(new_n10327_1, new_n10325, new_n10330);
nand_1 g09954(new_n10330, new_n10329, new_n10331);
nand_1 g09955(n2515, n1512, new_n10332);
nand_1 g09956(n1564, n1199, new_n10333);
nand_1 g09957(n4828, n533, new_n10334);
nand_1 g09958(new_n10334, new_n10333, new_n10335);
not_4  g09959(new_n10333, new_n10336);
not_4  g09960(new_n10334, new_n10337);
nand_1 g09961(new_n10337, new_n10336, new_n10338);
nand_1 g09962(new_n10338, new_n10335, new_n10339);
xnor_1 g09963(new_n10339, new_n10332, new_n10340);
not_4  g09964(new_n10340, new_n10341);
xnor_1 g09965(new_n10341, new_n10331, new_n10342);
nand_1 g09966(new_n10099, new_n10095, new_n10343);
nand_1 g09967(new_n10105, new_n10343, new_n10344);
nand_1 g09968(n12391, n5069, new_n10345);
not_4  g09969(new_n10345, new_n10346);
nand_1 g09970(n7891, n6806, new_n10347);
nand_1 g09971(n12069, n12044, new_n10348);
not_4  g09972(new_n10348, new_n10349);
xnor_1 g09973(new_n10349, new_n10347, new_n10350);
xnor_1 g09974(new_n10350, new_n10346, new_n10351);
xnor_1 g09975(new_n10351, new_n10344, new_n10352);
xnor_1 g09976(new_n10352, new_n10342, new_n10353);
xnor_1 g09977(new_n10353, new_n10323, new_n10354);
xnor_1 g09978(new_n10354, new_n10118, new_n10355);
nand_1 g09979(new_n10122, new_n10092, new_n10356);
nand_1 g09980(new_n10356, new_n10127, new_n10357);
xnor_1 g09981(new_n10357, new_n10355, new_n10358);
nor_1  g09982(new_n10139, new_n10136, new_n10359);
nor_1  g09983(new_n10134, new_n10012, new_n10360);
nor_1  g09984(new_n10360, new_n10359, new_n10361);
nand_1 g09985(new_n10180, new_n10361, new_n10362);
nand_1 g09986(new_n10362, new_n10135, new_n10363);
nand_1 g09987(new_n10363, new_n10358, new_n10364);
not_4  g09988(new_n10358, new_n10365);
not_4  g09989(new_n10180, new_n10366);
nor_1  g09990(new_n10366, new_n10141, new_n10367);
nor_1  g09991(new_n10367, new_n10359, new_n10368);
nand_1 g09992(new_n10368, new_n10365, new_n10369);
nand_1 g09993(new_n10369, new_n10364, new_n10370);
nor_1  g09994(new_n10370, new_n10316, new_n10371);
nor_1  g09995(new_n10368, new_n10365, new_n10372);
nor_1  g09996(new_n10363, new_n10358, new_n10373);
nor_1  g09997(new_n10373, new_n10372, new_n10374);
nor_1  g09998(new_n10374, new_n10315, new_n10375);
nor_1  g09999(new_n10375, new_n10371, new_n10376);
nand_1 g10000(new_n10376, new_n10273, new_n10377);
nand_1 g10001(new_n10374, new_n10315, new_n10378);
nand_1 g10002(new_n10370, new_n10316, new_n10379);
nand_1 g10003(new_n10379, new_n10378, new_n10380);
nand_1 g10004(new_n10380, new_n10272, new_n10381);
nand_1 g10005(new_n10381, new_n10377, new_n10382);
nor_1  g10006(new_n10382, new_n10230, new_n10383);
not_4  g10007(new_n10230, new_n10384);
nor_1  g10008(new_n10380, new_n10272, new_n10385);
nor_1  g10009(new_n10376, new_n10273, new_n10386);
nor_1  g10010(new_n10386, new_n10385, new_n10387);
nor_1  g10011(new_n10387, new_n10384, new_n10388);
nor_1  g10012(new_n10388, new_n10383, new_n10389);
nand_1 g10013(new_n10389, new_n9820_1, new_n10390);
not_4  g10014(new_n9782, new_n10391_1);
nand_1 g10015(new_n9781, new_n9780, new_n10392);
nand_1 g10016(new_n10392, new_n10391_1, new_n10393);
not_4  g10017(new_n10393, new_n10394);
not_4  g10018(new_n9779, new_n10395);
xnor_1 g10019(new_n10395, new_n9778, new_n10396);
xnor_1 g10020(new_n10224, new_n10190, new_n10397);
nor_1  g10021(new_n10397, new_n10396, new_n10398);
xnor_1 g10022(new_n9776, new_n9767_1, new_n10399);
xnor_1 g10023(new_n10221, new_n10197, new_n10400);
nor_1  g10024(new_n10400, new_n10399, new_n10401);
not_4  g10025(new_n10401, new_n10402);
not_4  g10026(new_n10400, new_n10403);
xnor_1 g10027(new_n10403, new_n10399, new_n10404);
xnor_1 g10028(new_n10218, new_n10206, new_n10405);
nand_1 g10029(new_n9747, new_n377, new_n10406);
nand_1 g10030(new_n10406, new_n9769, new_n10407);
not_4  g10031(new_n10406, new_n10408);
nand_1 g10032(new_n10408, new_n9745, new_n10409);
nand_1 g10033(new_n10409, new_n10407, new_n10410);
nand_1 g10034(new_n10410, new_n10405, new_n10411);
xnor_1 g10035(new_n10410, new_n10405, new_n10412);
nand_1 g10036(new_n387, new_n9741, new_n10413);
nand_1 g10037(new_n9773, new_n9771, new_n10414);
nand_1 g10038(new_n10414, new_n9775, new_n10415);
nand_1 g10039(new_n10415, new_n10413, new_n10416);
xnor_1 g10040(new_n10216, new_n10214, new_n10417);
xnor_1 g10041(new_n10415, new_n10413, new_n10418);
nor_1  g10042(new_n10418, new_n10417, new_n10419);
not_4  g10043(new_n10419, new_n10420);
nand_1 g10044(new_n10420, new_n10416, new_n10421);
not_4  g10045(new_n10421, new_n10422);
nor_1  g10046(new_n10422, new_n10412, new_n10423);
not_4  g10047(new_n10423, new_n10424);
nand_1 g10048(new_n10424, new_n10411, new_n10425);
nand_1 g10049(new_n10425, new_n10404, new_n10426);
nand_1 g10050(new_n10426, new_n10402, new_n10427);
not_4  g10051(new_n10427, new_n10428);
not_4  g10052(new_n10398, new_n10429);
nand_1 g10053(new_n10397, new_n10396, new_n10430);
nand_1 g10054(new_n10430, new_n10429, new_n10431);
nor_1  g10055(new_n10431, new_n10428, new_n10432);
nor_1  g10056(new_n10432, new_n10398, new_n10433);
nor_1  g10057(new_n10433, new_n10394, new_n10434);
not_4  g10058(new_n10434, new_n10435);
xnor_1 g10059(new_n10227, new_n10185, new_n10436);
nand_1 g10060(new_n10433, new_n10394, new_n10437);
nand_1 g10061(new_n10437, new_n10435, new_n10438);
nor_1  g10062(new_n10438, new_n10436, new_n10439_1);
not_4  g10063(new_n10439_1, new_n10440);
nand_1 g10064(new_n10440, new_n10435, new_n10441);
nand_1 g10065(new_n10387, new_n10384, new_n10442);
nand_1 g10066(new_n10382, new_n10230, new_n10443);
nand_1 g10067(new_n10443, new_n10442, new_n10444);
nor_1  g10068(new_n10444, new_n9819, new_n10445);
nor_1  g10069(new_n10389, new_n9820_1, new_n10446);
nor_1  g10070(new_n10446, new_n10445, new_n10447);
nand_1 g10071(new_n10447, new_n10441, new_n10448);
nand_1 g10072(new_n10448, new_n10390, new_n10449);
nand_1 g10073(new_n10378, new_n10364, new_n10450);
not_4  g10074(new_n10450, new_n10451_1);
nor_1  g10075(new_n10383, new_n10385, new_n10452);
nand_1 g10076(new_n10452, new_n10451_1, new_n10453);
nand_1 g10077(new_n10442, new_n10377, new_n10454);
nand_1 g10078(new_n10454, new_n10450, new_n10455);
nand_1 g10079(new_n10455, new_n10453, new_n10456);
not_4  g10080(new_n10231, new_n10457);
nand_1 g10081(new_n10266, new_n10457, new_n10458);
not_4  g10082(new_n10267, new_n10459);
nor_1  g10083(new_n10271, new_n10459, new_n10460);
not_4  g10084(new_n10460, new_n10461);
nand_1 g10085(new_n10461, new_n10458, new_n10462);
nand_1 g10086(new_n10321, new_n10319, new_n10463);
not_4  g10087(new_n10353, new_n10464);
nand_1 g10088(new_n10464, new_n10323, new_n10465);
nand_1 g10089(new_n10465, new_n10463, new_n10466);
nand_1 g10090(new_n10298, new_n10292, new_n10467);
nand_1 g10091(new_n10467, new_n10289, new_n10468);
not_4  g10092(new_n10332, new_n10469);
nand_1 g10093(new_n10335, new_n10469, new_n10470);
nand_1 g10094(new_n10470, new_n10338, new_n10471);
xnor_1 g10095(new_n10471, new_n10468, new_n10472);
nand_1 g10096(n8028, n4817, new_n10473);
nand_1 g10097(n7523, n7354, new_n10474);
xnor_1 g10098(new_n10474, new_n10473, new_n10475);
nand_1 g10099(n10848, n9457, new_n10476_1);
nand_1 g10100(n11222, n1906, new_n10477);
xnor_1 g10101(new_n10477, new_n10476_1, new_n10478);
nand_1 g10102(n6986, n4928, new_n10479);
nand_1 g10103(n4141, n2226, new_n10480);
not_4  g10104(new_n10480, new_n10481);
xnor_1 g10105(new_n10481, new_n10479, new_n10482);
xnor_1 g10106(new_n10482, new_n10478, new_n10483);
xnor_1 g10107(new_n10483, new_n10475, new_n10484);
not_4  g10108(new_n9797, new_n10485);
nand_1 g10109(new_n9803, new_n10485, new_n10486);
nand_1 g10110(new_n10486, new_n9802, new_n10487);
nand_1 g10111(n4516, n2509, new_n10488);
nand_1 g10112(n12704, n996, new_n10489);
nand_1 g10113(n12720, n3627, new_n10490);
not_4  g10114(new_n10490, new_n10491);
xnor_1 g10115(new_n10491, new_n10489, new_n10492);
xnor_1 g10116(new_n10492, new_n10488, new_n10493);
xnor_1 g10117(new_n10493, new_n10487, new_n10494);
xnor_1 g10118(new_n10494, new_n10484, new_n10495);
nand_1 g10119(n2515, n533, new_n10496);
nand_1 g10120(n1512, n1199, new_n10497);
nand_1 g10121(n12391, n12044, new_n10498);
xnor_1 g10122(new_n10498, new_n10497, new_n10499);
xnor_1 g10123(new_n10499, new_n10496, new_n10500);
xnor_1 g10124(new_n10500, new_n10495, new_n10501);
xnor_1 g10125(new_n10501, new_n10472, new_n10502);
not_4  g10126(new_n10275, new_n10503);
nand_1 g10127(new_n10282, new_n10503, new_n10504);
not_4  g10128(new_n10300, new_n10505);
nand_1 g10129(new_n10505, new_n10283, new_n10506);
nand_1 g10130(new_n10506, new_n10504, new_n10507);
nand_1 g10131(new_n10295, new_n10294, new_n10508);
nand_1 g10132(new_n10297, new_n10293, new_n10509);
nand_1 g10133(new_n10509, new_n10508, new_n10510_1);
nand_1 g10134(n12069, n5694, new_n10511);
nand_1 g10135(n11153, n4903, new_n10512);
xnor_1 g10136(new_n10512, new_n10511, new_n10513);
nand_1 g10137(n7294, n5767, new_n10514);
nand_1 g10138(n8336, n783, new_n10515);
xnor_1 g10139(new_n10515, new_n10514, new_n10516);
xnor_1 g10140(new_n10516, new_n10513, new_n10517);
xnor_1 g10141(new_n10517, new_n10510_1, new_n10518);
nand_1 g10142(n4189, n4005, new_n10519);
nand_1 g10143(n5814, n5314, new_n10520);
xnor_1 g10144(new_n10520, new_n10519, new_n10521);
xnor_1 g10145(new_n10521, new_n10518, new_n10522);
xnor_1 g10146(new_n10522, new_n10507, new_n10523);
xnor_1 g10147(new_n10523, new_n10502, new_n10524);
xnor_1 g10148(new_n10524, new_n10466, new_n10525);
xnor_1 g10149(new_n10525, new_n10462, new_n10526);
nand_1 g10150(new_n10354, new_n10124, new_n10527);
nand_1 g10151(new_n10357, new_n10355, new_n10528);
nand_1 g10152(new_n10528, new_n10527, new_n10529);
not_4  g10153(new_n10004, new_n10530);
nand_1 g10154(new_n10309, new_n10530, new_n10531);
nand_1 g10155(new_n10314, new_n10310, new_n10532);
nand_1 g10156(new_n10532, new_n10531, new_n10533);
nand_1 g10157(new_n9793, new_n9788, new_n10534);
not_4  g10158(new_n9794, new_n10535);
nand_1 g10159(new_n9806, new_n10535, new_n10536);
nand_1 g10160(new_n10536, new_n10534, new_n10537);
nand_1 g10161(new_n9791, new_n9790, new_n10538);
not_4  g10162(new_n9792, new_n10539);
nand_1 g10163(new_n10539, new_n9789, new_n10540);
nand_1 g10164(new_n10540, new_n10538, new_n10541);
xnor_1 g10165(new_n10541, new_n10537, new_n10542);
nand_1 g10166(new_n10279, new_n10278_1, new_n10543);
nand_1 g10167(new_n10281, new_n10276, new_n10544);
nand_1 g10168(new_n10544, new_n10543, new_n10545_1);
nand_1 g10169(new_n10348, new_n10347, new_n10546);
nand_1 g10170(new_n10350, new_n10345, new_n10547_1);
nand_1 g10171(new_n10547_1, new_n10546, new_n10548);
xnor_1 g10172(new_n10548, new_n10545_1, new_n10549);
xnor_1 g10173(new_n10549, new_n10542, new_n10550);
xnor_1 g10174(new_n10550, new_n10533, new_n10551);
not_4  g10175(new_n10551, new_n10552);
not_4  g10176(new_n9814, new_n10553);
nor_1  g10177(new_n9818, new_n9783, new_n10554);
nor_1  g10178(new_n10554, new_n10553, new_n10555);
not_4  g10179(new_n10344, new_n10556);
nand_1 g10180(new_n10351, new_n10556, new_n10557);
not_4  g10181(new_n10342, new_n10558);
nand_1 g10182(new_n10352, new_n10558, new_n10559);
nand_1 g10183(new_n10559, new_n10557, new_n10560);
nand_1 g10184(n6578, n1564, new_n10561);
xnor_1 g10185(new_n10561, new_n10560, new_n10562);
xnor_1 g10186(new_n10562, new_n10555, new_n10563);
nand_1 g10187(new_n10563, new_n10552, new_n10564);
not_4  g10188(new_n10562, new_n10565);
xnor_1 g10189(new_n10565, new_n10555, new_n10566);
nand_1 g10190(new_n10566, new_n10551, new_n10567);
nand_1 g10191(new_n10567, new_n10564, new_n10568);
nand_1 g10192(new_n10306, new_n10304, new_n10569);
not_4  g10193(new_n10301, new_n10570);
nand_1 g10194(new_n10308, new_n10570, new_n10571);
nand_1 g10195(new_n10571, new_n10569, new_n10572);
not_4  g10196(new_n10250, new_n10573);
nand_1 g10197(new_n10256, new_n10573, new_n10574);
nand_1 g10198(new_n10574, new_n10248, new_n10575);
nand_1 g10199(new_n10240, new_n10239, new_n10576);
nand_1 g10200(new_n10242, new_n10238, new_n10577);
nand_1 g10201(new_n10577, new_n10576, new_n10578);
nand_1 g10202(n5319, n1980, new_n10579);
nand_1 g10203(n9920, n2508, new_n10580);
nand_1 g10204(n10678, n1209, new_n10581);
xnor_1 g10205(new_n10581, new_n10580, new_n10582);
xnor_1 g10206(new_n10582, new_n10579, new_n10583);
xnor_1 g10207(new_n10583, new_n10578, new_n10584);
xnor_1 g10208(new_n10584, new_n10575, new_n10585);
xnor_1 g10209(new_n10585, new_n10572, new_n10586);
nor_1  g10210(new_n10243, new_n10236, new_n10587);
not_4  g10211(new_n10244, new_n10588);
nor_1  g10212(new_n10257, new_n10588, new_n10589_1);
nor_1  g10213(new_n10589_1, new_n10587, new_n10590);
nand_1 g10214(new_n10253, new_n10252, new_n10591);
nand_1 g10215(new_n10255, new_n10251, new_n10592);
nand_1 g10216(new_n10592, new_n10591, new_n10593);
nand_1 g10217(n4828, n2802, new_n10594);
nand_1 g10218(n10928, n8236, new_n10595);
nand_1 g10219(n5105, n1094, new_n10596);
xnor_1 g10220(new_n10596, new_n10595, new_n10597);
xnor_1 g10221(new_n10597, new_n10594, new_n10598);
xnor_1 g10222(new_n10598, new_n10593, new_n10599);
xnor_1 g10223(new_n10599, new_n10590, new_n10600);
xnor_1 g10224(new_n10600, new_n10586, new_n10601);
not_4  g10225(new_n10601, new_n10602);
not_4  g10226(new_n10331, new_n10603);
nand_1 g10227(new_n10341, new_n10603, new_n10604);
nand_1 g10228(new_n10604, new_n10329, new_n10605);
nand_1 g10229(n7891, n5069, new_n10606);
nand_1 g10230(n6038, n2087, new_n10607);
xnor_1 g10231(new_n10607, new_n10606, new_n10608);
xnor_1 g10232(new_n10608, new_n10605, new_n10609);
nand_1 g10233(n7160, n6806, new_n10610);
nand_1 g10234(n6687, n615, new_n10611);
xnor_1 g10235(new_n10611, new_n10610, new_n10612);
xnor_1 g10236(new_n10612, new_n10609, new_n10613);
xnor_1 g10237(new_n10613, new_n10602, new_n10614);
nand_1 g10238(new_n9810, new_n9809, new_n10615);
nand_1 g10239(new_n9812, new_n9815, new_n10616);
nand_1 g10240(new_n10616, new_n10615, new_n10617);
nand_1 g10241(new_n10263, new_n10260, new_n10618);
not_4  g10242(new_n10258, new_n10619);
nand_1 g10243(new_n10265, new_n10619, new_n10620);
nand_1 g10244(new_n10620, new_n10618, new_n10621);
nand_1 g10245(new_n9795, new_n9702, new_n10622);
not_4  g10246(new_n9796, new_n10623);
nand_1 g10247(new_n9805, new_n10623, new_n10624);
nand_1 g10248(new_n10624, new_n10622, new_n10625);
nand_1 g10249(n7500, n7320, new_n10626);
not_4  g10250(new_n10626, new_n10627);
nand_1 g10251(n12706, n2564, new_n10628);
nand_1 g10252(n6770, n2585, new_n10629);
xnor_1 g10253(new_n10629, new_n10628, new_n10630);
xnor_1 g10254(new_n10630, new_n10627, new_n10631);
xnor_1 g10255(new_n10631, new_n10625, new_n10632);
xnor_1 g10256(new_n10632, new_n10621, new_n10633);
xnor_1 g10257(new_n10633, new_n10617, new_n10634);
xnor_1 g10258(new_n10634, new_n10614, new_n10635);
nand_1 g10259(new_n10635, new_n10568, new_n10636);
nor_1  g10260(new_n10566, new_n10551, new_n10637);
nor_1  g10261(new_n10563, new_n10552, new_n10638);
nor_1  g10262(new_n10638, new_n10637, new_n10639);
not_4  g10263(new_n10635, new_n10640);
nand_1 g10264(new_n10640, new_n10639, new_n10641);
nand_1 g10265(new_n10641, new_n10636, new_n10642);
nor_1  g10266(new_n10642, new_n10529, new_n10643);
not_4  g10267(new_n10529, new_n10644_1);
nor_1  g10268(new_n10640, new_n10639, new_n10645);
nor_1  g10269(new_n10635, new_n10568, new_n10646);
nor_1  g10270(new_n10646, new_n10645, new_n10647);
nor_1  g10271(new_n10647, new_n10644_1, new_n10648);
nor_1  g10272(new_n10648, new_n10643, new_n10649);
nor_1  g10273(new_n10649, new_n10526, new_n10650);
not_4  g10274(new_n10526, new_n10651);
nand_1 g10275(new_n10647, new_n10644_1, new_n10652);
nand_1 g10276(new_n10642, new_n10529, new_n10653);
nand_1 g10277(new_n10653, new_n10652, new_n10654);
nor_1  g10278(new_n10654, new_n10651, new_n10655);
nor_1  g10279(new_n10655, new_n10650, new_n10656);
nand_1 g10280(new_n10656, new_n10456, new_n10657);
nor_1  g10281(new_n10454, new_n10450, new_n10658);
nor_1  g10282(new_n10452, new_n10451_1, new_n10659);
nor_1  g10283(new_n10659, new_n10658, new_n10660);
nand_1 g10284(new_n10654, new_n10651, new_n10661);
nand_1 g10285(new_n10649, new_n10526, new_n10662);
nand_1 g10286(new_n10662, new_n10661, new_n10663);
nand_1 g10287(new_n10663, new_n10660, new_n10664);
nand_1 g10288(new_n10664, new_n10657, new_n10665);
nor_1  g10289(new_n10665, new_n10449, new_n10666);
not_4  g10290(new_n10441, new_n10667);
nand_1 g10291(new_n10444, new_n9819, new_n10668);
nand_1 g10292(new_n10668, new_n10390, new_n10669);
nor_1  g10293(new_n10669, new_n10667, new_n10670);
nor_1  g10294(new_n10670, new_n10445, new_n10671);
nor_1  g10295(new_n10663, new_n10660, new_n10672);
nor_1  g10296(new_n10656, new_n10456, new_n10673);
nor_1  g10297(new_n10673, new_n10672, new_n10674);
nor_1  g10298(new_n10674, new_n10671, new_n10675);
nor_1  g10299(new_n10675, new_n10666, n3654);
nand_1 g10300(new_n10438, new_n10436, new_n10677);
nand_1 g10301(new_n10677, new_n10440, n3661);
nand_1 g10302(n7456, n5305, new_n10679);
nand_1 g10303(n5964, n3932, new_n10680);
not_4  g10304(new_n10680, new_n10681);
nand_1 g10305(n1798, n1097, new_n10682);
nand_1 g10306(n12591, n5305, new_n10683);
nand_1 g10307(new_n10683, new_n10682, new_n10684);
nand_1 g10308(new_n10684, new_n10681, new_n10685_1);
nor_1  g10309(new_n10683, new_n10682, new_n10686);
not_4  g10310(new_n10686, new_n10687);
nand_1 g10311(new_n10687, new_n10685_1, new_n10688);
xnor_1 g10312(new_n10688, new_n10679, new_n10689);
nand_1 g10313(n3932, n1097, new_n10690);
nand_1 g10314(n4312, n1798, new_n10691);
nand_1 g10315(n12591, n5964, new_n10692);
xnor_1 g10316(new_n10692, new_n10691, new_n10693);
xnor_1 g10317(new_n10693, new_n10690, new_n10694);
xnor_1 g10318(new_n10694, new_n10689, new_n10695_1);
nand_1 g10319(new_n10687, new_n10684, new_n10696);
not_4  g10320(new_n10696, new_n10697);
nor_1  g10321(new_n10697, new_n6819, new_n10698);
nand_1 g10322(new_n10698, new_n10695_1, new_n10699);
nand_1 g10323(n11662, n5305, new_n10700);
not_4  g10324(new_n10700, new_n10701);
nand_1 g10325(n7456, n5964, new_n10702);
nand_1 g10326(n4312, n3932, new_n10703);
nand_1 g10327(n12591, n1097, new_n10704);
nand_1 g10328(n12705, n1798, new_n10705);
not_4  g10329(new_n10705, new_n10706);
xnor_1 g10330(new_n10706, new_n10704, new_n10707);
not_4  g10331(new_n10707, new_n10708);
xnor_1 g10332(new_n10708, new_n10703, new_n10709);
nor_1  g10333(new_n10709, new_n10702, new_n10710);
not_4  g10334(new_n10710, new_n10711);
nand_1 g10335(new_n10709, new_n10702, new_n10712);
nand_1 g10336(new_n10712, new_n10711, new_n10713);
nand_1 g10337(new_n10692, new_n10691, new_n10714);
not_4  g10338(new_n10693, new_n10715);
nand_1 g10339(new_n10715, new_n10690, new_n10716);
nand_1 g10340(new_n10716, new_n10714, new_n10717);
nor_1  g10341(new_n10717, new_n10713, new_n10718);
not_4  g10342(new_n10718, new_n10719);
nand_1 g10343(new_n10717, new_n10713, new_n10720);
nand_1 g10344(new_n10720, new_n10719, new_n10721);
not_4  g10345(new_n10721, new_n10722);
nand_1 g10346(new_n10722, new_n10701, new_n10723);
nand_1 g10347(new_n10721, new_n10700, new_n10724);
nand_1 g10348(new_n10724, new_n10723, new_n10725);
not_4  g10349(new_n10679, new_n10726);
nand_1 g10350(new_n10688, new_n10726, new_n10727);
not_4  g10351(new_n10689, new_n10728);
nor_1  g10352(new_n10694, new_n10728, new_n10729);
not_4  g10353(new_n10729, new_n10730);
nand_1 g10354(new_n10730, new_n10727, new_n10731);
xnor_1 g10355(new_n10731, new_n10725, new_n10732);
xnor_1 g10356(new_n10732, new_n10699, new_n10733);
not_4  g10357(new_n10733, new_n10734);
xnor_1 g10358(new_n10698, new_n10695_1, new_n10735);
nand_1 g10359(n11023, n8759, new_n10736);
nand_1 g10360(n8759, n3022, new_n10737);
nand_1 g10361(n12299, n6703, new_n10738);
nand_1 g10362(new_n10738, new_n10737, new_n10739);
nand_1 g10363(n12299, n3022, new_n10740);
not_4  g10364(new_n10740, new_n10741);
nand_1 g10365(new_n10741, new_n6822_1, new_n10742);
nand_1 g10366(n9640, n6776, new_n10743);
nand_1 g10367(new_n10743, new_n10742, new_n10744);
nand_1 g10368(new_n10744, new_n10739, new_n10745);
nor_1  g10369(new_n10745, new_n10736, new_n10746);
not_4  g10370(new_n10746, new_n10747);
nand_1 g10371(new_n10745, new_n10736, new_n10748);
nand_1 g10372(new_n10748, new_n10747, new_n10749);
nand_1 g10373(n12299, n9640, new_n10750);
not_4  g10374(new_n10750, new_n10751);
nand_1 g10375(n6776, n3022, new_n10752);
nand_1 g10376(n7436, n6703, new_n10753);
nand_1 g10377(new_n10753, new_n10752, new_n10754);
not_4  g10378(new_n10752, new_n10755);
not_4  g10379(new_n10753, new_n10756);
nand_1 g10380(new_n10756, new_n10755, new_n10757);
nand_1 g10381(new_n10757, new_n10754, new_n10758);
xnor_1 g10382(new_n10758, new_n10751, new_n10759);
xnor_1 g10383(new_n10759, new_n10749, new_n10760);
not_4  g10384(new_n10743, new_n10761);
nand_1 g10385(new_n10761, new_n6802, new_n10762);
nand_1 g10386(new_n10742, new_n10739, new_n10763);
nand_1 g10387(new_n10763, new_n10762, new_n10764);
not_4  g10388(new_n10764, new_n10765);
nand_1 g10389(new_n10765, new_n10761, new_n10766);
xnor_1 g10390(new_n10766, new_n10760, new_n10767);
not_4  g10391(new_n10767, new_n10768);
nand_1 g10392(n11922, n5331, new_n10769);
nand_1 g10393(n2530, n1067, new_n10770);
not_4  g10394(new_n10770, new_n10771);
nand_1 g10395(n8665, n8476, new_n10772);
nand_1 g10396(n12648, n5645, new_n10773);
nand_1 g10397(new_n10773, new_n10772, new_n10774);
not_4  g10398(new_n10772, new_n10775);
not_4  g10399(new_n10773, new_n10776);
nand_1 g10400(new_n10776, new_n10775, new_n10777);
nand_1 g10401(new_n10777, new_n10774, new_n10778);
xnor_1 g10402(new_n10778, new_n10771, new_n10779);
xnor_1 g10403(new_n10779, new_n10769, new_n10780);
nand_1 g10404(n8665, n5331, new_n10781);
nand_1 g10405(n5645, n2530, new_n10782);
nand_1 g10406(new_n10782, new_n10781, new_n10783);
nand_1 g10407(n8476, n1067, new_n10784);
nand_1 g10408(n8665, n2530, new_n10785);
not_4  g10409(new_n10785, new_n10786);
nand_1 g10410(new_n10786, new_n6804, new_n10787);
nand_1 g10411(new_n10787, new_n10784, new_n10788);
nand_1 g10412(new_n10788, new_n10783, new_n10789_1);
not_4  g10413(new_n10789_1, new_n10790);
xnor_1 g10414(new_n10790, new_n10780, new_n10791);
nand_1 g10415(new_n10787, new_n10783, new_n10792);
not_4  g10416(new_n10792, new_n10793);
nor_1  g10417(new_n10793, new_n6840, new_n10794);
xnor_1 g10418(new_n10794, new_n10791, new_n10795);
nand_1 g10419(n7965, n2749, new_n10796);
nand_1 g10420(n7965, n3754, new_n10797);
nand_1 g10421(n11892, n11876, new_n10798);
nand_1 g10422(new_n10798, new_n10797, new_n10799);
nand_1 g10423(n11892, n3754, new_n10800);
not_4  g10424(new_n10800, new_n10801);
nand_1 g10425(new_n10801, new_n6806_1, new_n10802);
nand_1 g10426(n10898, n7388, new_n10803);
nand_1 g10427(new_n10803, new_n10802, new_n10804);
nand_1 g10428(new_n10804, new_n10799, new_n10805);
xnor_1 g10429(new_n10805, new_n10796, new_n10806);
nand_1 g10430(n11892, n10898, new_n10807);
nand_1 g10431(n7388, n3754, new_n10808);
nand_1 g10432(n11876, n2393, new_n10809);
nand_1 g10433(new_n10809, new_n10808, new_n10810);
not_4  g10434(new_n10810, new_n10811);
nor_1  g10435(new_n10809, new_n10808, new_n10812);
nor_1  g10436(new_n10812, new_n10811, new_n10813);
nor_1  g10437(new_n10813, new_n10807, new_n10814);
nand_1 g10438(new_n10813, new_n10807, new_n10815);
not_4  g10439(new_n10815, new_n10816);
nor_1  g10440(new_n10816, new_n10814, new_n10817);
nor_1  g10441(new_n10817, new_n10806, new_n10818);
not_4  g10442(new_n10818, new_n10819);
nand_1 g10443(new_n10817, new_n10806, new_n10820);
nand_1 g10444(new_n10820, new_n10819, new_n10821);
not_4  g10445(new_n10803, new_n10822);
nand_1 g10446(new_n10822, new_n6805, new_n10823);
nand_1 g10447(new_n10802, new_n10799, new_n10824);
nand_1 g10448(new_n10824, new_n10823, new_n10825);
not_4  g10449(new_n10825, new_n10826);
nand_1 g10450(new_n10826, new_n10822, new_n10827);
not_4  g10451(new_n10827, new_n10828);
xnor_1 g10452(new_n10828, new_n10821, new_n10829);
nand_1 g10453(new_n10829, new_n10795, new_n10830);
nor_1  g10454(new_n10829, new_n10795, new_n10831);
not_4  g10455(new_n10831, new_n10832);
nand_1 g10456(new_n10832, new_n10830, new_n10833);
not_4  g10457(new_n10823, new_n10834);
nand_1 g10458(new_n10834, new_n10799, new_n10835);
nand_1 g10459(new_n10835, new_n10825, new_n10836);
not_4  g10460(new_n6807, new_n10837);
nand_1 g10461(new_n6832, new_n10837, new_n10838);
nand_1 g10462(new_n6844, new_n10838, new_n10839);
not_4  g10463(new_n10839, new_n10840);
nand_1 g10464(new_n10840, new_n10836, new_n10841);
xnor_1 g10465(new_n10839, new_n10836, new_n10842);
nor_1  g10466(new_n10784, new_n6804, new_n10843);
not_4  g10467(new_n10843, new_n10844);
nor_1  g10468(new_n10844, new_n10783, new_n10845);
not_4  g10469(new_n10845, new_n10846);
nand_1 g10470(new_n10844, new_n10793, new_n10847);
nand_1 g10471(new_n10847, new_n10846, new_n10848_1);
not_4  g10472(new_n10848_1, new_n10849);
nand_1 g10473(new_n10849, new_n10842, new_n10850);
nand_1 g10474(new_n10850, new_n10841, new_n10851_1);
xnor_1 g10475(new_n10851_1, new_n10833, new_n10852);
xnor_1 g10476(new_n10852, new_n10768, new_n10853);
not_4  g10477(new_n10762, new_n10854);
nand_1 g10478(new_n10854, new_n10739, new_n10855);
nand_1 g10479(new_n10855, new_n10764, new_n10856);
not_4  g10480(new_n6823, new_n10857);
nand_1 g10481(new_n6827, new_n10857, new_n10858);
not_4  g10482(new_n6845, new_n10859);
nand_1 g10483(new_n10859, new_n6828, new_n10860);
nand_1 g10484(new_n10860, new_n10858, new_n10861);
not_4  g10485(new_n10861, new_n10862);
nand_1 g10486(new_n10862, new_n10856, new_n10863);
xnor_1 g10487(new_n10848_1, new_n10842, new_n10864);
xnor_1 g10488(new_n10861, new_n10856, new_n10865);
nand_1 g10489(new_n10865, new_n10864, new_n10866);
nand_1 g10490(new_n10866, new_n10863, new_n10867);
xnor_1 g10491(new_n10867, new_n10853, new_n10868);
nor_1  g10492(new_n10868, new_n10735, new_n10869);
xnor_1 g10493(new_n10868, new_n10735, new_n10870);
xnor_1 g10494(new_n10865, new_n10864, new_n10871);
nand_1 g10495(new_n10681, new_n6800, new_n10872);
nor_1  g10496(new_n10872, new_n10684, new_n10873);
not_4  g10497(new_n10873, new_n10874);
nand_1 g10498(new_n10872, new_n10697, new_n10875);
nand_1 g10499(new_n10875, new_n10874, new_n10876);
nor_1  g10500(new_n10876, new_n10871, new_n10877);
not_4  g10501(new_n6820, new_n10878);
nand_1 g10502(new_n10878, new_n6813, new_n10879);
nand_1 g10503(new_n6846, new_n6821, new_n10880);
nand_1 g10504(new_n10880, new_n10879, new_n10881);
xnor_1 g10505(new_n10876, new_n10871, new_n10882);
nor_1  g10506(new_n10882, new_n10881, new_n10883);
nor_1  g10507(new_n10883, new_n10877, new_n10884);
not_4  g10508(new_n10884, new_n10885);
nor_1  g10509(new_n10885, new_n10870, new_n10886);
nor_1  g10510(new_n10886, new_n10869, new_n10887);
nand_1 g10511(new_n10887, new_n10734, new_n10888);
nor_1  g10512(new_n10887, new_n10734, new_n10889);
not_4  g10513(new_n10889, new_n10890);
nand_1 g10514(new_n10890, new_n10888, new_n10891);
not_4  g10515(new_n10766, new_n10892);
nand_1 g10516(new_n10892, new_n10760, new_n10893);
nand_1 g10517(n10451, n8759, new_n10894);
nand_1 g10518(n11023, n6776, new_n10895);
nand_1 g10519(new_n10757, new_n10750, new_n10896);
nand_1 g10520(new_n10896, new_n10754, new_n10897);
not_4  g10521(new_n10897, new_n10898_1);
xnor_1 g10522(new_n10898_1, new_n10895, new_n10899);
nand_1 g10523(n9640, n7436, new_n10900);
not_4  g10524(new_n10900, new_n10901);
nand_1 g10525(n8276, n6703, new_n10902);
nand_1 g10526(new_n10902, new_n10740, new_n10903);
not_4  g10527(new_n10902, new_n10904);
nand_1 g10528(new_n10904, new_n10741, new_n10905);
nand_1 g10529(new_n10905, new_n10903, new_n10906);
xnor_1 g10530(new_n10906, new_n10901, new_n10907);
xnor_1 g10531(new_n10907, new_n10899, new_n10908);
not_4  g10532(new_n10908, new_n10909);
xnor_1 g10533(new_n10909, new_n10894, new_n10910);
not_4  g10534(new_n10749, new_n10911);
nand_1 g10535(new_n10759, new_n10911, new_n10912);
nand_1 g10536(new_n10912, new_n10747, new_n10913_1);
xnor_1 g10537(new_n10913_1, new_n10910, new_n10914);
not_4  g10538(new_n10914, new_n10915);
xnor_1 g10539(new_n10915, new_n10893, new_n10916);
not_4  g10540(new_n10916, new_n10917);
not_4  g10541(new_n10821, new_n10918);
nand_1 g10542(new_n10828, new_n10918, new_n10919);
nand_1 g10543(n7965, n159, new_n10920);
nor_1  g10544(new_n10805, new_n10796, new_n10921);
nor_1  g10545(new_n10818, new_n10921, new_n10922);
not_4  g10546(new_n10922, new_n10923);
xnor_1 g10547(new_n10923, new_n10920, new_n10924);
nand_1 g10548(n7388, n2749, new_n10925);
nand_1 g10549(new_n10815, new_n10810, new_n10926);
not_4  g10550(new_n10926, new_n10927);
xnor_1 g10551(new_n10927, new_n10925, new_n10928_1);
nand_1 g10552(n11876, n5860, new_n10929);
nand_1 g10553(n10898, n2393, new_n10930);
xnor_1 g10554(new_n10930, new_n10929, new_n10931);
not_4  g10555(new_n10931, new_n10932);
xnor_1 g10556(new_n10932, new_n10800, new_n10933);
nand_1 g10557(new_n10933, new_n10928_1, new_n10934);
not_4  g10558(new_n10934, new_n10935);
nor_1  g10559(new_n10933, new_n10928_1, new_n10936);
nor_1  g10560(new_n10936, new_n10935, new_n10937);
xnor_1 g10561(new_n10937, new_n10924, new_n10938);
not_4  g10562(new_n10938, new_n10939);
xnor_1 g10563(new_n10939, new_n10919, new_n10940);
not_4  g10564(new_n10791, new_n10941);
nand_1 g10565(new_n10794, new_n10941, new_n10942);
nand_1 g10566(n5331, n2551, new_n10943);
nand_1 g10567(n11922, n8476, new_n10944);
nand_1 g10568(new_n10777, new_n10770, new_n10945);
nand_1 g10569(new_n10945, new_n10774, new_n10946);
not_4  g10570(new_n10946, new_n10947);
xnor_1 g10571(new_n10947, new_n10944, new_n10948);
nand_1 g10572(n12648, n1067, new_n10949_1);
not_4  g10573(new_n10949_1, new_n10950);
nand_1 g10574(n10545, n5645, new_n10951);
nand_1 g10575(new_n10951, new_n10785, new_n10952);
nor_1  g10576(new_n10951, new_n10785, new_n10953);
not_4  g10577(new_n10953, new_n10954);
nand_1 g10578(new_n10954, new_n10952, new_n10955);
xnor_1 g10579(new_n10955, new_n10950, new_n10956);
not_4  g10580(new_n10956, new_n10957);
xnor_1 g10581(new_n10957, new_n10948, new_n10958);
xnor_1 g10582(new_n10958, new_n10943, new_n10959);
not_4  g10583(new_n10769, new_n10960);
nand_1 g10584(new_n10779, new_n10960, new_n10961);
nand_1 g10585(new_n10790, new_n10780, new_n10962);
nand_1 g10586(new_n10962, new_n10961, new_n10963);
xnor_1 g10587(new_n10963, new_n10959, new_n10964);
not_4  g10588(new_n10964, new_n10965_1);
xnor_1 g10589(new_n10965_1, new_n10942, new_n10966);
nand_1 g10590(new_n10966, new_n10940, new_n10967);
nor_1  g10591(new_n10966, new_n10940, new_n10968);
not_4  g10592(new_n10968, new_n10969);
nand_1 g10593(new_n10969, new_n10967, new_n10970);
not_4  g10594(new_n10833, new_n10971);
nand_1 g10595(new_n10851_1, new_n10971, new_n10972);
nand_1 g10596(new_n10972, new_n10832, new_n10973);
xnor_1 g10597(new_n10973, new_n10970, new_n10974);
nor_1  g10598(new_n10974, new_n10917, new_n10975);
not_4  g10599(new_n10975, new_n10976);
nand_1 g10600(new_n10974, new_n10917, new_n10977);
nand_1 g10601(new_n10977, new_n10976, new_n10978);
nand_1 g10602(new_n10852, new_n10768, new_n10979);
not_4  g10603(new_n10853, new_n10980);
nand_1 g10604(new_n10867, new_n10980, new_n10981);
nand_1 g10605(new_n10981, new_n10979, new_n10982);
nor_1  g10606(new_n10982, new_n10978, new_n10983);
not_4  g10607(new_n10983, new_n10984);
nand_1 g10608(new_n10982, new_n10978, new_n10985);
nand_1 g10609(new_n10985, new_n10984, new_n10986);
not_4  g10610(new_n10986, new_n10987);
xnor_1 g10611(new_n10987, new_n10891, n3677);
xnor_1 g10612(new_n9491, new_n9490, n3849);
not_4  g10613(new_n6795, new_n10990_1);
xnor_1 g10614(new_n10990_1, new_n6794, n4088);
xnor_1 g10615(new_n1225, new_n1101, n4155);
xnor_1 g10616(new_n3172_1, new_n3171, n4159);
xnor_1 g10617(new_n6784, new_n6587, n4226);
nand_1 g10618(n12591, n4312, new_n10995);
nand_1 g10619(new_n10705, new_n10704, new_n10996);
nand_1 g10620(new_n10707, new_n10703, new_n10997);
nand_1 g10621(new_n10997, new_n10996, new_n10998);
not_4  g10622(new_n10998, new_n10999);
xnor_1 g10623(new_n10999, new_n10995, new_n11000);
nand_1 g10624(n12705, n3932, new_n11001);
nand_1 g10625(n12025, n1798, new_n11002);
nand_1 g10626(new_n11002, new_n11001, new_n11003);
not_4  g10627(new_n11001, new_n11004);
not_4  g10628(new_n11002, new_n11005);
nand_1 g10629(new_n11005, new_n11004, new_n11006);
nand_1 g10630(new_n11006, new_n11003, new_n11007);
xnor_1 g10631(new_n11007, new_n11000, new_n11008);
not_4  g10632(new_n11008, new_n11009);
nand_1 g10633(n11662, n5964, new_n11010);
not_4  g10634(new_n11010, new_n11011);
nand_1 g10635(n7456, n1097, new_n11012);
not_4  g10636(new_n11012, new_n11013);
nand_1 g10637(new_n11013, new_n11011, new_n11014);
nand_1 g10638(new_n11012, new_n11010, new_n11015);
nand_1 g10639(new_n11015, new_n11014, new_n11016);
nand_1 g10640(new_n11016, new_n11009, new_n11017);
not_4  g10641(new_n11016, new_n11018);
nand_1 g10642(new_n11018, new_n11008, new_n11019);
nand_1 g10643(new_n11019, new_n11017, new_n11020);
not_4  g10644(new_n11020, new_n11021);
nand_1 g10645(new_n10719, new_n10711, new_n11022);
nand_1 g10646(new_n11022, new_n11021, new_n11023_1);
not_4  g10647(new_n11022, new_n11024);
nand_1 g10648(new_n11024, new_n11020, new_n11025);
nand_1 g10649(new_n11025, new_n11023_1, new_n11026);
not_4  g10650(new_n11026, new_n11027);
not_4  g10651(new_n10725, new_n11028);
nand_1 g10652(new_n10731, new_n11028, new_n11029);
nand_1 g10653(new_n11029, new_n10723, new_n11030);
nand_1 g10654(new_n11030, new_n11027, new_n11031);
nand_1 g10655(new_n10998, new_n10995, new_n11032);
nand_1 g10656(new_n11007, new_n11000, new_n11033);
nand_1 g10657(new_n11033, new_n11032, new_n11034);
nand_1 g10658(n10327, n5964, new_n11035);
nand_1 g10659(n11662, n1097, new_n11036);
nand_1 g10660(n9583, n5305, new_n11037);
not_4  g10661(new_n11037, new_n11038);
xnor_1 g10662(new_n11038, new_n11036, new_n11039);
xnor_1 g10663(new_n11039, new_n11035, new_n11040);
xnor_1 g10664(new_n11040, new_n11034, new_n11041);
nand_1 g10665(n7456, n4312, new_n11042);
xnor_1 g10666(new_n11042, new_n11006, new_n11043);
nand_1 g10667(n12025, n3932, new_n11044);
not_4  g10668(new_n11044, new_n11045);
nand_1 g10669(n12705, n12591, new_n11046);
nand_1 g10670(n11257, n1798, new_n11047);
not_4  g10671(new_n11047, new_n11048);
xnor_1 g10672(new_n11048, new_n11046, new_n11049);
xnor_1 g10673(new_n11049, new_n11045, new_n11050);
xnor_1 g10674(new_n11050, new_n11043, new_n11051);
xnor_1 g10675(new_n11051, new_n11041, new_n11052);
not_4  g10676(new_n11052, new_n11053);
nor_1  g10677(new_n11023_1, new_n11014, new_n11054);
not_4  g10678(new_n11054, new_n11055);
nand_1 g10679(new_n11023_1, new_n11014, new_n11056);
nand_1 g10680(new_n11056, new_n11055, new_n11057);
nand_1 g10681(new_n11057, new_n11019, new_n11058);
xnor_1 g10682(new_n11058, new_n11053, new_n11059);
xnor_1 g10683(new_n11059, new_n11031, new_n11060);
nand_1 g10684(n10327, n5305, new_n11061);
not_4  g10685(new_n11061, new_n11062);
xnor_1 g10686(new_n11030, new_n11026, new_n11063);
nor_1  g10687(new_n11063, new_n11062, new_n11064);
not_4  g10688(new_n11064, new_n11065);
not_4  g10689(new_n10699, new_n11066);
nand_1 g10690(new_n10732, new_n11066, new_n11067);
nand_1 g10691(new_n11063, new_n11062, new_n11068);
nand_1 g10692(new_n11068, new_n11065, new_n11069);
not_4  g10693(new_n11069, new_n11070);
nand_1 g10694(new_n11070, new_n11067, new_n11071);
nand_1 g10695(new_n11071, new_n11065, new_n11072);
xnor_1 g10696(new_n11072, new_n11060, new_n11073);
not_4  g10697(new_n11073, new_n11074);
nor_1  g10698(new_n10897, new_n10895, new_n11075);
not_4  g10699(new_n11075, new_n11076);
nand_1 g10700(new_n10907, new_n10899, new_n11077);
nand_1 g10701(new_n11077, new_n11076, new_n11078);
nand_1 g10702(n10451, n6776, new_n11079);
nand_1 g10703(n12299, n11023, new_n11080);
not_4  g10704(new_n11080, new_n11081);
xnor_1 g10705(new_n11081, new_n11079, new_n11082);
xnor_1 g10706(new_n11082, new_n11078, new_n11083);
nand_1 g10707(n7436, n3022, new_n11084);
nand_1 g10708(n9640, n8276, new_n11085);
nand_1 g10709(n9241, n6703, new_n11086);
nand_1 g10710(new_n11086, new_n11085, new_n11087);
not_4  g10711(new_n11085, new_n11088);
not_4  g10712(new_n11086, new_n11089);
nand_1 g10713(new_n11089, new_n11088, new_n11090);
nand_1 g10714(new_n11090, new_n11087, new_n11091);
xnor_1 g10715(new_n11091, new_n11084, new_n11092);
nand_1 g10716(new_n10905, new_n10900, new_n11093);
nand_1 g10717(new_n11093, new_n10903, new_n11094);
xnor_1 g10718(new_n11094, new_n11092, new_n11095);
xnor_1 g10719(new_n11095, new_n11083, new_n11096);
not_4  g10720(new_n11096, new_n11097);
not_4  g10721(new_n10894, new_n11098);
nand_1 g10722(new_n10909, new_n11098, new_n11099);
nand_1 g10723(new_n10913_1, new_n10910, new_n11100);
nand_1 g10724(new_n11100, new_n11099, new_n11101);
nand_1 g10725(new_n11101, new_n11097, new_n11102);
nand_1 g10726(new_n11091, new_n11084, new_n11103);
not_4  g10727(new_n11092, new_n11104);
nand_1 g10728(new_n11094, new_n11104, new_n11105);
nand_1 g10729(new_n11105, new_n11103, new_n11106);
nand_1 g10730(n10278, n6776, new_n11107);
nand_1 g10731(n12299, n10451, new_n11108);
nand_1 g10732(n11423, n8759, new_n11109);
not_4  g10733(new_n11109, new_n11110);
xnor_1 g10734(new_n11110, new_n11108, new_n11111);
xnor_1 g10735(new_n11111, new_n11107, new_n11112);
xnor_1 g10736(new_n11112, new_n11106, new_n11113);
nand_1 g10737(n11023, n7436, new_n11114);
not_4  g10738(new_n11114, new_n11115);
xnor_1 g10739(new_n11115, new_n11090, new_n11116);
nand_1 g10740(n9640, n9241, new_n11117);
nand_1 g10741(n8276, n3022, new_n11118);
nand_1 g10742(n10510, n6703, new_n11119);
not_4  g10743(new_n11119, new_n11120);
xnor_1 g10744(new_n11120, new_n11118, new_n11121);
xnor_1 g10745(new_n11121, new_n11117, new_n11122);
not_4  g10746(new_n11122, new_n11123);
xnor_1 g10747(new_n11123, new_n11116, new_n11124);
xnor_1 g10748(new_n11124, new_n11113, new_n11125);
nand_1 g10749(new_n11082, new_n11078, new_n11126);
nor_1  g10750(new_n11080, new_n11079, new_n11127);
nor_1  g10751(new_n11095, new_n11083, new_n11128);
xnor_1 g10752(new_n11128, new_n11127, new_n11129);
nand_1 g10753(new_n11129, new_n11126, new_n11130);
xnor_1 g10754(new_n11130, new_n11125, new_n11131);
xnor_1 g10755(new_n11131, new_n11102, new_n11132);
nand_1 g10756(n10278, n8759, new_n11133);
not_4  g10757(new_n11133, new_n11134);
xnor_1 g10758(new_n11101, new_n11096, new_n11135);
nand_1 g10759(new_n11135, new_n11134, new_n11136);
not_4  g10760(new_n10893, new_n11137);
nand_1 g10761(new_n10915, new_n11137, new_n11138);
not_4  g10762(new_n11138, new_n11139);
xnor_1 g10763(new_n11135, new_n11133, new_n11140);
nand_1 g10764(new_n11140, new_n11139, new_n11141);
nand_1 g10765(new_n11141, new_n11136, new_n11142);
xnor_1 g10766(new_n11142, new_n11132, new_n11143);
nand_1 g10767(n12648, n8665, new_n11144);
nand_1 g10768(n10545, n1067, new_n11145);
nand_1 g10769(n7690, n5645, new_n11146);
not_4  g10770(new_n11146, new_n11147);
xnor_1 g10771(new_n11147, new_n11145, new_n11148);
xnor_1 g10772(new_n11148, new_n11144, new_n11149);
not_4  g10773(new_n11149, new_n11150);
nand_1 g10774(new_n10954, new_n10949_1, new_n11151);
nand_1 g10775(new_n11151, new_n10952, new_n11152);
not_4  g10776(new_n11152, new_n11153_1);
xnor_1 g10777(new_n11153_1, new_n11150, new_n11154);
not_4  g10778(new_n11154, new_n11155);
nand_1 g10779(n8476, n2551, new_n11156);
nand_1 g10780(n11922, n2530, new_n11157);
not_4  g10781(new_n11157, new_n11158);
xnor_1 g10782(new_n11158, new_n11156, new_n11159);
xnor_1 g10783(new_n11159, new_n11155, new_n11160);
nor_1  g10784(new_n10946, new_n10944, new_n11161);
not_4  g10785(new_n11161, new_n11162);
nand_1 g10786(new_n10956, new_n10948, new_n11163);
nand_1 g10787(new_n11163, new_n11162, new_n11164);
xnor_1 g10788(new_n11164, new_n11160, new_n11165);
not_4  g10789(new_n11165, new_n11166);
not_4  g10790(new_n10943, new_n11167);
nand_1 g10791(new_n10958, new_n11167, new_n11168);
nand_1 g10792(new_n10963, new_n10959, new_n11169);
nand_1 g10793(new_n11169, new_n11168, new_n11170);
nand_1 g10794(new_n11170, new_n11166, new_n11171);
not_4  g10795(new_n11145, new_n11172);
nand_1 g10796(new_n11147, new_n11172, new_n11173);
not_4  g10797(new_n11173, new_n11174);
nand_1 g10798(n12648, n11922, new_n11175);
not_4  g10799(new_n11175, new_n11176);
nand_1 g10800(new_n11176, new_n11174, new_n11177);
nand_1 g10801(new_n11175, new_n11173, new_n11178);
nand_1 g10802(new_n11178, new_n11177, new_n11179);
nand_1 g10803(n7690, n1067, new_n11180);
nand_1 g10804(n10545, n8665, new_n11181);
nand_1 g10805(n5645, n3616, new_n11182);
not_4  g10806(new_n11182, new_n11183);
xnor_1 g10807(new_n11183, new_n11181, new_n11184);
xnor_1 g10808(new_n11184, new_n11180, new_n11185);
not_4  g10809(new_n11185, new_n11186);
xnor_1 g10810(new_n11186, new_n11179, new_n11187);
not_4  g10811(new_n11144, new_n11188);
nand_1 g10812(new_n11148, new_n11188, new_n11189);
nand_1 g10813(new_n11153_1, new_n11149, new_n11190);
nand_1 g10814(new_n11190, new_n11189, new_n11191);
nand_1 g10815(n12826, n8476, new_n11192);
nand_1 g10816(n2551, n2530, new_n11193);
nand_1 g10817(n5331, n4094, new_n11194);
not_4  g10818(new_n11194, new_n11195);
xnor_1 g10819(new_n11195, new_n11193, new_n11196);
not_4  g10820(new_n11196, new_n11197);
xnor_1 g10821(new_n11197, new_n11192, new_n11198);
xnor_1 g10822(new_n11198, new_n11191, new_n11199);
xnor_1 g10823(new_n11199, new_n11187, new_n11200);
nand_1 g10824(new_n11159, new_n11154, new_n11201);
nor_1  g10825(new_n11157, new_n11156, new_n11202);
nand_1 g10826(new_n11164, new_n11160, new_n11203);
not_4  g10827(new_n11203, new_n11204);
xnor_1 g10828(new_n11204, new_n11202, new_n11205);
nand_1 g10829(new_n11205, new_n11201, new_n11206);
xnor_1 g10830(new_n11206, new_n11200, new_n11207);
xnor_1 g10831(new_n11207, new_n11171, new_n11208);
nand_1 g10832(n12826, n5331, new_n11209);
not_4  g10833(new_n11209, new_n11210);
xnor_1 g10834(new_n11170, new_n11165, new_n11211);
nor_1  g10835(new_n11211, new_n11210, new_n11212);
not_4  g10836(new_n11212, new_n11213);
not_4  g10837(new_n10942, new_n11214);
nand_1 g10838(new_n10965_1, new_n11214, new_n11215);
xnor_1 g10839(new_n11211, new_n11209, new_n11216_1);
nand_1 g10840(new_n11216_1, new_n11215, new_n11217);
nand_1 g10841(new_n11217, new_n11213, new_n11218);
xnor_1 g10842(new_n11218, new_n11208, new_n11219);
nand_1 g10843(n7965, n1510, new_n11220);
not_4  g10844(new_n11220, new_n11221);
not_4  g10845(new_n10925, new_n11222_1);
nand_1 g10846(new_n10927, new_n11222_1, new_n11223);
nand_1 g10847(new_n10934, new_n11223, new_n11224);
nand_1 g10848(n7388, n159, new_n11225);
not_4  g10849(new_n11225, new_n11226);
nand_1 g10850(n11892, n2749, new_n11227);
not_4  g10851(new_n11227, new_n11228);
nand_1 g10852(new_n11228, new_n11226, new_n11229);
nand_1 g10853(new_n11227, new_n11225, new_n11230);
nand_1 g10854(new_n11230, new_n11229, new_n11231);
xnor_1 g10855(new_n11231, new_n11224, new_n11232);
nand_1 g10856(n3754, n2393, new_n11233);
nand_1 g10857(n10898, n5860, new_n11234);
nand_1 g10858(n11876, n3986, new_n11235);
not_4  g10859(new_n11235, new_n11236);
xnor_1 g10860(new_n11236, new_n11234, new_n11237);
xnor_1 g10861(new_n11237, new_n11233, new_n11238);
nand_1 g10862(new_n10930, new_n10929, new_n11239);
not_4  g10863(new_n11239, new_n11240);
nor_1  g10864(new_n10931, new_n10801, new_n11241);
nor_1  g10865(new_n11241, new_n11240, new_n11242);
xnor_1 g10866(new_n11242, new_n11238, new_n11243);
xnor_1 g10867(new_n11243, new_n11232, new_n11244);
nor_1  g10868(new_n10922, new_n10920, new_n11245);
not_4  g10869(new_n11245, new_n11246);
nand_1 g10870(new_n10937, new_n10924, new_n11247);
nand_1 g10871(new_n11247, new_n11246, new_n11248);
nand_1 g10872(new_n11248, new_n11244, new_n11249);
not_4  g10873(new_n11249, new_n11250);
nor_1  g10874(new_n11248, new_n11244, new_n11251);
nor_1  g10875(new_n11251, new_n11250, new_n11252);
nand_1 g10876(new_n11252, new_n11221, new_n11253);
not_4  g10877(new_n10919, new_n11254);
nand_1 g10878(new_n10939, new_n11254, new_n11255);
xnor_1 g10879(new_n11252, new_n11220, new_n11256);
not_4  g10880(new_n11256, new_n11257_1);
nor_1  g10881(new_n11257_1, new_n11255, new_n11258);
not_4  g10882(new_n11258, new_n11259);
nand_1 g10883(new_n11259, new_n11253, new_n11260);
not_4  g10884(new_n11224, new_n11261);
nand_1 g10885(new_n11231, new_n11261, new_n11262);
nand_1 g10886(new_n11243, new_n11232, new_n11263);
nand_1 g10887(new_n11263, new_n11262, new_n11264);
xnor_1 g10888(new_n11264, new_n11229, new_n11265);
nand_1 g10889(n7388, n1510, new_n11266);
nand_1 g10890(n11892, n159, new_n11267);
not_4  g10891(new_n11267, new_n11268);
nand_1 g10892(n12247, n7965, new_n11269);
xnor_1 g10893(new_n11269, new_n11268, new_n11270);
xnor_1 g10894(new_n11270, new_n11266, new_n11271);
not_4  g10895(new_n11233, new_n11272);
nand_1 g10896(new_n11237, new_n11272, new_n11273);
nand_1 g10897(new_n11242, new_n11238, new_n11274);
nand_1 g10898(new_n11274, new_n11273, new_n11275);
not_4  g10899(new_n11275, new_n11276);
xnor_1 g10900(new_n11276, new_n11271, new_n11277);
not_4  g10901(new_n11234, new_n11278);
nand_1 g10902(new_n11236, new_n11278, new_n11279);
not_4  g10903(new_n11279, new_n11280);
nand_1 g10904(n2749, n2393, new_n11281);
not_4  g10905(new_n11281, new_n11282);
nand_1 g10906(new_n11282, new_n11280, new_n11283);
nand_1 g10907(new_n11281, new_n11279, new_n11284);
nand_1 g10908(new_n11284, new_n11283, new_n11285);
not_4  g10909(new_n11285, new_n11286);
nand_1 g10910(n10898, n3986, new_n11287);
nand_1 g10911(n11876, n5857, new_n11288);
nand_1 g10912(n5860, n3754, new_n11289);
not_4  g10913(new_n11289, new_n11290);
xnor_1 g10914(new_n11290, new_n11288, new_n11291);
xnor_1 g10915(new_n11291, new_n11287, new_n11292);
not_4  g10916(new_n11292, new_n11293);
xnor_1 g10917(new_n11293, new_n11286, new_n11294);
xnor_1 g10918(new_n11294, new_n11277, new_n11295);
xnor_1 g10919(new_n11295, new_n11265, new_n11296_1);
not_4  g10920(new_n11296_1, new_n11297);
xnor_1 g10921(new_n11297, new_n11249, new_n11298);
xnor_1 g10922(new_n11298, new_n11260, new_n11299);
xnor_1 g10923(new_n11299, new_n11219, new_n11300);
xnor_1 g10924(new_n11256, new_n11255, new_n11301);
xnor_1 g10925(new_n11216_1, new_n11215, new_n11302);
nor_1  g10926(new_n11302, new_n11301, new_n11303);
not_4  g10927(new_n11303, new_n11304);
not_4  g10928(new_n10970, new_n11305);
nand_1 g10929(new_n10973, new_n11305, new_n11306);
nand_1 g10930(new_n11306, new_n10969, new_n11307);
nand_1 g10931(new_n11302, new_n11301, new_n11308);
nand_1 g10932(new_n11308, new_n11304, new_n11309);
not_4  g10933(new_n11309, new_n11310);
nand_1 g10934(new_n11310, new_n11307, new_n11311_1);
nand_1 g10935(new_n11311_1, new_n11304, new_n11312);
xnor_1 g10936(new_n11312, new_n11300, new_n11313);
xnor_1 g10937(new_n11313, new_n11143, new_n11314);
xnor_1 g10938(new_n11140, new_n11138, new_n11315);
not_4  g10939(new_n11307, new_n11316);
nand_1 g10940(new_n11309, new_n11316, new_n11317);
nand_1 g10941(new_n11317, new_n11311_1, new_n11318);
nor_1  g10942(new_n11318, new_n11315, new_n11319);
not_4  g10943(new_n11319, new_n11320);
nand_1 g10944(new_n10984, new_n10976, new_n11321);
nand_1 g10945(new_n11318, new_n11315, new_n11322);
nand_1 g10946(new_n11322, new_n11320, new_n11323);
nor_1  g10947(new_n11323, new_n11321, new_n11324);
not_4  g10948(new_n11324, new_n11325);
nand_1 g10949(new_n11325, new_n11320, new_n11326_1);
not_4  g10950(new_n11326_1, new_n11327);
nor_1  g10951(new_n11327, new_n11314, new_n11328);
not_4  g10952(new_n11328, new_n11329);
nand_1 g10953(new_n11327, new_n11314, new_n11330);
nand_1 g10954(new_n11330, new_n11329, new_n11331);
not_4  g10955(new_n11331, new_n11332);
nand_1 g10956(new_n11332, new_n11074, new_n11333);
nand_1 g10957(new_n11331, new_n11073, new_n11334);
nand_1 g10958(new_n11334, new_n11333, new_n11335);
not_4  g10959(new_n11067, new_n11336);
nand_1 g10960(new_n11069, new_n11336, new_n11337);
nand_1 g10961(new_n11337, new_n11071, new_n11338);
nand_1 g10962(new_n11323, new_n11321, new_n11339);
nand_1 g10963(new_n11339, new_n11325, new_n11340);
nor_1  g10964(new_n11340, new_n11338, new_n11341);
not_4  g10965(new_n11341, new_n11342);
nand_1 g10966(new_n11340, new_n11338, new_n11343);
nand_1 g10967(new_n11343, new_n11342, new_n11344);
nor_1  g10968(new_n10986, new_n10891, new_n11345);
nor_1  g10969(new_n11345, new_n10889, new_n11346);
not_4  g10970(new_n11346, new_n11347);
nor_1  g10971(new_n11347, new_n11344, new_n11348);
not_4  g10972(new_n11348, new_n11349);
nand_1 g10973(new_n11349, new_n11342, new_n11350);
not_4  g10974(new_n11350, new_n11351);
nor_1  g10975(new_n11351, new_n11335, new_n11352);
not_4  g10976(new_n11352, new_n11353);
nand_1 g10977(new_n11353, new_n11333, new_n11354);
not_4  g10978(new_n11354, new_n11355);
not_4  g10979(new_n11102, new_n11356);
nand_1 g10980(new_n11131, new_n11356, new_n11357);
nand_1 g10981(new_n11142, new_n11132, new_n11358);
nand_1 g10982(new_n11358, new_n11357, new_n11359);
not_4  g10983(new_n11359, new_n11360);
nand_1 g10984(new_n11313, new_n11143, new_n11361);
nand_1 g10985(new_n11329, new_n11361, new_n11362);
nand_1 g10986(new_n11042, new_n11006, new_n11363);
not_4  g10987(new_n11043, new_n11364);
nand_1 g10988(new_n11050, new_n11364, new_n11365);
nand_1 g10989(new_n11365, new_n11363, new_n11366);
nand_1 g10990(n11662, n4312, new_n11367);
xnor_1 g10991(new_n11367, new_n11366, new_n11368);
not_4  g10992(new_n11090, new_n11369);
nand_1 g10993(new_n11115, new_n11369, new_n11370);
nand_1 g10994(new_n11122, new_n11116, new_n11371);
nand_1 g10995(new_n11371, new_n11370, new_n11372);
nand_1 g10996(n12299, n10278, new_n11373);
xnor_1 g10997(new_n11373, new_n11372, new_n11374);
nand_1 g10998(new_n11109, new_n11108, new_n11375);
nand_1 g10999(new_n11111, new_n11107, new_n11376);
nand_1 g11000(new_n11376, new_n11375, new_n11377);
nand_1 g11001(n10451, n7436, new_n11378);
nand_1 g11002(n9241, n3022, new_n11379);
xnor_1 g11003(new_n11379, new_n11378, new_n11380);
nand_1 g11004(n11257, n3932, new_n11381);
nand_1 g11005(n10327, n1097, new_n11382);
xnor_1 g11006(new_n11382, new_n11381, new_n11383);
xnor_1 g11007(new_n11383, new_n11380, new_n11384);
xnor_1 g11008(new_n11384, new_n11377, new_n11385);
nand_1 g11009(new_n11289, new_n11288, new_n11386);
nand_1 g11010(new_n11291, new_n11287, new_n11387);
nand_1 g11011(new_n11387, new_n11386, new_n11388);
nand_1 g11012(n2393, n159, new_n11389);
nand_1 g11013(n5860, n2749, new_n11390);
xnor_1 g11014(new_n11390, new_n11389, new_n11391);
xnor_1 g11015(new_n11391, new_n11388, new_n11392);
xnor_1 g11016(new_n11392, new_n11385, new_n11393);
xnor_1 g11017(new_n11393, new_n11374, new_n11394);
xnor_1 g11018(new_n11394, new_n11368, new_n11395);
nor_1  g11019(new_n11207, new_n11171, new_n11396);
nor_1  g11020(new_n11218, new_n11208, new_n11397);
nor_1  g11021(new_n11397, new_n11396, new_n11398);
xnor_1 g11022(new_n11398, new_n11395, new_n11399);
nor_1  g11023(new_n11264, new_n11229, new_n11400);
nor_1  g11024(new_n11295, new_n11265, new_n11401);
nor_1  g11025(new_n11401, new_n11400, new_n11402);
nand_1 g11026(new_n11270, new_n11266, new_n11403);
nand_1 g11027(new_n11403, new_n11268, new_n11404);
not_4  g11028(new_n11404, new_n11405);
nand_1 g11029(n12247, n7388, new_n11406);
not_4  g11030(new_n11406, new_n11407_1);
nand_1 g11031(new_n11407_1, new_n11405, new_n11408);
nand_1 g11032(new_n11407_1, new_n11220, new_n11409);
nand_1 g11033(new_n11409, new_n11404, new_n11410);
nand_1 g11034(new_n11410, new_n11408, new_n11411);
nand_1 g11035(n10898, n5857, new_n11412);
nand_1 g11036(n12591, n12025, new_n11413);
nand_1 g11037(n11876, n45, new_n11414);
xnor_1 g11038(new_n11414, new_n11413, new_n11415);
xnor_1 g11039(new_n11415, new_n11412, new_n11416);
xnor_1 g11040(new_n11416, new_n11411, new_n11417);
xnor_1 g11041(new_n11417, new_n11402, new_n11418);
nand_1 g11042(new_n11119, new_n11118, new_n11419);
nand_1 g11043(new_n11121, new_n11117, new_n11420);
nand_1 g11044(new_n11420, new_n11419, new_n11421);
nand_1 g11045(n12705, n7456, new_n11422);
nand_1 g11046(n11023, n8276, new_n11423_1);
xnor_1 g11047(new_n11423_1, new_n11422, new_n11424);
xnor_1 g11048(new_n11424, new_n11421, new_n11425);
nand_1 g11049(n9583, n5964, new_n11426);
nand_1 g11050(n12511, n7965, new_n11427);
xnor_1 g11051(new_n11427, new_n11426, new_n11428);
xnor_1 g11052(new_n11428, new_n11425, new_n11429);
nand_1 g11053(new_n11128, new_n11127, new_n11430);
not_4  g11054(new_n11125, new_n11431);
nand_1 g11055(new_n11130, new_n11431, new_n11432);
nand_1 g11056(new_n11432, new_n11430, new_n11433);
not_4  g11057(new_n11106, new_n11434);
nor_1  g11058(new_n11112, new_n11434, new_n11435);
not_4  g11059(new_n11113, new_n11436);
nor_1  g11060(new_n11124, new_n11436, new_n11437);
nor_1  g11061(new_n11437, new_n11435, new_n11438);
xnor_1 g11062(new_n11438, new_n11433, new_n11439);
xnor_1 g11063(new_n11439, new_n11429, new_n11440);
xnor_1 g11064(new_n11440, new_n11418, new_n11441);
not_4  g11065(new_n11441, new_n11442);
nand_1 g11066(new_n11297, new_n11250, new_n11443);
nand_1 g11067(new_n11298, new_n11260, new_n11444);
nand_1 g11068(new_n11444, new_n11443, new_n11445);
nand_1 g11069(new_n11204, new_n11202, new_n11446);
nand_1 g11070(new_n11206, new_n11200, new_n11447);
nand_1 g11071(new_n11447, new_n11446, new_n11448);
not_4  g11072(new_n11040, new_n11449);
nand_1 g11073(new_n11449, new_n11034, new_n11450);
nand_1 g11074(new_n11051, new_n11041, new_n11451);
nand_1 g11075(new_n11451, new_n11450, new_n11452);
xnor_1 g11076(new_n11452, new_n11448, new_n11453);
nand_1 g11077(n3986, n3754, new_n11454);
nand_1 g11078(n11423, n6776, new_n11455);
xnor_1 g11079(new_n11455, new_n11454, new_n11456);
nand_1 g11080(n8759, n2278, new_n11457);
nand_1 g11081(n10510, n9640, new_n11458);
xnor_1 g11082(new_n11458, new_n11457, new_n11459);
xnor_1 g11083(new_n11459, new_n11456, new_n11460);
nand_1 g11084(n8476, n4094, new_n11461);
nand_1 g11085(n5305, n753, new_n11462);
xnor_1 g11086(new_n11462, new_n11461, new_n11463);
nand_1 g11087(n3616, n1067, new_n11464);
nand_1 g11088(n10644, n6703, new_n11465);
not_4  g11089(new_n11465, new_n11466);
xnor_1 g11090(new_n11466, new_n11464, new_n11467);
xnor_1 g11091(new_n11467, new_n11463, new_n11468);
xnor_1 g11092(new_n11468, new_n11460, new_n11469);
nand_1 g11093(new_n11037, new_n11036, new_n11470);
nand_1 g11094(new_n11039, new_n11035, new_n11471);
nand_1 g11095(new_n11471, new_n11470, new_n11472);
nand_1 g11096(new_n11047, new_n11046, new_n11473);
nand_1 g11097(new_n11049, new_n11044, new_n11474);
nand_1 g11098(new_n11474, new_n11473, new_n11475);
xnor_1 g11099(new_n11475, new_n11472, new_n11476);
xnor_1 g11100(new_n11476, new_n11469, new_n11477);
xnor_1 g11101(new_n11477, new_n11453, new_n11478_1);
nand_1 g11102(new_n11058, new_n11052, new_n11479);
nand_1 g11103(new_n11479, new_n11055, new_n11480);
not_4  g11104(new_n11271, new_n11481);
nand_1 g11105(new_n11276, new_n11481, new_n11482);
not_4  g11106(new_n11294, new_n11483);
nand_1 g11107(new_n11483, new_n11277, new_n11484);
nand_1 g11108(new_n11484, new_n11482, new_n11485);
nand_1 g11109(new_n11292, new_n11286, new_n11486);
nand_1 g11110(new_n11486, new_n11283, new_n11487);
nand_1 g11111(new_n11182, new_n11181, new_n11488);
nand_1 g11112(new_n11184, new_n11180, new_n11489);
nand_1 g11113(new_n11489, new_n11488, new_n11490);
nand_1 g11114(n10547, n1798, new_n11491);
nand_1 g11115(n8665, n7690, new_n11492);
xnor_1 g11116(new_n11492, new_n11491, new_n11493);
nand_1 g11117(n12826, n2530, new_n11494);
nand_1 g11118(n11892, n1510, new_n11495);
xnor_1 g11119(new_n11495, new_n11494, new_n11496);
xnor_1 g11120(new_n11496, new_n11493, new_n11497);
xnor_1 g11121(new_n11497, new_n11490, new_n11498);
xnor_1 g11122(new_n11498, new_n11487, new_n11499);
xnor_1 g11123(new_n11499, new_n11485, new_n11500);
not_4  g11124(new_n11500, new_n11501);
nand_1 g11125(n11922, n10545, new_n11502);
not_4  g11126(new_n11191, new_n11503);
nand_1 g11127(new_n11198, new_n11503, new_n11504);
nand_1 g11128(new_n11199, new_n11187, new_n11505);
nand_1 g11129(new_n11505, new_n11504, new_n11506);
xnor_1 g11130(new_n11506, new_n11502, new_n11507);
not_4  g11131(new_n11179, new_n11508);
nand_1 g11132(new_n11185, new_n11508, new_n11509);
nand_1 g11133(new_n11509, new_n11177, new_n11510);
nand_1 g11134(new_n11194, new_n11193, new_n11511);
nand_1 g11135(new_n11196, new_n11192, new_n11512);
nand_1 g11136(new_n11512, new_n11511, new_n11513);
xnor_1 g11137(new_n11513, new_n11510, new_n11514);
nand_1 g11138(n12648, n2551, new_n11515);
nand_1 g11139(n10685, n5331, new_n11516);
nand_1 g11140(n5645, n4499, new_n11517);
xnor_1 g11141(new_n11517, new_n11516, new_n11518);
xnor_1 g11142(new_n11518, new_n11515, new_n11519);
xnor_1 g11143(new_n11519, new_n11514, new_n11520);
xnor_1 g11144(new_n11520, new_n11507, new_n11521);
xnor_1 g11145(new_n11521, new_n11501, new_n11522);
nor_1  g11146(new_n11522, new_n11480, new_n11523);
not_4  g11147(new_n11480, new_n11524);
xnor_1 g11148(new_n11521, new_n11500, new_n11525);
nor_1  g11149(new_n11525, new_n11524, new_n11526);
nor_1  g11150(new_n11526, new_n11523, new_n11527);
nand_1 g11151(new_n11527, new_n11478_1, new_n11528);
not_4  g11152(new_n11478_1, new_n11529);
nand_1 g11153(new_n11525, new_n11524, new_n11530);
nand_1 g11154(new_n11522, new_n11480, new_n11531);
nand_1 g11155(new_n11531, new_n11530, new_n11532);
nand_1 g11156(new_n11532, new_n11529, new_n11533);
nand_1 g11157(new_n11533, new_n11528, new_n11534);
nor_1  g11158(new_n11534, new_n11445, new_n11535);
not_4  g11159(new_n11445, new_n11536_1);
nor_1  g11160(new_n11532, new_n11529, new_n11537);
nor_1  g11161(new_n11527, new_n11478_1, new_n11538);
nor_1  g11162(new_n11538, new_n11537, new_n11539);
nor_1  g11163(new_n11539, new_n11536_1, new_n11540);
nor_1  g11164(new_n11540, new_n11535, new_n11541);
nand_1 g11165(new_n11541, new_n11442, new_n11542);
nand_1 g11166(new_n11539, new_n11536_1, new_n11543);
nand_1 g11167(new_n11534, new_n11445, new_n11544);
nand_1 g11168(new_n11544, new_n11543, new_n11545);
nand_1 g11169(new_n11545, new_n11441, new_n11546);
nand_1 g11170(new_n11546, new_n11542, new_n11547);
nor_1  g11171(new_n11547, new_n11399, new_n11548);
not_4  g11172(new_n11399, new_n11549);
nor_1  g11173(new_n11545, new_n11441, new_n11550);
nor_1  g11174(new_n11541, new_n11442, new_n11551);
nor_1  g11175(new_n11551, new_n11550, new_n11552);
nor_1  g11176(new_n11552, new_n11549, new_n11553);
nor_1  g11177(new_n11553, new_n11548, new_n11554);
not_4  g11178(new_n11059, new_n11555);
nor_1  g11179(new_n11555, new_n11031, new_n11556);
not_4  g11180(new_n11060, new_n11557);
nor_1  g11181(new_n11072, new_n11557, new_n11558);
nor_1  g11182(new_n11558, new_n11556, new_n11559);
nand_1 g11183(new_n11299, new_n11219, new_n11560);
not_4  g11184(new_n11560, new_n11561);
not_4  g11185(new_n11312, new_n11562);
nor_1  g11186(new_n11562, new_n11300, new_n11563);
nor_1  g11187(new_n11563, new_n11561, new_n11564);
xnor_1 g11188(new_n11564, new_n11559, new_n11565);
not_4  g11189(new_n11565, new_n11566);
nand_1 g11190(new_n11566, new_n11554, new_n11567);
nand_1 g11191(new_n11552, new_n11549, new_n11568);
nand_1 g11192(new_n11547, new_n11399, new_n11569);
nand_1 g11193(new_n11569, new_n11568, new_n11570);
nand_1 g11194(new_n11565, new_n11570, new_n11571);
nand_1 g11195(new_n11571, new_n11567, new_n11572);
nor_1  g11196(new_n11572, new_n11362, new_n11573);
not_4  g11197(new_n11362, new_n11574);
nor_1  g11198(new_n11565, new_n11570, new_n11575);
nor_1  g11199(new_n11566, new_n11554, new_n11576);
nor_1  g11200(new_n11576, new_n11575, new_n11577);
nor_1  g11201(new_n11577, new_n11574, new_n11578);
nor_1  g11202(new_n11578, new_n11573, new_n11579);
nand_1 g11203(new_n11579, new_n11360, new_n11580);
nand_1 g11204(new_n11577, new_n11574, new_n11581);
nand_1 g11205(new_n11572, new_n11362, new_n11582);
nand_1 g11206(new_n11582, new_n11581, new_n11583);
nand_1 g11207(new_n11583, new_n11359, new_n11584);
nand_1 g11208(new_n11584, new_n11580, new_n11585);
nor_1  g11209(new_n11585, new_n11355, new_n11586);
nor_1  g11210(new_n11583, new_n11359, new_n11587);
nor_1  g11211(new_n11579, new_n11360, new_n11588);
nor_1  g11212(new_n11588, new_n11587, new_n11589);
nor_1  g11213(new_n11589, new_n11354, new_n11590);
nor_1  g11214(new_n11590, new_n11586, n4230);
nand_1 g11215(new_n6574, new_n6573, new_n11592);
nand_1 g11216(new_n11592, new_n6576, n4300);
nand_1 g11217(new_n3913, new_n3912, new_n11594);
nand_1 g11218(new_n11594, new_n3915, n4326);
nand_1 g11219(n6687, n5320, new_n11596);
nor_1  g11220(new_n1347, new_n1338, new_n11597);
nor_1  g11221(new_n1353_1, new_n1348, new_n11598);
nor_1  g11222(new_n11598, new_n11597, new_n11599);
not_4  g11223(new_n11599, new_n11600);
xnor_1 g11224(new_n11600, new_n11596, new_n11601);
nand_1 g11225(n4370, n2564, new_n11602);
not_4  g11226(new_n11602, new_n11603);
nand_1 g11227(new_n1351, new_n1350, new_n11604);
not_4  g11228(new_n1352, new_n11605);
nand_1 g11229(new_n11605, new_n1349, new_n11606);
nand_1 g11230(new_n11606, new_n11604, new_n11607);
xnor_1 g11231(new_n11607, new_n11603, new_n11608);
nand_1 g11232(n6770, n5212, new_n11609);
nand_1 g11233(n11877, n4189, new_n11610);
nand_1 g11234(n11407, n9920, new_n11611);
not_4  g11235(new_n11611, new_n11612);
xnor_1 g11236(new_n11612, new_n11610, new_n11613);
xnor_1 g11237(new_n11613, new_n11609, new_n11614);
not_4  g11238(new_n11614, new_n11615);
xnor_1 g11239(new_n11615, new_n11608, new_n11616);
xnor_1 g11240(new_n11616, new_n11601, new_n11617);
not_4  g11241(new_n11617, new_n11618);
xnor_1 g11242(new_n11618, new_n1363, new_n11619);
not_4  g11243(new_n11619, new_n11620);
not_4  g11244(new_n1488, new_n11621);
nand_1 g11245(new_n11621, new_n1487, new_n11622);
nand_1 g11246(n8336, n2433, new_n11623);
nand_1 g11247(n10928, n8819, new_n11624);
nand_1 g11248(new_n1480, new_n1473, new_n11625);
nand_1 g11249(new_n11625, new_n1477, new_n11626);
nor_1  g11250(new_n11626, new_n11624, new_n11627);
not_4  g11251(new_n11627, new_n11628);
nand_1 g11252(new_n11626, new_n11624, new_n11629);
nand_1 g11253(new_n11629, new_n11628, new_n11630);
nand_1 g11254(n11728, n2226, new_n11631);
not_4  g11255(new_n11631, new_n11632);
nand_1 g11256(n12709, n1094, new_n11633);
nand_1 g11257(new_n11633, new_n1400, new_n11634);
not_4  g11258(new_n11633, new_n11635);
nand_1 g11259(new_n11635, new_n1401, new_n11636);
nand_1 g11260(new_n11636, new_n11634, new_n11637);
xnor_1 g11261(new_n11637, new_n11632, new_n11638);
xnor_1 g11262(new_n11638, new_n11630, new_n11639);
xnor_1 g11263(new_n11639, new_n11623, new_n11640);
not_4  g11264(new_n1472, new_n11641);
nand_1 g11265(new_n1482, new_n11641, new_n11642);
nand_1 g11266(new_n1485, new_n1483, new_n11643);
nand_1 g11267(new_n11643, new_n11642, new_n11644);
xnor_1 g11268(new_n11644, new_n11640, new_n11645);
not_4  g11269(new_n11645, new_n11646);
xnor_1 g11270(new_n11646, new_n11622, new_n11647);
nand_1 g11271(new_n1551, new_n1489, new_n11648);
nor_1  g11272(new_n1558, new_n1552, new_n11649);
not_4  g11273(new_n11649, new_n11650);
nand_1 g11274(new_n11650, new_n11648, new_n11651);
xnor_1 g11275(new_n11651, new_n11647, new_n11652);
nand_1 g11276(n12069, n11967, new_n11653);
nand_1 g11277(n12391, n6254, new_n11654);
nand_1 g11278(new_n1499, new_n1498, new_n11655);
nand_1 g11279(new_n1501, new_n1497, new_n11656);
nand_1 g11280(new_n11656, new_n11655, new_n11657);
not_4  g11281(new_n11657, new_n11658);
xnor_1 g11282(new_n11658, new_n11654, new_n11659);
nand_1 g11283(n7160, n7159, new_n11660);
not_4  g11284(new_n11660, new_n11661);
nand_1 g11285(n12777, n7891, new_n11662_1);
nand_1 g11286(n12489, n4828, new_n11663);
nand_1 g11287(new_n11663, new_n11662_1, new_n11664);
not_4  g11288(new_n11662_1, new_n11665);
not_4  g11289(new_n11663, new_n11666);
nand_1 g11290(new_n11666, new_n11665, new_n11667);
nand_1 g11291(new_n11667, new_n11664, new_n11668);
xnor_1 g11292(new_n11668, new_n11661, new_n11669);
nand_1 g11293(new_n11669, new_n11659, new_n11670);
not_4  g11294(new_n11670, new_n11671);
nor_1  g11295(new_n11669, new_n11659, new_n11672);
nor_1  g11296(new_n11672, new_n11671, new_n11673);
xnor_1 g11297(new_n11673, new_n11653, new_n11674);
nand_1 g11298(new_n1505, new_n1494, new_n11675);
xnor_1 g11299(new_n11675, new_n11674, new_n11676);
not_4  g11300(new_n11676, new_n11677);
xnor_1 g11301(new_n11677, new_n1511, new_n11678);
nand_1 g11302(n12947, n11222, new_n11679);
nand_1 g11303(n11791, n11153, new_n11680);
nand_1 g11304(new_n1528, new_n1521, new_n11681);
nand_1 g11305(new_n11681, new_n1525, new_n11682);
not_4  g11306(new_n11682, new_n11683);
xnor_1 g11307(new_n11683, new_n11680, new_n11684);
not_4  g11308(new_n11684, new_n11685);
nand_1 g11309(n5760, n996, new_n11686);
not_4  g11310(new_n11686, new_n11687);
nand_1 g11311(n5314, n1478, new_n11688);
nand_1 g11312(n10990, n5767, new_n11689);
nand_1 g11313(new_n11689, new_n11688, new_n11690);
not_4  g11314(new_n11688, new_n11691);
not_4  g11315(new_n11689, new_n11692);
nand_1 g11316(new_n11692, new_n11691, new_n11693);
nand_1 g11317(new_n11693, new_n11690, new_n11694);
xnor_1 g11318(new_n11694, new_n11687, new_n11695);
xnor_1 g11319(new_n11695, new_n11685, new_n11696);
xnor_1 g11320(new_n11696, new_n11679, new_n11697);
not_4  g11321(new_n11697, new_n11698);
nand_1 g11322(new_n1531, new_n1518, new_n11699);
xnor_1 g11323(new_n11699, new_n11698, new_n11700);
xnor_1 g11324(new_n11700, new_n1537, new_n11701);
nand_1 g11325(new_n1549, new_n1542, new_n11702);
xnor_1 g11326(new_n11702, new_n11701, new_n11703);
xnor_1 g11327(new_n11703, new_n11678, new_n11704);
nor_1  g11328(new_n11704, new_n11652, new_n11705);
not_4  g11329(new_n11705, new_n11706);
nand_1 g11330(new_n11704, new_n11652, new_n11707_1);
nand_1 g11331(new_n11707_1, new_n11706, new_n11708);
xnor_1 g11332(new_n11708, new_n11620, new_n11709);
not_4  g11333(new_n1365, new_n11710);
nand_1 g11334(new_n1469, new_n11710, new_n11711);
nand_1 g11335(new_n1559, new_n1470, new_n11712);
nand_1 g11336(new_n11712, new_n11711, new_n11713);
xnor_1 g11337(new_n11713, new_n11709, n4333);
nand_1 g11338(n11877, n11757, new_n11715);
nand_1 g11339(n5240, n5212, new_n11716);
not_4  g11340(new_n11716, new_n11717);
nand_1 g11341(n11821, n11407, new_n11718);
not_4  g11342(new_n11718, new_n11719);
nand_1 g11343(new_n11719, new_n11717, new_n11720);
nand_1 g11344(new_n11718, new_n11716, new_n11721);
nand_1 g11345(new_n11721, new_n11720, new_n11722);
xnor_1 g11346(new_n11722, new_n11715, new_n11723);
nand_1 g11347(n11407, n5240, new_n11724);
nand_1 g11348(n11877, n3172, new_n11725);
nand_1 g11349(new_n11725, new_n11724, new_n11726);
nand_1 g11350(n11757, n5212, new_n11727);
not_4  g11351(new_n11725, new_n11728_1);
xnor_1 g11352(new_n11728_1, new_n11724, new_n11729);
nand_1 g11353(new_n11729, new_n11727, new_n11730);
nand_1 g11354(new_n11730, new_n11726, new_n11731);
xnor_1 g11355(new_n11731, new_n11723, new_n11732);
nand_1 g11356(n5320, n1333, new_n11733);
nand_1 g11357(n4370, n3172, new_n11734);
not_4  g11358(new_n11734, new_n11735);
xnor_1 g11359(new_n11735, new_n11733, new_n11736);
xnor_1 g11360(new_n11736, new_n11732, new_n11737);
nand_1 g11361(n4370, n1333, new_n11738);
nand_1 g11362(n11877, n1333, new_n11739);
nand_1 g11363(n11757, n11407, new_n11740);
nand_1 g11364(new_n11740, new_n11739, new_n11741);
nand_1 g11365(n5212, n3172, new_n11742);
xnor_1 g11366(new_n11740, new_n11739, new_n11743);
not_4  g11367(new_n11743, new_n11744);
nand_1 g11368(new_n11744, new_n11742, new_n11745);
nand_1 g11369(new_n11745, new_n11741, new_n11746);
nor_1  g11370(new_n11746, new_n11738, new_n11747);
not_4  g11371(new_n11747, new_n11748);
xnor_1 g11372(new_n11746, new_n11738, new_n11749);
not_4  g11373(new_n11749, new_n11750);
xnor_1 g11374(new_n11729, new_n11727, new_n11751);
nand_1 g11375(new_n11751, new_n11750, new_n11752);
nand_1 g11376(new_n11752, new_n11748, new_n11753);
xnor_1 g11377(new_n11753, new_n11737, new_n11754);
nand_1 g11378(n7862, n5320, new_n11755_1);
not_4  g11379(new_n11751, new_n11756);
nand_1 g11380(new_n11756, new_n11749, new_n11757_1);
nand_1 g11381(new_n11757_1, new_n11752, new_n11758);
nand_1 g11382(new_n11758, new_n11755_1, new_n11759);
xnor_1 g11383(new_n11758, new_n11755_1, new_n11760);
not_4  g11384(new_n11760, new_n11761);
nand_1 g11385(n7862, n4370, new_n11762);
nand_1 g11386(n11407, n3172, new_n11763);
nand_1 g11387(n11877, n7862, new_n11764);
nand_1 g11388(new_n11764, new_n11763, new_n11765);
nand_1 g11389(n11407, n7862, new_n11766);
not_4  g11390(new_n11766, new_n11767);
nand_1 g11391(new_n11767, new_n11728_1, new_n11768);
nand_1 g11392(n5212, n1333, new_n11769);
nand_1 g11393(new_n11769, new_n11768, new_n11770);
nand_1 g11394(new_n11770, new_n11765, new_n11771);
nor_1  g11395(new_n11771, new_n11762, new_n11772);
xnor_1 g11396(new_n11771, new_n11762, new_n11773);
xnor_1 g11397(new_n11743, new_n11742, new_n11774);
nor_1  g11398(new_n11774, new_n11773, new_n11775);
nor_1  g11399(new_n11775, new_n11772, new_n11776);
nand_1 g11400(new_n11776, new_n11761, new_n11777);
nand_1 g11401(new_n11777, new_n11759, new_n11778);
nor_1  g11402(new_n11778, new_n11754, new_n11779);
not_4  g11403(new_n11732, new_n11780_1);
nand_1 g11404(new_n11736, new_n11780_1, new_n11781);
nor_1  g11405(new_n11734, new_n11733, new_n11782);
nand_1 g11406(new_n11753, new_n11737, new_n11783);
not_4  g11407(new_n11783, new_n11784);
xnor_1 g11408(new_n11784, new_n11782, new_n11785);
nand_1 g11409(new_n11785, new_n11781, new_n11786);
nand_1 g11410(n11757, n4370, new_n11787);
not_4  g11411(new_n11787, new_n11788);
xnor_1 g11412(new_n11788, new_n11720, new_n11789);
nand_1 g11413(n11821, n5212, new_n11790);
nand_1 g11414(n11877, n5240, new_n11791_1);
nand_1 g11415(n11407, n9080, new_n11792);
not_4  g11416(new_n11792, new_n11793);
xnor_1 g11417(new_n11793, new_n11791_1, new_n11794);
xnor_1 g11418(new_n11794, new_n11790, new_n11795);
xnor_1 g11419(new_n11795, new_n11789, new_n11796);
nand_1 g11420(new_n11722, new_n11715, new_n11797);
not_4  g11421(new_n11723, new_n11798);
nand_1 g11422(new_n11731, new_n11798, new_n11799);
nand_1 g11423(new_n11799, new_n11797, new_n11800);
nand_1 g11424(n12000, n1333, new_n11801);
nand_1 g11425(n5320, n3172, new_n11802);
nand_1 g11426(n9725, n7862, new_n11803);
not_4  g11427(new_n11803, new_n11804);
xnor_1 g11428(new_n11804, new_n11802, new_n11805);
xnor_1 g11429(new_n11805, new_n11801, new_n11806);
xnor_1 g11430(new_n11806, new_n11800, new_n11807);
xnor_1 g11431(new_n11807, new_n11796, new_n11808);
not_4  g11432(new_n11808, new_n11809);
xnor_1 g11433(new_n11809, new_n11786, new_n11810);
xnor_1 g11434(new_n11810, new_n11779, new_n11811);
not_4  g11435(new_n11811, new_n11812);
nand_1 g11436(n12000, n7862, new_n11813);
xnor_1 g11437(new_n11778, new_n11754, new_n11814);
nand_1 g11438(new_n11814, new_n11813, new_n11815);
xnor_1 g11439(new_n11774, new_n11773, new_n11816);
not_4  g11440(new_n11816, new_n11817);
nand_1 g11441(new_n11768, new_n11765, new_n11818);
not_4  g11442(new_n11818, new_n11819);
nand_1 g11443(n11407, n1333, new_n11820);
not_4  g11444(new_n11820, new_n11821_1);
nand_1 g11445(n7862, n5212, new_n11822);
not_4  g11446(new_n11822, new_n11823);
nand_1 g11447(new_n11823, new_n11821_1, new_n11824);
nor_1  g11448(new_n11824, new_n11819, new_n11825);
nand_1 g11449(new_n11825, new_n11817, new_n11826);
xnor_1 g11450(new_n11776, new_n11760, new_n11827);
nor_1  g11451(new_n11827, new_n11826, new_n11828);
not_4  g11452(new_n11828, new_n11829);
xnor_1 g11453(new_n11814, new_n11813, new_n11830);
not_4  g11454(new_n11830, new_n11831);
nand_1 g11455(new_n11831, new_n11829, new_n11832);
nand_1 g11456(new_n11832, new_n11815, new_n11833);
xnor_1 g11457(new_n11833, new_n11812, new_n11834);
nand_1 g11458(n8819, n6877, new_n11835);
nand_1 g11459(n12709, n2464, new_n11836);
not_4  g11460(new_n11836, new_n11837);
nand_1 g11461(n6877, n6429, new_n11838);
not_4  g11462(new_n11838, new_n11839);
nand_1 g11463(new_n11839, new_n11837, new_n11840);
nand_1 g11464(new_n11838, new_n11836, new_n11841);
nand_1 g11465(n11728, n9400, new_n11842);
not_4  g11466(new_n11842, new_n11843);
nand_1 g11467(new_n11843, new_n11841, new_n11844);
nand_1 g11468(new_n11844, new_n11840, new_n11845);
xnor_1 g11469(new_n11845, new_n11835, new_n11846);
nand_1 g11470(n11728, n2464, new_n11847);
not_4  g11471(new_n11847, new_n11848);
nand_1 g11472(n12709, n11311, new_n11849);
nand_1 g11473(n9400, n6429, new_n11850);
nand_1 g11474(new_n11850, new_n11849, new_n11851);
nor_1  g11475(new_n11850, new_n11849, new_n11852);
not_4  g11476(new_n11852, new_n11853);
nand_1 g11477(new_n11853, new_n11851, new_n11854);
xnor_1 g11478(new_n11854, new_n11848, new_n11855);
xnor_1 g11479(new_n11855, new_n11846, new_n11856);
not_4  g11480(new_n11856, new_n11857);
nand_1 g11481(new_n11841, new_n11840, new_n11858);
not_4  g11482(new_n11858, new_n11859);
nand_1 g11483(n12709, n9400, new_n11860);
not_4  g11484(new_n11860, new_n11861);
nand_1 g11485(n11728, n6877, new_n11862);
not_4  g11486(new_n11862, new_n11863);
nand_1 g11487(new_n11863, new_n11861, new_n11864);
nor_1  g11488(new_n11864, new_n11859, new_n11865);
nand_1 g11489(new_n11865, new_n11857, new_n11866);
not_4  g11490(new_n11866, new_n11867);
nand_1 g11491(n6877, n2433, new_n11868);
not_4  g11492(new_n11868, new_n11869);
nand_1 g11493(n9400, n8819, new_n11870);
nand_1 g11494(new_n11853, new_n11847, new_n11871);
nand_1 g11495(new_n11871, new_n11851, new_n11872);
nor_1  g11496(new_n11872, new_n11870, new_n11873);
not_4  g11497(new_n11873, new_n11874);
nand_1 g11498(new_n11872, new_n11870, new_n11875);
nand_1 g11499(new_n11875, new_n11874, new_n11876_1);
nand_1 g11500(n11728, n11311, new_n11877_1);
nand_1 g11501(n6429, n2464, new_n11878);
nand_1 g11502(n12709, n4187, new_n11879);
xnor_1 g11503(new_n11879, new_n11878, new_n11880);
xnor_1 g11504(new_n11880, new_n11877_1, new_n11881);
nor_1  g11505(new_n11881, new_n11876_1, new_n11882);
not_4  g11506(new_n11882, new_n11883);
nand_1 g11507(new_n11881, new_n11876_1, new_n11884);
nand_1 g11508(new_n11884, new_n11883, new_n11885);
not_4  g11509(new_n11885, new_n11886);
nand_1 g11510(new_n11886, new_n11869, new_n11887);
nand_1 g11511(new_n11885, new_n11868, new_n11888);
nand_1 g11512(new_n11888, new_n11887, new_n11889);
not_4  g11513(new_n11835, new_n11890);
nand_1 g11514(new_n11845, new_n11890, new_n11891);
nand_1 g11515(new_n11855, new_n11846, new_n11892_1);
nand_1 g11516(new_n11892_1, new_n11891, new_n11893);
xnor_1 g11517(new_n11893, new_n11889, new_n11894);
nand_1 g11518(new_n11894, new_n11867, new_n11895);
nand_1 g11519(n8717, n6877, new_n11896);
nand_1 g11520(n11311, n6429, new_n11897);
nand_1 g11521(n12709, n4203, new_n11898);
nand_1 g11522(n11728, n4187, new_n11899);
not_4  g11523(new_n11899, new_n11900);
xnor_1 g11524(new_n11900, new_n11898, new_n11901);
xnor_1 g11525(new_n11901, new_n11897, new_n11902);
nand_1 g11526(new_n11879, new_n11878, new_n11903);
not_4  g11527(new_n11880, new_n11904);
nand_1 g11528(new_n11904, new_n11877_1, new_n11905);
nand_1 g11529(new_n11905, new_n11903, new_n11906);
xnor_1 g11530(new_n11906, new_n11902, new_n11907);
nand_1 g11531(n9400, n2433, new_n11908);
nand_1 g11532(n8819, n2464, new_n11909);
not_4  g11533(new_n11909, new_n11910);
xnor_1 g11534(new_n11910, new_n11908, new_n11911);
xnor_1 g11535(new_n11911, new_n11907, new_n11912);
nand_1 g11536(new_n11883, new_n11874, new_n11913);
xnor_1 g11537(new_n11913, new_n11912, new_n11914);
not_4  g11538(new_n11889, new_n11915);
nand_1 g11539(new_n11893, new_n11915, new_n11916);
nand_1 g11540(new_n11916, new_n11887, new_n11917_1);
nand_1 g11541(new_n11917_1, new_n11914, new_n11918);
not_4  g11542(new_n11918, new_n11919_1);
nor_1  g11543(new_n11917_1, new_n11914, new_n11920);
nor_1  g11544(new_n11920, new_n11919_1, new_n11921);
xnor_1 g11545(new_n11921, new_n11896, new_n11922_1);
xnor_1 g11546(new_n11922_1, new_n11895, new_n11923);
xnor_1 g11547(new_n11894, new_n11866, new_n11924);
xnor_1 g11548(new_n11865, new_n11856, new_n11925);
nand_1 g11549(n12489, n4805, new_n11926);
not_4  g11550(new_n11926, new_n11927);
nand_1 g11551(n10990, n7236, new_n11928);
not_4  g11552(new_n11928, new_n11929);
nand_1 g11553(new_n11929, new_n11927, new_n11930);
not_4  g11554(new_n11930, new_n11931);
nand_1 g11555(n12489, n11478, new_n11932);
nand_1 g11556(n7159, n4805, new_n11933);
not_4  g11557(new_n11933, new_n11934);
xnor_1 g11558(new_n11934, new_n11932, new_n11935);
nor_1  g11559(new_n11935, new_n11931, new_n11936);
not_4  g11560(new_n11936, new_n11937);
xnor_1 g11561(new_n11935, new_n11930, new_n11938);
nand_1 g11562(n10990, n3992, new_n11939);
nand_1 g11563(n7236, n5760, new_n11940);
xnor_1 g11564(new_n11940, new_n11939, new_n11941);
nand_1 g11565(new_n11941, new_n11938, new_n11942);
nand_1 g11566(new_n11942, new_n11937, new_n11943);
nand_1 g11567(n10990, n8384, new_n11944);
not_4  g11568(new_n11944, new_n11945);
nand_1 g11569(n7236, n1478, new_n11946);
not_4  g11570(new_n11946, new_n11947);
nand_1 g11571(new_n11947, new_n11945, new_n11948);
nand_1 g11572(n5760, n3992, new_n11949);
not_4  g11573(new_n11949, new_n11950);
nand_1 g11574(new_n11950, new_n11928, new_n11951);
nand_1 g11575(new_n11946, new_n11944, new_n11952);
not_4  g11576(new_n11952, new_n11953);
nand_1 g11577(new_n11953, new_n11951, new_n11954);
nand_1 g11578(new_n11954, new_n11948, new_n11955);
nor_1  g11579(new_n11953, new_n11951, new_n11956);
nor_1  g11580(new_n11956, new_n11955, new_n11957);
not_4  g11581(new_n11957, new_n11958);
nand_1 g11582(new_n11958, new_n11943, new_n11959);
xnor_1 g11583(new_n11957, new_n11943, new_n11960);
nand_1 g11584(n11478, n7159, new_n11961);
not_4  g11585(new_n11961, new_n11962);
nand_1 g11586(new_n11962, new_n11926, new_n11963);
nand_1 g11587(n12489, n5283, new_n11964);
nand_1 g11588(n12777, n4805, new_n11965);
nand_1 g11589(new_n11965, new_n11964, new_n11966);
not_4  g11590(new_n11964, new_n11967_1);
not_4  g11591(new_n11965, new_n11968);
nand_1 g11592(new_n11968, new_n11967_1, new_n11969);
nand_1 g11593(new_n11969, new_n11966, new_n11970);
nand_1 g11594(new_n11970, new_n11963, new_n11971);
not_4  g11595(new_n11966, new_n11972);
nor_1  g11596(new_n11972, new_n11963, new_n11973);
not_4  g11597(new_n11973, new_n11974);
nand_1 g11598(new_n11974, new_n11971, new_n11975);
nand_1 g11599(new_n11975, new_n11960, new_n11976);
nand_1 g11600(new_n11976, new_n11959, new_n11977);
nand_1 g11601(n6254, n4805, new_n11978);
nand_1 g11602(new_n11966, new_n11962, new_n11979);
nand_1 g11603(new_n11979, new_n11969, new_n11980);
xnor_1 g11604(new_n11980, new_n11978, new_n11981);
nand_1 g11605(n7159, n5283, new_n11982);
not_4  g11606(new_n11982, new_n11983);
nand_1 g11607(n12489, n137, new_n11984);
nand_1 g11608(n12777, n11478, new_n11985);
xnor_1 g11609(new_n11985, new_n11984, new_n11986);
xnor_1 g11610(new_n11986, new_n11983, new_n11987);
nand_1 g11611(new_n11987, new_n11981, new_n11988);
not_4  g11612(new_n11988, new_n11989);
nor_1  g11613(new_n11987, new_n11981, new_n11990);
nor_1  g11614(new_n11990, new_n11989, new_n11991);
not_4  g11615(new_n11932, new_n11992);
nand_1 g11616(new_n11934, new_n11992, new_n11993);
not_4  g11617(new_n11993, new_n11994);
nand_1 g11618(new_n11970, new_n11994, new_n11995);
xnor_1 g11619(new_n11995, new_n11991, new_n11996);
nand_1 g11620(n11791, n7236, new_n11997);
nand_1 g11621(new_n11949, new_n11948, new_n11998);
nand_1 g11622(new_n11998, new_n11952, new_n11999_1);
xnor_1 g11623(new_n11999_1, new_n11997, new_n12000_1);
nand_1 g11624(n8384, n5760, new_n12001);
not_4  g11625(new_n12001, new_n12002);
nand_1 g11626(n10990, n6358, new_n12003);
nand_1 g11627(n3992, n1478, new_n12004);
xnor_1 g11628(new_n12004, new_n12003, new_n12005_1);
not_4  g11629(new_n12005_1, new_n12006);
xnor_1 g11630(new_n12006, new_n12002, new_n12007);
not_4  g11631(new_n12007, new_n12008);
xnor_1 g11632(new_n12008, new_n12000_1, new_n12009);
nand_1 g11633(new_n11955, new_n11950, new_n12010);
xnor_1 g11634(new_n12010, new_n12009, new_n12011);
not_4  g11635(new_n12011, new_n12012);
xnor_1 g11636(new_n12012, new_n11996, new_n12013);
xnor_1 g11637(new_n12013, new_n11977, new_n12014_1);
nand_1 g11638(new_n12014_1, new_n11925, new_n12015);
not_4  g11639(new_n11925, new_n12016);
xnor_1 g11640(new_n12014_1, new_n12016, new_n12017);
xnor_1 g11641(new_n11975, new_n11960, new_n12018);
not_4  g11642(new_n12018, new_n12019);
nand_1 g11643(n12709, n6877, new_n12020_1);
nand_1 g11644(new_n12020_1, new_n11843, new_n12021);
nand_1 g11645(new_n12021, new_n11858, new_n12022);
not_4  g11646(new_n12021, new_n12023);
nand_1 g11647(new_n12023, new_n11841, new_n12024);
nand_1 g11648(new_n12024, new_n12022, new_n12025_1);
nor_1  g11649(new_n12025_1, new_n12019, new_n12026);
not_4  g11650(new_n12026, new_n12027);
xnor_1 g11651(new_n12025_1, new_n12018, new_n12028);
xnor_1 g11652(new_n11941, new_n11938, new_n12029);
nand_1 g11653(new_n11862, new_n11860, new_n12030);
nand_1 g11654(new_n12030, new_n11864, new_n12031);
not_4  g11655(new_n12031, new_n12032);
nand_1 g11656(new_n12032, new_n12029, new_n12033);
not_4  g11657(new_n12020_1, new_n12034);
nand_1 g11658(new_n11928, new_n11926, new_n12035);
nand_1 g11659(new_n12035, new_n11930, new_n12036);
not_4  g11660(new_n12036, new_n12037);
nand_1 g11661(new_n12037, new_n12034, new_n12038);
not_4  g11662(new_n12038, new_n12039);
xnor_1 g11663(new_n12031, new_n12029, new_n12040);
nand_1 g11664(new_n12040, new_n12039, new_n12041);
nand_1 g11665(new_n12041, new_n12033, new_n12042);
nand_1 g11666(new_n12042, new_n12028, new_n12043);
nand_1 g11667(new_n12043, new_n12027, new_n12044_1);
nand_1 g11668(new_n12044_1, new_n12017, new_n12045);
nand_1 g11669(new_n12045, new_n12015, new_n12046);
nor_1  g11670(new_n12046, new_n11924, new_n12047);
xnor_1 g11671(new_n12046, new_n11924, new_n12048);
not_4  g11672(new_n11995, new_n12049);
nand_1 g11673(new_n12049, new_n11991, new_n12050);
nand_1 g11674(n7159, n137, new_n12051);
nand_1 g11675(n12777, n5283, new_n12052);
nand_1 g11676(n12489, n6294, new_n12053);
not_4  g11677(new_n12053, new_n12054);
xnor_1 g11678(new_n12054, new_n12052, new_n12055);
xnor_1 g11679(new_n12055, new_n12051, new_n12056);
not_4  g11680(new_n12056, new_n12057);
nand_1 g11681(n11478, n6254, new_n12058);
nand_1 g11682(new_n11985, new_n11984, new_n12059);
not_4  g11683(new_n12059, new_n12060);
nor_1  g11684(new_n11986, new_n11983, new_n12061);
nor_1  g11685(new_n12061, new_n12060, new_n12062);
xnor_1 g11686(new_n12062, new_n12058, new_n12063);
xnor_1 g11687(new_n12063, new_n12057, new_n12064);
not_4  g11688(new_n12064, new_n12065);
nand_1 g11689(n11967, n4805, new_n12066);
not_4  g11690(new_n12066, new_n12067);
not_4  g11691(new_n11978, new_n12068);
nand_1 g11692(new_n11980, new_n12068, new_n12069_1);
nand_1 g11693(new_n11988, new_n12069_1, new_n12070);
xnor_1 g11694(new_n12070, new_n12067, new_n12071);
xnor_1 g11695(new_n12071, new_n12065, new_n12072);
not_4  g11696(new_n12072, new_n12073);
xnor_1 g11697(new_n12073, new_n12050, new_n12074);
not_4  g11698(new_n12009, new_n12075);
nor_1  g11699(new_n12010, new_n12075, new_n12076_1);
nand_1 g11700(n6358, n5760, new_n12077);
nand_1 g11701(n8384, n1478, new_n12078);
nand_1 g11702(n10990, n5198, new_n12079);
not_4  g11703(new_n12079, new_n12080);
xnor_1 g11704(new_n12080, new_n12078, new_n12081);
xnor_1 g11705(new_n12081, new_n12077, new_n12082);
nand_1 g11706(n11791, n3992, new_n12083);
nand_1 g11707(new_n12004, new_n12003, new_n12084);
not_4  g11708(new_n12084, new_n12085);
nor_1  g11709(new_n12005_1, new_n12002, new_n12086);
nor_1  g11710(new_n12086, new_n12085, new_n12087);
xnor_1 g11711(new_n12087, new_n12083, new_n12088);
xnor_1 g11712(new_n12088, new_n12082, new_n12089);
nand_1 g11713(n12947, n7236, new_n12090);
nor_1  g11714(new_n11999_1, new_n11997, new_n12091);
nor_1  g11715(new_n12007, new_n12000_1, new_n12092);
nor_1  g11716(new_n12092, new_n12091, new_n12093);
not_4  g11717(new_n12093, new_n12094);
xnor_1 g11718(new_n12094, new_n12090, new_n12095);
not_4  g11719(new_n12095, new_n12096);
xnor_1 g11720(new_n12096, new_n12089, new_n12097);
xnor_1 g11721(new_n12097, new_n12076_1, new_n12098);
xnor_1 g11722(new_n12098, new_n12074, new_n12099);
not_4  g11723(new_n12099, new_n12100);
nor_1  g11724(new_n12011, new_n11996, new_n12101);
not_4  g11725(new_n12101, new_n12102);
nand_1 g11726(new_n12013, new_n11977, new_n12103);
nand_1 g11727(new_n12103, new_n12102, new_n12104);
xnor_1 g11728(new_n12104, new_n12100, new_n12105);
nor_1  g11729(new_n12105, new_n12048, new_n12106);
nor_1  g11730(new_n12106, new_n12047, new_n12107);
nor_1  g11731(new_n12107, new_n11923, new_n12108);
not_4  g11732(new_n12108, new_n12109);
not_4  g11733(new_n12076_1, new_n12110);
nor_1  g11734(new_n12097, new_n12110, new_n12111_1);
nand_1 g11735(n7236, n6441, new_n12112);
not_4  g11736(new_n12083, new_n12113);
nand_1 g11737(new_n12087, new_n12113, new_n12114);
nand_1 g11738(new_n12088, new_n12082, new_n12115);
nand_1 g11739(new_n12115, new_n12114, new_n12116);
nand_1 g11740(n12947, n3992, new_n12117);
nand_1 g11741(n11791, n8384, new_n12118);
xnor_1 g11742(new_n12118, new_n12117, new_n12119);
not_4  g11743(new_n12119, new_n12120);
xnor_1 g11744(new_n12120, new_n12116, new_n12121);
nand_1 g11745(n6358, n1478, new_n12122);
nand_1 g11746(n5760, n5198, new_n12123);
nand_1 g11747(n10990, n1471, new_n12124);
nand_1 g11748(new_n12124, new_n12123, new_n12125);
not_4  g11749(new_n12123, new_n12126);
not_4  g11750(new_n12124, new_n12127);
nand_1 g11751(new_n12127, new_n12126, new_n12128);
nand_1 g11752(new_n12128, new_n12125, new_n12129);
not_4  g11753(new_n12129, new_n12130);
xnor_1 g11754(new_n12130, new_n12122, new_n12131);
not_4  g11755(new_n12131, new_n12132);
nand_1 g11756(new_n12079, new_n12078, new_n12133);
nand_1 g11757(new_n12081, new_n12077, new_n12134);
nand_1 g11758(new_n12134, new_n12133, new_n12135);
nor_1  g11759(new_n12135, new_n12132, new_n12136);
not_4  g11760(new_n12136, new_n12137);
nand_1 g11761(new_n12135, new_n12132, new_n12138);
nand_1 g11762(new_n12138, new_n12137, new_n12139);
xnor_1 g11763(new_n12139, new_n12121, new_n12140);
nand_1 g11764(new_n12093, new_n12090, new_n12141);
nand_1 g11765(new_n12095, new_n12089, new_n12142);
nand_1 g11766(new_n12142, new_n12141, new_n12143);
nor_1  g11767(new_n12143, new_n12140, new_n12144);
not_4  g11768(new_n12144, new_n12145_1);
nand_1 g11769(new_n12143, new_n12140, new_n12146);
nand_1 g11770(new_n12146, new_n12145_1, new_n12147);
nor_1  g11771(new_n12147, new_n12112, new_n12148);
not_4  g11772(new_n12148, new_n12149);
nand_1 g11773(new_n12147, new_n12112, new_n12150);
nand_1 g11774(new_n12150, new_n12149, new_n12151);
not_4  g11775(new_n12151, new_n12152);
nand_1 g11776(new_n12152, new_n12111_1, new_n12153);
not_4  g11777(new_n12111_1, new_n12154);
nand_1 g11778(new_n12151, new_n12154, new_n12155);
nand_1 g11779(new_n12155, new_n12153, new_n12156);
nor_1  g11780(new_n12072, new_n12050, new_n12157);
nand_1 g11781(n4805, n447, new_n12158);
not_4  g11782(new_n12058, new_n12159);
nand_1 g11783(new_n12062, new_n12159, new_n12160);
nand_1 g11784(new_n12063, new_n12056, new_n12161);
nand_1 g11785(new_n12161, new_n12160, new_n12162);
nand_1 g11786(n11967, n11478, new_n12163);
nand_1 g11787(n6254, n5283, new_n12164);
xnor_1 g11788(new_n12164, new_n12163, new_n12165);
not_4  g11789(new_n12165, new_n12166);
xnor_1 g11790(new_n12166, new_n12162, new_n12167);
nand_1 g11791(n12777, n137, new_n12168);
nand_1 g11792(n7159, n6294, new_n12169);
nand_1 g11793(n12489, n6797, new_n12170);
nand_1 g11794(new_n12170, new_n12169, new_n12171);
not_4  g11795(new_n12169, new_n12172);
not_4  g11796(new_n12170, new_n12173);
nand_1 g11797(new_n12173, new_n12172, new_n12174);
nand_1 g11798(new_n12174, new_n12171, new_n12175);
not_4  g11799(new_n12175, new_n12176);
xnor_1 g11800(new_n12176, new_n12168, new_n12177);
not_4  g11801(new_n12177, new_n12178);
nand_1 g11802(new_n12053, new_n12052, new_n12179);
nand_1 g11803(new_n12055, new_n12051, new_n12180);
nand_1 g11804(new_n12180, new_n12179, new_n12181);
nor_1  g11805(new_n12181, new_n12178, new_n12182);
not_4  g11806(new_n12182, new_n12183);
nand_1 g11807(new_n12181, new_n12178, new_n12184);
nand_1 g11808(new_n12184, new_n12183, new_n12185);
not_4  g11809(new_n12185, new_n12186);
xnor_1 g11810(new_n12186, new_n12167, new_n12187);
nor_1  g11811(new_n12070, new_n12067, new_n12188);
nor_1  g11812(new_n12071, new_n12064, new_n12189);
nor_1  g11813(new_n12189, new_n12188, new_n12190);
nand_1 g11814(new_n12190, new_n12187, new_n12191);
not_4  g11815(new_n12191, new_n12192);
nor_1  g11816(new_n12190, new_n12187, new_n12193);
nor_1  g11817(new_n12193, new_n12192, new_n12194);
xnor_1 g11818(new_n12194, new_n12158, new_n12195);
nand_1 g11819(new_n12195, new_n12157, new_n12196);
not_4  g11820(new_n12157, new_n12197);
not_4  g11821(new_n12158, new_n12198);
xnor_1 g11822(new_n12194, new_n12198, new_n12199);
nand_1 g11823(new_n12199, new_n12197, new_n12200);
nand_1 g11824(new_n12200, new_n12196, new_n12201);
not_4  g11825(new_n12201, new_n12202);
nand_1 g11826(new_n12098, new_n12074, new_n12203);
nor_1  g11827(new_n12104, new_n12099, new_n12204);
not_4  g11828(new_n12204, new_n12205);
nand_1 g11829(new_n12205, new_n12203, new_n12206);
xnor_1 g11830(new_n12206, new_n12202, new_n12207);
xnor_1 g11831(new_n12207, new_n12156, new_n12208);
nand_1 g11832(new_n12107, new_n11923, new_n12209);
nand_1 g11833(new_n12209, new_n12109, new_n12210);
not_4  g11834(new_n12210, new_n12211);
nand_1 g11835(new_n12211, new_n12208, new_n12212);
nand_1 g11836(new_n12212, new_n12109, new_n12213);
nand_1 g11837(new_n11911, new_n11907, new_n12214);
nor_1  g11838(new_n11909, new_n11908, new_n12215);
not_4  g11839(new_n11912, new_n12216);
nand_1 g11840(new_n11913, new_n12216, new_n12217);
not_4  g11841(new_n12217, new_n12218);
xnor_1 g11842(new_n12218, new_n12215, new_n12219);
nand_1 g11843(new_n12219, new_n12214, new_n12220);
not_4  g11844(new_n11897, new_n12221_1);
nand_1 g11845(new_n11901, new_n12221_1, new_n12222);
not_4  g11846(new_n11906, new_n12223);
nand_1 g11847(new_n12223, new_n11902, new_n12224);
nand_1 g11848(new_n12224, new_n12222, new_n12225);
nand_1 g11849(n9400, n8717, new_n12226);
nand_1 g11850(n2464, n2433, new_n12227);
nand_1 g11851(n7730, n6877, new_n12228);
not_4  g11852(new_n12228, new_n12229);
xnor_1 g11853(new_n12229, new_n12227, new_n12230);
xnor_1 g11854(new_n12230, new_n12226, new_n12231);
xnor_1 g11855(new_n12231, new_n12225, new_n12232);
nor_1  g11856(new_n11899, new_n11898, new_n12233);
nand_1 g11857(n11311, n8819, new_n12234);
xnor_1 g11858(new_n12234, new_n12233, new_n12235);
nand_1 g11859(n11728, n4203, new_n12236);
nand_1 g11860(n6429, n4187, new_n12237);
nand_1 g11861(n12753, n12709, new_n12238);
not_4  g11862(new_n12238, new_n12239);
xnor_1 g11863(new_n12239, new_n12237, new_n12240);
xnor_1 g11864(new_n12240, new_n12236, new_n12241);
not_4  g11865(new_n12241, new_n12242);
xnor_1 g11866(new_n12242, new_n12235, new_n12243);
xnor_1 g11867(new_n12243, new_n12232, new_n12244);
xnor_1 g11868(new_n12244, new_n12220, new_n12245);
not_4  g11869(new_n12245, new_n12246);
xnor_1 g11870(new_n12246, new_n11918, new_n12247_1);
not_4  g11871(new_n11896, new_n12248);
nand_1 g11872(new_n11921, new_n12248, new_n12249);
not_4  g11873(new_n11895, new_n12250);
nand_1 g11874(new_n11922_1, new_n12250, new_n12251);
nand_1 g11875(new_n12251, new_n12249, new_n12252);
xnor_1 g11876(new_n12252, new_n12247_1, new_n12253);
not_4  g11877(new_n12253, new_n12254);
nand_1 g11878(n11478, n447, new_n12255);
nand_1 g11879(n11967, n5283, new_n12256);
not_4  g11880(new_n12256, new_n12257);
nand_1 g11881(n4805, n1353, new_n12258);
xnor_1 g11882(new_n12258, new_n12257, new_n12259);
xnor_1 g11883(new_n12259, new_n12255, new_n12260);
not_4  g11884(new_n12260, new_n12261);
not_4  g11885(new_n12168, new_n12262);
nand_1 g11886(new_n12176, new_n12262, new_n12263);
nand_1 g11887(new_n12183, new_n12263, new_n12264);
xnor_1 g11888(new_n12264, new_n12261, new_n12265);
nand_1 g11889(n6254, n137, new_n12266);
xnor_1 g11890(new_n12266, new_n12174, new_n12267);
nand_1 g11891(n7159, n6797, new_n12268);
nand_1 g11892(n12777, n6294, new_n12269);
nand_1 g11893(n12489, n3146, new_n12270);
nand_1 g11894(new_n12270, new_n12269, new_n12271);
not_4  g11895(new_n12269, new_n12272);
not_4  g11896(new_n12270, new_n12273);
nand_1 g11897(new_n12273, new_n12272, new_n12274);
nand_1 g11898(new_n12274, new_n12271, new_n12275);
xnor_1 g11899(new_n12275, new_n12268, new_n12276);
not_4  g11900(new_n12276, new_n12277);
xnor_1 g11901(new_n12277, new_n12267, new_n12278);
xnor_1 g11902(new_n12278, new_n12265, new_n12279);
nand_1 g11903(new_n12166, new_n12162, new_n12280);
nor_1  g11904(new_n12164, new_n12163, new_n12281);
nor_1  g11905(new_n12185, new_n12167, new_n12282);
xnor_1 g11906(new_n12282, new_n12281, new_n12283);
nand_1 g11907(new_n12283, new_n12280, new_n12284);
xnor_1 g11908(new_n12284, new_n12279, new_n12285);
xnor_1 g11909(new_n12285, new_n12192, new_n12286);
nand_1 g11910(new_n12194, new_n12198, new_n12287);
nand_1 g11911(new_n12196, new_n12287, new_n12288);
not_4  g11912(new_n12288, new_n12289);
nor_1  g11913(new_n12289, new_n12286, new_n12290);
xnor_1 g11914(new_n12285, new_n12191, new_n12291);
nor_1  g11915(new_n12288, new_n12291, new_n12292);
nor_1  g11916(new_n12292, new_n12290, new_n12293);
not_4  g11917(new_n12122, new_n12294);
nand_1 g11918(new_n12130, new_n12294, new_n12295);
nand_1 g11919(new_n12137, new_n12295, new_n12296);
nand_1 g11920(n6441, n3992, new_n12297);
nand_1 g11921(n12947, n8384, new_n12298);
nand_1 g11922(n11999, n7236, new_n12299_1);
not_4  g11923(new_n12299_1, new_n12300);
xnor_1 g11924(new_n12300, new_n12298, new_n12301);
xnor_1 g11925(new_n12301, new_n12297, new_n12302);
not_4  g11926(new_n12302, new_n12303);
xnor_1 g11927(new_n12303, new_n12296, new_n12304);
not_4  g11928(new_n12128, new_n12305);
nand_1 g11929(n11791, n6358, new_n12306);
not_4  g11930(new_n12306, new_n12307);
nand_1 g11931(new_n12307, new_n12305, new_n12308);
nand_1 g11932(new_n12306, new_n12128, new_n12309);
nand_1 g11933(new_n12309, new_n12308, new_n12310);
nand_1 g11934(n5760, n1471, new_n12311);
nand_1 g11935(n5198, n1478, new_n12312);
nand_1 g11936(n10990, n7646, new_n12313);
not_4  g11937(new_n12313, new_n12314);
xnor_1 g11938(new_n12314, new_n12312, new_n12315);
xnor_1 g11939(new_n12315, new_n12311, new_n12316);
xnor_1 g11940(new_n12316, new_n12310, new_n12317);
xnor_1 g11941(new_n12317, new_n12304, new_n12318);
nand_1 g11942(new_n12120, new_n12116, new_n12319);
nor_1  g11943(new_n12118, new_n12117, new_n12320);
nor_1  g11944(new_n12139, new_n12121, new_n12321);
xnor_1 g11945(new_n12321, new_n12320, new_n12322);
nand_1 g11946(new_n12322, new_n12319, new_n12323);
xnor_1 g11947(new_n12323, new_n12318, new_n12324);
xnor_1 g11948(new_n12324, new_n12145_1, new_n12325);
nand_1 g11949(new_n12153, new_n12149, new_n12326);
nor_1  g11950(new_n12326, new_n12325, new_n12327);
xnor_1 g11951(new_n12324, new_n12144, new_n12328);
not_4  g11952(new_n12326, new_n12329);
nor_1  g11953(new_n12329, new_n12328, new_n12330);
nor_1  g11954(new_n12330, new_n12327, new_n12331);
nand_1 g11955(new_n12331, new_n12293, new_n12332);
nand_1 g11956(new_n12288, new_n12291, new_n12333);
nand_1 g11957(new_n12289, new_n12286, new_n12334);
nand_1 g11958(new_n12334, new_n12333, new_n12335);
nand_1 g11959(new_n12329, new_n12328, new_n12336);
nand_1 g11960(new_n12326, new_n12325, new_n12337);
nand_1 g11961(new_n12337, new_n12336, new_n12338);
nand_1 g11962(new_n12338, new_n12335, new_n12339);
nand_1 g11963(new_n12339, new_n12332, new_n12340);
nor_1  g11964(new_n12206, new_n12202, new_n12341);
not_4  g11965(new_n12156, new_n12342);
nor_1  g11966(new_n12207, new_n12342, new_n12343);
nor_1  g11967(new_n12343, new_n12341, new_n12344);
not_4  g11968(new_n12344, new_n12345);
nor_1  g11969(new_n12345, new_n12340, new_n12346);
nor_1  g11970(new_n12338, new_n12335, new_n12347);
nor_1  g11971(new_n12331, new_n12293, new_n12348);
nor_1  g11972(new_n12348, new_n12347, new_n12349);
nor_1  g11973(new_n12344, new_n12349, new_n12350);
nor_1  g11974(new_n12350, new_n12346, new_n12351);
nor_1  g11975(new_n12351, new_n12254, new_n12352);
nand_1 g11976(new_n12344, new_n12349, new_n12353);
nand_1 g11977(new_n12345, new_n12340, new_n12354);
nand_1 g11978(new_n12354, new_n12353, new_n12355);
nor_1  g11979(new_n12355, new_n12253, new_n12356);
nor_1  g11980(new_n12356, new_n12352, new_n12357);
nand_1 g11981(new_n12357, new_n12213, new_n12358);
not_4  g11982(new_n12213, new_n12359);
nand_1 g11983(new_n12355, new_n12253, new_n12360);
nand_1 g11984(new_n12351, new_n12254, new_n12361);
nand_1 g11985(new_n12361, new_n12360, new_n12362);
nand_1 g11986(new_n12362, new_n12359, new_n12363);
nand_1 g11987(new_n12363, new_n12358, new_n12364);
nor_1  g11988(new_n12364, new_n11834, new_n12365);
not_4  g11989(new_n11834, new_n12366);
nor_1  g11990(new_n12362, new_n12359, new_n12367);
nor_1  g11991(new_n12357, new_n12213, new_n12368);
nor_1  g11992(new_n12368, new_n12367, new_n12369);
nand_1 g11993(new_n12369, new_n12366, new_n12370);
nand_1 g11994(new_n12364, new_n11834, new_n12371);
nand_1 g11995(new_n12371, new_n12370, new_n12372);
xnor_1 g11996(new_n11831, new_n11828, new_n12373);
nand_1 g11997(new_n11827, new_n11826, new_n12374);
nand_1 g11998(new_n12374, new_n11829, new_n12375);
not_4  g11999(new_n12105, new_n12376);
xnor_1 g12000(new_n12376, new_n12048, new_n12377);
nand_1 g12001(new_n12377, new_n12375, new_n12378);
not_4  g12002(new_n12378, new_n12379);
nor_1  g12003(new_n12377, new_n12375, new_n12380);
nor_1  g12004(new_n12380, new_n12379, new_n12381);
xnor_1 g12005(new_n11825, new_n11816, new_n12382);
not_4  g12006(new_n12017, new_n12383);
xnor_1 g12007(new_n12044_1, new_n12383, new_n12384);
nor_1  g12008(new_n12384, new_n12382, new_n12385);
xnor_1 g12009(new_n12042, new_n12028, new_n12386);
not_4  g12010(new_n12386, new_n12387);
nor_1  g12011(new_n11769, new_n11767, new_n12388);
not_4  g12012(new_n12388, new_n12389);
nor_1  g12013(new_n12389, new_n11765, new_n12390);
not_4  g12014(new_n12390, new_n12391_1);
nand_1 g12015(new_n12389, new_n11819, new_n12392);
nand_1 g12016(new_n12392, new_n12391_1, new_n12393);
nor_1  g12017(new_n12393, new_n12387, new_n12394);
not_4  g12018(new_n12394, new_n12395);
xnor_1 g12019(new_n12393, new_n12386, new_n12396);
xnor_1 g12020(new_n12037, new_n12020_1, new_n12397);
nand_1 g12021(new_n12397, new_n11767, new_n12398);
nand_1 g12022(new_n11822, new_n11820, new_n12399);
nand_1 g12023(new_n12399, new_n11824, new_n12400);
nand_1 g12024(new_n12400, new_n12398, new_n12401);
xnor_1 g12025(new_n12040, new_n12038, new_n12402);
xnor_1 g12026(new_n12400, new_n12398, new_n12403);
nor_1  g12027(new_n12403, new_n12402, new_n12404);
not_4  g12028(new_n12404, new_n12405);
nand_1 g12029(new_n12405, new_n12401, new_n12406);
nand_1 g12030(new_n12406, new_n12396, new_n12407);
nand_1 g12031(new_n12407, new_n12395, new_n12408);
not_4  g12032(new_n12408, new_n12409);
xnor_1 g12033(new_n12384, new_n12382, new_n12410);
nor_1  g12034(new_n12410, new_n12409, new_n12411);
nor_1  g12035(new_n12411, new_n12385, new_n12412);
not_4  g12036(new_n12412, new_n12413);
nand_1 g12037(new_n12413, new_n12381, new_n12414);
nand_1 g12038(new_n12414, new_n12378, new_n12415);
nand_1 g12039(new_n12415, new_n12373, new_n12416);
xnor_1 g12040(new_n12210, new_n12208, new_n12417);
not_4  g12041(new_n12417, new_n12418);
xnor_1 g12042(new_n12415, new_n12373, new_n12419);
nor_1  g12043(new_n12419, new_n12418, new_n12420);
not_4  g12044(new_n12420, new_n12421);
nand_1 g12045(new_n12421, new_n12416, new_n12422);
not_4  g12046(new_n12422, new_n12423);
nor_1  g12047(new_n12423, new_n12372, new_n12424);
nor_1  g12048(new_n12424, new_n12365, new_n12425);
nand_1 g12049(new_n12360, new_n12359, new_n12426);
nand_1 g12050(new_n12426, new_n12361, new_n12427);
nand_1 g12051(new_n11810, new_n11779, new_n12428);
not_4  g12052(new_n11833, new_n12429);
nand_1 g12053(new_n12429, new_n11812, new_n12430);
nand_1 g12054(new_n12430, new_n12428, new_n12431);
nand_1 g12055(new_n12282, new_n12281, new_n12432);
not_4  g12056(new_n12279, new_n12433);
nand_1 g12057(new_n12284, new_n12433, new_n12434);
nand_1 g12058(new_n12434, new_n12432, new_n12435);
nand_1 g12059(new_n12299_1, new_n12298, new_n12436);
nand_1 g12060(new_n12301, new_n12297, new_n12437);
nand_1 g12061(new_n12437, new_n12436, new_n12438);
nand_1 g12062(n4805, n4436, new_n12439);
nand_1 g12063(n8384, n6441, new_n12440);
nand_1 g12064(n11791, n5198, new_n12441);
xnor_1 g12065(new_n12441, new_n12440, new_n12442);
xnor_1 g12066(new_n12442, new_n12439, new_n12443);
xnor_1 g12067(new_n12443, new_n12438, new_n12444_1);
nand_1 g12068(n7159, n3146, new_n12445);
nand_1 g12069(n11967, n137, new_n12446);
xnor_1 g12070(new_n12446, new_n12445, new_n12447);
nand_1 g12071(n6294, n6254, new_n12448);
nand_1 g12072(n12947, n6358, new_n12449);
xnor_1 g12073(new_n12449, new_n12448, new_n12450);
nand_1 g12074(n11407, n6826, new_n12451);
nand_1 g12075(n7862, n6604, new_n12452);
xnor_1 g12076(new_n12452, new_n12451, new_n12453);
xnor_1 g12077(new_n12453, new_n12450, new_n12454);
xnor_1 g12078(new_n12454, new_n12447, new_n12455);
xnor_1 g12079(new_n12455, new_n12444_1, new_n12456);
nand_1 g12080(n6429, n4203, new_n12457);
nor_1  g12081(new_n12266, new_n12174, new_n12458);
nor_1  g12082(new_n12276, new_n12267, new_n12459);
nor_1  g12083(new_n12459, new_n12458, new_n12460);
xnor_1 g12084(new_n12460, new_n12457, new_n12461);
xnor_1 g12085(new_n12461, new_n12456, new_n12462);
nor_1  g12086(new_n12264, new_n12260, new_n12463);
not_4  g12087(new_n12265, new_n12464);
nor_1  g12088(new_n12278, new_n12464, new_n12465);
nor_1  g12089(new_n12465, new_n12463, new_n12466);
nor_1  g12090(new_n12302, new_n12296, new_n12467);
not_4  g12091(new_n12304, new_n12468);
nor_1  g12092(new_n12317, new_n12468, new_n12469);
nor_1  g12093(new_n12469, new_n12467, new_n12470);
nand_1 g12094(n11478, n1353, new_n12471);
not_4  g12095(new_n12471, new_n12472);
nand_1 g12096(new_n12259, new_n12255, new_n12473);
nand_1 g12097(new_n12473, new_n12257, new_n12474);
not_4  g12098(new_n12474, new_n12475);
nand_1 g12099(new_n12475, new_n12472, new_n12476);
nand_1 g12100(new_n12472, new_n12158, new_n12477);
nand_1 g12101(new_n12477, new_n12474, new_n12478);
nand_1 g12102(new_n12478, new_n12476, new_n12479);
not_4  g12103(new_n12268, new_n12480);
nand_1 g12104(new_n12271, new_n12480, new_n12481);
nand_1 g12105(new_n12481, new_n12274, new_n12482);
xnor_1 g12106(new_n12482, new_n12479, new_n12483);
xnor_1 g12107(new_n12483, new_n12470, new_n12484);
xnor_1 g12108(new_n12484, new_n12466, new_n12485);
xnor_1 g12109(new_n12485, new_n12462, new_n12486);
not_4  g12110(new_n12486, new_n12487);
nand_1 g12111(new_n11784, new_n11782, new_n12488);
nand_1 g12112(new_n11808, new_n11786, new_n12489_1);
nand_1 g12113(new_n12489_1, new_n12488, new_n12490);
nand_1 g12114(n12777, n6797, new_n12491);
xnor_1 g12115(new_n12491, new_n12490, new_n12492);
xnor_1 g12116(new_n12492, new_n12487, new_n12493);
xnor_1 g12117(new_n12493, new_n12435, new_n12494);
xnor_1 g12118(new_n12494, new_n12431, new_n12495);
xnor_1 g12119(new_n12495, new_n12427, new_n12496);
nand_1 g12120(new_n12246, new_n11919_1, new_n12497);
nand_1 g12121(new_n12252, new_n12247_1, new_n12498);
nand_1 g12122(new_n12498, new_n12497, new_n12499);
nand_1 g12123(new_n12285, new_n12192, new_n12500);
nand_1 g12124(new_n12333, new_n12500, new_n12501);
xnor_1 g12125(new_n12501, new_n12499, new_n12502);
nand_1 g12126(new_n12324, new_n12144, new_n12503);
nand_1 g12127(new_n12337, new_n12503, new_n12504);
nand_1 g12128(new_n12231, new_n12225, new_n12505);
not_4  g12129(new_n12232, new_n12506);
nand_1 g12130(new_n12243, new_n12506, new_n12507);
nand_1 g12131(new_n12507, new_n12505, new_n12508);
nand_1 g12132(new_n12228, new_n12227, new_n12509);
nand_1 g12133(new_n12230, new_n12226, new_n12510);
nand_1 g12134(new_n12510, new_n12509, new_n12511_1);
nand_1 g12135(n5283, n447, new_n12512);
nand_1 g12136(n11999, n3992, new_n12513);
not_4  g12137(new_n12513, new_n12514);
xnor_1 g12138(new_n12514, new_n12512, new_n12515);
xnor_1 g12139(new_n12515, new_n12511_1, new_n12516);
xnor_1 g12140(new_n12516, new_n12508, new_n12517);
nand_1 g12141(n7646, n5760, new_n12518);
nand_1 g12142(n10990, n4722, new_n12519);
xnor_1 g12143(new_n12519, new_n12518, new_n12520);
xnor_1 g12144(new_n12520, new_n12517, new_n12521);
xnor_1 g12145(new_n12521, new_n12504, new_n12522);
xnor_1 g12146(new_n12522, new_n12502, new_n12523);
nor_1  g12147(new_n12346, new_n12347, new_n12524);
nand_1 g12148(new_n12218, new_n12215, new_n12525);
nand_1 g12149(new_n12244, new_n12220, new_n12526);
nand_1 g12150(new_n12526, new_n12525, new_n12527);
not_4  g12151(new_n11806, new_n12528);
nand_1 g12152(new_n12528, new_n11800, new_n12529);
nand_1 g12153(new_n11807, new_n11796, new_n12530);
nand_1 g12154(new_n12530, new_n12529, new_n12531);
nand_1 g12155(new_n12238, new_n12237, new_n12532);
nand_1 g12156(new_n12240, new_n12236, new_n12533);
nand_1 g12157(new_n12533, new_n12532, new_n12534);
nand_1 g12158(n12000, n3172, new_n12535);
nand_1 g12159(n9725, n1333, new_n12536);
nand_1 g12160(n12709, n10174, new_n12537);
xnor_1 g12161(new_n12537, new_n12536, new_n12538);
xnor_1 g12162(new_n12538, new_n12535, new_n12539);
xnor_1 g12163(new_n12539, new_n12534, new_n12540);
not_4  g12164(new_n12234, new_n12541);
nand_1 g12165(new_n12541, new_n12233, new_n12542);
nand_1 g12166(new_n12241, new_n12235, new_n12543);
nand_1 g12167(new_n12543, new_n12542, new_n12544);
nand_1 g12168(new_n12313, new_n12312, new_n12545);
nand_1 g12169(new_n12315, new_n12311, new_n12546);
nand_1 g12170(new_n12546, new_n12545, new_n12547);
nand_1 g12171(n6877, n1198, new_n12548);
nand_1 g12172(n12753, n11728, new_n12549);
not_4  g12173(new_n12549, new_n12550);
xnor_1 g12174(new_n12550, new_n12548, new_n12551);
xnor_1 g12175(new_n12551, new_n12547, new_n12552);
xnor_1 g12176(new_n12552, new_n12544, new_n12553);
xnor_1 g12177(new_n12553, new_n12540, new_n12554);
xnor_1 g12178(new_n12554, new_n12531, new_n12555);
nand_1 g12179(n12489, n4938, new_n12556);
nand_1 g12180(new_n11803, new_n11802, new_n12557);
nand_1 g12181(new_n11805, new_n11801, new_n12558);
nand_1 g12182(new_n12558, new_n12557, new_n12559);
nand_1 g12183(n11757, n5320, new_n12560);
nand_1 g12184(n9080, n5212, new_n12561);
xnor_1 g12185(new_n12561, new_n12560, new_n12562);
nand_1 g12186(n11877, n11821, new_n12563);
nand_1 g12187(n5240, n4370, new_n12564);
xnor_1 g12188(new_n12564, new_n12563, new_n12565);
xnor_1 g12189(new_n12565, new_n12562, new_n12566);
xnor_1 g12190(new_n12566, new_n12559, new_n12567);
nand_1 g12191(n9400, n7730, new_n12568);
nand_1 g12192(n11311, n2433, new_n12569);
not_4  g12193(new_n12569, new_n12570);
xnor_1 g12194(new_n12570, new_n12568, new_n12571);
xnor_1 g12195(new_n12571, new_n12567, new_n12572);
nand_1 g12196(new_n11792, new_n11791_1, new_n12573);
nand_1 g12197(new_n11794, new_n11790, new_n12574);
nand_1 g12198(new_n12574, new_n12573, new_n12575);
nand_1 g12199(new_n11787, new_n11720, new_n12576);
not_4  g12200(new_n11795, new_n12577);
nand_1 g12201(new_n12577, new_n11789, new_n12578);
nand_1 g12202(new_n12578, new_n12576, new_n12579);
xnor_1 g12203(new_n12579, new_n12575, new_n12580);
xnor_1 g12204(new_n12580, new_n12572, new_n12581);
xnor_1 g12205(new_n12581, new_n12556, new_n12582);
xnor_1 g12206(new_n12582, new_n12555, new_n12583);
xnor_1 g12207(new_n12583, new_n12527, new_n12584);
nand_1 g12208(new_n12321, new_n12320, new_n12585);
not_4  g12209(new_n12318, new_n12586);
nand_1 g12210(new_n12323, new_n12586, new_n12587);
nand_1 g12211(new_n12587, new_n12585, new_n12588);
nand_1 g12212(n8819, n4187, new_n12589);
nand_1 g12213(n1478, n1471, new_n12590);
xnor_1 g12214(new_n12590, new_n12589, new_n12591_1);
nand_1 g12215(n8717, n2464, new_n12592);
nand_1 g12216(n10022, n7236, new_n12593);
xnor_1 g12217(new_n12593, new_n12592, new_n12594);
xnor_1 g12218(new_n12594, new_n12591_1, new_n12595);
not_4  g12219(new_n12310, new_n12596);
nand_1 g12220(new_n12316, new_n12596, new_n12597);
nand_1 g12221(new_n12597, new_n12308, new_n12598);
xnor_1 g12222(new_n12598, new_n12595, new_n12599);
xnor_1 g12223(new_n12599, new_n12588, new_n12600);
xnor_1 g12224(new_n12600, new_n12584, new_n12601);
xnor_1 g12225(new_n12601, new_n12524, new_n12602);
xnor_1 g12226(new_n12602, new_n12523, new_n12603);
xnor_1 g12227(new_n12603, new_n12496, new_n12604);
not_4  g12228(new_n12604, new_n12605);
nand_1 g12229(new_n12605, new_n12425, new_n12606);
nor_1  g12230(new_n12369, new_n12366, new_n12607);
nor_1  g12231(new_n12607, new_n12365, new_n12608);
nand_1 g12232(new_n12422, new_n12608, new_n12609);
nand_1 g12233(new_n12609, new_n12370, new_n12610);
nand_1 g12234(new_n12604, new_n12610, new_n12611);
nand_1 g12235(new_n12611, new_n12606, n4378);
xnor_1 g12236(new_n4203_1, new_n4086_1, n4397);
xnor_1 g12237(new_n4533, new_n4300_1, n4553);
xnor_1 g12238(new_n927, new_n918, n4686);
xnor_1 g12239(new_n10425, new_n10404, n4689);
xnor_1 g12240(new_n5627, new_n5489, n4733);
nand_1 g12241(new_n2278_1, new_n2268, new_n12618);
nand_1 g12242(new_n12618, new_n2280, n4757);
xnor_1 g12243(new_n5484, new_n5483, n4971);
xnor_1 g12244(new_n7331, new_n7330, n5030);
xnor_1 g12245(new_n3169, new_n3136, n5034);
nand_1 g12246(new_n3160, new_n3148, new_n12623);
nand_1 g12247(new_n12623, new_n3162, n5094);
not_4  g12248(new_n11607, new_n12625);
nand_1 g12249(new_n12625, new_n11603, new_n12626);
nand_1 g12250(new_n11614, new_n11608, new_n12627);
nand_1 g12251(new_n12627, new_n12626, new_n12628);
nand_1 g12252(n5320, n2564, new_n12629);
nand_1 g12253(n4370, n4189, new_n12630);
xnor_1 g12254(new_n12630, new_n12629, new_n12631);
not_4  g12255(new_n12631, new_n12632);
xnor_1 g12256(new_n12632, new_n12628, new_n12633);
nand_1 g12257(n11877, n6770, new_n12634);
nand_1 g12258(new_n11611, new_n11610, new_n12635);
nand_1 g12259(new_n11613, new_n11609, new_n12636);
nand_1 g12260(new_n12636, new_n12635, new_n12637);
not_4  g12261(new_n12637, new_n12638);
xnor_1 g12262(new_n12638, new_n12634, new_n12639);
nand_1 g12263(n9920, n5212, new_n12640);
nand_1 g12264(n11407, n3627, new_n12641);
nand_1 g12265(new_n12641, new_n12640, new_n12642);
not_4  g12266(new_n12640, new_n12643);
not_4  g12267(new_n12641, new_n12644);
nand_1 g12268(new_n12644, new_n12643, new_n12645);
nand_1 g12269(new_n12645, new_n12642, new_n12646);
xnor_1 g12270(new_n12646, new_n12639, new_n12647);
xnor_1 g12271(new_n12647, new_n12633, new_n12648_1);
nor_1  g12272(new_n11599, new_n11596, new_n12649);
not_4  g12273(new_n12649, new_n12650);
nand_1 g12274(new_n11616, new_n11601, new_n12651);
nand_1 g12275(new_n12651, new_n12650, new_n12652);
nand_1 g12276(new_n12652, new_n12648_1, new_n12653);
nor_1  g12277(new_n12637, new_n12634, new_n12654);
not_4  g12278(new_n12654, new_n12655);
not_4  g12279(new_n12646, new_n12656);
nand_1 g12280(new_n12656, new_n12639, new_n12657);
nand_1 g12281(new_n12657, new_n12655, new_n12658);
nand_1 g12282(n12000, n2564, new_n12659);
nand_1 g12283(n5320, n4189, new_n12660);
nand_1 g12284(n9725, n6687, new_n12661);
nand_1 g12285(new_n12661, new_n12660, new_n12662);
not_4  g12286(new_n12660, new_n12663);
not_4  g12287(new_n12661, new_n12664);
nand_1 g12288(new_n12664, new_n12663, new_n12665);
nand_1 g12289(new_n12665, new_n12662, new_n12666);
xnor_1 g12290(new_n12666, new_n12659, new_n12667);
xnor_1 g12291(new_n12667, new_n12658, new_n12668);
nand_1 g12292(n6770, n4370, new_n12669);
nand_1 g12293(new_n12669, new_n12645, new_n12670);
not_4  g12294(new_n12645, new_n12671);
not_4  g12295(new_n12669, new_n12672);
nand_1 g12296(new_n12672, new_n12671, new_n12673);
nand_1 g12297(new_n12673, new_n12670, new_n12674);
nand_1 g12298(n5212, n3627, new_n12675);
nand_1 g12299(n11877, n9920, new_n12676);
nand_1 g12300(n11407, n4516, new_n12677);
nand_1 g12301(new_n12677, new_n12676, new_n12678);
not_4  g12302(new_n12676, new_n12679);
not_4  g12303(new_n12677, new_n12680);
nand_1 g12304(new_n12680, new_n12679, new_n12681);
nand_1 g12305(new_n12681, new_n12678, new_n12682);
xnor_1 g12306(new_n12682, new_n12675, new_n12683);
not_4  g12307(new_n12683, new_n12684);
xnor_1 g12308(new_n12684, new_n12674, new_n12685);
xnor_1 g12309(new_n12685, new_n12668, new_n12686);
not_4  g12310(new_n12686, new_n12687);
nand_1 g12311(new_n12632, new_n12628, new_n12688);
nor_1  g12312(new_n12630, new_n12629, new_n12689);
not_4  g12313(new_n12647, new_n12690);
nor_1  g12314(new_n12690, new_n12633, new_n12691);
xnor_1 g12315(new_n12691, new_n12689, new_n12692);
nand_1 g12316(new_n12692, new_n12688, new_n12693);
xnor_1 g12317(new_n12693, new_n12687, new_n12694);
xnor_1 g12318(new_n12694, new_n12653, new_n12695);
nand_1 g12319(n12000, n6687, new_n12696);
xnor_1 g12320(new_n12652, new_n12648_1, new_n12697);
nor_1  g12321(new_n12697, new_n12696, new_n12698);
nand_1 g12322(new_n11618, new_n1362, new_n12699);
xnor_1 g12323(new_n12697, new_n12696, new_n12700);
nor_1  g12324(new_n12700, new_n12699, new_n12701);
nor_1  g12325(new_n12701, new_n12698, new_n12702);
xnor_1 g12326(new_n12702, new_n12695, new_n12703);
nand_1 g12327(n8717, n8336, new_n12704_1);
not_4  g12328(new_n12704_1, new_n12705_1);
nand_1 g12329(n6429, n2226, new_n12706_1);
not_4  g12330(new_n12706_1, new_n12707);
nand_1 g12331(n11728, n1094, new_n12708);
nand_1 g12332(n12709, n10678, new_n12709_1);
not_4  g12333(new_n12709_1, new_n12710);
xnor_1 g12334(new_n12710, new_n12708, new_n12711);
xnor_1 g12335(new_n12711, new_n12707, new_n12712);
nand_1 g12336(new_n11636, new_n11631, new_n12713);
nand_1 g12337(new_n12713, new_n11634, new_n12714);
nor_1  g12338(new_n12714, new_n12712, new_n12715);
not_4  g12339(new_n12715, new_n12716);
nand_1 g12340(new_n12714, new_n12712, new_n12717);
nand_1 g12341(new_n12717, new_n12716, new_n12718);
nand_1 g12342(n10928, n2433, new_n12719);
nand_1 g12343(n8819, n6986, new_n12720_1);
not_4  g12344(new_n12720_1, new_n12721);
xnor_1 g12345(new_n12721, new_n12719, new_n12722);
xnor_1 g12346(new_n12722, new_n12718, new_n12723);
not_4  g12347(new_n11630, new_n12724);
nand_1 g12348(new_n11638, new_n12724, new_n12725);
nand_1 g12349(new_n12725, new_n11628, new_n12726);
xnor_1 g12350(new_n12726, new_n12723, new_n12727);
not_4  g12351(new_n11623, new_n12728);
nand_1 g12352(new_n11639, new_n12728, new_n12729);
nand_1 g12353(new_n11644, new_n11640, new_n12730);
nand_1 g12354(new_n12730, new_n12729, new_n12731);
xnor_1 g12355(new_n12731, new_n12727, new_n12732);
nand_1 g12356(new_n12732, new_n12705_1, new_n12733);
not_4  g12357(new_n11622, new_n12734);
nand_1 g12358(new_n11646, new_n12734, new_n12735);
not_4  g12359(new_n12735, new_n12736);
xnor_1 g12360(new_n12732, new_n12704_1, new_n12737);
nand_1 g12361(new_n12737, new_n12736, new_n12738);
nand_1 g12362(new_n12738, new_n12733, new_n12739);
not_4  g12363(new_n12727, new_n12740);
nand_1 g12364(new_n12731, new_n12740, new_n12741);
nand_1 g12365(new_n12711, new_n12707, new_n12742);
nand_1 g12366(new_n12716, new_n12742, new_n12743);
nand_1 g12367(n10928, n8717, new_n12744);
not_4  g12368(new_n12744, new_n12745);
nand_1 g12369(n6986, n2433, new_n12746);
nand_1 g12370(n8336, n7730, new_n12747);
not_4  g12371(new_n12747, new_n12748);
xnor_1 g12372(new_n12748, new_n12746, new_n12749);
xnor_1 g12373(new_n12749, new_n12745, new_n12750);
xnor_1 g12374(new_n12750, new_n12743, new_n12751);
not_4  g12375(new_n12708, new_n12752);
nand_1 g12376(new_n12710, new_n12752, new_n12753_1);
nand_1 g12377(n8819, n2226, new_n12754);
nand_1 g12378(new_n12754, new_n12753_1, new_n12755);
not_4  g12379(new_n12753_1, new_n12756);
not_4  g12380(new_n12754, new_n12757);
nand_1 g12381(new_n12757, new_n12756, new_n12758);
nand_1 g12382(new_n12758, new_n12755, new_n12759);
not_4  g12383(new_n12759, new_n12760);
nand_1 g12384(n11728, n10678, new_n12761);
nand_1 g12385(n6429, n1094, new_n12762);
nand_1 g12386(n12709, n7320, new_n12763);
not_4  g12387(new_n12763, new_n12764);
xnor_1 g12388(new_n12764, new_n12762, new_n12765);
xnor_1 g12389(new_n12765, new_n12761, new_n12766);
not_4  g12390(new_n12766, new_n12767);
xnor_1 g12391(new_n12767, new_n12760, new_n12768);
xnor_1 g12392(new_n12768, new_n12751, new_n12769);
not_4  g12393(new_n12718, new_n12770);
nand_1 g12394(new_n12722, new_n12770, new_n12771);
nor_1  g12395(new_n12720_1, new_n12719, new_n12772);
nand_1 g12396(new_n12726, new_n12723, new_n12773);
not_4  g12397(new_n12773, new_n12774);
xnor_1 g12398(new_n12774, new_n12772, new_n12775);
nand_1 g12399(new_n12775, new_n12771, new_n12776);
xnor_1 g12400(new_n12776, new_n12769, new_n12777_1);
xnor_1 g12401(new_n12777_1, new_n12741, new_n12778);
xnor_1 g12402(new_n12778, new_n12739, new_n12779);
xnor_1 g12403(new_n12737, new_n12735, new_n12780);
not_4  g12404(new_n12780, new_n12781);
nand_1 g12405(new_n11651, new_n11647, new_n12782);
nand_1 g12406(new_n11706, new_n12782, new_n12783);
not_4  g12407(new_n12783, new_n12784);
nand_1 g12408(new_n12784, new_n12781, new_n12785);
not_4  g12409(new_n1537, new_n12786);
nand_1 g12410(new_n11700, new_n12786, new_n12787);
nand_1 g12411(n11222, n6441, new_n12788);
not_4  g12412(new_n11680, new_n12789);
nand_1 g12413(new_n11683, new_n12789, new_n12790);
nand_1 g12414(new_n11695, new_n11684, new_n12791);
nand_1 g12415(new_n12791, new_n12790, new_n12792);
nand_1 g12416(n12947, n11153, new_n12793);
nand_1 g12417(n11791, n5314, new_n12794);
xnor_1 g12418(new_n12794, new_n12793, new_n12795);
not_4  g12419(new_n12795, new_n12796);
xnor_1 g12420(new_n12796, new_n12792, new_n12797);
nand_1 g12421(n1478, n996, new_n12798);
nand_1 g12422(n10990, n5319, new_n12799);
nand_1 g12423(n5767, n5760, new_n12800);
nand_1 g12424(new_n12800, new_n12799, new_n12801);
not_4  g12425(new_n12799, new_n12802);
not_4  g12426(new_n12800, new_n12803);
nand_1 g12427(new_n12803, new_n12802, new_n12804);
nand_1 g12428(new_n12804, new_n12801, new_n12805);
not_4  g12429(new_n12805, new_n12806);
xnor_1 g12430(new_n12806, new_n12798, new_n12807_1);
nand_1 g12431(new_n11693, new_n11686, new_n12808);
nand_1 g12432(new_n12808, new_n11690, new_n12809);
xnor_1 g12433(new_n12809, new_n12807_1, new_n12810);
not_4  g12434(new_n12810, new_n12811);
xnor_1 g12435(new_n12811, new_n12797, new_n12812);
not_4  g12436(new_n11679, new_n12813);
nand_1 g12437(new_n11696, new_n12813, new_n12814);
nand_1 g12438(new_n11699, new_n11697, new_n12815);
nand_1 g12439(new_n12815, new_n12814, new_n12816);
xnor_1 g12440(new_n12816, new_n12812, new_n12817);
xnor_1 g12441(new_n12817, new_n12788, new_n12818);
xnor_1 g12442(new_n12818, new_n12787, new_n12819);
nand_1 g12443(new_n11677, new_n1510_1, new_n12820);
not_4  g12444(new_n12820, new_n12821);
nand_1 g12445(n12069, n447, new_n12822);
not_4  g12446(new_n12822, new_n12823);
nand_1 g12447(n12777, n7160, new_n12824);
not_4  g12448(new_n12824, new_n12825);
nand_1 g12449(n7159, n4828, new_n12826_1);
nand_1 g12450(n12489, n2515, new_n12827);
not_4  g12451(new_n12827, new_n12828);
xnor_1 g12452(new_n12828, new_n12826_1, new_n12829);
xnor_1 g12453(new_n12829, new_n12825, new_n12830);
nand_1 g12454(new_n11667, new_n11660, new_n12831);
nand_1 g12455(new_n12831, new_n11664, new_n12832);
nor_1  g12456(new_n12832, new_n12830, new_n12833);
not_4  g12457(new_n12833, new_n12834);
nand_1 g12458(new_n12832, new_n12830, new_n12835);
nand_1 g12459(new_n12835, new_n12834, new_n12836);
nand_1 g12460(n12391, n11967, new_n12837);
nand_1 g12461(n7891, n6254, new_n12838);
not_4  g12462(new_n12838, new_n12839);
xnor_1 g12463(new_n12839, new_n12837, new_n12840);
xnor_1 g12464(new_n12840, new_n12836, new_n12841);
nor_1  g12465(new_n11657, new_n11654, new_n12842);
nor_1  g12466(new_n11671, new_n12842, new_n12843);
xnor_1 g12467(new_n12843, new_n12841, new_n12844);
not_4  g12468(new_n11653, new_n12845);
nand_1 g12469(new_n11673, new_n12845, new_n12846);
nand_1 g12470(new_n11675, new_n11674, new_n12847);
nand_1 g12471(new_n12847, new_n12846, new_n12848);
nand_1 g12472(new_n12848, new_n12844, new_n12849);
not_4  g12473(new_n12849, new_n12850);
nor_1  g12474(new_n12848, new_n12844, new_n12851);
nor_1  g12475(new_n12851, new_n12850, new_n12852);
nand_1 g12476(new_n12852, new_n12823, new_n12853);
nor_1  g12477(new_n12852, new_n12823, new_n12854);
not_4  g12478(new_n12854, new_n12855);
nand_1 g12479(new_n12855, new_n12853, new_n12856);
nand_1 g12480(new_n12856, new_n12821, new_n12857);
nor_1  g12481(new_n12856, new_n12821, new_n12858);
not_4  g12482(new_n12858, new_n12859);
nand_1 g12483(new_n12859, new_n12857, new_n12860);
not_4  g12484(new_n11702, new_n12861);
nand_1 g12485(new_n12861, new_n11701, new_n12862);
nand_1 g12486(new_n11703, new_n11678, new_n12863);
nand_1 g12487(new_n12863, new_n12862, new_n12864);
xnor_1 g12488(new_n12864, new_n12860, new_n12865);
xnor_1 g12489(new_n12865, new_n12819, new_n12866);
nand_1 g12490(new_n12783, new_n12780, new_n12867);
nand_1 g12491(new_n12867, new_n12785, new_n12868);
nor_1  g12492(new_n12868, new_n12866, new_n12869);
not_4  g12493(new_n12869, new_n12870);
nand_1 g12494(new_n12870, new_n12785, new_n12871);
nand_1 g12495(new_n12871, new_n12779, new_n12872);
nor_1  g12496(new_n12871, new_n12779, new_n12873);
not_4  g12497(new_n12873, new_n12874);
nand_1 g12498(new_n12874, new_n12872, new_n12875);
not_4  g12499(new_n12875, new_n12876);
not_4  g12500(new_n12812, new_n12877);
nand_1 g12501(new_n12816, new_n12877, new_n12878);
not_4  g12502(new_n12798, new_n12879);
nand_1 g12503(new_n12806, new_n12879, new_n12880);
not_4  g12504(new_n12807_1, new_n12881);
nor_1  g12505(new_n12809, new_n12881, new_n12882);
not_4  g12506(new_n12882, new_n12883);
nand_1 g12507(new_n12883, new_n12880, new_n12884);
nand_1 g12508(n11153, n6441, new_n12885);
not_4  g12509(new_n12885, new_n12886);
nand_1 g12510(n12947, n5314, new_n12887);
nand_1 g12511(n11999, n11222, new_n12888);
not_4  g12512(new_n12888, new_n12889);
xnor_1 g12513(new_n12889, new_n12887, new_n12890);
xnor_1 g12514(new_n12890, new_n12886, new_n12891);
xnor_1 g12515(new_n12891, new_n12884, new_n12892);
nand_1 g12516(n11791, n996, new_n12893);
nand_1 g12517(new_n12893, new_n12804, new_n12894);
not_4  g12518(new_n12804, new_n12895);
not_4  g12519(new_n12893, new_n12896);
nand_1 g12520(new_n12896, new_n12895, new_n12897);
nand_1 g12521(new_n12897, new_n12894, new_n12898);
not_4  g12522(new_n12898, new_n12899);
nand_1 g12523(n5760, n5319, new_n12900);
nand_1 g12524(n5767, n1478, new_n12901);
nand_1 g12525(n10990, n9457, new_n12902);
not_4  g12526(new_n12902, new_n12903);
xnor_1 g12527(new_n12903, new_n12901, new_n12904);
xnor_1 g12528(new_n12904, new_n12900, new_n12905);
not_4  g12529(new_n12905, new_n12906);
xnor_1 g12530(new_n12906, new_n12899, new_n12907);
xnor_1 g12531(new_n12907, new_n12892, new_n12908);
nand_1 g12532(new_n12796, new_n12792, new_n12909);
nor_1  g12533(new_n12794, new_n12793, new_n12910);
nor_1  g12534(new_n12811, new_n12797, new_n12911);
xnor_1 g12535(new_n12911, new_n12910, new_n12912);
nand_1 g12536(new_n12912, new_n12909, new_n12913);
xnor_1 g12537(new_n12913, new_n12908, new_n12914);
xnor_1 g12538(new_n12914, new_n12878, new_n12915);
not_4  g12539(new_n12788, new_n12916);
nand_1 g12540(new_n12817, new_n12916, new_n12917);
not_4  g12541(new_n12787, new_n12918);
nand_1 g12542(new_n12818, new_n12918, new_n12919);
nand_1 g12543(new_n12919, new_n12917, new_n12920);
xnor_1 g12544(new_n12920, new_n12915, new_n12921);
nand_1 g12545(new_n12829, new_n12825, new_n12922);
nand_1 g12546(new_n12834, new_n12922, new_n12923);
nand_1 g12547(n12391, n447, new_n12924);
nand_1 g12548(n11967, n7891, new_n12925_1);
nand_1 g12549(n12069, n1353, new_n12926);
nand_1 g12550(new_n12926, new_n12925_1, new_n12927);
not_4  g12551(new_n12925_1, new_n12928);
not_4  g12552(new_n12926, new_n12929);
nand_1 g12553(new_n12929, new_n12928, new_n12930);
nand_1 g12554(new_n12930, new_n12927, new_n12931);
xnor_1 g12555(new_n12931, new_n12924, new_n12932);
xnor_1 g12556(new_n12932, new_n12923, new_n12933);
not_4  g12557(new_n12826_1, new_n12934);
nand_1 g12558(new_n12828, new_n12934, new_n12935);
not_4  g12559(new_n12935, new_n12936);
nand_1 g12560(n7160, n6254, new_n12937);
not_4  g12561(new_n12937, new_n12938);
nand_1 g12562(new_n12938, new_n12936, new_n12939);
nand_1 g12563(new_n12937, new_n12935, new_n12940);
nand_1 g12564(new_n12940, new_n12939, new_n12941);
nand_1 g12565(n7159, n2515, new_n12942);
nand_1 g12566(n12777, n4828, new_n12943);
nand_1 g12567(n12489, n1199, new_n12944);
nand_1 g12568(new_n12944, new_n12943, new_n12945);
not_4  g12569(new_n12943, new_n12946);
not_4  g12570(new_n12944, new_n12947_1);
nand_1 g12571(new_n12947_1, new_n12946, new_n12948);
nand_1 g12572(new_n12948, new_n12945, new_n12949);
xnor_1 g12573(new_n12949, new_n12942, new_n12950);
not_4  g12574(new_n12950, new_n12951);
xnor_1 g12575(new_n12951, new_n12941, new_n12952);
xnor_1 g12576(new_n12952, new_n12933, new_n12953);
not_4  g12577(new_n12836, new_n12954);
nand_1 g12578(new_n12840, new_n12954, new_n12955);
nor_1  g12579(new_n12838, new_n12837, new_n12956);
not_4  g12580(new_n12843, new_n12957);
nand_1 g12581(new_n12957, new_n12841, new_n12958);
not_4  g12582(new_n12958, new_n12959);
xnor_1 g12583(new_n12959, new_n12956, new_n12960);
nand_1 g12584(new_n12960, new_n12955, new_n12961);
xnor_1 g12585(new_n12961, new_n12953, new_n12962);
xnor_1 g12586(new_n12962, new_n12849, new_n12963);
nand_1 g12587(new_n12859, new_n12855, new_n12964);
xnor_1 g12588(new_n12964, new_n12963, new_n12965);
xnor_1 g12589(new_n12965, new_n12921, new_n12966);
nand_1 g12590(new_n12864, new_n12860, new_n12967);
not_4  g12591(new_n12865, new_n12968);
nand_1 g12592(new_n12968, new_n12819, new_n12969);
nand_1 g12593(new_n12969, new_n12967, new_n12970);
xnor_1 g12594(new_n12970, new_n12966, new_n12971);
not_4  g12595(new_n12971, new_n12972);
nand_1 g12596(new_n12972, new_n12876, new_n12973);
nand_1 g12597(new_n12971, new_n12875, new_n12974);
nand_1 g12598(new_n12974, new_n12973, new_n12975);
nand_1 g12599(new_n12975, new_n12703, new_n12976);
not_4  g12600(new_n12976, new_n12977);
nor_1  g12601(new_n12975, new_n12703, new_n12978);
nor_1  g12602(new_n12978, new_n12977, new_n12979);
xnor_1 g12603(new_n12700, new_n12699, new_n12980);
nor_1  g12604(new_n11708, new_n11620, new_n12981);
not_4  g12605(new_n11713, new_n12982);
nor_1  g12606(new_n12982, new_n11709, new_n12983);
nor_1  g12607(new_n12983, new_n12981, new_n12984);
nand_1 g12608(new_n12984, new_n12980, new_n12985);
xnor_1 g12609(new_n12984, new_n12980, new_n12986);
not_4  g12610(new_n12986, new_n12987);
nand_1 g12611(new_n12868, new_n12866, new_n12988);
nand_1 g12612(new_n12988, new_n12870, new_n12989);
not_4  g12613(new_n12989, new_n12990);
nand_1 g12614(new_n12990, new_n12987, new_n12991);
nand_1 g12615(new_n12991, new_n12985, new_n12992);
xnor_1 g12616(new_n12992, new_n12979, n5132);
xnor_1 g12617(new_n12397, new_n11766, n5191);
not_4  g12618(new_n4080, new_n12995);
nand_1 g12619(new_n12995, new_n3934, new_n12996);
nand_1 g12620(new_n12996, new_n3931, new_n12997);
nand_1 g12621(new_n4078, new_n4073, new_n12998);
not_4  g12622(new_n3449, new_n12999);
nand_1 g12623(new_n3485, new_n12999, new_n13000);
nand_1 g12624(new_n3508, new_n3486, new_n13001);
nand_1 g12625(new_n13001, new_n13000, new_n13002);
nand_1 g12626(new_n3482, new_n3480, new_n13003);
not_4  g12627(new_n3478, new_n13004);
nand_1 g12628(new_n3484, new_n13004, new_n13005);
nand_1 g12629(new_n13005, new_n13003, new_n13006);
nand_1 g12630(n11478, n10965, new_n13007);
not_4  g12631(new_n3959, new_n13008);
nand_1 g12632(new_n3965, new_n13008, new_n13009);
nand_1 g12633(new_n13009, new_n3957, new_n13010);
nand_1 g12634(n8433, n4722, new_n13011);
nand_1 g12635(n8065, n2464, new_n13012);
nand_1 g12636(n7646, n405, new_n13013);
xnor_1 g12637(new_n13013, new_n13012, new_n13014);
xnor_1 g12638(new_n13014, new_n13011, new_n13015);
xnor_1 g12639(new_n13015, new_n13010, new_n13016);
xnor_1 g12640(new_n13016, new_n13007, new_n13017);
xnor_1 g12641(new_n13017, new_n13006, new_n13018);
nor_1  g12642(new_n4036, new_n4032, new_n13019);
nor_1  g12643(new_n4050, new_n4037, new_n13020);
nor_1  g12644(new_n13020, new_n13019, new_n13021);
not_4  g12645(new_n4001, new_n13022);
nand_1 g12646(new_n4011, new_n13022, new_n13023);
nand_1 g12647(new_n13023, new_n4000, new_n13024);
not_4  g12648(new_n4039, new_n13025);
nand_1 g12649(new_n13025, new_n4038, new_n13026);
not_4  g12650(new_n4049, new_n13027);
nand_1 g12651(new_n13027, new_n4040, new_n13028);
nand_1 g12652(new_n13028, new_n13026, new_n13029);
xnor_1 g12653(new_n13029, new_n13024, new_n13030);
nand_1 g12654(n8384, n6359, new_n13031);
nand_1 g12655(n7546, n4805, new_n13032);
xnor_1 g12656(new_n13032, new_n13031, new_n13033);
nand_1 g12657(n12925, n4938, new_n13034);
nand_1 g12658(n11536, n7862, new_n13035);
xnor_1 g12659(new_n13035, new_n13034, new_n13036);
not_4  g12660(new_n4041, new_n13037);
nand_1 g12661(new_n4044, new_n13037, new_n13038);
nand_1 g12662(new_n13038, new_n4047, new_n13039);
xnor_1 g12663(new_n13039, new_n13036, new_n13040);
xnor_1 g12664(new_n13040, new_n13033, new_n13041);
xnor_1 g12665(new_n13041, new_n13030, new_n13042);
xnor_1 g12666(new_n13042, new_n13021, new_n13043);
not_4  g12667(new_n3992_1, new_n13044);
nand_1 g12668(new_n13044, new_n3990, new_n13045);
not_4  g12669(new_n4012, new_n13046);
nand_1 g12670(new_n13046, new_n3993, new_n13047);
nand_1 g12671(new_n13047, new_n13045, new_n13048);
nand_1 g12672(new_n4029, new_n4028, new_n13049);
nand_1 g12673(new_n4031, new_n4027, new_n13050);
nand_1 g12674(new_n13050, new_n13049, new_n13051);
nand_1 g12675(n9956, n6826, new_n13052);
nand_1 g12676(n6797, n4826, new_n13053);
xnor_1 g12677(new_n13053, new_n13052, new_n13054);
nand_1 g12678(n7610, n6294, new_n13055);
nand_1 g12679(n6611, n6358, new_n13056);
xnor_1 g12680(new_n13056, new_n13055, new_n13057);
xnor_1 g12681(new_n13057, new_n13054, new_n13058);
xnor_1 g12682(new_n13058, new_n13051, new_n13059);
nand_1 g12683(n7733, n3146, new_n13060);
nand_1 g12684(new_n3986_1, new_n3985, new_n13061);
nand_1 g12685(new_n3988, new_n3984, new_n13062);
nand_1 g12686(new_n13062, new_n13061, new_n13063);
xnor_1 g12687(new_n13063, new_n13060, new_n13064);
xnor_1 g12688(new_n13064, new_n13059, new_n13065);
nand_1 g12689(n5198, n217, new_n13066);
nand_1 g12690(n5283, n503, new_n13067);
xnor_1 g12691(new_n13067, new_n13066, new_n13068);
nand_1 g12692(n4970, n137, new_n13069);
nand_1 g12693(n11296, n3992, new_n13070);
not_4  g12694(new_n13070, new_n13071);
xnor_1 g12695(new_n13071, new_n13069, new_n13072);
xnor_1 g12696(new_n13072, new_n13068, new_n13073);
not_4  g12697(new_n4002, new_n13074);
nand_1 g12698(new_n4005_1, new_n13074, new_n13075);
nand_1 g12699(new_n13075, new_n4008, new_n13076);
nand_1 g12700(n11311, n10439, new_n13077);
nand_1 g12701(n6126, n4203, new_n13078);
xnor_1 g12702(new_n13078, new_n13077, new_n13079);
xnor_1 g12703(new_n13079, new_n13076, new_n13080);
xnor_1 g12704(new_n13080, new_n13073, new_n13081);
xnor_1 g12705(new_n13081, new_n13065, new_n13082);
xnor_1 g12706(new_n13082, new_n13048, new_n13083);
xnor_1 g12707(new_n13083, new_n13043, new_n13084);
nand_1 g12708(new_n3972, new_n3970, new_n13085);
not_4  g12709(new_n3967, new_n13086);
nand_1 g12710(new_n3974, new_n13086, new_n13087);
nand_1 g12711(new_n13087, new_n13085, new_n13088);
nor_1  g12712(new_n3862, new_n3851, new_n13089);
nor_1  g12713(new_n4017, new_n4013, new_n13090);
nor_1  g12714(new_n13090, new_n13089, new_n13091);
xnor_1 g12715(new_n13091, new_n13088, new_n13092);
xnor_1 g12716(new_n13092, new_n13084, new_n13093);
xnor_1 g12717(new_n13093, new_n13018, new_n13094);
xnor_1 g12718(new_n13094, new_n13002, new_n13095);
not_4  g12719(new_n3937, new_n13096);
nand_1 g12720(new_n3975, new_n13096, new_n13097);
nand_1 g12721(new_n3979, new_n3976, new_n13098);
nand_1 g12722(new_n13098, new_n13097, new_n13099);
nor_1  g12723(new_n3950, new_n3947, new_n13100);
not_4  g12724(new_n3951, new_n13101);
nor_1  g12725(new_n3966, new_n13101, new_n13102);
nor_1  g12726(new_n13102, new_n13100, new_n13103);
nand_1 g12727(n4086, n1471, new_n13104);
nand_1 g12728(n10391, n9400, new_n13105);
not_4  g12729(new_n13105, new_n13106);
not_4  g12730(new_n3940, new_n13107);
nand_1 g12731(new_n3946, new_n13107, new_n13108);
not_4  g12732(new_n13108, new_n13109);
nand_1 g12733(new_n13109, new_n13106, new_n13110);
nand_1 g12734(new_n13106, new_n3568, new_n13111);
nand_1 g12735(new_n13111, new_n13108, new_n13112);
nand_1 g12736(new_n13112, new_n13110, new_n13113);
nand_1 g12737(n11757, n2577, new_n13114);
nand_1 g12738(n9637, n3172, new_n13115);
nand_1 g12739(n5240, n3842, new_n13116);
xnor_1 g12740(new_n13116, new_n13115, new_n13117);
xnor_1 g12741(new_n13117, new_n13114, new_n13118);
not_4  g12742(new_n3453, new_n13119);
nand_1 g12743(new_n3456_1, new_n13119, new_n13120);
nand_1 g12744(new_n13120, new_n3459, new_n13121);
xnor_1 g12745(new_n13121, new_n13118, new_n13122);
xnor_1 g12746(new_n13122, new_n13113, new_n13123);
xnor_1 g12747(new_n13123, new_n13104, new_n13124);
nand_1 g12748(n7236, n1357, new_n13125);
nand_1 g12749(new_n3475, new_n3469, new_n13126);
nand_1 g12750(new_n13126, new_n3466, new_n13127);
xnor_1 g12751(new_n13127, new_n13125, new_n13128);
xnor_1 g12752(new_n13128, new_n13124, new_n13129);
xnor_1 g12753(new_n13129, new_n13103, new_n13130);
nand_1 g12754(n1835, n1333, new_n13131);
nand_1 g12755(n11917, n11821, new_n13132);
xnor_1 g12756(new_n13132, new_n13131, new_n13133);
nand_1 g12757(n12753, n3602, new_n13134);
nand_1 g12758(n8595, n4187, new_n13135);
xnor_1 g12759(new_n13135, new_n13134, new_n13136);
nand_1 g12760(n6877, n4190, new_n13137);
nand_1 g12761(n10174, n3719, new_n13138);
xnor_1 g12762(new_n13138, new_n13137, new_n13139);
xnor_1 g12763(new_n13139, new_n13136, new_n13140);
xnor_1 g12764(new_n13140, new_n13133, new_n13141);
nand_1 g12765(new_n3962, new_n3961, new_n13142);
nand_1 g12766(new_n3964, new_n3960, new_n13143);
nand_1 g12767(new_n13143, new_n13142, new_n13144);
nand_1 g12768(n9080, n4921, new_n13145);
xnor_1 g12769(new_n13145, new_n13144, new_n13146);
xnor_1 g12770(new_n13146, new_n13141, new_n13147);
not_4  g12771(new_n3452, new_n13148);
nand_1 g12772(new_n3461, new_n13148, new_n13149);
not_4  g12773(new_n3477, new_n13150);
nand_1 g12774(new_n13150, new_n3462, new_n13151);
nand_1 g12775(new_n13151, new_n13149, new_n13152);
xnor_1 g12776(new_n13152, new_n13147, new_n13153);
xnor_1 g12777(new_n13153, new_n13130, new_n13154);
nand_1 g12778(new_n4058, new_n4055, new_n13155);
nand_1 g12779(new_n4060, new_n4051, new_n13156);
nand_1 g12780(new_n13156, new_n13155, new_n13157);
xnor_1 g12781(new_n13157, new_n13154, new_n13158);
xnor_1 g12782(new_n13158, new_n13099, new_n13159);
not_4  g12783(new_n3983, new_n13160);
nand_1 g12784(new_n4018, new_n13160, new_n13161);
nand_1 g12785(new_n4025, new_n4019, new_n13162);
nand_1 g12786(new_n13162, new_n13161, new_n13163);
xnor_1 g12787(new_n13163, new_n13159, new_n13164);
xnor_1 g12788(new_n13164, new_n13095, new_n13165);
not_4  g12789(new_n4064, new_n13166);
nor_1  g12790(new_n13166, new_n4026, new_n13167);
not_4  g12791(new_n4065, new_n13168);
nor_1  g12792(new_n4069, new_n13168, new_n13169);
nor_1  g12793(new_n13169, new_n13167, new_n13170);
nand_1 g12794(new_n4061, new_n3817, new_n13171);
not_4  g12795(new_n4063, new_n13172);
nand_1 g12796(new_n13172, new_n4062, new_n13173);
nand_1 g12797(new_n13173, new_n13171, new_n13174);
nand_1 g12798(new_n3472, new_n3471, new_n13175);
nand_1 g12799(new_n3474, new_n3470, new_n13176);
nand_1 g12800(new_n13176, new_n13175, new_n13177);
xnor_1 g12801(new_n13177, new_n13174, new_n13178);
xnor_1 g12802(new_n13178, new_n13170, new_n13179);
xnor_1 g12803(new_n13179, new_n13165, new_n13180);
xnor_1 g12804(new_n13180, new_n12998, new_n13181);
xnor_1 g12805(new_n13181, new_n12997, n5257);
xnor_1 g12806(new_n12406, new_n12396, n5411);
nand_1 g12807(new_n3917, new_n3905, new_n13184);
nand_1 g12808(new_n13184, new_n3919, n5435);
xnor_1 g12809(new_n6811, new_n6800, n5641);
xnor_1 g12810(new_n9493, new_n9483, n5670);
nand_1 g12811(new_n5486, new_n5453, new_n13188);
nand_1 g12812(new_n13188, new_n5488, n5693);
xnor_1 g12813(new_n1467, new_n1453, n5934);
xnor_1 g12814(new_n12410, new_n12409, n6089);
not_4  g12815(new_n8665_1, new_n13192);
nand_1 g12816(new_n8669, new_n13192, new_n13193);
not_4  g12817(new_n8644, new_n13194);
nand_1 g12818(new_n8648, new_n13194, new_n13195);
nand_1 g12819(new_n8653, new_n8649, new_n13196);
nand_1 g12820(new_n13196, new_n13195, new_n13197);
nand_1 g12821(n2564, n2253, new_n13198);
nand_1 g12822(n9195, n4189, new_n13199);
nand_1 g12823(n6687, n3865, new_n13200);
nand_1 g12824(new_n13200, new_n13199, new_n13201);
not_4  g12825(new_n13199, new_n13202);
not_4  g12826(new_n13200, new_n13203);
nand_1 g12827(new_n13203, new_n13202, new_n13204);
nand_1 g12828(new_n13204, new_n13201, new_n13205);
xnor_1 g12829(new_n13205, new_n13198, new_n13206);
xnor_1 g12830(new_n13206, new_n13197, new_n13207);
not_4  g12831(new_n8645, new_n13208);
nand_1 g12832(new_n8647, new_n13208, new_n13209);
nand_1 g12833(n6770, n4634, new_n13210);
xnor_1 g12834(new_n13210, new_n13209, new_n13211);
nand_1 g12835(n3627, n2879, new_n13212);
not_4  g12836(new_n13212, new_n13213);
nand_1 g12837(n10223, n9920, new_n13214);
nand_1 g12838(n7265, n4516, new_n13215);
not_4  g12839(new_n13215, new_n13216);
xnor_1 g12840(new_n13216, new_n13214, new_n13217);
xnor_1 g12841(new_n13217, new_n13213, new_n13218);
xnor_1 g12842(new_n13218, new_n13211, new_n13219);
xnor_1 g12843(new_n13219, new_n13207, new_n13220);
not_4  g12844(new_n8654, new_n13221);
nand_1 g12845(new_n8658, new_n13221, new_n13222);
nor_1  g12846(new_n8656, new_n8655, new_n13223);
nand_1 g12847(new_n8664, new_n8659, new_n13224);
not_4  g12848(new_n13224, new_n13225);
xnor_1 g12849(new_n13225, new_n13223, new_n13226);
nand_1 g12850(new_n13226, new_n13222, new_n13227);
xnor_1 g12851(new_n13227, new_n13220, new_n13228);
not_4  g12852(new_n13228, new_n13229);
xnor_1 g12853(new_n13229, new_n13193, new_n13230);
nand_1 g12854(new_n8677, new_n8673, new_n13231);
xnor_1 g12855(new_n13231, new_n13230, new_n13232);
not_4  g12856(new_n13232, new_n13233);
nand_1 g12857(new_n8717_1, new_n8714, new_n13234);
nand_1 g12858(new_n8821, new_n13234, new_n13235);
not_4  g12859(new_n13235, new_n13236);
not_4  g12860(new_n8683, new_n13237);
nand_1 g12861(new_n8712, new_n13237, new_n13238);
not_4  g12862(new_n8682, new_n13239);
nand_1 g12863(new_n8713, new_n13239, new_n13240);
nand_1 g12864(new_n13240, new_n13238, new_n13241);
not_4  g12865(new_n8707, new_n13242);
nand_1 g12866(new_n8711, new_n13242, new_n13243);
not_4  g12867(new_n8684, new_n13244);
nand_1 g12868(new_n8688, new_n13244, new_n13245);
nand_1 g12869(new_n8694, new_n13245, new_n13246);
not_4  g12870(new_n13246, new_n13247);
nand_1 g12871(n12221, n10928, new_n13248);
nand_1 g12872(n12145, n6986, new_n13249);
nand_1 g12873(n10217, n8336, new_n13250);
nand_1 g12874(new_n13250, new_n13249, new_n13251);
not_4  g12875(new_n13249, new_n13252);
not_4  g12876(new_n13250, new_n13253);
nand_1 g12877(new_n13253, new_n13252, new_n13254);
nand_1 g12878(new_n13254, new_n13251, new_n13255);
xnor_1 g12879(new_n13255, new_n13248, new_n13256);
xnor_1 g12880(new_n13256, new_n13247, new_n13257);
nor_1  g12881(new_n8686, new_n8685, new_n13258);
nand_1 g12882(n2522, n2226, new_n13259);
not_4  g12883(new_n13259, new_n13260);
xnor_1 g12884(new_n13260, new_n13258, new_n13261);
nand_1 g12885(n10678, n2024, new_n13262);
nand_1 g12886(n9189, n1094, new_n13263);
nand_1 g12887(n7946, n7320, new_n13264);
not_4  g12888(new_n13264, new_n13265);
xnor_1 g12889(new_n13265, new_n13263, new_n13266);
xnor_1 g12890(new_n13266, new_n13262, new_n13267);
not_4  g12891(new_n13267, new_n13268);
xnor_1 g12892(new_n13268, new_n13261, new_n13269);
xnor_1 g12893(new_n13269, new_n13257, new_n13270);
not_4  g12894(new_n8700, new_n13271);
nand_1 g12895(new_n13271, new_n8697, new_n13272);
nor_1  g12896(new_n8699, new_n8698, new_n13273);
nand_1 g12897(new_n8706, new_n8701, new_n13274);
not_4  g12898(new_n13274, new_n13275);
xnor_1 g12899(new_n13275, new_n13273, new_n13276);
nand_1 g12900(new_n13276, new_n13272, new_n13277);
xnor_1 g12901(new_n13277, new_n13270, new_n13278);
xnor_1 g12902(new_n13278, new_n13243, new_n13279);
xnor_1 g12903(new_n13279, new_n13241, new_n13280);
nand_1 g12904(n7160, n521, new_n13281);
not_4  g12905(new_n13281, new_n13282);
xnor_1 g12906(new_n13282, new_n8736, new_n13283);
nand_1 g12907(n2515, n2498, new_n13284);
not_4  g12908(new_n13284, new_n13285);
nand_1 g12909(n2558, n1199, new_n13286);
nand_1 g12910(n5579, n4828, new_n13287);
nand_1 g12911(new_n13287, new_n13286, new_n13288);
not_4  g12912(new_n13286, new_n13289);
not_4  g12913(new_n13287, new_n13290);
nand_1 g12914(new_n13290, new_n13289, new_n13291);
nand_1 g12915(new_n13291, new_n13288, new_n13292);
xnor_1 g12916(new_n13292, new_n13285, new_n13293);
xnor_1 g12917(new_n13293, new_n13283, new_n13294);
nand_1 g12918(new_n8747, new_n8729, new_n13295);
nand_1 g12919(n12391, n5798, new_n13296);
not_4  g12920(new_n13296, new_n13297);
nand_1 g12921(n7891, n6016, new_n13298);
nand_1 g12922(n12069, n2347, new_n13299);
not_4  g12923(new_n13299, new_n13300);
xnor_1 g12924(new_n13300, new_n13298, new_n13301);
xnor_1 g12925(new_n13301, new_n13297, new_n13302);
xnor_1 g12926(new_n13302, new_n13295, new_n13303);
xnor_1 g12927(new_n13303, new_n13294, new_n13304);
not_4  g12928(new_n8756, new_n13305);
nand_1 g12929(new_n13305, new_n8749, new_n13306);
not_4  g12930(new_n8755, new_n13307);
xnor_1 g12931(new_n8764, new_n13307, new_n13308);
not_4  g12932(new_n13308, new_n13309);
nand_1 g12933(new_n13309, new_n13306, new_n13310);
xnor_1 g12934(new_n13310, new_n13304, new_n13311);
not_4  g12935(new_n13311, new_n13312);
nand_1 g12936(new_n13312, new_n8771, new_n13313);
nand_1 g12937(new_n13311, new_n8772, new_n13314);
nand_1 g12938(new_n13314, new_n13313, new_n13315);
not_4  g12939(new_n13315, new_n13316);
nand_1 g12940(new_n8780, new_n8776, new_n13317);
nand_1 g12941(new_n13317, new_n13316, new_n13318);
nor_1  g12942(new_n13317, new_n13316, new_n13319);
not_4  g12943(new_n13319, new_n13320);
nand_1 g12944(new_n13320, new_n13318, new_n13321);
not_4  g12945(new_n8803, new_n13322);
nand_1 g12946(new_n8807, new_n13322, new_n13323);
not_4  g12947(new_n8785, new_n13324);
nand_1 g12948(new_n8789, new_n13324, new_n13325);
not_4  g12949(new_n8790, new_n13326);
nor_1  g12950(new_n8792, new_n13326, new_n13327);
not_4  g12951(new_n13327, new_n13328);
nand_1 g12952(new_n13328, new_n13325, new_n13329);
nand_1 g12953(n11153, n5153, new_n13330);
not_4  g12954(new_n13330, new_n13331);
nand_1 g12955(n7270, n5314, new_n13332);
nand_1 g12956(n11222, n2507, new_n13333);
not_4  g12957(new_n13333, new_n13334);
xnor_1 g12958(new_n13334, new_n13332, new_n13335);
xnor_1 g12959(new_n13335, new_n13331, new_n13336);
xnor_1 g12960(new_n13336, new_n13329, new_n13337);
not_4  g12961(new_n8786, new_n13338);
nand_1 g12962(new_n8788, new_n13338, new_n13339);
nand_1 g12963(n996, n806, new_n13340);
xnor_1 g12964(new_n13340, new_n13339, new_n13341);
nand_1 g12965(n9111, n5319, new_n13342);
not_4  g12966(new_n13342, new_n13343);
nand_1 g12967(n5767, n3342, new_n13344);
nand_1 g12968(n9763, n9457, new_n13345);
not_4  g12969(new_n13345, new_n13346);
xnor_1 g12970(new_n13346, new_n13344, new_n13347);
xnor_1 g12971(new_n13347, new_n13343, new_n13348);
xnor_1 g12972(new_n13348, new_n13341, new_n13349);
xnor_1 g12973(new_n13349, new_n13337, new_n13350);
nand_1 g12974(new_n8798, new_n8793, new_n13351);
nor_1  g12975(new_n8796, new_n8795, new_n13352);
nand_1 g12976(new_n8802, new_n8799, new_n13353);
not_4  g12977(new_n13353, new_n13354);
xnor_1 g12978(new_n13354, new_n13352, new_n13355);
nand_1 g12979(new_n13355, new_n13351, new_n13356);
xnor_1 g12980(new_n13356, new_n13350, new_n13357);
xnor_1 g12981(new_n13357, new_n13323, new_n13358);
not_4  g12982(new_n8808, new_n13359);
nand_1 g12983(new_n13359, new_n8784, new_n13360);
nand_1 g12984(new_n8809, new_n6528, new_n13361);
nand_1 g12985(new_n13361, new_n13360, new_n13362);
xnor_1 g12986(new_n13362, new_n13358, new_n13363);
nand_1 g12987(new_n13363, new_n13321, new_n13364);
not_4  g12988(new_n13364, new_n13365);
nor_1  g12989(new_n13363, new_n13321, new_n13366);
nor_1  g12990(new_n13366, new_n13365, new_n13367);
nand_1 g12991(new_n8817, new_n8812, new_n13368);
not_4  g12992(new_n13368, new_n13369);
nand_1 g12993(new_n13369, new_n13367, new_n13370);
not_4  g12994(new_n13370, new_n13371);
nor_1  g12995(new_n13369, new_n13367, new_n13372);
nor_1  g12996(new_n13372, new_n13371, new_n13373);
nand_1 g12997(new_n13373, new_n13280, new_n13374);
not_4  g12998(new_n13374, new_n13375);
nor_1  g12999(new_n13373, new_n13280, new_n13376);
nor_1  g13000(new_n13376, new_n13375, new_n13377);
nand_1 g13001(new_n13377, new_n13236, new_n13378);
not_4  g13002(new_n13378, new_n13379);
nor_1  g13003(new_n13377, new_n13236, new_n13380);
nor_1  g13004(new_n13380, new_n13379, new_n13381);
nand_1 g13005(new_n13381, new_n13233, new_n13382);
not_4  g13006(new_n8679, new_n13383);
nand_1 g13007(new_n13383, new_n8678, new_n13384);
not_4  g13008(new_n8823, new_n13385);
nand_1 g13009(new_n13385, new_n8680, new_n13386);
nand_1 g13010(new_n13386, new_n13384, new_n13387);
not_4  g13011(new_n13382, new_n13388);
nor_1  g13012(new_n13381, new_n13233, new_n13389);
nor_1  g13013(new_n13389, new_n13388, new_n13390);
not_4  g13014(new_n13390, new_n13391);
nor_1  g13015(new_n13391, new_n13387, new_n13392);
not_4  g13016(new_n13392, new_n13393);
nand_1 g13017(new_n13393, new_n13382, new_n13394);
not_4  g13018(new_n13394, new_n13395);
nand_1 g13019(new_n13378, new_n13374, new_n13396);
not_4  g13020(new_n13396, new_n13397);
nand_1 g13021(new_n13370, new_n13364, new_n13398);
not_4  g13022(new_n13398, new_n13399);
nand_1 g13023(new_n13275, new_n13273, new_n13400);
not_4  g13024(new_n13270, new_n13401);
nand_1 g13025(new_n13277, new_n13401, new_n13402);
nand_1 g13026(new_n13402, new_n13400, new_n13403);
not_4  g13027(new_n13197, new_n13404);
nand_1 g13028(new_n13206, new_n13404, new_n13405);
nand_1 g13029(new_n13219, new_n13207, new_n13406);
nand_1 g13030(new_n13406, new_n13405, new_n13407);
nand_1 g13031(n2522, n1094, new_n13408);
nand_1 g13032(new_n13333, new_n13332, new_n13409);
nand_1 g13033(new_n13335, new_n13330, new_n13410);
nand_1 g13034(new_n13410, new_n13409, new_n13411);
xnor_1 g13035(new_n13411, new_n13408, new_n13412);
xnor_1 g13036(new_n13412, new_n13407, new_n13413);
xnor_1 g13037(new_n13413, new_n13403, new_n13414);
nand_1 g13038(new_n13256, new_n13247, new_n13415);
not_4  g13039(new_n13257, new_n13416);
nand_1 g13040(new_n13269, new_n13416, new_n13417);
nand_1 g13041(new_n13417, new_n13415, new_n13418);
nand_1 g13042(n10678, n9189, new_n13419);
xnor_1 g13043(new_n13419, new_n13418, new_n13420);
nand_1 g13044(new_n13264, new_n13263, new_n13421);
nand_1 g13045(new_n13266, new_n13262, new_n13422);
nand_1 g13046(new_n13422, new_n13421, new_n13423);
nand_1 g13047(n7946, n7523, new_n13424);
nand_1 g13048(n10223, n3627, new_n13425);
nand_1 g13049(n3865, n2564, new_n13426);
xnor_1 g13050(new_n13426, new_n13425, new_n13427);
xnor_1 g13051(new_n13427, new_n13424, new_n13428);
xnor_1 g13052(new_n13428, new_n13423, new_n13429);
nand_1 g13053(n12221, n6986, new_n13430);
nand_1 g13054(n8336, n7823, new_n13431);
xnor_1 g13055(new_n13431, new_n13430, new_n13432);
xnor_1 g13056(new_n13432, new_n13429, new_n13433);
nand_1 g13057(new_n13215, new_n13214, new_n13434);
nand_1 g13058(new_n13217, new_n13212, new_n13435);
nand_1 g13059(new_n13435, new_n13434, new_n13436);
nor_1  g13060(new_n13260, new_n13258, new_n13437);
nor_1  g13061(new_n13267, new_n13261, new_n13438);
nor_1  g13062(new_n13438, new_n13437, new_n13439);
xnor_1 g13063(new_n13439, new_n13436, new_n13440);
nand_1 g13064(new_n13299, new_n13298, new_n13441);
nand_1 g13065(new_n13301, new_n13296, new_n13442);
nand_1 g13066(new_n13442, new_n13441, new_n13443);
nand_1 g13067(n6687, n2512, new_n13444);
nand_1 g13068(new_n13288, new_n13285, new_n13445);
nand_1 g13069(new_n13445, new_n13291, new_n13446);
xnor_1 g13070(new_n13446, new_n13444, new_n13447);
xnor_1 g13071(new_n13447, new_n13443, new_n13448);
xnor_1 g13072(new_n13448, new_n13440, new_n13449);
xnor_1 g13073(new_n13449, new_n13433, new_n13450);
nand_1 g13074(n11153, n2507, new_n13451);
nand_1 g13075(n7270, n996, new_n13452);
xnor_1 g13076(new_n13452, new_n13451, new_n13453);
nand_1 g13077(n7160, n6016, new_n13454);
nand_1 g13078(n5767, n806, new_n13455);
xnor_1 g13079(new_n13455, new_n13454, new_n13456);
xnor_1 g13080(new_n13456, new_n13453, new_n13457);
nand_1 g13081(n4828, n521, new_n13458);
nand_1 g13082(n5579, n2515, new_n13459);
xnor_1 g13083(new_n13459, new_n13458, new_n13460);
nand_1 g13084(n12069, n1576, new_n13461);
nand_1 g13085(n5314, n5153, new_n13462);
xnor_1 g13086(new_n13462, new_n13461, new_n13463);
xnor_1 g13087(new_n13463, new_n13460, new_n13464);
xnor_1 g13088(new_n13464, new_n13457, new_n13465);
not_4  g13089(new_n13198, new_n13466);
nand_1 g13090(new_n13201, new_n13466, new_n13467);
nand_1 g13091(new_n13467, new_n13204, new_n13468);
nand_1 g13092(n4516, n2879, new_n13469);
not_4  g13093(new_n13469, new_n13470);
nand_1 g13094(n4189, n2253, new_n13471);
nand_1 g13095(n9920, n4634, new_n13472);
xnor_1 g13096(new_n13472, new_n13471, new_n13473);
xnor_1 g13097(new_n13473, new_n13470, new_n13474);
xnor_1 g13098(new_n13474, new_n13468, new_n13475);
xnor_1 g13099(new_n13475, new_n13465, new_n13476);
nand_1 g13100(new_n13210, new_n13209, new_n13477);
not_4  g13101(new_n13211, new_n13478);
nand_1 g13102(new_n13218, new_n13478, new_n13479);
nand_1 g13103(new_n13479, new_n13477, new_n13480);
nor_1  g13104(new_n13340, new_n13339, new_n13481);
nor_1  g13105(new_n13348, new_n13341, new_n13482);
nor_1  g13106(new_n13482, new_n13481, new_n13483);
xnor_1 g13107(new_n13483, new_n13480, new_n13484);
xnor_1 g13108(new_n13484, new_n13476, new_n13485);
xnor_1 g13109(new_n13485, new_n13450, new_n13486);
xnor_1 g13110(new_n13486, new_n13420, new_n13487);
xnor_1 g13111(new_n13487, new_n13414, new_n13488);
nand_1 g13112(new_n13354, new_n13352, new_n13489);
nand_1 g13113(new_n13356, new_n13350, new_n13490);
nand_1 g13114(new_n13490, new_n13489, new_n13491);
nand_1 g13115(n12145, n2226, new_n13492);
not_4  g13116(new_n13248, new_n13493);
nand_1 g13117(new_n13251, new_n13493, new_n13494);
nand_1 g13118(new_n13494, new_n13254, new_n13495);
nand_1 g13119(n9195, n6770, new_n13496);
nand_1 g13120(n11222, n6431, new_n13497);
xnor_1 g13121(new_n13497, new_n13496, new_n13498);
nand_1 g13122(n10928, n10217, new_n13499);
nand_1 g13123(n7320, n2024, new_n13500);
xnor_1 g13124(new_n13500, new_n13499, new_n13501);
xnor_1 g13125(new_n13501, new_n13498, new_n13502);
nand_1 g13126(n5319, n3342, new_n13503);
nand_1 g13127(n9457, n9111, new_n13504);
nand_1 g13128(n9763, n4817, new_n13505);
not_4  g13129(new_n13505, new_n13506);
xnor_1 g13130(new_n13506, new_n13504, new_n13507);
xnor_1 g13131(new_n13507, new_n13503, new_n13508);
xnor_1 g13132(new_n13508, new_n13502, new_n13509);
xnor_1 g13133(new_n13509, new_n13495, new_n13510);
xnor_1 g13134(new_n13510, new_n13492, new_n13511);
xnor_1 g13135(new_n13511, new_n13491, new_n13512);
xnor_1 g13136(new_n13512, new_n13488, new_n13513);
not_4  g13137(new_n13243, new_n13514);
nand_1 g13138(new_n13278, new_n13514, new_n13515);
nand_1 g13139(new_n13279, new_n13241, new_n13516);
nand_1 g13140(new_n13516, new_n13515, new_n13517);
nand_1 g13141(new_n8763, new_n13307, new_n13518);
nand_1 g13142(new_n13310, new_n13304, new_n13519);
nand_1 g13143(new_n13519, new_n13518, new_n13520);
nand_1 g13144(new_n13225, new_n13223, new_n13521);
nand_1 g13145(new_n13227, new_n13220, new_n13522);
nand_1 g13146(new_n13522, new_n13521, new_n13523);
not_4  g13147(new_n13329, new_n13524);
nand_1 g13148(new_n13336, new_n13524, new_n13525);
nand_1 g13149(new_n13349, new_n13337, new_n13526);
nand_1 g13150(new_n13526, new_n13525, new_n13527);
not_4  g13151(new_n8736, new_n13528);
nand_1 g13152(new_n13282, new_n13528, new_n13529);
nand_1 g13153(new_n13293, new_n13283, new_n13530);
nand_1 g13154(new_n13530, new_n13529, new_n13531);
nand_1 g13155(n7891, n5798, new_n13532);
xnor_1 g13156(new_n13532, new_n13531, new_n13533);
nand_1 g13157(n12391, n2347, new_n13534);
nand_1 g13158(n7265, n2087, new_n13535);
xnor_1 g13159(new_n13535, new_n13534, new_n13536);
xnor_1 g13160(new_n13536, new_n13533, new_n13537);
xnor_1 g13161(new_n13537, new_n13527, new_n13538);
nand_1 g13162(n2498, n1199, new_n13539);
nand_1 g13163(n6578, n2558, new_n13540);
xnor_1 g13164(new_n13540, new_n13539, new_n13541);
xnor_1 g13165(new_n13541, new_n13538, new_n13542);
xnor_1 g13166(new_n13542, new_n13523, new_n13543);
xnor_1 g13167(new_n13543, new_n13520, new_n13544);
xnor_1 g13168(new_n13544, new_n13517, new_n13545);
xnor_1 g13169(new_n13545, new_n13513, new_n13546);
nor_1  g13170(new_n13357, new_n13323, new_n13547);
nor_1  g13171(new_n13362, new_n13358, new_n13548);
nor_1  g13172(new_n13548, new_n13547, new_n13549);
nand_1 g13173(new_n13345, new_n13344, new_n13550);
nand_1 g13174(new_n13347, new_n13342, new_n13551);
nand_1 g13175(new_n13551, new_n13550, new_n13552);
not_4  g13176(new_n13295, new_n13553);
nand_1 g13177(new_n13302, new_n13553, new_n13554);
nand_1 g13178(new_n13303, new_n13294, new_n13555);
nand_1 g13179(new_n13555, new_n13554, new_n13556);
xnor_1 g13180(new_n13556, new_n13552, new_n13557);
xnor_1 g13181(new_n13557, new_n13549, new_n13558);
xnor_1 g13182(new_n13558, new_n13546, new_n13559);
xnor_1 g13183(new_n13559, new_n13399, new_n13560);
not_4  g13184(new_n13193, new_n13561);
nand_1 g13185(new_n13229, new_n13561, new_n13562);
not_4  g13186(new_n13231, new_n13563);
nand_1 g13187(new_n13563, new_n13230, new_n13564);
nand_1 g13188(new_n13564, new_n13562, new_n13565);
nand_1 g13189(new_n13318, new_n13313, new_n13566);
xnor_1 g13190(new_n13566, new_n13565, new_n13567);
nand_1 g13191(new_n13567, new_n13560, new_n13568);
xnor_1 g13192(new_n13559, new_n13398, new_n13569);
not_4  g13193(new_n13567, new_n13570);
nand_1 g13194(new_n13570, new_n13569, new_n13571);
nand_1 g13195(new_n13571, new_n13568, new_n13572);
nand_1 g13196(new_n13572, new_n13397, new_n13573);
nor_1  g13197(new_n13570, new_n13569, new_n13574);
nor_1  g13198(new_n13567, new_n13560, new_n13575);
nor_1  g13199(new_n13575, new_n13574, new_n13576);
nand_1 g13200(new_n13576, new_n13396, new_n13577);
nand_1 g13201(new_n13577, new_n13573, new_n13578);
nand_1 g13202(new_n13578, new_n13395, new_n13579);
nor_1  g13203(new_n13576, new_n13396, new_n13580);
nor_1  g13204(new_n13572, new_n13397, new_n13581);
nor_1  g13205(new_n13581, new_n13580, new_n13582);
nand_1 g13206(new_n13582, new_n13394, new_n13583);
nand_1 g13207(new_n13583, new_n13579, n6192);
xnor_1 g13208(new_n941, new_n911_1, n6273);
nand_1 g13209(new_n8419, new_n8417, new_n13586);
nand_1 g13210(new_n13586, new_n8421, n6445);
xnor_1 g13211(new_n10431, new_n10428, n6645);
nand_1 g13212(new_n8870, new_n8869, new_n13589);
nand_1 g13213(new_n13589, new_n8872, n6689);
xnor_1 g13214(new_n1455, new_n1357_1, n6742);
xnor_1 g13215(new_n2295, new_n2474, n6809);
xnor_1 g13216(new_n7536, new_n7532, n6822);
nand_1 g13217(new_n12403, new_n12402, new_n13594);
nand_1 g13218(new_n13594, new_n12405, n6860);
nand_1 g13219(new_n10422, new_n10412, new_n13596);
nand_1 g13220(new_n13596, new_n10424, n7193);
xnor_1 g13221(new_n8631, new_n8422, n7568);
nand_1 g13222(new_n1463, new_n1462, new_n13599);
nand_1 g13223(new_n13599, new_n1465, n7676);
not_4  g13224(new_n954, new_n13601);
nand_1 g13225(new_n1095, new_n13601, new_n13602);
nand_1 g13226(new_n13602, new_n953, new_n13603);
nor_1  g13227(new_n1089, new_n1000, new_n13604);
not_4  g13228(new_n13604, new_n13605);
not_4  g13229(new_n1094_1, new_n13606);
nand_1 g13230(new_n13606, new_n1091, new_n13607);
nand_1 g13231(new_n13607, new_n13605, new_n13608);
not_4  g13232(new_n1086, new_n13609);
nand_1 g13233(new_n1088, new_n13609, new_n13610);
nand_1 g13234(new_n13610, new_n1085, new_n13611);
nand_1 g13235(n9241, n1209, new_n13612);
nand_1 g13236(new_n1078, new_n891, new_n13613);
not_4  g13237(new_n1081, new_n13614);
nand_1 g13238(new_n13614, new_n1079, new_n13615);
nand_1 g13239(new_n13615, new_n13613, new_n13616);
nand_1 g13240(new_n1075, new_n1073, new_n13617);
nand_1 g13241(new_n1077, new_n1069, new_n13618);
nand_1 g13242(new_n13618, new_n13617, new_n13619);
not_4  g13243(new_n468, new_n13620);
nand_1 g13244(new_n477, new_n13620, new_n13621);
nand_1 g13245(new_n494, new_n478, new_n13622);
nand_1 g13246(new_n13622, new_n13621, new_n13623);
not_4  g13247(new_n486, new_n13624);
nand_1 g13248(new_n492, new_n13624, new_n13625);
nand_1 g13249(new_n13625, new_n484, new_n13626);
nand_1 g13250(n12705, n2508, new_n13627);
not_4  g13251(new_n469, new_n13628);
nand_1 g13252(new_n472, new_n13628, new_n13629);
nand_1 g13253(new_n13629, new_n475, new_n13630);
xnor_1 g13254(new_n13630, new_n13627, new_n13631);
nand_1 g13255(n3986, n1980, new_n13632);
nand_1 g13256(n10848, n5857, new_n13633);
xnor_1 g13257(new_n13633, new_n13632, new_n13634);
nand_1 g13258(n11257, n2509, new_n13635);
nand_1 g13259(n4005, n1097, new_n13636);
not_4  g13260(new_n13636, new_n13637);
xnor_1 g13261(new_n13637, new_n13635, new_n13638);
xnor_1 g13262(new_n13638, new_n13634, new_n13639);
xnor_1 g13263(new_n13639, new_n13631, new_n13640);
xnor_1 g13264(new_n13640, new_n13626, new_n13641);
nand_1 g13265(n8028, n45, new_n13642);
not_4  g13266(new_n13642, new_n13643);
nand_1 g13267(new_n959, new_n958, new_n13644);
nand_1 g13268(new_n961, new_n957, new_n13645);
nand_1 g13269(new_n13645, new_n13644, new_n13646);
xnor_1 g13270(new_n13646, new_n13643, new_n13647);
not_4  g13271(new_n973, new_n13648);
nand_1 g13272(new_n976, new_n13648, new_n13649);
nand_1 g13273(new_n13649, new_n979, new_n13650);
xnor_1 g13274(new_n13650, new_n13647, new_n13651);
nand_1 g13275(n4312, n2585, new_n13652);
nand_1 g13276(new_n489, new_n488, new_n13653);
nand_1 g13277(new_n491, new_n487, new_n13654);
nand_1 g13278(new_n13654, new_n13653, new_n13655);
nand_1 g13279(n10644, n7354, new_n13656);
not_4  g13280(new_n13656, new_n13657);
nand_1 g13281(n12706, n5964, new_n13658);
nand_1 g13282(n12720, n12025, new_n13659);
xnor_1 g13283(new_n13659, new_n13658, new_n13660);
xnor_1 g13284(new_n13660, new_n13657, new_n13661);
xnor_1 g13285(new_n13661, new_n13655, new_n13662);
xnor_1 g13286(new_n13662, new_n13652, new_n13663);
xnor_1 g13287(new_n13663, new_n13651, new_n13664);
xnor_1 g13288(new_n13664, new_n13641, new_n13665);
xnor_1 g13289(new_n13665, new_n13623, new_n13666);
nand_1 g13290(n7436, n4141, new_n13667);
not_4  g13291(new_n972, new_n13668);
nand_1 g13292(new_n982, new_n13668, new_n13669);
nand_1 g13293(new_n13669, new_n970, new_n13670);
xnor_1 g13294(new_n13670, new_n13667, new_n13671);
xnor_1 g13295(new_n13671, new_n13666, new_n13672);
xnor_1 g13296(new_n13672, new_n13619, new_n13673);
xnor_1 g13297(new_n13673, new_n13616, new_n13674);
xnor_1 g13298(new_n13674, new_n13612, new_n13675);
xnor_1 g13299(new_n13675, new_n13611, new_n13676);
nand_1 g13300(n10547, n6038, new_n13677);
nand_1 g13301(new_n1008, new_n1007, new_n13678);
nand_1 g13302(new_n1010, new_n1005, new_n13679);
nand_1 g13303(new_n13679, new_n13678, new_n13680);
xnor_1 g13304(new_n13680, new_n13677, new_n13681);
nand_1 g13305(new_n1024, new_n1023, new_n13682);
nand_1 g13306(new_n1026, new_n1022, new_n13683);
nand_1 g13307(new_n13683, new_n13682, new_n13684);
nand_1 g13308(n12044, n8476, new_n13685);
nand_1 g13309(n11892, n5814, new_n13686);
nand_1 g13310(n3616, n1512, new_n13687);
xnor_1 g13311(new_n13687, new_n13686, new_n13688);
xnor_1 g13312(new_n13688, new_n13685, new_n13689);
xnor_1 g13313(new_n13689, new_n13684, new_n13690);
xnor_1 g13314(new_n13690, new_n13681, new_n13691);
nand_1 g13315(n12299, n4928, new_n13692);
nand_1 g13316(new_n1063, new_n1062, new_n13693);
nand_1 g13317(new_n1065, new_n1061, new_n13694);
nand_1 g13318(new_n13694, new_n13693, new_n13695);
xnor_1 g13319(new_n13695, new_n13692, new_n13696);
nand_1 g13320(n5069, n2530, new_n13697);
nand_1 g13321(n10545, n2802, new_n13698);
xnor_1 g13322(new_n13698, new_n13697, new_n13699);
xnor_1 g13323(new_n13699, new_n13696, new_n13700);
xnor_1 g13324(new_n13700, new_n13691, new_n13701);
not_4  g13325(new_n1004, new_n13702);
nand_1 g13326(new_n1011, new_n13702, new_n13703);
not_4  g13327(new_n1029, new_n13704);
nand_1 g13328(new_n13704, new_n1012, new_n13705);
nand_1 g13329(new_n13705, new_n13703, new_n13706);
not_4  g13330(new_n1057, new_n13707);
nand_1 g13331(new_n1059, new_n13707, new_n13708);
nand_1 g13332(new_n1066, new_n1060, new_n13709);
nand_1 g13333(new_n13709, new_n13708, new_n13710);
nand_1 g13334(new_n1027, new_n1021, new_n13711);
nand_1 g13335(new_n13711, new_n1019, new_n13712);
nand_1 g13336(n7690, n533, new_n13713);
not_4  g13337(new_n13713, new_n13714);
xnor_1 g13338(new_n13714, new_n13712, new_n13715);
xnor_1 g13339(new_n13715, new_n13710, new_n13716);
xnor_1 g13340(new_n13716, new_n13706, new_n13717);
xnor_1 g13341(new_n13717, new_n13701, new_n13718);
nand_1 g13342(n12704, n2393, new_n13719);
nand_1 g13343(n7294, n5860, new_n13720);
xnor_1 g13344(new_n13720, new_n13719, new_n13721);
nand_1 g13345(n12648, n6806, new_n13722);
nand_1 g13346(n4499, n1564, new_n13723);
xnor_1 g13347(new_n13723, new_n13722, new_n13724);
xnor_1 g13348(new_n13724, new_n13721, new_n13725);
nand_1 g13349(new_n1051, new_n1050, new_n13726);
nand_1 g13350(new_n1053, new_n1049, new_n13727);
nand_1 g13351(new_n13727, new_n13726, new_n13728);
nand_1 g13352(n5694, n5331, new_n13729);
nand_1 g13353(n7388, n4903, new_n13730);
xnor_1 g13354(new_n13730, new_n13729, new_n13731);
xnor_1 g13355(new_n13731, new_n13728, new_n13732);
xnor_1 g13356(new_n13732, new_n13725, new_n13733);
nand_1 g13357(n8276, n5105, new_n13734);
nand_1 g13358(n5305, n615, new_n13735);
xnor_1 g13359(new_n13735, new_n13734, new_n13736);
xnor_1 g13360(new_n13736, new_n13733, new_n13737);
xnor_1 g13361(new_n13737, new_n13718, new_n13738);
nand_1 g13362(new_n990, new_n987, new_n13739);
not_4  g13363(new_n984, new_n13740);
nand_1 g13364(new_n992_1, new_n13740, new_n13741);
nand_1 g13365(new_n13741, new_n13739, new_n13742);
nor_1  g13366(new_n1036, new_n839, new_n13743);
nor_1  g13367(new_n1039, new_n1030, new_n13744);
nor_1  g13368(new_n13744, new_n13743, new_n13745);
xnor_1 g13369(new_n13745, new_n13742, new_n13746);
xnor_1 g13370(new_n13746, new_n13738, new_n13747);
nand_1 g13371(n8759, n783, new_n13748);
nand_1 g13372(n10510, n7500, new_n13749);
not_4  g13373(new_n13749, new_n13750);
xnor_1 g13374(new_n13750, new_n13748, new_n13751);
nand_1 g13375(new_n499, new_n497, new_n13752);
nand_1 g13376(new_n501, new_n495, new_n13753);
nand_1 g13377(new_n13753, new_n13752, new_n13754);
nor_1  g13378(new_n1054, new_n1048, new_n13755);
nor_1  g13379(new_n1068, new_n1055, new_n13756);
nor_1  g13380(new_n13756, new_n13755, new_n13757);
xnor_1 g13381(new_n13757, new_n13754, new_n13758);
xnor_1 g13382(new_n13758, new_n13751, new_n13759);
xnor_1 g13383(new_n13759, new_n13747, new_n13760);
not_4  g13384(new_n1001, new_n13761);
nand_1 g13385(new_n1040, new_n13761, new_n13762);
nand_1 g13386(new_n1045, new_n1041, new_n13763);
nand_1 g13387(new_n13763, new_n13762, new_n13764);
nand_1 g13388(n7965, n1906, new_n13765);
xnor_1 g13389(new_n13765, new_n13764, new_n13766);
xnor_1 g13390(new_n13766, new_n13760, new_n13767);
not_4  g13391(new_n462, new_n13768);
nand_1 g13392(new_n503_1, new_n13768, new_n13769);
nand_1 g13393(new_n524, new_n504, new_n13770);
nand_1 g13394(new_n13770, new_n13769, new_n13771);
nand_1 g13395(new_n993, new_n607, new_n13772);
nand_1 g13396(new_n999, new_n994, new_n13773);
nand_1 g13397(new_n13773, new_n13772, new_n13774);
nor_1  g13398(new_n962, new_n956, new_n13775);
not_4  g13399(new_n964, new_n13776);
nor_1  g13400(new_n983, new_n13776, new_n13777);
nor_1  g13401(new_n13777, new_n13775, new_n13778);
nand_1 g13402(n8236, n6776, new_n13779);
xnor_1 g13403(new_n13779, new_n13778, new_n13780);
xnor_1 g13404(new_n13780, new_n13774, new_n13781);
xnor_1 g13405(new_n13781, new_n13771, new_n13782);
xnor_1 g13406(new_n13782, new_n13767, new_n13783);
xnor_1 g13407(new_n13783, new_n13676, new_n13784);
xnor_1 g13408(new_n13784, new_n13608, new_n13785);
not_4  g13409(new_n13785, new_n13786);
xnor_1 g13410(new_n13786, new_n13603, n7966);
nand_1 g13411(new_n13391, new_n13387, new_n13788);
nand_1 g13412(new_n13788, new_n13393, n7981);
nand_1 g13413(new_n12992, new_n12979, new_n13790);
nand_1 g13414(new_n13790, new_n12976, new_n13791);
nand_1 g13415(new_n12973, new_n12874, new_n13792);
not_4  g13416(new_n12921, new_n13793);
nand_1 g13417(new_n12965, new_n13793, new_n13794);
nand_1 g13418(new_n12970, new_n12966, new_n13795);
nand_1 g13419(new_n13795, new_n13794, new_n13796);
nand_1 g13420(new_n12962, new_n12850, new_n13797);
not_4  g13421(new_n12964, new_n13798);
nand_1 g13422(new_n13798, new_n12963, new_n13799);
nand_1 g13423(new_n13799, new_n13797, new_n13800);
nand_1 g13424(new_n12691, new_n12689, new_n13801);
nand_1 g13425(new_n12693, new_n12687, new_n13802);
nand_1 g13426(new_n13802, new_n13801, new_n13803);
not_4  g13427(new_n12942, new_n13804);
nand_1 g13428(new_n12945, new_n13804, new_n13805);
nand_1 g13429(new_n13805, new_n12948, new_n13806);
nand_1 g13430(n8717, n6986, new_n13807);
not_4  g13431(new_n13807, new_n13808);
nand_1 g13432(n11222, n10022, new_n13809);
nand_1 g13433(n12391, n1353, new_n13810);
xnor_1 g13434(new_n13810, new_n13809, new_n13811);
xnor_1 g13435(new_n13811, new_n13808, new_n13812);
xnor_1 g13436(new_n13812, new_n13806, new_n13813);
xnor_1 g13437(new_n13813, new_n13803, new_n13814);
xnor_1 g13438(new_n13814, new_n13800, new_n13815);
xnor_1 g13439(new_n13815, new_n13796, new_n13816);
nand_1 g13440(new_n12959, new_n12956, new_n13817);
not_4  g13441(new_n12953, new_n13818);
nand_1 g13442(new_n12961, new_n13818, new_n13819);
nand_1 g13443(new_n13819, new_n13817, new_n13820);
not_4  g13444(new_n12923, new_n13821);
nand_1 g13445(new_n12932, new_n13821, new_n13822);
not_4  g13446(new_n12952, new_n13823);
nand_1 g13447(new_n13823, new_n12933, new_n13824);
nand_1 g13448(new_n13824, new_n13822, new_n13825);
nand_1 g13449(n12069, n4436, new_n13826);
nand_1 g13450(n11999, n11153, new_n13827);
xnor_1 g13451(new_n13827, new_n13826, new_n13828);
nand_1 g13452(n7159, n1199, new_n13829);
nand_1 g13453(n11967, n7160, new_n13830);
not_4  g13454(new_n13830, new_n13831);
xnor_1 g13455(new_n13831, new_n13829, new_n13832);
xnor_1 g13456(new_n13832, new_n13828, new_n13833);
not_4  g13457(new_n12924, new_n13834);
nand_1 g13458(new_n12927, new_n13834, new_n13835);
nand_1 g13459(new_n13835, new_n12930, new_n13836);
nand_1 g13460(n6254, n4828, new_n13837);
nand_1 g13461(n11407, n2087, new_n13838);
xnor_1 g13462(new_n13838, new_n13837, new_n13839);
xnor_1 g13463(new_n13839, new_n13836, new_n13840);
xnor_1 g13464(new_n13840, new_n13833, new_n13841);
xnor_1 g13465(new_n13841, new_n13825, new_n13842);
xnor_1 g13466(new_n13842, new_n13820, new_n13843);
not_4  g13467(new_n12884, new_n13844);
nand_1 g13468(new_n12891, new_n13844, new_n13845);
not_4  g13469(new_n12907, new_n13846);
nand_1 g13470(new_n13846, new_n12892, new_n13847);
nand_1 g13471(new_n13847, new_n13845, new_n13848);
nand_1 g13472(n12489, n6578, new_n13849);
nand_1 g13473(n12947, n996, new_n13850);
nand_1 g13474(n9457, n5760, new_n13851);
xnor_1 g13475(new_n13851, new_n13850, new_n13852);
xnor_1 g13476(new_n13852, new_n13849, new_n13853);
xnor_1 g13477(new_n13853, new_n13848, new_n13854);
not_4  g13478(new_n12941, new_n13855);
nand_1 g13479(new_n12951, new_n13855, new_n13856);
nand_1 g13480(new_n13856, new_n12939, new_n13857);
nand_1 g13481(n7891, n447, new_n13858);
xnor_1 g13482(new_n13858, new_n13857, new_n13859);
nand_1 g13483(n12777, n2515, new_n13860);
nand_1 g13484(new_n12902, new_n12901, new_n13861);
nand_1 g13485(new_n12904, new_n12900, new_n13862);
nand_1 g13486(new_n13862, new_n13861, new_n13863);
nand_1 g13487(new_n12888, new_n12887, new_n13864);
nand_1 g13488(new_n12890, new_n12885, new_n13865);
nand_1 g13489(new_n13865, new_n13864, new_n13866);
xnor_1 g13490(new_n13866, new_n13863, new_n13867);
xnor_1 g13491(new_n13867, new_n13860, new_n13868);
xnor_1 g13492(new_n13868, new_n13859, new_n13869);
nand_1 g13493(n6441, n5314, new_n13870);
nand_1 g13494(n11791, n5767, new_n13871);
xnor_1 g13495(new_n13871, new_n13870, new_n13872);
nand_1 g13496(new_n12905, new_n12899, new_n13873);
nand_1 g13497(new_n13873, new_n12897, new_n13874);
nand_1 g13498(n6687, n6604, new_n13875);
xnor_1 g13499(new_n13875, new_n13874, new_n13876);
xnor_1 g13500(new_n13876, new_n13872, new_n13877);
xnor_1 g13501(new_n13877, new_n13869, new_n13878);
xnor_1 g13502(new_n13878, new_n13854, new_n13879);
xnor_1 g13503(new_n13879, new_n13843, new_n13880);
nand_1 g13504(new_n12774, new_n12772, new_n13881);
not_4  g13505(new_n12769, new_n13882);
nand_1 g13506(new_n12776, new_n13882, new_n13883);
nand_1 g13507(new_n13883, new_n13881, new_n13884);
not_4  g13508(new_n12743, new_n13885);
nand_1 g13509(new_n12750, new_n13885, new_n13886);
not_4  g13510(new_n12768, new_n13887);
nand_1 g13511(new_n13887, new_n12751, new_n13888);
nand_1 g13512(new_n13888, new_n13886, new_n13889);
nand_1 g13513(n10678, n6429, new_n13890);
xnor_1 g13514(new_n13890, new_n13889, new_n13891);
nand_1 g13515(new_n12766, new_n12760, new_n13892);
nand_1 g13516(new_n13892, new_n12758, new_n13893);
nand_1 g13517(n2433, n2226, new_n13894);
nand_1 g13518(n8819, n1094, new_n13895);
nand_1 g13519(n10928, n7730, new_n13896);
xnor_1 g13520(new_n13896, new_n13895, new_n13897);
xnor_1 g13521(new_n13897, new_n13894, new_n13898);
xnor_1 g13522(new_n13898, new_n13893, new_n13899);
xnor_1 g13523(new_n13899, new_n13891, new_n13900);
xnor_1 g13524(new_n13900, new_n13884, new_n13901);
xnor_1 g13525(new_n13901, new_n13880, new_n13902);
nand_1 g13526(new_n12911, new_n12910, new_n13903);
not_4  g13527(new_n12908, new_n13904);
nand_1 g13528(new_n12913, new_n13904, new_n13905);
nand_1 g13529(new_n13905, new_n13903, new_n13906);
nor_1  g13530(new_n12694, new_n12653, new_n13907);
nor_1  g13531(new_n12702, new_n12695, new_n13908);
nor_1  g13532(new_n13908, new_n13907, new_n13909);
xnor_1 g13533(new_n13909, new_n13906, new_n13910);
xnor_1 g13534(new_n13910, new_n13902, new_n13911);
not_4  g13535(new_n12878, new_n13912);
nand_1 g13536(new_n12914, new_n13912, new_n13913);
nand_1 g13537(new_n12920, new_n12915, new_n13914);
nand_1 g13538(new_n13914, new_n13913, new_n13915);
not_4  g13539(new_n12741, new_n13916);
nand_1 g13540(new_n12777_1, new_n13916, new_n13917);
nand_1 g13541(new_n12778, new_n12739, new_n13918);
nand_1 g13542(new_n13918, new_n13917, new_n13919);
not_4  g13543(new_n12667, new_n13920);
nor_1  g13544(new_n13920, new_n12658, new_n13921);
not_4  g13545(new_n12668, new_n13922);
nor_1  g13546(new_n12685, new_n13922, new_n13923);
nor_1  g13547(new_n13923, new_n13921, new_n13924);
not_4  g13548(new_n12659, new_n13925);
nand_1 g13549(new_n12662, new_n13925, new_n13926);
nand_1 g13550(new_n13926, new_n12665, new_n13927);
nand_1 g13551(n12709, n7523, new_n13928);
nand_1 g13552(n12000, n4189, new_n13929);
xnor_1 g13553(new_n13929, new_n13928, new_n13930);
xnor_1 g13554(new_n13930, new_n13927, new_n13931);
nand_1 g13555(n9725, n2564, new_n13932);
nand_1 g13556(n9920, n4370, new_n13933);
xnor_1 g13557(new_n13933, new_n13932, new_n13934);
nand_1 g13558(n5212, n4516, new_n13935);
nand_1 g13559(n6770, n5320, new_n13936);
nand_1 g13560(n5319, n1478, new_n13937);
xnor_1 g13561(new_n13937, new_n13936, new_n13938);
xnor_1 g13562(new_n13938, new_n13935, new_n13939);
xnor_1 g13563(new_n13939, new_n13934, new_n13940);
nand_1 g13564(n11728, n7320, new_n13941);
nand_1 g13565(new_n12763, new_n12762, new_n13942);
nand_1 g13566(new_n12765, new_n12761, new_n13943);
nand_1 g13567(new_n13943, new_n13942, new_n13944);
xnor_1 g13568(new_n13944, new_n13941, new_n13945);
xnor_1 g13569(new_n13945, new_n13940, new_n13946);
xnor_1 g13570(new_n13946, new_n13931, new_n13947);
not_4  g13571(new_n12675, new_n13948);
nand_1 g13572(new_n12678, new_n13948, new_n13949);
nand_1 g13573(new_n13949, new_n12681, new_n13950);
nand_1 g13574(n10990, n4817, new_n13951);
nand_1 g13575(n11877, n3627, new_n13952);
nand_1 g13576(n8336, n1198, new_n13953);
not_4  g13577(new_n13953, new_n13954);
xnor_1 g13578(new_n13954, new_n13952, new_n13955);
xnor_1 g13579(new_n13955, new_n13951, new_n13956);
xnor_1 g13580(new_n13956, new_n13950, new_n13957);
not_4  g13581(new_n12674, new_n13958);
nand_1 g13582(new_n12684, new_n13958, new_n13959);
nand_1 g13583(new_n13959, new_n12673, new_n13960);
nand_1 g13584(new_n12747, new_n12746, new_n13961);
nand_1 g13585(new_n12749, new_n12744, new_n13962);
nand_1 g13586(new_n13962, new_n13961, new_n13963);
xnor_1 g13587(new_n13963, new_n13960, new_n13964);
xnor_1 g13588(new_n13964, new_n13957, new_n13965);
xnor_1 g13589(new_n13965, new_n13947, new_n13966);
xnor_1 g13590(new_n13966, new_n13924, new_n13967);
xnor_1 g13591(new_n13967, new_n13919, new_n13968);
xnor_1 g13592(new_n13968, new_n13915, new_n13969);
xnor_1 g13593(new_n13969, new_n13911, new_n13970);
xnor_1 g13594(new_n13970, new_n13816, new_n13971);
xnor_1 g13595(new_n13971, new_n13792, new_n13972);
xnor_1 g13596(new_n13972, new_n13791, n8100);
nand_1 g13597(new_n10418, new_n10417, new_n13974);
nand_1 g13598(new_n13974, new_n10420, n8138);
nand_1 g13599(new_n6565, new_n6564, new_n13976);
nand_1 g13600(new_n13976, new_n6567, n8202);
xnor_1 g13601(new_n3907, new_n3898, n8303);
nand_1 g13602(new_n3156, new_n3155, new_n13979);
nand_1 g13603(new_n13979, new_n3158, n8398);
nand_1 g13604(new_n4539, new_n4538, new_n13981);
nand_1 g13605(new_n13981, new_n4541, n9137);
nand_1 g13606(new_n7670, new_n7668, new_n13983);
nand_1 g13607(new_n13983, new_n7672, n9387);
nand_1 g13608(new_n12419, new_n12418, new_n13985);
nand_1 g13609(new_n13985, new_n12421, n9571);
not_4  g13610(new_n944, new_n13987);
xnor_1 g13611(new_n947, new_n13987, n9578);
xnor_1 g13612(new_n1238, new_n1236, n9706);
xnor_1 g13613(new_n4542, new_n4532, n9756);
nand_1 g13614(new_n7335, new_n7315, new_n13991);
nand_1 g13615(new_n13991, new_n7314, new_n13992);
nand_1 g13616(n12826, n7891, new_n13993);
nand_1 g13617(new_n7021, new_n7019, new_n13994);
not_4  g13618(new_n7017, new_n13995);
nand_1 g13619(new_n7023, new_n13995, new_n13996);
nand_1 g13620(new_n13996, new_n13994, new_n13997);
xnor_1 g13621(new_n13997, new_n13993, new_n13998);
nand_1 g13622(new_n7310, new_n7284, new_n13999);
nand_1 g13623(n8336, n2278, new_n14000);
not_4  g13624(new_n6896, new_n14001);
nand_1 g13625(new_n6930, new_n14001, new_n14002);
nand_1 g13626(new_n6942, new_n6931, new_n14003);
nand_1 g13627(new_n14003, new_n14002, new_n14004);
xnor_1 g13628(new_n14004, new_n14000, new_n14005);
not_4  g13629(new_n14005, new_n14006);
not_4  g13630(new_n7135, new_n14007);
nor_1  g13631(new_n14007, new_n7091, new_n14008);
not_4  g13632(new_n7136, new_n14009);
nor_1  g13633(new_n7149, new_n14009, new_n14010);
nor_1  g13634(new_n14010, new_n14008, new_n14011);
nor_1  g13635(new_n6911, new_n6910, new_n14012);
nor_1  g13636(new_n6921, new_n6912, new_n14013);
nor_1  g13637(new_n14013, new_n14012, new_n14014);
not_4  g13638(new_n6995, new_n14015);
nand_1 g13639(new_n7002, new_n14015, new_n14016);
nand_1 g13640(new_n7016, new_n7003, new_n14017);
nand_1 g13641(new_n14017, new_n14016, new_n14018);
nand_1 g13642(n11662, n6770, new_n14019);
nand_1 g13643(n10451, n2226, new_n14020);
nand_1 g13644(n5319, n3754, new_n14021);
xnor_1 g13645(new_n14021, new_n14020, new_n14022);
xnor_1 g13646(new_n14022, new_n14019, new_n14023);
nand_1 g13647(new_n7012, new_n7011, new_n14024);
nand_1 g13648(new_n7014, new_n7010, new_n14025);
nand_1 g13649(new_n14025, new_n14024, new_n14026);
xnor_1 g13650(new_n14026, new_n14023, new_n14027);
not_4  g13651(new_n6913, new_n14028);
nand_1 g13652(new_n6916, new_n14028, new_n14029);
nand_1 g13653(new_n14029, new_n6919, new_n14030);
nand_1 g13654(n10278, n6986, new_n14031);
nand_1 g13655(n10678, n3022, new_n14032);
xnor_1 g13656(new_n14032, new_n14031, new_n14033);
xnor_1 g13657(new_n14033, new_n14030, new_n14034);
xnor_1 g13658(new_n14034, new_n14027, new_n14035);
not_4  g13659(new_n7006, new_n14036);
nand_1 g13660(new_n7008, new_n14036, new_n14037);
nand_1 g13661(new_n7015, new_n7009, new_n14038);
nand_1 g13662(new_n14038, new_n14037, new_n14039);
nor_1  g13663(new_n7000, new_n6998, new_n14040);
not_4  g13664(new_n6996, new_n14041);
nor_1  g13665(new_n7001, new_n14041, new_n14042);
nor_1  g13666(new_n14042, new_n14040, new_n14043);
xnor_1 g13667(new_n14043, new_n14039, new_n14044);
xnor_1 g13668(new_n14044, new_n14035, new_n14045);
xnor_1 g13669(new_n14045, new_n14018, new_n14046);
xnor_1 g13670(new_n14046, new_n14014, new_n14047);
nand_1 g13671(new_n6903, new_n6902, new_n14048);
nand_1 g13672(new_n6905, new_n6901, new_n14049);
nand_1 g13673(new_n14049, new_n14048, new_n14050);
nand_1 g13674(n8665, n2515, new_n14051);
nand_1 g13675(n10898, n9457, new_n14052);
nand_1 g13676(n12511, n11222, new_n14053);
xnor_1 g13677(new_n14053, new_n14052, new_n14054);
xnor_1 g13678(new_n14054, new_n14051, new_n14055);
xnor_1 g13679(new_n14055, new_n14050, new_n14056);
xnor_1 g13680(new_n14056, new_n14047, new_n14057);
nand_1 g13681(n12391, n4094, new_n14058);
nor_1  g13682(new_n6906, new_n6900, new_n14059);
not_4  g13683(new_n6908, new_n14060);
nor_1  g13684(new_n6923, new_n14060, new_n14061);
nor_1  g13685(new_n14061, new_n14059, new_n14062);
nand_1 g13686(n4516, n3932, new_n14063);
nand_1 g13687(n7523, n6703, new_n14064);
xnor_1 g13688(new_n14064, new_n14063, new_n14065);
nand_1 g13689(n11423, n10928, new_n14066);
nand_1 g13690(n12591, n3627, new_n14067);
xnor_1 g13691(new_n14067, new_n14066, new_n14068);
xnor_1 g13692(new_n14068, new_n14065, new_n14069);
xnor_1 g13693(new_n14069, new_n14062, new_n14070);
nand_1 g13694(n11876, n4817, new_n14071);
not_4  g13695(new_n7116, new_n14072);
nand_1 g13696(new_n7119, new_n14072, new_n14073);
nand_1 g13697(new_n14073, new_n7122, new_n14074);
nand_1 g13698(n10327, n4189, new_n14075);
nand_1 g13699(n9920, n7456, new_n14076);
xnor_1 g13700(new_n14076, new_n14075, new_n14077);
xnor_1 g13701(new_n14077, new_n14074, new_n14078);
xnor_1 g13702(new_n14078, new_n14071, new_n14079);
xnor_1 g13703(new_n14079, new_n14070, new_n14080);
xnor_1 g13704(new_n14080, new_n14058, new_n14081);
xnor_1 g13705(new_n14081, new_n14057, new_n14082);
xnor_1 g13706(new_n14082, new_n14011, new_n14083);
xnor_1 g13707(new_n14083, new_n14006, new_n14084);
nand_1 g13708(new_n6927, new_n6926, new_n14085);
not_4  g13709(new_n6924, new_n14086);
nand_1 g13710(new_n6929, new_n14086, new_n14087);
nand_1 g13711(new_n14087, new_n14085, new_n14088);
nor_1  g13712(new_n7131, new_n7062, new_n14089);
not_4  g13713(new_n7128, new_n14090);
nor_1  g13714(new_n7134, new_n14090, new_n14091);
nor_1  g13715(new_n14091, new_n14089, new_n14092);
xnor_1 g13716(new_n14092, new_n14088, new_n14093);
nand_1 g13717(new_n7204, new_n7202, new_n14094);
nand_1 g13718(new_n7231, new_n7206, new_n14095);
nand_1 g13719(new_n14095, new_n14094, new_n14096);
nand_1 g13720(n11023, n1094, new_n14097);
xnor_1 g13721(new_n14097, new_n14096, new_n14098);
nand_1 g13722(new_n7216, new_n7210, new_n14099);
not_4  g13723(new_n7217, new_n14100);
nand_1 g13724(new_n7230, new_n14100, new_n14101);
nand_1 g13725(new_n14101, new_n14099, new_n14102);
not_4  g13726(new_n7115, new_n14103);
nand_1 g13727(new_n7125, new_n14103, new_n14104);
nand_1 g13728(new_n14104, new_n7114, new_n14105);
nand_1 g13729(new_n7213, new_n7212, new_n14106);
nand_1 g13730(new_n7215, new_n7211, new_n14107);
nand_1 g13731(new_n14107, new_n14106, new_n14108);
nand_1 g13732(new_n7225, new_n7224, new_n14109);
nand_1 g13733(new_n7227, new_n7223, new_n14110);
nand_1 g13734(new_n14110, new_n14109, new_n14111);
xnor_1 g13735(new_n14111, new_n14108, new_n14112);
nand_1 g13736(n12069, n10685, new_n14113);
nand_1 g13737(n6578, n5645, new_n14114);
xnor_1 g13738(new_n14114, new_n14113, new_n14115);
nand_1 g13739(n5767, n2749, new_n14116);
nand_1 g13740(n996, n159, new_n14117);
nand_1 g13741(n5314, n1510, new_n14118);
xnor_1 g13742(new_n14118, new_n14117, new_n14119);
xnor_1 g13743(new_n14119, new_n14116, new_n14120);
xnor_1 g13744(new_n14120, new_n14115, new_n14121);
xnor_1 g13745(new_n14121, new_n14112, new_n14122);
not_4  g13746(new_n7219, new_n14123);
nand_1 g13747(new_n7221, new_n14123, new_n14124);
nand_1 g13748(new_n7228, new_n7222, new_n14125);
nand_1 g13749(new_n14125, new_n14124, new_n14126);
nand_1 g13750(n7160, n2551, new_n14127);
nand_1 g13751(n9583, n2564, new_n14128);
nand_1 g13752(n9640, n7320, new_n14129);
xnor_1 g13753(new_n14129, new_n14128, new_n14130);
xnor_1 g13754(new_n14130, new_n14127, new_n14131);
nand_1 g13755(n1199, n1067, new_n14132);
nand_1 g13756(n12247, n11153, new_n14133);
xnor_1 g13757(new_n14133, new_n14132, new_n14134);
xnor_1 g13758(new_n14134, new_n14131, new_n14135);
xnor_1 g13759(new_n14135, new_n14126, new_n14136);
xnor_1 g13760(new_n14136, new_n14122, new_n14137);
xnor_1 g13761(new_n14137, new_n14105, new_n14138);
nand_1 g13762(new_n7105, new_n7098, new_n14139);
nand_1 g13763(new_n7127, new_n7107, new_n14140);
nand_1 g13764(new_n14140, new_n14139, new_n14141);
nand_1 g13765(new_n7102, new_n7101, new_n14142);
nand_1 g13766(new_n7104, new_n7099, new_n14143);
nand_1 g13767(new_n14143, new_n14142, new_n14144);
nand_1 g13768(n6687, n753, new_n14145);
nand_1 g13769(n2087, n1798, new_n14146);
xnor_1 g13770(new_n14146, new_n14145, new_n14147);
xnor_1 g13771(new_n14147, new_n14144, new_n14148);
xnor_1 g13772(new_n14148, new_n14141, new_n14149);
xnor_1 g13773(new_n14149, new_n14138, new_n14150);
xnor_1 g13774(new_n14150, new_n14102, new_n14151);
xnor_1 g13775(new_n14151, new_n14098, new_n14152);
xnor_1 g13776(new_n14152, new_n14093, new_n14153);
not_4  g13777(new_n7199, new_n14154);
nand_1 g13778(new_n7233, new_n14154, new_n14155);
nand_1 g13779(new_n7249, new_n7234, new_n14156);
nand_1 g13780(new_n14156, new_n14155, new_n14157);
not_4  g13781(new_n6989, new_n14158);
nand_1 g13782(new_n7024, new_n14158, new_n14159);
not_4  g13783(new_n7038, new_n14160);
nand_1 g13784(new_n14160, new_n7025, new_n14161);
nand_1 g13785(new_n14161, new_n14159, new_n14162);
xnor_1 g13786(new_n14162, new_n14157, new_n14163);
xnor_1 g13787(new_n14163, new_n14153, new_n14164);
xnor_1 g13788(new_n14164, new_n14084, new_n14165);
nand_1 g13789(n11922, n4828, new_n14166);
not_4  g13790(new_n7279, new_n14167);
nor_1  g13791(new_n7280, new_n7150, new_n14168);
nor_1  g13792(new_n14168, new_n14167, new_n14169);
xnor_1 g13793(new_n14169, new_n14166, new_n14170);
not_4  g13794(new_n14170, new_n14171);
nor_1  g13795(new_n14171, new_n14165, new_n14172);
xnor_1 g13796(new_n14083, new_n14005, new_n14173);
xnor_1 g13797(new_n14164, new_n14173, new_n14174);
nor_1  g13798(new_n14170, new_n14174, new_n14175);
nor_1  g13799(new_n14175, new_n14172, new_n14176);
nor_1  g13800(new_n14176, new_n13999, new_n14177);
not_4  g13801(new_n13999, new_n14178);
nand_1 g13802(new_n14170, new_n14174, new_n14179);
nand_1 g13803(new_n14171, new_n14165, new_n14180);
nand_1 g13804(new_n14180, new_n14179, new_n14181);
nor_1  g13805(new_n14181, new_n14178, new_n14182);
nor_1  g13806(new_n14182, new_n14177, new_n14183);
nand_1 g13807(new_n14183, new_n13998, new_n14184);
not_4  g13808(new_n13998, new_n14185);
nand_1 g13809(new_n14181, new_n14178, new_n14186);
nand_1 g13810(new_n14176, new_n13999, new_n14187);
nand_1 g13811(new_n14187, new_n14186, new_n14188);
nand_1 g13812(new_n14188, new_n14185, new_n14189);
nand_1 g13813(new_n14189, new_n14184, new_n14190);
nand_1 g13814(new_n14190, new_n13992, new_n14191);
not_4  g13815(new_n13992, new_n14192);
nor_1  g13816(new_n14188, new_n14185, new_n14193);
nor_1  g13817(new_n14183, new_n13998, new_n14194);
nor_1  g13818(new_n14194, new_n14193, new_n14195);
nand_1 g13819(new_n14195, new_n14192, new_n14196);
nand_1 g13820(new_n14196, new_n14191, n9767);
nand_1 g13821(new_n2274, new_n2273, new_n14198);
nand_1 g13822(new_n14198, new_n2276, n9820);
nand_1 g13823(new_n10669, new_n10667, new_n14200);
nand_1 g13824(new_n14200, new_n10448, n9938);
not_4  g13825(new_n939, new_n14202);
xnor_1 g13826(new_n14202, new_n938, n10476);
xnor_1 g13827(new_n936, new_n926, n10589);
xnor_1 g13828(new_n1233, new_n1232, n10695);
not_4  g13829(new_n3928, new_n14206);
nand_1 g13830(new_n3887, new_n3885, new_n14207);
xnor_1 g13831(new_n14207, new_n14206, n10789);
xnor_1 g13832(new_n3150, new_n3141, n10851);
nand_1 g13833(new_n5479, new_n5467, new_n14210);
nand_1 g13834(new_n14210, new_n5481, n10913);
xnor_1 g13835(new_n7816, new_n7677, n10949);
nand_1 g13836(new_n12423, new_n12372, new_n14213);
nand_1 g13837(new_n14213, new_n12609, n11216);
xnor_1 g13838(new_n5469, new_n5460, n11326);
nor_1  g13839(new_n6237, new_n6242, new_n14216);
nor_1  g13840(new_n14216, new_n6093, new_n14217);
not_4  g13841(new_n6141, new_n14218);
nand_1 g13842(new_n6142, new_n14218, new_n14219);
nand_1 g13843(new_n6236, new_n6143, new_n14220);
nand_1 g13844(new_n14220, new_n14219, new_n14221);
not_4  g13845(new_n14221, new_n14222);
not_4  g13846(new_n6101, new_n14223);
nand_1 g13847(new_n6139, new_n14223, new_n14224);
nand_1 g13848(new_n6140, new_n6099, new_n14225);
nand_1 g13849(new_n14225, new_n14224, new_n14226);
nand_1 g13850(new_n6136, new_n6135, new_n14227);
not_4  g13851(new_n6133, new_n14228);
nand_1 g13852(new_n6138, new_n14228, new_n14229);
nand_1 g13853(new_n14229, new_n14227, new_n14230);
nand_1 g13854(n9763, n45, new_n14231);
nand_1 g13855(n8759, n7823, new_n14232);
xnor_1 g13856(new_n14232, new_n14231, new_n14233);
xnor_1 g13857(new_n14233, new_n14230, new_n14234);
nand_1 g13858(new_n5764, new_n5763, new_n14235);
nand_1 g13859(new_n5766, new_n5762, new_n14236);
nand_1 g13860(new_n14236, new_n14235, new_n14237);
nand_1 g13861(n9241, n9189, new_n14238);
xnor_1 g13862(new_n14238, new_n14237, new_n14239);
nand_1 g13863(n12705, n4634, new_n14240);
nand_1 g13864(n12145, n7436, new_n14241);
xnor_1 g13865(new_n14241, new_n14240, new_n14242);
nand_1 g13866(n9195, n4312, new_n14243);
nand_1 g13867(n10217, n6776, new_n14244);
not_4  g13868(new_n14244, new_n14245);
xnor_1 g13869(new_n14245, new_n14243, new_n14246);
xnor_1 g13870(new_n14246, new_n14242, new_n14247);
xnor_1 g13871(new_n14247, new_n14239, new_n14248);
nand_1 g13872(new_n6129, new_n6119, new_n14249);
nand_1 g13873(new_n14249, new_n6116, new_n14250);
nand_1 g13874(new_n6106, new_n6105, new_n14251);
nand_1 g13875(new_n6108, new_n6104, new_n14252);
nand_1 g13876(new_n14252, new_n14251, new_n14253);
xnor_1 g13877(new_n14253, new_n14250, new_n14254);
xnor_1 g13878(new_n14254, new_n14248, new_n14255);
nand_1 g13879(new_n6124, new_n6121, new_n14256);
nand_1 g13880(new_n14256, new_n6127, new_n14257);
xnor_1 g13881(new_n14257, new_n14255, new_n14258);
nand_1 g13882(n3986, n3342, new_n14259);
nand_1 g13883(n8276, n2522, new_n14260);
nand_1 g13884(n12299, n12221, new_n14261);
xnor_1 g13885(new_n14261, new_n14260, new_n14262);
xnor_1 g13886(new_n14262, new_n14259, new_n14263);
xnor_1 g13887(new_n14263, new_n14258, new_n14264);
nor_1  g13888(new_n6111, new_n6103, new_n14265);
nor_1  g13889(new_n6131, new_n6112, new_n14266);
nor_1  g13890(new_n14266, new_n14265, new_n14267);
not_4  g13891(new_n6219, new_n14268);
nor_1  g13892(new_n14268, new_n6038_1, new_n14269);
nor_1  g13893(new_n6221, new_n6216, new_n14270);
nor_1  g13894(new_n14270, new_n14269, new_n14271);
xnor_1 g13895(new_n14271, new_n14267, new_n14272);
xnor_1 g13896(new_n14272, new_n14264, new_n14273);
xnor_1 g13897(new_n14273, new_n14234, new_n14274);
xnor_1 g13898(new_n14274, new_n14226, new_n14275);
nand_1 g13899(n12025, n10223, new_n14276);
not_4  g13900(new_n14276, new_n14277);
nand_1 g13901(new_n5767_1, new_n5761, new_n14278);
nand_1 g13902(new_n14278, new_n5759, new_n14279);
xnor_1 g13903(new_n14279, new_n14277, new_n14280);
xnor_1 g13904(new_n14280, new_n14275, new_n14281);
not_4  g13905(new_n6190, new_n14282);
nand_1 g13906(new_n6197, new_n14282, new_n14283);
not_4  g13907(new_n6215, new_n14284);
nand_1 g13908(new_n14284, new_n6198, new_n14285);
nand_1 g13909(new_n14285, new_n14283, new_n14286);
nand_1 g13910(n7690, n5579, new_n14287);
nand_1 g13911(n7388, n2507, new_n14288);
xnor_1 g13912(new_n14288, new_n14287, new_n14289);
nand_1 g13913(n7270, n2393, new_n14290);
nand_1 g13914(n5331, n1576, new_n14291);
xnor_1 g13915(new_n14291, new_n14290, new_n14292);
xnor_1 g13916(new_n14292, new_n14289, new_n14293);
nand_1 g13917(n3616, n2498, new_n14294);
nand_1 g13918(n12648, n6016, new_n14295);
xnor_1 g13919(new_n14295, new_n14294, new_n14296);
xnor_1 g13920(new_n14296, new_n14293, new_n14297);
nand_1 g13921(n5798, n2530, new_n14298);
nand_1 g13922(n10644, n7946, new_n14299);
not_4  g13923(new_n14299, new_n14300);
xnor_1 g13924(new_n14300, new_n14298, new_n14301);
nand_1 g13925(new_n6194, new_n6193, new_n14302);
nand_1 g13926(new_n6196, new_n6191, new_n14303);
nand_1 g13927(new_n14303, new_n14302, new_n14304);
nand_1 g13928(new_n5749, new_n5748, new_n14305);
nand_1 g13929(new_n5751, new_n5747, new_n14306);
nand_1 g13930(new_n14306, new_n14305, new_n14307);
xnor_1 g13931(new_n14307, new_n14304, new_n14308);
xnor_1 g13932(new_n14308, new_n14301, new_n14309);
xnor_1 g13933(new_n14309, new_n14297, new_n14310);
xnor_1 g13934(new_n14310, new_n14286, new_n14311);
nand_1 g13935(new_n6175, new_n6173, new_n14312);
nand_1 g13936(new_n6177, new_n6169, new_n14313);
nand_1 g13937(new_n14313, new_n14312, new_n14314);
nand_1 g13938(new_n6210, new_n6209, new_n14315);
nand_1 g13939(new_n6212, new_n6208, new_n14316);
nand_1 g13940(new_n14316, new_n14315, new_n14317);
nand_1 g13941(new_n6213, new_n6207, new_n14318);
nand_1 g13942(new_n14318, new_n6204, new_n14319);
nand_1 g13943(n7965, n6431, new_n14320);
nand_1 g13944(n9111, n5857, new_n14321);
xnor_1 g13945(new_n14321, new_n14320, new_n14322);
nand_1 g13946(n11892, n5153, new_n14323);
nand_1 g13947(n5860, n806, new_n14324);
xnor_1 g13948(new_n14324, new_n14323, new_n14325);
nand_1 g13949(n10545, n521, new_n14326);
nand_1 g13950(n10547, n7265, new_n14327);
xnor_1 g13951(new_n14327, new_n14326, new_n14328);
xnor_1 g13952(new_n14328, new_n14325, new_n14329);
xnor_1 g13953(new_n14329, new_n14322, new_n14330);
xnor_1 g13954(new_n14330, new_n14319, new_n14331);
xnor_1 g13955(new_n14331, new_n14317, new_n14332);
xnor_1 g13956(new_n14332, new_n14314, new_n14333);
not_4  g13957(new_n5746, new_n14334);
nand_1 g13958(new_n5753, new_n14334, new_n14335);
not_4  g13959(new_n5769, new_n14336);
nand_1 g13960(new_n14336, new_n5754, new_n14337);
nand_1 g13961(new_n14337, new_n14335, new_n14338);
nor_1  g13962(new_n6159, new_n6158, new_n14339);
nor_1  g13963(new_n6167, new_n6160, new_n14340);
nor_1  g13964(new_n14340, new_n14339, new_n14341);
xnor_1 g13965(new_n14341, new_n14338, new_n14342);
xnor_1 g13966(new_n14342, new_n14333, new_n14343);
xnor_1 g13967(new_n14343, new_n14311, new_n14344);
not_4  g13968(new_n6146, new_n14345);
nand_1 g13969(new_n6178, new_n14345, new_n14346);
nand_1 g13970(new_n6183, new_n6179, new_n14347);
nand_1 g13971(new_n14347, new_n14346, new_n14348);
nand_1 g13972(new_n5729, new_n5773, new_n14349);
not_4  g13973(new_n5770, new_n14350);
nand_1 g13974(new_n5775, new_n14350, new_n14351);
nand_1 g13975(new_n14351, new_n14349, new_n14352);
not_4  g13976(new_n6152, new_n14353);
nand_1 g13977(new_n6155, new_n14353, new_n14354);
nand_1 g13978(new_n6168, new_n6156, new_n14355);
nand_1 g13979(new_n14355, new_n14354, new_n14356);
nand_1 g13980(new_n6164, new_n6163, new_n14357);
nand_1 g13981(new_n6166, new_n6161, new_n14358);
nand_1 g13982(new_n14358, new_n14357, new_n14359);
nand_1 g13983(n4499, n2558, new_n14360);
nand_1 g13984(n5305, n2512, new_n14361);
not_4  g13985(new_n14361, new_n14362);
xnor_1 g13986(new_n14362, new_n14360, new_n14363);
xnor_1 g13987(new_n14363, new_n14359, new_n14364);
nand_1 g13988(new_n6151, new_n6147, new_n14365);
nand_1 g13989(new_n14365, new_n6149, new_n14366);
not_4  g13990(new_n14366, new_n14367);
nand_1 g13991(n8476, n2347, new_n14368);
not_4  g13992(new_n14368, new_n14369);
nand_1 g13993(new_n14369, new_n14367, new_n14370);
nand_1 g13994(new_n14369, new_n6001, new_n14371);
nand_1 g13995(new_n14371, new_n14366, new_n14372);
nand_1 g13996(new_n14372, new_n14370, new_n14373);
nand_1 g13997(n2253, n1097, new_n14374);
nand_1 g13998(n5964, n3865, new_n14375);
xnor_1 g13999(new_n14375, new_n14374, new_n14376);
xnor_1 g14000(new_n14376, new_n14373, new_n14377);
xnor_1 g14001(new_n14377, new_n14364, new_n14378);
xnor_1 g14002(new_n14378, new_n14356, new_n14379);
nand_1 g14003(n10510, n2024, new_n14380);
nand_1 g14004(n11257, n2879, new_n14381);
xnor_1 g14005(new_n14381, new_n14380, new_n14382);
xnor_1 g14006(new_n14382, new_n14379, new_n14383);
xnor_1 g14007(new_n14383, new_n14352, new_n14384);
xnor_1 g14008(new_n14384, new_n14348, new_n14385);
xnor_1 g14009(new_n14385, new_n14344, new_n14386);
xnor_1 g14010(new_n14386, new_n14281, new_n14387);
not_4  g14011(new_n6230, new_n14388);
nand_1 g14012(new_n14388, new_n6184, new_n14389);
nand_1 g14013(new_n6235, new_n6231, new_n14390);
nand_1 g14014(new_n14390, new_n14389, new_n14391);
not_4  g14015(new_n5745, new_n14392);
nand_1 g14016(new_n5776, new_n14392, new_n14393);
nand_1 g14017(new_n5788, new_n5777, new_n14394);
nand_1 g14018(new_n14394, new_n14393, new_n14395);
nand_1 g14019(new_n6222, new_n6186, new_n14396);
not_4  g14020(new_n6229, new_n14397);
nand_1 g14021(new_n14397, new_n6224, new_n14398);
nand_1 g14022(new_n14398, new_n14396, new_n14399);
xnor_1 g14023(new_n14399, new_n14395, new_n14400);
xnor_1 g14024(new_n14400, new_n14391, new_n14401);
xnor_1 g14025(new_n14401, new_n14387, new_n14402);
xnor_1 g14026(new_n14402, new_n14222, new_n14403);
nand_1 g14027(new_n14403, new_n14217, new_n14404);
nand_1 g14028(new_n6239, new_n6241, new_n14405);
xnor_1 g14029(new_n14402, new_n14221, new_n14406);
nand_1 g14030(new_n14406, new_n14405, new_n14407);
nand_1 g14031(new_n14407, new_n14404, n11707);
nand_1 g14032(new_n6791, new_n6790, new_n14409);
nand_1 g14033(new_n14409, new_n6793, n11755);
not_4  g14034(new_n3921, new_n14411);
xnor_1 g14035(new_n14411, new_n3920, n11780);
xnor_1 g14036(new_n10882, new_n10881, n11919);
xnor_1 g14037(new_n10884, new_n10870, n12005);
xnor_1 g14038(new_n11347, new_n11344, n12014);
xnor_1 g14039(new_n9498, new_n9472, n12020);
xnor_1 g14040(new_n12413, new_n12381, n12076);
xnor_1 g14041(new_n12990, new_n12987, n12111);
nand_1 g14042(new_n11351, new_n11335, new_n14419);
nand_1 g14043(new_n14419, new_n11353, n12444);
nand_1 g14044(new_n6083, new_n6090, new_n14421);
nand_1 g14045(new_n14421, new_n6085, n12807);
endmodule


